.SUBCKT icecap c0
*.PININFO c0:B
.ENDS
.SUBCKT sky130_fd_io__amuxsplitv2_switch_levelshifter fbk fbk_n hold reset 
+ switch_lv switch_lv_n vgnd vpwr_hv vpwr_lv
*.PININFO hold:I reset:I switch_lv:I switch_lv_n:I fbk:O fbk_n:O vgnd:B 
*.PININFO vpwr_hv:B vpwr_lv:B
XICEnet97 net97 / icecap
XICEhold hold / icecap
XICEnet105 net105 / icecap
XICEfbk fbk / icecap
XICEfbk_n fbk_n / icecap
XICEreset reset / icecap
XICEnet109 net109 / icecap
XICEnet117 net117 / icecap
XICEswitch_lv_n switch_lv_n / icecap
XICEswitch_lv switch_lv / icecap
mI184 fbk reset vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI183 net97 vpwr_lv net109 vgnd sky130_fd_pr__nfet_05v0_nvt m=4 w=1.00 l=0.90 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI18 fbk hold net105 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI182 net105 vpwr_lv net117 vgnd sky130_fd_pr__nfet_05v0_nvt m=4 w=1.00 l=0.90 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI16 net109 switch_lv vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=4 w=1.00 l=0.15 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI15 fbk_n hold net97 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI19 net117 switch_lv_n vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=4 w=1.00 l=0.15 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI185 fbk_n fbk vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI20 fbk fbk_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__amuxsplitv2_switch_s0 hold in_lv out_h reset vccd vdda vssa 
+ vssd
*.PININFO hold:I in_lv:I reset:I out_h:O vccd:B vdda:B vssa:B vssd:B
XICEnet17 net17 / icecap
XICEout_h out_h / icecap
XICEreset reset / icecap
XICEin_lv_n in_lv_n / icecap
XICEin_lv_i in_lv_i / icecap
XICEnet13 net13 / icecap
XICEhold hold / icecap
XICEin_lv in_lv / icecap
XI0 net17 net13 hold reset in_lv_i in_lv_n vssa vdda vccd / 
+ sky130_fd_io__amuxsplitv2_switch_levelshifter
mI22 in_lv_n in_lv vssd vssd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.25 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI21 in_lv_i in_lv_n vssd vssd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.25 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI16 out_h net13 vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI20 in_lv_n in_lv vccd vccd sky130_fd_pr__pfet_01v8_hvt m=1 w=1.00 l=0.25 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI19 in_lv_i in_lv_n vccd vccd sky130_fd_pr__pfet_01v8_hvt m=1 w=1.00 l=0.25 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI15 out_h net13 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__amuxsplitv2_switch_sl hold in_lv out_h out_h_n reset vccd 
+ vdda vssa vssd vswitch
*.PININFO hold:I in_lv:I reset:I out_h:O out_h_n:O vccd:B vdda:B vssa:B vssd:B 
*.PININFO vswitch:B
XICEin_lv_i in_lv_i / icecap
XICEin_lv_n in_lv_n / icecap
XICEnet39 net39 / icecap
XICEhold hold / icecap
XICEout_h_n out_h_n / icecap
XICEout_h out_h / icecap
XICEnet48 net48 / icecap
XICEnet44 net44 / icecap
XICEin_lv in_lv / icecap
XICEnet35 net35 / icecap
XICEreset reset / icecap
mI14 out_h net44 vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI15 out_h_n net39 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI19 in_lv_i in_lv_n vccd vccd sky130_fd_pr__pfet_01v8_hvt m=1 w=1.00 l=0.25 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI20 in_lv_n in_lv vccd vccd sky130_fd_pr__pfet_01v8_hvt m=1 w=1.00 l=0.25 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI13 out_h net44 vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI16 out_h_n net39 vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI21 in_lv_i in_lv_n vssd vssd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.25 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI22 in_lv_n in_lv vssd vssd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.25 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
XI0 net39 net35 hold reset in_lv_i in_lv_n vssa vdda vccd / 
+ sky130_fd_io__amuxsplitv2_switch_levelshifter
XI1 net48 net44 hold reset in_lv_i in_lv_n vssa vswitch vccd / 
+ sky130_fd_io__amuxsplitv2_switch_levelshifter
.ENDS
* .SUBCKT s8_esd_res75only_small pad rout
* *.PININFO pad:B rout:B
* rI175 pad rout sky130_fd_pr__res_generic_po m=1 w=2 l=3.15
* .ENDS
.SUBCKT sky130_fd_io__amuxsplitv2_switch amuxbus_l amuxbus_r ngate_sl_h ngate_sr_h 
+ nmid_h pgate_sl_h_n pgate_sr_h_n vdda vssa
*.PININFO ngate_sl_h:I ngate_sr_h:I nmid_h:I pgate_sl_h_n:I pgate_sr_h_n:I 
*.PININFO amuxbus_l:B amuxbus_r:B vdda:B vssa:B
XICEpgate_sl_h_n pgate_sl_h_n / icecap
XICEpgate_sr_h_n pgate_sr_h_n / icecap
XICEnmid_h nmid_h / icecap
XICEngate_sl_h ngate_sl_h / icecap
XICEamuxbus_l amuxbus_l / icecap
XICEngate_sr_h ngate_sr_h / icecap
XICEnmid_h_s nmid_h_s / icecap
XICEamuxbus_r amuxbus_r / icecap
XICEmid mid / icecap
xI20 mid vdda condiode
xI19 vssa vdda condiode
XI18 vssa nmid_h_s / s8_esd_res75only_small
mI1 amuxbus_l ngate_sl_h mid mid sky130_fd_pr__nfet_g5v0d10v5 m=30 w=10.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI2 mid ngate_sr_h amuxbus_r mid sky130_fd_pr__nfet_g5v0d10v5 m=30 w=10.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI4 mid nmid_h nmid_h_s vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI0 mid pgate_sl_h_n amuxbus_l vdda sky130_fd_pr__pfet_g5v0d10v5 m=14 w=10.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI3 amuxbus_r pgate_sr_h_n mid vdda sky130_fd_pr__pfet_g5v0d10v5 m=14 w=10.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
* .SUBCKT sky130_fd_io__hvsbt_nand2 in0 in1 out vgnd vpwr
* *.PININFO in0:I in1:I vgnd:I vpwr:I out:O
* XICEout out / icecap
* XICEin0 in0 / icecap
* XICEin1 in1 / icecap
* mI3 out in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI5 out in1 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI1 out in1 net25 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI6 net25 in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
.SUBCKT sky130_fd_io__amuxsplitv2_delay enable_vdda_h hld_vdda_h_n hold reset 
+ vcc_io vgnd
*.PININFO enable_vdda_h:I hld_vdda_h_n:I hold:O reset:O vcc_io:B vgnd:B
XICEhold hold / icecap
XICEhld_vdda_h hld_vdda_h / icecap
XICEreset reset / icecap
XICEenable_vdda_h_n enable_vdda_h_n / icecap
XICEenable_vdda_h enable_vdda_h / icecap
XICEhld_vdda_h_n_switch hld_vdda_h_n_switch / icecap
XICEhld_vdda_h_n hld_vdda_h_n / icecap
XICEenable_vdda_switch enable_vdda_switch / icecap
XI33 enable_vdda_switch hld_vdda_h_n_switch reset vgnd vcc_io / 
+ sky130_fd_io__hvsbt_nand2
mI29 hld_vdda_h_n_switch hld_vdda_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.60 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI28 hld_vdda_h hld_vdda_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI12 enable_vdda_switch enable_vdda_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.60 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI13 enable_vdda_h_n enable_vdda_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI36 hold reset vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI31 hld_vdda_h_n_switch hld_vdda_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.60 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI30 hld_vdda_h hld_vdda_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI14 enable_vdda_switch enable_vdda_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.60 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI15 enable_vdda_h_n enable_vdda_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI37 hold reset vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__top_amuxsplitv2 amuxbus_a_l amuxbus_a_r amuxbus_b_l 
+ amuxbus_b_r enable_vdda_h hld_vdda_h_n switch_aa_s0 switch_aa_sl 
+ switch_aa_sr switch_bb_s0 switch_bb_sl switch_bb_sr vccd vcchib vdda vddio 
+ vddio_q vssa vssd vssio vssio_q vswitch
*.PININFO enable_vdda_h:I hld_vdda_h_n:I switch_aa_s0:I switch_aa_sl:I 
*.PININFO switch_aa_sr:I switch_bb_s0:I switch_bb_sl:I switch_bb_sr:I 
*.PININFO amuxbus_a_l:B amuxbus_a_r:B amuxbus_b_l:B amuxbus_b_r:B vccd:B 
*.PININFO vcchib:B vdda:B vddio:B vddio_q:B vssa:B vssd:B vssio:B vssio_q:B 
*.PININFO vswitch:B
xI22 vssa vdda condiode
XI18 hold switch_aa_s0 ng_vdda_aa_s0_h reset vccd vdda vssa vssd / 
+ sky130_fd_io__amuxsplitv2_switch_s0
XI348 hold switch_bb_s0 ng_vdda_bb_s0_h reset vccd vdda vssa vssd / 
+ sky130_fd_io__amuxsplitv2_switch_s0
XI347 hold switch_aa_sl ng_vswitch_aa_sl_h pg_vdda_aa_sl_h_n reset vccd vdda 
+ vssa vssd vswitch / sky130_fd_io__amuxsplitv2_switch_sl
XI24 hold switch_aa_sr ng_vswitch_aa_sr_h pg_vdda_aa_sr_h_n reset vccd vdda 
+ vssa vssd vswitch / sky130_fd_io__amuxsplitv2_switch_sl
XI349 hold switch_bb_sr ng_vswitch_bb_sr_h pg_vdda_bb_sr_h_n reset vccd vdda 
+ vssa vssd vswitch / sky130_fd_io__amuxsplitv2_switch_sl
XI350 hold switch_bb_sl ng_vswitch_bb_sl_h pg_vdda_bb_sl_h_n reset vccd vdda 
+ vssa vssd vswitch / sky130_fd_io__amuxsplitv2_switch_sl
XI6 amuxbus_a_l amuxbus_a_r ng_vswitch_aa_sl_h ng_vswitch_aa_sr_h 
+ ng_vdda_aa_s0_h pg_vdda_aa_sl_h_n pg_vdda_aa_sr_h_n vdda vssa / 
+ sky130_fd_io__amuxsplitv2_switch
XI8 amuxbus_b_l amuxbus_b_r ng_vswitch_bb_sl_h ng_vswitch_bb_sr_h 
+ ng_vdda_bb_s0_h pg_vdda_bb_sl_h_n pg_vdda_bb_sr_h_n vdda vssa / 
+ sky130_fd_io__amuxsplitv2_switch
XI342 enable_vdda_h hld_vdda_h_n hold reset vdda vssa / 
+ sky130_fd_io__amuxsplitv2_delay
XICEnet27 enable_vdda_h / icecap
XICEamuxbus_b_r amuxbus_b_r / icecap
XICEswitch_aa_sl_h ng_vswitch_aa_sl_h / icecap
XICEamuxbus_a_l amuxbus_a_l / icecap
XICEswitch_bb_sl_h_n pg_vdda_bb_sl_h_n / icecap
XICEswitch_bb_sr_h ng_vswitch_bb_sr_h / icecap
XICEswitch_aa_s0_h ng_vdda_aa_s0_h / icecap
XICEswitch_aa_s0 hold / icecap
XICEswitch_aa_sr_h ng_vswitch_aa_sr_h / icecap
XICEswitch_aa_sl_h_n pg_vdda_aa_sl_h_n / icecap
XICEswitch_bb_sl_h ng_vswitch_bb_sl_h / icecap
XICEswitch_bb_s0_h ng_vdda_bb_s0_h / icecap
XICEswitch_bb_sr_h_n pg_vdda_bb_sr_h_n / icecap
XICEswitch_aa_sr_h_n pg_vdda_aa_sr_h_n / icecap
XI355 hold / icecap
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_nonoverlap_leak_fix p1g p1gb p2g padlo 
+ vgnd vpwr
*.PININFO padlo:I vgnd:I vpwr:I p1g:O p1gb:O p2g:O
XICEpadlo_bar padlo_bar / icecap
XICEp2gb p2gb / icecap
XICEp1gb p1gb / icecap
XICEp2g p2g / icecap
XICEp1g_new p1g_new / icecap
XICEp1g p1g / icecap
XICEpadlo padlo / icecap
XICEp2g_new p2g_new / icecap
mI76 p1g p1gb vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI64 p1g_new padlo vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=1.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI53 padlo_bar padlo vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI50 p2g_new p1g_new vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=1.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI49 p2g_new padlo_bar vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=1.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI65 p1g_new p2g_new vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=1.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI77 p2g p2gb vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI70 p2gb p2g_new vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI72 p1gb p1g_new vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI54 padlo_bar padlo vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI69 p1g_new padlo net140 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=4.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI78 p2g p2gb vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=0.42 l=2.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI67 net140 p2g_new vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=8.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI71 p2gb p2g_new vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI79 p1g p1gb vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=2.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI51 p2g_new padlo_bar net124 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=4.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI73 p1gb p1g_new vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI52 net124 p1g_new vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=8.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_pug_ovtfix padlo pug4_h pug7_h tie_hi 
+ vpb_drvr
*.PININFO padlo:I tie_hi:I vpb_drvr:I pug4_h:O pug7_h:O
mI52 pug4_h padlo tie_hi vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.50 sa=1.825 
+ sb=1.825 sd=280e-3 topography=normal perim=1.14
mI53 pug7_h padlo tie_hi vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__sio_hvsbt_nand2 in0 in1 out vgnd vnb vpb vpwr
*.PININFO in0:I in1:I vgnd:I vnb:I vpb:I vpwr:I out:O
XICEout out / icecap
XICEin1 in1 / icecap
XICEin0 in0 / icecap
mI3 out in0 vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI5 out in1 vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI1 out in1 net25 vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI6 net25 in0 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__sio_hvsbt_inv_x1 in out vgnd vnb vpb vpwr
*.PININFO in:I vgnd:I vnb:I vpb:I vpwr:I out:O
XICEout out / icecap
XICEin in / icecap
mI2 out in vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal perim=1.14
mI1 out in vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__sio_hvsbt_nor in0 in1 out vgnd vnb vpb vpwr
*.PININFO in0:I in1:I vgnd:I vnb:I vpb:I vpwr:I out:O
XICEin0 in0 / icecap
XICEin1 in1 / icecap
XICEout out / icecap
mI3 net17 in0 vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI12 out in1 net17 vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI1 out in0 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI6 out in1 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
* .SUBCKT sky130_fd_io__tk_em1o a b
* *.PININFO a:B b:B
* rI1 a net11 short
* rI2 b net7 short
* .ENDS
* .SUBCKT sky130_fd_io__tk_em1s a b
* *.PININFO a:B b:B
* rI1 a net8 short
* rI2 b net8 short
* .ENDS
.SUBCKT sky130_fd_io__sio_hotswap_dly in out out_n vcc_io vgnd
*.PININFO in:I vcc_io:I vgnd:I out:O out_n:O
XICEa5 a5 / icecap
XICEa3 a3 / icecap
XICEout out / icecap
XICEa2 a2 / icecap
XICEa7 a7 / icecap
XICEout_n out_n / icecap
XICEa4 a4 / icecap
XICEa6 a6 / icecap
XICEa1 a1 / icecap
XICEin in / icecap
XI228 out_n a5 / sky130_fd_io__tk_em1o
XI229 out_n a7 / sky130_fd_io__tk_em1o
XI227 a6 out / sky130_fd_io__tk_em1o
XI214 out_n a1 / sky130_fd_io__tk_em1o
XI215 a2 out / sky130_fd_io__tk_em1o
XEdly0 in out / sky130_fd_io__tk_em1o
XI217 out_n a3 / sky130_fd_io__tk_em1s
XEdly2 a4 out / sky130_fd_io__tk_em1s
mI196 a1 in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI204 a4 a3 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI199 a2 a1 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI198 a3 a2 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI232 a5 a4 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI231 a6 a5 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI230 a7 a6 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI197 a1 in vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI202 a4 a3 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI201 a2 a1 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI200 a3 a2 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI235 a5 a4 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI234 a6 a5 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI233 a7 a6 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__sio_hotswap_log_i2c_fix dishs_h dishs_h_n en_h enhs_h 
+ enhs_h_n enhs_lat_h_n exiths_h forcehi_h<1> od_i_h_n vcc_io vgnd
*.PININFO en_h:I enhs_lat_h_n:I forcehi_h<1>:I od_i_h_n:I vcc_io:I vgnd:I 
*.PININFO dishs_h:O dishs_h_n:O enhs_h:O enhs_h_n:O exiths_h:O
XICEdishs_h_n dishs_h_n / icecap
XICEnet39 net39 / icecap
XICEdishs_h dishs_h / icecap
XICEnet74 net74 / icecap
XICEod_i_h_n od_i_h_n / icecap
XICEen_h en_h / icecap
XICEenhs_dly_h_n enhs_dly_h_n / icecap
XICEenhs_h_n enhs_h_n / icecap
XICEnet46 net46 / icecap
XICEnet80 net80 / icecap
XICEforcehi_h<1> forcehi_h<1> / icecap
XICEenhs_dly_h enhs_dly_h / icecap
XICEexiths_h exiths_h / icecap
XICEenhs_lat_h_n enhs_lat_h_n / icecap
XICEenhs_h enhs_h / icecap
XI664 net39 net46 dishs_h vgnd vgnd vcc_io vcc_io / sky130_fd_io__sio_hvsbt_nand2
XI663 net80 forcehi_h<1> net46 vgnd vgnd vcc_io vcc_io / 
+ sky130_fd_io__sio_hvsbt_nand2
XI662 od_i_h_n en_h net39 vgnd vgnd vcc_io vcc_io / sky130_fd_io__sio_hvsbt_nand2
XI658 od_i_h_n net80 vgnd vgnd vcc_io vcc_io / sky130_fd_io__sio_hvsbt_inv_x1
XI666 enhs_lat_h_n net74 vgnd vgnd vcc_io vcc_io / sky130_fd_io__sio_hvsbt_inv_x1
XI565 net74 enhs_h_n vgnd vgnd vcc_io vcc_io / sky130_fd_io__sio_hvsbt_inv_x1
XI667 dishs_h dishs_h_n vgnd vgnd vcc_io vcc_io / sky130_fd_io__sio_hvsbt_inv_x1
XI637 enhs_h_n enhs_h vgnd vgnd vcc_io vcc_io / sky130_fd_io__sio_hvsbt_inv_x1
XI553 net74 enhs_dly_h_n exiths_h vgnd vgnd vcc_io vcc_io / 
+ sky130_fd_io__sio_hvsbt_nor
XI521 net74 enhs_dly_h enhs_dly_h_n vcc_io vgnd / sky130_fd_io__sio_hotswap_dly
.ENDS
.SUBCKT sky130_fd_io__sio_hotswap_hys in out vcc_io vgnd
*.PININFO in:I vcc_io:I vgnd:I out:O
XICEvcc_io_buf vcc_io_buf / icecap
XICEout out / icecap
XICEvgnd_buf vgnd_buf / icecap
XICEin in / icecap
XICEint_p int_p / icecap
XICEint_n int_n / icecap
mI650 vcc_io_buf out int_n vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI649 int_n in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI648 out in int_n vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=0.42 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI655 vgnd_buf vcc_io vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI647 vgnd_buf out int_p vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI656 vcc_io_buf vgnd vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI646 out in int_p vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI645 int_p in vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__sio_hotswap_pghspd in1 in2 out vgnd
*.PININFO in1:I in2:I vgnd:I out:O
XICEin2 in2 / icecap
XICEnet25 net25 / icecap
XICEnet34 net34 / icecap
XICEnet27 net27 / icecap
XICEnet30 net30 / icecap
XICEnet42 net42 / icecap
XICEin1 in1 / icecap
XICEout out / icecap
XICEnet38 net38 / icecap
XEin2b vgnd net25 / sky130_fd_io__tk_em1o
XEoutb net38 out / sky130_fd_io__tk_em1o
XEin1b vgnd net27 / sky130_fd_io__tk_em1o
XEin1a in1 net27 / sky130_fd_io__tk_em1s
XEouta net42 out / sky130_fd_io__tk_em1s
XEin2a in2 net25 / sky130_fd_io__tk_em1s
mI481 net50 in2 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI507 out in1 net50 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI651 net42 net27 net34 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=6 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI654 net38 net27 net30 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI652 net34 net25 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=6 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI653 net30 net25 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__sio_hotswap_wpd en out vgnd
*.PININFO en:I vgnd:I out:O
XICEout out / icecap
XICEnpd<17> sky130_fd_pr__special_nfet_latch<17> / icecap
XICEen en / icecap
XICEnpd<14> sky130_fd_pr__special_nfet_latch<14> / icecap
XICEnpd<15> sky130_fd_pr__special_nfet_latch<15> / icecap
XICEnpd<18> sky130_fd_pr__special_nfet_latch<18> / icecap
XICEnpd<16> sky130_fd_pr__special_nfet_latch<16> / icecap
XI198 sky130_fd_pr__special_nfet_latch<15> sky130_fd_pr__special_nfet_latch<16> / sky130_fd_io__tk_em1o
XI209 vgnd sky130_fd_pr__special_nfet_latch<14> / sky130_fd_io__tk_em1o
XI196 sky130_fd_pr__special_nfet_latch<17> sky130_fd_pr__special_nfet_latch<18> / sky130_fd_io__tk_em1o
XI197 sky130_fd_pr__special_nfet_latch<16> sky130_fd_pr__special_nfet_latch<17> / sky130_fd_io__tk_em1o
XE20 sky130_fd_pr__special_nfet_latch<18> out / sky130_fd_io__tk_em1o
XI208 sky130_fd_pr__special_nfet_latch<14> sky130_fd_pr__special_nfet_latch<15> / sky130_fd_io__tk_em1o
mnen17 sky130_fd_pr__special_nfet_latch<17> en sky130_fd_pr__special_nfet_latch<16> vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mnen15 sky130_fd_pr__special_nfet_latch<15> en sky130_fd_pr__special_nfet_latch<14> vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mnen14 sky130_fd_pr__special_nfet_latch<14> en vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mnen16 sky130_fd_pr__special_nfet_latch<16> en sky130_fd_pr__special_nfet_latch<15> vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mnen19 out en sky130_fd_pr__special_nfet_latch<18> vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mnen18 sky130_fd_pr__special_nfet_latch<18> en sky130_fd_pr__special_nfet_latch<17> vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_latch dishs_h dishs_h_n enhs_h enhs_h_n 
+ enhs_lat_h_n enhs_lathys_h_n exiths_h p3out pad_esd pghs_h vcc_io vgnd 
+ vpb_drvr vpwr_ka
*.PININFO dishs_h:I dishs_h_n:I enhs_h:I enhs_h_n:I exiths_h:I pad_esd:I 
*.PININFO vcc_io:I vgnd:I vpb_drvr:I vpwr_ka:I enhs_lat_h_n:O 
*.PININFO enhs_lathys_h_n:O p3out:O pghs_h:B
XI660 vgnd net102 vgnd vgnd vcc_io vcc_io / sky130_fd_io__sio_hvsbt_inv_x1
XI528 n6 net96 vgnd vgnd vcc_io vcc_io / sky130_fd_io__sio_hvsbt_inv_x1
XEhys2 enhs_lathys_h_n enhs_lat_h_n / sky130_fd_io__tk_em1o
XI658 net96 enhs_lat_h_n / sky130_fd_io__tk_em1s
XEhys1 net117 enhs_lathys_h_n / sky130_fd_io__tk_em1s
Xhys n6 net117 vcc_io vgnd / sky130_fd_io__sio_hotswap_hys
Xpghspd enhs_h n2 pghs_h vgnd / sky130_fd_io__sio_hotswap_pghspd
Xwpdenhs vpwr_ka net127 vgnd / sky130_fd_io__sio_hotswap_wpd
Xwpdexhs vpwr_ka net124 vgnd / sky130_fd_io__sio_hotswap_wpd
mI502 net186 pghs_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI484 net161 enhs_h pghs_h vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI491 n5 n6 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI498 n2 n6 net124 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI500 net170 enhs_h_n n2 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mnexiths pghs_h exiths_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI485 n3 n2 net161 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI499 n4 pghs_h net170 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI497 n6 n5 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mndishs pghs_h dishs_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI508 n2 enhs_h_n net186 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI696 vgnd exiths_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI487 pghs_h n5 net127 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI697 vgnd dishs_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI492 n5 n6 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI503 n4 vgnd vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=2.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI488 n3 vgnd vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=2.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI505 n6 n5 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI493 n5 n3 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI323 n2 dishs_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI279 n2 pad_esd vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI504 n6 n4 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI689 p3out pad_esd vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=12 w=10.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_ctl_i2c_fix en_h enhs_lat_h_n forcehi_h<1> 
+ od_i_h_n p3out pad_esd pghs_h vddio vpb_drvr vpwr_ka vssd
*.PININFO en_h:I forcehi_h<1>:I od_i_h_n:I pad_esd:I vddio:I vpb_drvr:I 
*.PININFO vpwr_ka:I vssd:I enhs_lat_h_n:O p3out:O pghs_h:B
XICEvpb_drvr vpb_drvr / icecap
XICEpghs_h pghs_h / icecap
XICEforcehi_h<1> forcehi_h<1> / icecap
XICEdishs_h dishs_h / icecap
XICEdishs_h_n dishs_h_n / icecap
XICEpad_esd pad_esd / icecap
XICEenhs_lathys_h_n enhs_lathys_h_n / icecap
XICEp3out p3out / icecap
XICEen_h en_h / icecap
XICEenhs_h_n enhs_h_n / icecap
XICEod_i_h_n od_i_h_n / icecap
XICEenhs_h enhs_h / icecap
XICEenhs_lat_h_n enhs_lat_h_n / icecap
XICEexiths_h exiths_h / icecap
Xhslog dishs_h dishs_h_n en_h enhs_h enhs_h_n enhs_lathys_h_n exiths_h 
+ forcehi_h<1> od_i_h_n vddio vssd / sky130_fd_io__sio_hotswap_log_i2c_fix
Xhslatch dishs_h dishs_h_n enhs_h enhs_h_n enhs_lat_h_n enhs_lathys_h_n 
+ exiths_h p3out pad_esd pghs_h vddio vssd vpb_drvr vpwr_ka / 
+ sky130_fd_io__gpio_ovtv2_hotswap_latch
.ENDS
.SUBCKT sky130_fd_io__sio_tk_em1s a b
*.PININFO a:B b:B
rI1 a net8 short
rI2 b net8 short
.ENDS
.SUBCKT sky130_fd_io__sio_tk_em1o a b
*.PININFO a:B b:B
rI1 a net11 short
rI2 b net7 short
.ENDS
.SUBCKT sky130_fd_io__sio_hvsbt_inv_x4 in out vgnd vnb vpb vpwr
*.PININFO in:I vgnd:I vnb:I vpb:I vpwr:I out:O
XICEout out / icecap
XICEin in / icecap
mI2 out in vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=4 w=1.00 l=0.60 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal perim=1.14
mI1 out in vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.00 l=0.60 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_pghspu pad pghs_h pghs_h_latch tie_hi 
+ vcc_io_soft vpb_drvr
*.PININFO pad:I tie_hi:I vcc_io_soft:I vpb_drvr:I pghs_h:O pghs_h_latch:O
XEg9 tie_hi pg8 / sky130_fd_io__sio_tk_em1o
XEg2 pg2 vcc_io_soft / sky130_fd_io__sio_tk_em1s
XEg5 pg6 pg4 / sky130_fd_io__sio_tk_em1s
XEg4 pg4 pg3 / sky130_fd_io__sio_tk_em1s
XEpghs3 padhi3 pghs_h_latch / sky130_fd_io__sio_tk_em1s
XEg3 pg3 pg2 / sky130_fd_io__sio_tk_em1s
XEpghs7 padhi7 net36 / sky130_fd_io__sio_tk_em1s
XEg7 pg7 pg6 / sky130_fd_io__sio_tk_em1s
XEg8 pg8 pg7 / sky130_fd_io__sio_tk_em1s
XEpghs2 padhi2 padhi3 / sky130_fd_io__sio_tk_em1s
XEpghs8 pghs_h padhi7 / sky130_fd_io__sio_tk_em1s
XICEpg2 pg2 / icecap
XICEpadhi7 padhi7 / icecap
XICEpg3 pg3 / icecap
XICEpadhi6 net36 / icecap
XICEpg7 pg7 / icecap
XICEpadhi4 pghs_h_latch / icecap
XICEpg8 pg8 / icecap
XICEpg4 pg4 / icecap
XICEpadhi3 padhi3 / icecap
XICEpadhi2 padhi2 / icecap
XICEpadhi8 pghs_h / icecap
XICEpg5 pg6 / icecap
XICEtie_hi tie_hi / icecap
mpghs8 pghs_h pg8 pad vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=20.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mpghs2 padhi2 pg2 pad vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=20.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mpghs3 padhi3 pg3 pad vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=20.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mpghs6 net36 pg6 pad vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mpghs4 pghs_h_latch pg4 pad vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mpghs7 padhi7 pg7 pad vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=20.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
* .SUBCKT s8_esd_signal_5_sym_hv_local_5term gate in nbody nwellRing vgnd
* *.PININFO gate:I in:B nbody:B nwellRing:B vgnd:B
* mI1 in gate vgnd nbody sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=5.40 l=0.60 sa=0.0 sb=0.0 sd=0.0 
* + topography=normal perim=0.94
* rI9 net18 nbody short
* rI8 net16 nwellRing short
* .ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_pghs_i2c_fix en_h force_h<1> od_i_h_n 
+ p3out pad padlo pghs_h tie_hi vcc_io_soft vddio vpb_drvr vpwr_ka vssd
*.PININFO en_h:I force_h<1>:I od_i_h_n:I pad:I tie_hi:I vcc_io_soft:I vddio:I 
*.PININFO vpb_drvr:I vpwr_ka:I vssd:I p3out:O padlo:O pghs_h:O
XICEtie_hi tie_hi / icecap
XICEen_h en_h / icecap
XICEenhs_latbuf_h_n enhs_latbuf_h_n / icecap
XICEpad pad / icecap
XICEvpb_drvr vpb_drvr / icecap
XICEp3out p3out / icecap
XICEenhs_lat_h enhs_lat_h / icecap
XICEnet54 net54 / icecap
XICEforce_h<1> force_h<1> / icecap
XICEvcc_io_soft vcc_io_soft / icecap
XICEod_i_h_n od_i_h_n / icecap
XICEenhs_lat_h_n enhs_lat_h_n / icecap
XICEnet50 net50 / icecap
XICEpadlo padlo / icecap
XICEpghs_h pghs_h / icecap
Xhsctl en_h enhs_lat_h_n force_h<1> od_i_h_n p3out pad net50 vddio vpb_drvr 
+ vpwr_ka vssd / sky130_fd_io__gpio_ovtv2_hotswap_ctl_i2c_fix
XI3 enhs_latbuf_h_n padlo / sky130_fd_io__sio_tk_em1s
XEpghs12 pghs_h net54 / sky130_fd_io__sio_tk_em1o
XI2 enhs_lat_h enhs_latbuf_h_n vssd vssd vddio vddio / 
+ sky130_fd_io__sio_hvsbt_inv_x4
XI1 enhs_lat_h_n enhs_lat_h vssd vssd vddio vddio / sky130_fd_io__sio_hvsbt_inv_x1
Xpghspu pad pghs_h net50 tie_hi vcc_io_soft vpb_drvr / 
+ sky130_fd_io__gpio_ovtv2_hotswap_pghspu
Xclamp vssd vddio vssd vddio pad / s8_esd_signal_5_sym_hv_local_5term
mpghs12 net54 padlo vpb_drvr vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__sio_tk_tie_r_out_esd a b
*.PININFO a:B b:B
resd_r a b sky130_fd_pr__res_generic_po m=1 w=0.5 l=10.2
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_pug pad padlo pug_h tie_hi vpb_drvr
*.PININFO pad:I padlo:I tie_hi:I vpb_drvr:I pug_h:O
XEg1 padlo net22 / sky130_fd_io__sio_tk_em1s
XI65 net24 tie_hi / sky130_fd_io__sio_tk_em1s
XEs2 net26 tie_hi / sky130_fd_io__sio_tk_em1s
XEs1 pad net26 / sky130_fd_io__sio_tk_em1o
XEg2 net22 net24 / sky130_fd_io__sio_tk_em1o
mI52 pug_h net22 net26 vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.50 sa=1.825 sb=1.825 
+ sd=280e-3 topography=normal perim=1.14
mI53 pug_h net24 net26 vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_bias pswg_h vcc_io vpb_drvr
*.PININFO pswg_h:I vcc_io:I vpb_drvr:O
XICEvpb_drvr vpb_drvr / icecap
XICEpswg_h pswg_h / icecap
mpsw_vccio vpb_drvr pswg_h vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=22 w=15.0 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI36 vpb_drvr pswg_h vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=9 w=10.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit pb pd pgin ps
*.PININFO pb:I pgin:I pd:B ps:B
XICEpd pd / icecap
XICEnet15 pgin / icecap
XICEpgin pgin / icecap
mpdrv pd pgin ps pb sky130_fd_pr__esd_pfet_g5v0d10v5 m=2 w=15.50 l=0.55 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias p2g pad soft_vcc_io tie_hi 
+ vpb_drvr
*.PININFO p2g:I pad:I soft_vcc_io:I tie_hi:I vpb_drvr:B
XICEsoft_vcc_io soft_vcc_io / icecap
XICEp2g p2g / icecap
XICEtie_hi tie_hi / icecap
Xpsw_pad4 vpb_drvr vpb_drvr p2g pad / sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
Xpsw_pad0 vpb_drvr vpb_drvr p2g pad / sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
Xpsw_pad3 vpb_drvr vpb_drvr p2g pad / sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
Xpsw_pad2 vpb_drvr vpb_drvr p2g pad / sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
Xpsw_pad5 vpb_drvr vpb_drvr soft_vcc_io pad / 
+ sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
Xpsw_pad1 vpb_drvr vpb_drvr p2g pad / sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
XI5 tie_hi soft_vcc_io / sky130_fd_io__tk_em1o
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_i2c_fix_leak_fix force_h<1> nghs_h 
+ od_i_h_n oe_hs_h p2g pad pad_esd pghs_h pug_h<7> pug_h<6> pug_h<5> pug_h<4> 
+ pug_h<3> pug_h<2> pug_h<1> pug_h<0> vcc_io_soft vddio vpb_drvr vpwr_ka vssd
*.PININFO force_h<1>:I od_i_h_n:I oe_hs_h:I pad:I pad_esd:I vddio:I vpwr_ka:I 
*.PININFO vssd:I nghs_h:O p2g:O pghs_h:O vcc_io_soft:O vpb_drvr:O pug_h<7>:B 
*.PININFO pug_h<6>:B pug_h<5>:B pug_h<4>:B pug_h<3>:B pug_h<2>:B pug_h<1>:B 
*.PININFO pug_h<0>:B
Xnon_overlap p1g nghs_h p2g padlo vssd vpb_drvr / 
+ sky130_fd_io__gpio_ovtv2_hotswap_nonoverlap_leak_fix
Xpug47 padlo pug_h<4> pug_h<7> tie_hi vpb_drvr / 
+ sky130_fd_io__gpio_ovtv2_hotswap_pug_ovtfix
Xpghs oe_hs_h force_h<1> od_i_h_n net74 pad_esd padlo p1g tie_hi vcc_io_soft 
+ vddio vpb_drvr vpwr_ka vssd / sky130_fd_io__gpio_ovtv2_hotswap_pghs_i2c_fix
Xresd_tiehi vpb_drvr tie_hi / sky130_fd_io__sio_tk_tie_r_out_esd
Xresd_vccio vddio vcc_io_soft / sky130_fd_io__sio_tk_tie_r_out_esd
Xpug<3> pad_esd padlo pug_h<3> tie_hi vpb_drvr / 
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xpug<2> pad_esd padlo pug_h<2> tie_hi vpb_drvr / 
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xpug<1> pad_esd padlo pug_h<1> tie_hi vpb_drvr / 
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xpug<0> pad_esd padlo pug_h<0> tie_hi vpb_drvr / 
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xpug<6> pad_esd padlo pug_h<6> tie_hi vpb_drvr / 
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xpug<5> pad_esd padlo pug_h<5> tie_hi vpb_drvr / 
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xp1_bias p1g vddio vpb_drvr / sky130_fd_io__gpio_ovtv2_hotswap_bias
Xp2p4_bias p2g pad vcc_io_soft vcc_io_soft vpb_drvr / 
+ sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias
XICEnet84 vpb_drvr / icecap
XICEnet135 vpb_drvr / icecap
XICEod_h od_i_h_n / icecap
XICEp1g p1g / icecap
XICEnet89 vpb_drvr / icecap
XICEp2g p2g / icecap
XICEoe_hs_h oe_hs_h / icecap
XICEnet136 vpb_drvr / icecap
XICEnet148 tie_hi / icecap
XICEnet152 padlo / icecap
XICEforce_h<1> force_h<1> / icecap
XICEpadlo padlo / icecap
XICEnet149 p1g / icecap
XICEvcc_io_soft vcc_io_soft / icecap
XICEnet142 vpb_drvr / icecap
XICEtie_hi tie_hi / icecap
XICEvpb_drvr vpb_drvr / icecap
rI26 p2g net137 short
rI39 p2g net74 short
rI49 pghs_h p1g short
.ENDS
* .SUBCKT sky130_fd_io__com_pad pad vgnd_io
* *.PININFO pad:B vgnd_io:B
* XICEpad pad / icecap
* .ENDS
* .SUBCKT sky130_fd_io__gpio_pddrvr_strong_slow pad pd_h vcc_io vgnd_io
* *.PININFO pd_h:I vcc_io:I vgnd_io:I pad:O
* XICEpd_h pd_h / icecap
* XICEpad pad / icecap
* XICEvcc_io vcc_io / icecap
* mndrv pad pd_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpio_pddrvr_weak pad pd_h vcc_io vgnd_io
* *.PININFO pd_h:I vcc_io:I vgnd_io:I pad:O
* XICEvcc_io vcc_io / icecap
* XICEpd_h pd_h / icecap
* XICEpad pad / icecap
* mndrv1 pad pd_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=6 w=5.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__com_res_strong_slow ra rb vgnd_io
* *.PININFO vgnd_io:I ra:B rb:B
* XICErb rb / icecap
* XICEnet30 net30 / icecap
* XICEra ra / icecap
* XICEnet34 net34 / icecap
* XI28 net34 net30 / sky130_fd_io__tk_em1s
* rI32 rb net30 sky130_fd_pr__res_generic_po m=1 w=2 l=2
* rI29 net30 net34 sky130_fd_pr__res_generic_po m=1 w=2 l=3
* rr1 net34 ra sky130_fd_pr__res_generic_po m=1 w=2 l=5
* .ENDS
* .SUBCKT sky130_fd_io__com_res_weak ra rb vgnd_io
* *.PININFO vgnd_io:I ra:B rb:B
* XICEn<3> n<3> / icecap
* XICEn<2> n<2> / icecap
* XICErb rb / icecap
* XICEn<0> n<0> / icecap
* XICEn<4> n<4> / icecap
* XICEra ra / icecap
* XICEnet64 net64 / icecap
* XICEn<1> n<1> / icecap
* XICEn<5> n<5> / icecap
* Xe9 n<0> n<1> / sky130_fd_io__tk_em1s
* Xe11 n<2> n<3> / sky130_fd_io__tk_em1s
* Xe10 n<1> n<2> / sky130_fd_io__tk_em1s
* Xe12 n<3> rb / sky130_fd_io__tk_em1s
* Xe13 n<4> n<0> / sky130_fd_io__tk_em1s
* Xe14 n<5> n<4> / sky130_fd_io__tk_em1o
* rI84 n<0> n<1> sky130_fd_pr__res_generic_po m=1 w=0.8 l=1.5
* rI62 n<3> rb sky130_fd_pr__res_generic_po m=1 w=0.8 l=1.5
* rI82 n<2> n<3> sky130_fd_pr__res_generic_po m=1 w=0.8 l=1.5
* rI85 ra net64 sky130_fd_pr__res_generic_po m=1 w=0.8 l=50
* rI83 n<1> n<2> sky130_fd_pr__res_generic_po m=1 w=0.8 l=1.5
* rI116 net64 n<5> sky130_fd_pr__res_generic_po m=1 w=0.8 l=12
* rI104 n<4> n<0> sky130_fd_pr__res_generic_po m=1 w=0.8 l=6
* rI134 n<5> n<4> sky130_fd_pr__res_generic_po m=1 w=0.8 l=6
* .ENDS
* .SUBCKT sky130_fd_io__tk_tie_r_out_esd a b
* *.PININFO a:B b:B
* resd_r a b sky130_fd_pr__res_generic_po m=1 w=0.5 l=10.2
* .ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pddrvr_unit nd ngin ns
*.PININFO ngin:I nd:B ns:B
XICEngin ngin / icecap
XICEnet13 ngin / icecap
XICEnd nd / icecap
mndrv nd ngin ns ns sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=40.31 l=0.55 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pddrvr pad pd_csd pd_h<3> pd_h<2> tie_lo_esd vddio 
+ vssio vssio_q
*.PININFO pd_csd:I pd_h<3>:I pd_h<2>:I tie_lo_esd:O pad:B vddio:B vssio:B 
*.PININFO vssio_q:B
XICEpd_csd pd_csd / icecap
XICEpd_h<2> pd_h<2> / icecap
XICEpd_h<3> pd_h<3> / icecap
XICEpad pad / icecap
XICEtie_lo_esd tie_lo_esd / icecap
XICEvssio_q vssio_q / icecap
XI26 vssio tie_lo_esd / sky130_fd_io__tk_tie_r_out_esd
Xn1 pad pd_h<2> vssio / sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn2 pad pd_h<2> vssio / sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn3 pad pd_h<2> vssio / sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn8 pad pd_h<3> vssio / sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn7 pad pd_h<3> vssio / sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn6 pad pd_h<3> vssio / sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn5 pad pd_h<3> vssio / sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn9 pad pd_h<3> vssio / sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn10 pad pd_h<3> vssio / sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn11 pad pd_h<3> vssio / sky130_fd_io__gpio_ovtv2_pddrvr_unit
rI8 vddio net96 short
mn14 pad pd_csd vssio_q vssio_q sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=40.31 l=0.55 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mn13 pad pd_csd vssio_q vssio_q sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=40.31 l=0.55 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
xI9 vssio vddio condiode
xI62 vssio_q vddio condiode
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pudrvr_weak nghs_h pad pghs_h pu_h_n pug_h vddio 
+ vpb_drvr vssd vssio
*.PININFO nghs_h:I pghs_h:I pu_h_n:I vddio:I vpb_drvr:I vssd:I vssio:I pad:B 
*.PININFO pug_h:B
XICEnet26 net26 / icecap
XICEpghs_h pghs_h / icecap
XICEnghs_h nghs_h / icecap
XICEpad pad / icecap
XICEpug_h pug_h / icecap
XICEpu_h_n pu_h_n / icecap
XI36 pad net26 / sky130_fd_io__tk_em1o
mI51 pug_h nghs_h pu_h_n vssio sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI50 pu_h_n pghs_h pug_h vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mpdrv pad pug_h vddio vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=3 w=10.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI35 net26 pug_h vddio vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=10.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI29 pad pug_h vddio vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=10.0 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pudrvr_strong_slow nghs_h pad pghs_h pu_h_n pug_h 
+ vddio vpb_drvr vssd vssio
*.PININFO nghs_h:I pghs_h:I pu_h_n:I vddio:I vpb_drvr:I vssd:I vssio:I pad:B 
*.PININFO pug_h:B
XICEvssio vssio / icecap
XICEpghs_h pghs_h / icecap
XICEnghs_h nghs_h / icecap
XICEpug_h pug_h / icecap
XICEpu_h_n pu_h_n / icecap
XICEpad pad / icecap
mI20 pug_h nghs_h pu_h_n vssio sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI30 pu_h_n pghs_h pug_h vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mpdrv pad pug_h vddio vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=12 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
* .SUBCKT sky130_fd_io__tk_em2o a b
* *.PININFO a:B b:B
* rI1 a net11 short
* rI2 b net7 short
* .ENDS
* .SUBCKT sky130_fd_io__tk_em2s a b
* *.PININFO a:B b:B
* rI1 a net8 short
* rI2 b net8 short
* .ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5 pb pd pgin ps
*.PININFO pgin:I pb:B pd:B ps:B
XICEnet15 pgin / icecap
XICEpgin pgin / icecap
XICEpd pd / icecap
mpdrv pd pgin ps pb sky130_fd_pr__esd_pfet_g5v0d10v5 m=1 w=15.50 l=0.55 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pudrvr_strong nghs_h<4> nghs_h<3> nghs_h<2> pad 
+ pghs_h<4> pghs_h<3> pghs_h<2> pu_csd_h pu_h_n<3> pu_h_n<2> pug_h<4> pug_h<3> 
+ pug_h<2> tie_hi_esd vddio vddio_amx vpb_drvr vssd vssio
*.PININFO nghs_h<4>:I nghs_h<3>:I nghs_h<2>:I pghs_h<4>:I pghs_h<3>:I 
*.PININFO pghs_h<2>:I pu_csd_h:I pu_h_n<3>:I pu_h_n<2>:I vddio:I vssd:I 
*.PININFO vssio:I tie_hi_esd:O pad:B pug_h<4>:B pug_h<3>:B pug_h<2>:B 
*.PININFO vddio_amx:B vpb_drvr:B
XI155<0> vpb_drvr / icecap
XI155<1> vpb_drvr / icecap
XICEtie_hi_vpbdrvr tie_hi_vpbdrvr / icecap
XICEpug_h<2> pug_h<2> / icecap
XICEnet83 net83 / icecap
XICEvddio_amx vddio_amx / icecap
XICEpu_h_n<3> pu_h_n<3> / icecap
XICEpug_h<3> pug_h<3> / icecap
XICEpghs_h<3> pghs_h<3> / icecap
XICEnet81 net81 / icecap
XICEpug_h<4> pug_h<4> / icecap
XICEpghs_h<4> pghs_h<4> / icecap
XICEnghs_h<4> nghs_h<4> / icecap
XICEpu_csd_h pu_csd_h / icecap
XICEtie_hi_esd tie_hi_esd / icecap
XICEpghs_h<2> pghs_h<2> / icecap
XICEnghs_h<2> nghs_h<2> / icecap
XICEnet079 net079 / icecap
XICEpu_h_n<2> pu_h_n<2> / icecap
XICEnghs_h<3> nghs_h<3> / icecap
XICEnet79 net79 / icecap
XICEpad pad / icecap
XI49 vddio tie_hi_esd / sky130_fd_io__tk_tie_r_out_esd
XI133 vpb_drvr tie_hi_vpbdrvr / sky130_fd_io__tk_tie_r_out_esd
XI112 pug_h<2> net83 / sky130_fd_io__tk_em2o
XI111 pug_h<4> net81 / sky130_fd_io__tk_em2o
XI141 pug_h<3> net79 / sky130_fd_io__tk_em2o
XI152 pug_h<4> net079 / sky130_fd_io__tk_em2o
XI142 tie_hi_vpbdrvr net79 / sky130_fd_io__tk_em2s
XI82 tie_hi_vpbdrvr net83 / sky130_fd_io__tk_em2s
XI109 tie_hi_vpbdrvr net81 / sky130_fd_io__tk_em2s
XI153 tie_hi_vpbdrvr net079 / sky130_fd_io__tk_em2s
Xn7 vpb_drvr pad pug_h<3> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn6 vpb_drvr pad pug_h<3> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn5<2> vpb_drvr pad pug_h<3> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn5<1> vpb_drvr pad pug_h<3> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn5<0> vpb_drvr pad pug_h<3> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn4 vpb_drvr pad pug_h<2> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn2<3> vpb_drvr pad net83 vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn2<2> vpb_drvr pad net83 vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn2<1> vpb_drvr pad net83 vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn2<0> vpb_drvr pad net83 vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn9<1> vpb_drvr pad net79 vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn9<0> vpb_drvr pad net79 vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn11<1> vpb_drvr pad pug_h<4> vddio_amx / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn11<0> vpb_drvr pad pug_h<4> vddio_amx / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn12<1> vpb_drvr pad net81 vddio_amx / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn12<0> vpb_drvr pad net81 vddio_amx / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn1<1> vpb_drvr pad pug_h<2> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn1<0> vpb_drvr pad pug_h<2> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn3<1> vpb_drvr pad pug_h<2> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn3<0> vpb_drvr pad pug_h<2> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn8<1> vpb_drvr pad pug_h<3> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn8<0> vpb_drvr pad pug_h<3> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn10<1> vpb_drvr pad net079 vddio_amx / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn10<0> vpb_drvr pad net079 vddio_amx / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
mI136 pug_h<4> nghs_h<4> pu_csd_h vssio sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI127 pug_h<2> nghs_h<2> pu_h_n<2> vssio sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI25 pug_h<3> nghs_h<3> pu_h_n<3> vssio sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI137 pu_csd_h pghs_h<4> pug_h<4> vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI128 pu_h_n<2> pghs_h<2> pug_h<2> vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI24 pu_h_n<3> pghs_h<3> pug_h<3> vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_odrvr_sub nghs_h pad pad_esd pd_csd_h pd_h<3> 
+ pd_h<2> pd_h<1> pd_h<0> pghs_h pu_csd_h pu_h_n<3> pu_h_n<2> pu_h_n<1> 
+ pu_h_n<0> pug_h<4> pug_h<3> pug_h<2> pug_h<1> pug_h<0> tie_hi_esd tie_lo_esd 
+ vddio vddio_amx vpb_drvr vssd vssio vssio_amx
*.PININFO nghs_h:I pd_csd_h:I pd_h<3>:I pd_h<2>:I pd_h<1>:I pd_h<0>:I pghs_h:I 
*.PININFO pu_csd_h:I pu_h_n<3>:I pu_h_n<2>:I pu_h_n<1>:I pu_h_n<0>:I vddio:I 
*.PININFO vssd:I vssio:I vssio_amx:I pad:B pad_esd:B pug_h<4>:B pug_h<3>:B 
*.PININFO pug_h<2>:B pug_h<1>:B pug_h<0>:B tie_hi_esd:B tie_lo_esd:B 
*.PININFO vddio_amx:B vpb_drvr:B
Xpddrvr_strong_slow strong_slow_pad pd_h<1> vddio vssio / 
+ sky130_fd_io__gpio_pddrvr_strong_slow
XI73 weak_pad pd_h<0> vddio vssio / sky130_fd_io__gpio_pddrvr_weak
Xres strong_slow_pad pad_esd vssio / sky130_fd_io__com_res_strong_slow
Xres_weak weak_pad pad_esd vssio / sky130_fd_io__com_res_weak
Xpd_drvr pad pd_csd_h pd_h<3> pd_h<2> tie_lo_esd vddio vssio vssio_amx / 
+ sky130_fd_io__gpio_ovtv2_pddrvr
Xpudrvr_weak nghs_h weak_pad pghs_h pu_h_n<0> pug_h<0> vddio vpb_drvr vssd 
+ vssio / sky130_fd_io__gpio_ovtv2_pudrvr_weak
Xstrong_slow_pudrvr nghs_h strong_slow_pad pghs_h pu_h_n<1> pug_h<1> vddio 
+ vpb_drvr vssd vssio / sky130_fd_io__gpio_ovtv2_pudrvr_strong_slow
Xpudrvr_strong nghs_h nghs_h nghs_h pad pghs_h pghs_h pghs_h pu_csd_h 
+ pu_h_n<3> pu_h_n<2> pug_h<4> pug_h<3> pug_h<2> tie_hi_esd vddio vddio_amx 
+ vpb_drvr vssd vssio / sky130_fd_io__gpio_ovtv2_pudrvr_strong
Xres_esd pad_esd pad / s8_esd_res75only_small
xI72 vssio vddio condiode
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_odrvr_i2c_fix_leak_fix force_h<1> nga_pad_vpmp_h 
+ ngb_pad_vpmp_h nghs_h od_i_h_n oe_hs_h pad pd_csd_h pd_h<3> pd_h<2> pd_h<1> 
+ pd_h<0> pghs_h pu_csd_h pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> pug_h<7> 
+ pug_h<6> pug_h<5> tie_hi_esd tie_lo_esd vddio vddio_amx vpb_drvr vssa vssd 
+ vssio vssio_amx
*.PININFO force_h<1>:I nga_pad_vpmp_h:I ngb_pad_vpmp_h:I od_i_h_n:I oe_hs_h:I 
*.PININFO pd_csd_h:I pd_h<3>:I pd_h<2>:I pd_h<1>:I pd_h<0>:I pu_csd_h:I 
*.PININFO pu_h_n<3>:I pu_h_n<2>:I pu_h_n<1>:I pu_h_n<0>:I vddio:I vssa:I 
*.PININFO vssd:I vssio:I vssio_amx:I nghs_h:O pad:O pghs_h:O tie_hi_esd:O 
*.PININFO tie_lo_esd:O pug_h<7>:B pug_h<6>:B pug_h<5>:B vddio_amx:B vpb_drvr:B
XICEnghs_h nghs_h / icecap
XICEtie_lo_esd tie_lo_esd / icecap
XICEpad_esd pad_esd / icecap
XICEpd_csd_h pd_csd_h / icecap
XICEpghs_h pghs_h / icecap
XICEoe_hs_h oe_hs_h / icecap
XICEvpb_drvr vpb_drvr / icecap
XICEod_i_h_n od_i_h_n / icecap
XICEpu_csd_h pu_csd_h / icecap
XICEnet74 net74 / icecap
XI196<0> pu_h_n<3> / icecap
XI196<1> pu_h_n<2> / icecap
XI196<2> pu_h_n<1> / icecap
XI196<3> pu_h_n<0> / icecap
XICEp2g p2g / icecap
XI195<0> pd_h<3> / icecap
XI195<1> pd_h<2> / icecap
XI195<2> pd_h<1> / icecap
XI199<0> pug_h<4> / icecap
XI199<1> pug_h<3> / icecap
XI199<2> pug_h<2> / icecap
XI199<3> pug_h<1> / icecap
XI199<4> pug_h<0> / icecap
XICEforce_h<1> force_h<1> / icecap
XICEpad pad / icecap
XI194<0> pd_h<3> / icecap
XI194<1> pd_h<2> / icecap
XI194<2> pd_h<1> / icecap
XI194<3> pd_h<0> / icecap
XI197<0> pd_csd_h / icecap
XI197<1> nga_pad_vpmp_h / icecap
XI197<2> ngb_pad_vpmp_h / icecap
XICEtie_hi_esd tie_hi_esd / icecap
XI198<0> pug_h<7> / icecap
XI198<1> pug_h<6> / icecap
XI198<2> pug_h<5> / icecap
XI198<3> pug_h<4> / icecap
XI198<4> pug_h<3> / icecap
XI198<5> pug_h<2> / icecap
XI198<6> pug_h<1> / icecap
XI198<7> pug_h<0> / icecap
Xhotswap force_h<1> nghs_h od_i_h_n oe_hs_h p2g pad pad_esd pghs_h pug_h<7> 
+ pug_h<6> pug_h<5> pug_h<4> pug_h<3> pug_h<2> pug_h<1> pug_h<0> net74 vddio 
+ vpb_drvr vddio vssd / sky130_fd_io__gpio_ovtv2_hotswap_i2c_fix_leak_fix
Xbondpad pad vssio / sky130_fd_io__com_pad
Xodrvr tie_hi_esd pad pad_esd pd_csd_h pd_h<3> pd_h<2> pd_h<1> pd_h<0> pghs_h 
+ pu_csd_h pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> pug_h<4> pug_h<3> pug_h<2> 
+ pug_h<1> pug_h<0> tie_hi_esd tie_lo_esd vddio vddio_amx vpb_drvr vssd vssio 
+ vssio_amx / sky130_fd_io__gpio_ovtv2_odrvr_sub
mI122<2> pd_h<3> pghs_h net106<0> vssio sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI122<1> pd_h<2> pghs_h net106<1> vssio sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI122<0> pd_h<1> pghs_h net106<2> vssio sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI85<2> net106<0> pghs_h vssio vssio sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI85<1> net106<1> pghs_h vssio vssio sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI85<0> net106<2> pghs_h vssio vssio sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI104<2> net102<0> pghs_h vssa vssio sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI104<1> net102<1> pghs_h vssa vssio sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI104<0> net102<2> pghs_h vssa vssio sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI103<2> pd_csd_h pghs_h net102<0> vssio sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI103<1> nga_pad_vpmp_h pghs_h net102<1> vssio sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI103<0> ngb_pad_vpmp_h pghs_h net102<2> vssio sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__nor3_dnw in0 in1 in2 out vgnd vpwr
*.PININFO in0:I in1:I in2:I vgnd:I vpwr:I out:O
XICEout out / icecap
XICEin0 in0 / icecap
XICEin1 in1 / icecap
XICEin2 in2 / icecap
mI3 net43 in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI12 net39 in1 net43 vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI16 out in2 net39 vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI1 out in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI6 out in1 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI18 out in2 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
* .SUBCKT sky130_fd_io__com_inv_x1_dnw in out vgnd vpwr
* *.PININFO in:I vgnd:I vpwr:I out:O
* XICEin in / icecap
* XICEout out / icecap
* mI1 out in vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI2 out in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__com_nand2_dnw in0 in1 out vgnd vpwr
* *.PININFO in0:I in1:I vgnd:I vpwr:I out:O
* XICEout out / icecap
* XICEin1 in1 / icecap
* XICEin0 in0 / icecap
* mI3 out in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI5 out in1 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI1 out in1 net25 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI6 net25 in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__com_nor2_dnw in0 in1 out vgnd vpwr
* *.PININFO in0:I in1:I vgnd:I vpwr:I out:O
* XICEin1 in1 / icecap
* XICEin0 in0 / icecap
* XICEout out / icecap
* mI3 net17 in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI12 out in1 net17 vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI1 out in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI6 out in1 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_predrvr_switch nmos_en pmos_en sig1 sig2 vcc_io 
+ vgnd_io
*.PININFO nmos_en:I pmos_en:I vcc_io:I vgnd_io:I sig1:B sig2:B
XICEpmos_en pmos_en / icecap
XICEsig1 sig1 / icecap
XICEnmos_en nmos_en / icecap
XICEsig2 sig2 / icecap
mI374 sig1 nmos_en sig2 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI375 sig2 pmos_en sig1 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_leak_fix drvlo_h_n en_cmos_b 
+ i2c_mode_h_n nghs_h nsw_en_int oe_i_h_n pad_cap pd_dis_h pd_h<3> pd_h<2> 
+ pden_h_n<1> pghs_h pug_h slew_ctl_h<1> slew_ctl_h<0> slew_ctl_h_n<1> 
+ slew_ctl_h_n<0> slow_h_n vcc_io vgnd_io vpb_drvr vssd
*.PININFO drvlo_h_n:I i2c_mode_h_n:I nghs_h:I oe_i_h_n:I pd_dis_h:I 
*.PININFO pden_h_n<1>:I pghs_h:I pug_h:I slew_ctl_h<1>:I slew_ctl_h<0>:I 
*.PININFO slew_ctl_h_n<1>:I slew_ctl_h_n<0>:I slow_h_n:I vcc_io:I vgnd_io:I 
*.PININFO vpb_drvr:I vssd:I en_cmos_b:O nsw_en_int:O pd_h<3>:O pd_h<2>:O 
*.PININFO pad_cap:B
XICEnsw_en_int nsw_en_int / icecap
XICEpug_h pug_h / icecap
XI319<0> cas3 / icecap
XI319<1> cas10 / icecap
XICEen_cmos_b en_cmos_b / icecap
XICEcas4 cas4 / icecap
XICEnet200 net200 / icecap
XICEna na / icecap
XICEnet519 net519 / icecap
XICEvdiode vdiode / icecap
XICEslew_ctl_h_n<1> slew_ctl_h_n<1> / icecap
XICEnet400 net400 / icecap
XICEpden_h_n<1> pden_h_n<1> / icecap
XICEcas2 cas2 / icecap
XICEslew_ctl_h<0> slew_ctl_h<0> / icecap
XICEne ne / icecap
XICEnet336 net336 / icecap
XICEpd_h<3> pd_h<3> / icecap
XICEdrvlo_h_n_i2c_4 drvlo_h_n_i2c_4 / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEcas5 cas5 / icecap
XICEslew_ctl_h<1> slew_ctl_h<1> / icecap
XICEnet278 net278 / icecap
XICEnet352 net352 / icecap
XICEnet404 net404 / icecap
XICEbiasp biasp / icecap
XI318<0> na / icecap
XI318<1> nb / icecap
XI318<2> nc / icecap
XI318<3> nd / icecap
XI318<4> ne / icecap
XI318<5> nf / icecap
XICEenb enb / icecap
XICEnet263 net263 / icecap
XICEcas10 cas10 / icecap
XICEnet303 net303 / icecap
XICEnet369 net369 / icecap
XICEnet288 net288 / icecap
XICEmode2b mode2b / icecap
XICEpad_cap pad_cap / icecap
XICEdrvlo_h_n_i2c_1 drvlo_h_n_i2c_1 / icecap
XICEnet313 net313 / icecap
XICEdrvlo_h_n_buf drvlo_h_n_buf / icecap
XICEen en / icecap
XICEnet531 net531 / icecap
XICEnet298 net298 / icecap
XICEnet193 net193 / icecap
XICEnet420 net420 / icecap
XICEvr vr / icecap
XICEnet388 net388 / icecap
XICEnc nc / icecap
XICEnet552 pd_h<3> / icecap
XICEnet318 net318 / icecap
XICEnet535 net535 / icecap
XICEslew_ctl_h_n<0> slew_ctl_h_n<0> / icecap
XICEpd_h<2> pd_h<2> / icecap
XICEnsw_en nsw_en / icecap
XICEdrvlo_h_n_i2c_2 drvlo_h_n_i2c_2 / icecap
XICEnet499 vcc_io / icecap
XICEnet283 net283 / icecap
XICEnghs_h nghs_h / icecap
XICEpd_dis_h pd_dis_h / icecap
XICE2vtn N0 / icecap
XICEvdelay vdelay / icecap
XICEnsw_enb nsw_enb / icecap
XICEoe_i_h_n oe_i_h_n / icecap
XICEdrvlo_h drvlo_h / icecap
XICEmode3b mode3b / icecap
XICEnet613 net352 / icecap
XICEnf nf / icecap
XICEpghs_h pghs_h / icecap
XICEnet190 net190 / icecap
XICEbiasp1 biasp1 / icecap
XICEpden_h<1> pden_h<1> / icecap
XICEmode1b mode1b / icecap
XICEnb nb / icecap
XICEi2c_mode_h_n i2c_mode_h_n / icecap
XICEdrvlo_h_n_i2c drvlo_h_n_i2c / icecap
XICEslow_h_n slow_h_n / icecap
XICEcas3 cas3 / icecap
XICEdrvlo_h_n_i2c_3 drvlo_h_n_i2c_3 / icecap
XICEnet293 net293 / icecap
XICEnd nd / icecap
rI288 N0 net193 sky130_fd_pr__res_generic_nd__hv m=1 w=0.5 l=113.375 isHV=TRUE
rI287 vdiode net190 sky130_fd_pr__res_generic_nd__hv m=1 w=0.5 l=113.375 isHV=TRUE
XI123 pd_dis_h nsw_enb oe_i_h_n net200 vgnd_io vcc_io / sky130_fd_io__nor3_dnw
xI208 vgnd_io vcc_io condiode
XI161 net293 drvlo_h_n_i2c_2 vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI159 net298 drvlo_h_n_i2c_1 vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI224 net288 net247 vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI605 en enb vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI176 net318 drvlo_h_n_i2c_4 vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI191 nsw_en nsw_enb vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI198 net303 drvlo_h_n_i2c vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI179 net283 nsw_en_int vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI168 net263 mode1b vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI122 drvlo_h drvlo_h_n_buf vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI170 net278 mode3b vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI715 pden_h_n<1> pden_h<1> vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI162 net313 drvlo_h_n_i2c_3 vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI254 drvlo_h_n drvlo_h vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI602 vdelay net200 en vgnd_io vcc_io / sky130_fd_io__com_nand2_dnw
XI112 pden_h<1> nsw_enb en_cmos_b vgnd_io vcc_io / sky130_fd_io__com_nand2_dnw
XI430 slew_ctl_h<1> slew_ctl_h_n<0> net263 vgnd_io vcc_io / 
+ sky130_fd_io__com_nand2_dnw
XI175 drvlo_h_n_i2c mode4b net318 vgnd_io vcc_io / sky130_fd_io__com_nor2_dnw
XI163 drvlo_h_n_i2c mode3b net313 vgnd_io vcc_io / sky130_fd_io__com_nor2_dnw
XI109 slow_h_n i2c_mode_h_n nsw_en vgnd_io vcc_io / sky130_fd_io__com_nor2_dnw
XI197 nsw_enb drvlo_h_n_buf net303 vgnd_io vcc_io / sky130_fd_io__com_nor2_dnw
XI158 drvlo_h_n_i2c mode1b net298 vgnd_io vcc_io / sky130_fd_io__com_nor2_dnw
XI160 drvlo_h_n_i2c mode2b net293 vgnd_io vcc_io / sky130_fd_io__com_nor2_dnw
XI225 slew_ctl_h<1> slew_ctl_h<0> net288 vgnd_io vcc_io / sky130_fd_io__com_nor2_dnw
XI181 pden_h_n<1> nsw_en net283 vgnd_io vcc_io / sky130_fd_io__com_nor2_dnw
XI169 slew_ctl_h<1> slew_ctl_h_n<0> net278 vgnd_io vcc_io / 
+ sky130_fd_io__com_nor2_dnw
xI99 net0101 net0100 net099 net098 sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3 m=18
mI206 N0 en vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI190 net531 en vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI220 net420 enb vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI153 pd_h<2> pden_h_n<1> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI182 vgnd_io vdelay vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.00 l=2.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI201 net352 N0 net190 vgnd_io sky130_fd_pr__nfet_05v0_nvt m=10 w=1.00 l=0.90 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI625 net404 pd_h<3> net348 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI339 net400 pden_h<1> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI125 pd_h<3> drvlo_h_n_buf net400 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI344 pd_h<3> pden_h_n<1> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI63 net388 vdiode pd_h<3> vgnd_io sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=0.90 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI189 net388 vgnd_io vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI10 biasp vdiode net336 vgnd_io sky130_fd_pr__nfet_05v0_nvt m=5 w=10.0 l=0.90 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI374 net519 nsw_en pd_h<3> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI137 biasp1 vdiode vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI13 net369 net369 vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=5 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI8 vdiode vdiode vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=5 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI165 vdiode en vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI14 N0 N0 net369 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=5 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI15 net352 N0 net190 vgnd_io sky130_fd_pr__nfet_05v0_nvt m=4 w=10.0 l=0.90 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI755 net348 pd_h<3> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI579 vdelay drvlo_h net404 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI192 net519 vgnd_io vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI219 net336 vdiode vr vgnd_io sky130_fd_pr__nfet_01v8_lvt m=5 w=7.00 l=0.15 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI232<1> cas3 pghs_h pd_h<3> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI232<0> cas10 pghs_h pd_h<3> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI278 vgnd_io vgnd_io vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI20 pug_h nghs_h nsw_enb vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI245 cas10 vcc_io cas4 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI196 nc biasp vcc_io vcc_io sky130_fd_pr__pfet_01v8 m=5 w=0.55 l=1.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI200 cas3 biasp1 nc vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI199 pd_h<3> drvlo_h_n_i2c_2 cas3 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI205 net352 en vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI156 cas5 biasp1 ne vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI580 vdelay drvlo_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI136 biasp biasp1 na vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI144 cas4 biasp1 nd vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI84 pd_h<3> drvlo_h_n_i2c cas2 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI230 nc vcc_io vcc_io vcc_io sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=1.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI79 nb biasp vcc_io vcc_io sky130_fd_pr__pfet_01v8 m=17 w=0.55 l=1.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI260 net535 enb vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI228 pd_h<3> drvlo_h_n_i2c net535 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI73 net388 drvlo_h_n_i2c net531 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI561 pd_h<3> drvlo_h_n_i2c_1 cas4 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI560 nd biasp vcc_io vcc_io sky130_fd_pr__pfet_01v8 m=14 w=0.55 l=1.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI375 pd_h<3> pug_h net519 vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI164 biasp enb vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI167 biasp1 enb vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI138 biasp1 biasp1 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI145 cas2 biasp1 nb vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI141 na biasp vcc_io vcc_io sky130_fd_pr__pfet_01v8 m=10 w=0.55 l=1.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI154 ne biasp vcc_io vcc_io sky130_fd_pr__pfet_01v8 m=14 w=0.55 l=1.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI178 net193 en vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI155 pd_h<3> drvlo_h_n_i2c_3 cas5 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI241 cas10 biasp1 nf vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI240 nf biasp vcc_io vcc_io sky130_fd_pr__pfet_01v8 m=8 w=0.55 l=1.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI229 ne vcc_io vcc_io vcc_io sky130_fd_pr__pfet_01v8 m=2 w=0.55 l=4.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI217 nb vcc_io vcc_io vcc_io sky130_fd_pr__pfet_01v8 m=3 w=0.55 l=1.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI216 nd vcc_io vcc_io vcc_io sky130_fd_pr__pfet_01v8 m=2 w=0.55 l=1.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI215 cas3 vcc_io cas2 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI214 cas5 vcc_io cas2 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI239 pd_h<3> drvlo_h_n_i2c_3 cas10 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI213 cas3 vcc_io cas4 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI212 na vcc_io vcc_io vcc_io sky130_fd_pr__pfet_01v8 m=2 w=0.55 l=1.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI211 vcc_io vcc_io vcc_io vcc_io sky130_fd_pr__pfet_01v8 m=4 w=0.55 l=1.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI210 vcc_io vcc_io vcc_io vcc_io sky130_fd_pr__pfet_01v8 m=6 w=0.55 l=4.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI248<5> na enb vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI248<4> nb enb vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI248<3> nc enb vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI248<2> nd enb vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI248<1> ne enb vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI248<0> nf enb vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI30 nsw_enb pghs_h pug_h vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI70 net531 en vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
XI94 nsw_en nsw_enb pd_h<2> pd_h<3> vcc_io vgnd_io / 
+ sky130_fd_io__gpio_ovtv2_predrvr_switch
rI221 net420 vr sky130_fd_pr__res_generic_po m=1 w=0.75 l=513.445
rI186 slew_ctl_h_n<0> mode4b short
rI157 net247 mode2b short
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_obpredrvr_new_leak_fix drvlo_h_n en_cmos_b 
+ i2c_mode_h_n nghs_h nsw_en oe_i_h_n pad pd_dis_h pd_h<3> pd_h<2> pden_h_n<1> 
+ pghs_h pug_h slew_ctl_h<1> slew_ctl_h<0> slew_ctl_h_n<1> slew_ctl_h_n<0> 
+ slow_h_n vcc_io vgnd_io vpb_drvr vssd
*.PININFO drvlo_h_n:I i2c_mode_h_n:I nghs_h:I oe_i_h_n:I pd_dis_h:I 
*.PININFO pden_h_n<1>:I pghs_h:I pug_h:I slew_ctl_h<1>:I slew_ctl_h<0>:I 
*.PININFO slew_ctl_h_n<1>:I slew_ctl_h_n<0>:I slow_h_n:I vcc_io:I vgnd_io:I 
*.PININFO vpb_drvr:I vssd:I en_cmos_b:O nsw_en:O pd_h<3>:O pd_h<2>:O pad:B
XICEpden_h_n<1> pden_h_n<1> / icecap
XICEpad pad / icecap
XICEvssd vssd / icecap
XICEoe_i_h_n oe_i_h_n / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEi2c_mode_h_n i2c_mode_h_n / icecap
XICEpug_h pug_h / icecap
XICEpghs_h pghs_h / icecap
XICEen_cmos_b en_cmos_b / icecap
XI89<0> slew_ctl_h<1> / icecap
XI89<1> slew_ctl_h<0> / icecap
XICEnghs_h nghs_h / icecap
XI88<0> pd_h<3> / icecap
XI88<1> pd_h<2> / icecap
XICEslow_h_n slow_h_n / icecap
XICEnsw_en nsw_en / icecap
XICEpd_dis_h pd_dis_h / icecap
XI90<0> slew_ctl_h_n<1> / icecap
XI90<1> slew_ctl_h_n<0> / icecap
XICEvpb_drvr vpb_drvr / icecap
Xpd_strong drvlo_h_n en_cmos_b i2c_mode_h_n nghs_h nsw_en oe_i_h_n pad 
+ pd_dis_h pd_h<3> pd_h<2> pden_h_n<1> pghs_h pug_h slew_ctl_h<1> 
+ slew_ctl_h<0> slew_ctl_h_n<1> slew_ctl_h_n<0> slow_h_n vcc_io vgnd_io 
+ vpb_drvr vssd / sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_leak_fix
.ENDS
* .SUBCKT sky130_fd_io__com_pupredrvr_strong_slow drvhi_h pu_h_n puen_h vcc_io vgnd_io
* *.PININFO drvhi_h:I puen_h:I vcc_io:I vgnd_io:I pu_h_n:O
* XICEnet17 net17 / icecap
* XICEdrvhi_h drvhi_h / icecap
* XICEpu_h_n pu_h_n / icecap
* XICEpuen_h puen_h / icecap
* mI3 pu_h_n drvhi_h net17 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI39 net17 puen_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI38 pu_h_n puen_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI37 pu_h_n drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=3 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__com_pupredrvr_weak drvhi_h pu_h_n puen_h vcc_io vgnd_io
* *.PININFO drvhi_h:I puen_h:I vcc_io:I vgnd_io:I pu_h_n:O
* XICEpu_h_n pu_h_n / icecap
* XICEpuen_h puen_h / icecap
* XICEdrvhi_h drvhi_h / icecap
* mI3 pu_h_n drvhi_h net21 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI39 net21 puen_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI38 pu_h_n puen_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI37 pu_h_n drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__com_pdpredrvr_weak drvlo_h_n pd_h pden_h_n vcc_io vgnd_io
* *.PININFO drvlo_h_n:I pden_h_n:I vcc_io:I vgnd_io:I pd_h:O
* XICEdrvlo_h_n drvlo_h_n / icecap
* XICEpd_h pd_h / icecap
* XICEnet25 net25 / icecap
* XICEpden_h_n pden_h_n / icecap
* mI26 pd_h pden_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI25 pd_h drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI24 net25 pden_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI23 pd_h drvlo_h_n net25 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__com_pdpredrvr_strong_slow drvlo_h_n pd_h pden_h_n vcc_io 
* + vgnd_io
* *.PININFO drvlo_h_n:I pden_h_n:I vcc_io:I vgnd_io:I pd_h:O
* XICEdrvlo_h_n drvlo_h_n / icecap
* XICEpd_h pd_h / icecap
* XICEnet25 net25 / icecap
* XICEpden_h_n pden_h_n / icecap
* mI26 pd_h pden_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI25 pd_h drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI24 net25 pden_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI23 pd_h drvlo_h_n net25 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__tk_opto out spd spu
* *.PININFO out:B spd:B spu:B
* Xe1 spu out / sky130_fd_io__tk_em1o
* Xe2 out spd / sky130_fd_io__tk_em1s
* .ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pdpredrvr_pbias drvlo_h_n en_h en_h_n pbias pd_h 
+ pden_h_n vcc_io vgnd_io
*.PININFO drvlo_h_n:I en_h:I en_h_n:I pd_h:I pden_h_n:I vcc_io:I vgnd_io:I 
*.PININFO pbias:O
XICEbias_g bias_g / icecap
XICEpbias pbias / icecap
XICEnet183 net183 / icecap
XICEpden_h_n pden_h_n / icecap
XICEen_h en_h / icecap
XICEn<101> n<101> / icecap
XICEnet157 net157 / icecap
XICEnet108 net108 / icecap
XICEnet171 net171 / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEdrvlo_i_h drvlo_i_h / icecap
XICEen_h_n en_h_n / icecap
XICEnet84 net84 / icecap
XICEpbias1 pbias1 / icecap
XICE2vtp N0 / icecap
XICEn<0> n<0> / icecap
XICEpd_h pd_h / icecap
XICEnet88 net88 / icecap
XICEn<1> n<1> / icecap
XICEnet161 net161 / icecap
XE1 n<1> n<0> / sky130_fd_io__tk_em1o
XE2 pbias pbias1 / sky130_fd_io__tk_em1o
XE3 pbias1 net88 / sky130_fd_io__tk_em1s
XE4 net108 pbias / sky130_fd_io__tk_em1s
XE6 pbias net84 / sky130_fd_io__tk_em1s
XE5 n<101> bias_g / sky130_fd_io__tk_em1s
XI27 n<0> pd_h en_h_n / sky130_fd_io__tk_opto
mI47 pbias bias_g vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=1.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI24 n<1> drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI18 bias_g drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI23 n<0> n<0> n<1> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI13 drvlo_i_h drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI20 bias_g n<1> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.60 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI19 bias_g en_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI34 net157 bias_g vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.60 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI36 net108 bias_g vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=1.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI38 n<1> pden_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI48 n<100> pd_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI41 n<101> pd_h n<100> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI44 pbias pbias pbias1 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI45 pbias1 pbias1 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI15 net183 en_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=10.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI16 net171 n<0> net183 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=10.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI6 pbias en_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI12 drvlo_i_h drvlo_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI17 bias_g drvlo_h_n net171 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=3 w=7.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI14 pbias drvlo_i_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI33 N0 vgnd_io vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=8.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI32 net161 net161 N0 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI31 net157 net157 net161 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI30 net88 N0 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI43 net84 bias_g vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI40 N0 drvlo_i_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr2 drvlo_h_n en_fast_n<1> 
+ en_fast_n<0> pd_h pden_h_n vcc_io vgnd_io
*.PININFO drvlo_h_n:I en_fast_n<1>:I en_fast_n<0>:I pden_h_n:I vcc_io:I 
*.PININFO vgnd_io:I pd_h:O
XICEpd_h pd_h / icecap
XICEen_fast_n<0> en_fast_n<0> / icecap
XICEpden_h_n pden_h_n / icecap
XICEint_nor<1> int_nor<1> / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEen_fast_n<1> en_fast_n<1> / icecap
XICEint_slow int_slow / icecap
XICEint_nor<0> int_nor<0> / icecap
XI373<0> int_nor<1> / icecap
XI373<1> int_nor<0> / icecap
mmnin pd_h drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=5 w=3.00 l=0.60 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI56 int_slow pden_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmpin_slow pd_h drvlo_h_n int_slow vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=4.00 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmpen_slow int_slow pden_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=4.00 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmpin_fast<1> pd_h drvlo_h_n int_nor<1> net19<0> sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmpin_fast<0> pd_h drvlo_h_n int_nor<0> net19<1> sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmpen_fast<1> int_nor<1> en_fast_n<1> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.00 l=1.00 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmpen_fast<0> int_nor<0> en_fast_n<0> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr3 drvlo_h_n en_fast_n<1> 
+ en_fast_n<0> pd_h pden_h_n vcc_io vgnd_io
*.PININFO drvlo_h_n:I en_fast_n<1>:I en_fast_n<0>:I pden_h_n:I vcc_io:I 
*.PININFO vgnd_io:I pd_h:O
XICEpd_h pd_h / icecap
XICEen_fast_n<0> en_fast_n<0> / icecap
XICEpden_h_n pden_h_n / icecap
XICEint_nor<1> int_nor<1> / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEen_fast_n<1> en_fast_n<1> / icecap
XICEint_slow int_slow / icecap
XICEint_nor<0> int_nor<0> / icecap
XI361<0> int_nor<1> / icecap
XI361<1> int_nor<0> / icecap
mmnin pd_h drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=5 w=3.00 l=0.60 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI56 int_slow pden_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmpin_slow pd_h drvlo_h_n int_slow vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=4.00 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmpen_slow int_slow pden_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=4.00 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmpin_fast<1> pd_h drvlo_h_n int_nor<1> net19<0> sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmpin_fast<0> pd_h drvlo_h_n int_nor<0> net19<1> sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmpen_fast<1> int_nor<1> en_fast_n<1> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.00 l=1.00 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmpen_fast<0> int_nor<0> en_fast_n<0> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
* .SUBCKT sky130_fd_io__tk_opti out spd spu
* *.PININFO out:B spd:B spu:B
* Xe2 spd out / sky130_fd_io__tk_em1o
* Xe1 out spu / sky130_fd_io__tk_em1s
* .ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_cmos drvhi_h drvlo_h_n en_cmos_b 
+ nsw_en_int pd_h<3> pd_h<2> pden_h_n slow_h vcc_io vgnd_io
*.PININFO drvhi_h:I drvlo_h_n:I en_cmos_b:I nsw_en_int:I pden_h_n:I slow_h:I 
*.PININFO vcc_io:I vgnd_io:I pd_h<3>:O pd_h<2>:O
Xbias drvhi_h en_fast_h en_fast_h_n pbias_out pd_h<2> pden_h_n vcc_io vgnd_io 
+ / sky130_fd_io__gpio_ovtv2_pdpredrvr_pbias
Xnr3 drvlo_h_n net76 net76 pd_h<2> nsw_en_int vcc_io vgnd_io / 
+ sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr2
Xnr2 drvlo_h_n en_fast2_n<1> en_fast2_n<0> pd_h<3> nsw_en_int vcc_io vgnd_io / 
+ sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr3
XI77 en_fast2_n<1> pbias_out en_fast_h_n / sky130_fd_io__tk_opto
XI76 net76 pbias_out en_fast_h_n / sky130_fd_io__tk_opto
XI79 en_fast2_n<0> en_fast2_n<1> vcc_io / sky130_fd_io__tk_opti
Xinv en_fast_h en_fast_h_n vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
Xnor slow_h en_cmos_b en_fast_h vgnd_io vcc_io / sky130_fd_io__com_nor2_dnw
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd3 drvhi_h en_fast<3> en_fast<2> 
+ en_fast<1> en_fast<0> pu_h_n puen_h vcc_io vgnd_io
*.PININFO drvhi_h:I en_fast<3>:I en_fast<2>:I en_fast<1>:I en_fast<0>:I 
*.PININFO puen_h:I vcc_io:I vgnd_io:I pu_h_n:O
XICEnet30 net30 / icecap
XICEint<0> int<0> / icecap
XICEdrvhi_h drvhi_h / icecap
XICEen_fast<0> en_fast<0> / icecap
XICEpu_h_n pu_h_n / icecap
XICEpuen_h puen_h / icecap
XI152<0> int<3> / icecap
XI152<1> int<2> / icecap
XI152<2> int<1> / icecap
XICEint_res int_res / icecap
XICEn<2> n<2> / icecap
XI150<0> en_fast<3> / icecap
XI150<1> en_fast<2> / icecap
XI150<2> en_fast<1> / icecap
XI151<0> int<3> / icecap
XI151<1> int<2> / icecap
XI151<2> int<1> / icecap
XI151<3> int<0> / icecap
XE1 net30 pu_h_n / sky130_fd_io__tk_em1s
rrespu1 int_res net30 sky130_fd_pr__res_generic_po m=1 w=0.33 l=11
rrespu2 pu_h_n int_res sky130_fd_pr__res_generic_po m=1 w=0.33 l=4
mmnin_fast<3> net30 drvhi_h int<3> net017<0> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmnin_fast<2> net30 drvhi_h int<2> net017<1> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmnin_fast<1> net30 drvhi_h int<1> net017<2> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmnin_fast<0> net30 drvhi_h int<0> net017<3> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmnen_slow1 n<2> puen_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=4.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmnin_slow pu_h_n drvhi_h n<2> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmnen_fast<3> int<3> en_fast<3> vgnd_io net018<0> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmnen_fast<2> int<2> en_fast<2> vgnd_io net018<1> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmnen_fast<1> int<1> en_fast<1> vgnd_io net018<2> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmnen_fast<0> int<0> en_fast<0> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmpen pu_h_n puen_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.60 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmpin pu_h_n drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=3 w=5.00 l=0.60 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd2 drvhi_h en_fast<3> en_fast<2> 
+ en_fast<1> en_fast<0> pu_h_n puen_h vcc_io vgnd_io
*.PININFO drvhi_h:I en_fast<3>:I en_fast<2>:I en_fast<1>:I en_fast<0>:I 
*.PININFO puen_h:I vcc_io:I vgnd_io:I pu_h_n:O
XI148<0> int<3> / icecap
XI148<1> int<2> / icecap
XI148<2> int<1> / icecap
XI148<3> int<0> / icecap
XI147<0> en_fast<3> / icecap
XI147<1> en_fast<2> / icecap
XI147<2> en_fast<1> / icecap
XICEn<2> n<2> / icecap
XICEpu_h_n pu_h_n / icecap
XICEnet30 net30 / icecap
XICEpuen_h puen_h / icecap
XICEint<0> int<0> / icecap
XICEdrvhi_h drvhi_h / icecap
XI149<0> int<3> / icecap
XI149<1> int<2> / icecap
XI149<2> int<1> / icecap
XICEen_fast<0> en_fast<0> / icecap
XICEint_res int_res / icecap
XE1 net30 pu_h_n / sky130_fd_io__tk_em1s
rrespu1 int_res net30 sky130_fd_pr__res_generic_po m=1 w=0.33 l=11
rrespu2 pu_h_n int_res sky130_fd_pr__res_generic_po m=1 w=0.33 l=4
mmnin_fast<3> net30 drvhi_h int<3> net017<0> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmnin_fast<2> net30 drvhi_h int<2> net017<1> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmnin_fast<1> net30 drvhi_h int<1> net017<2> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmnin_fast<0> net30 drvhi_h int<0> net017<3> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmnen_slow1 n<2> puen_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=4.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmnin_slow pu_h_n drvhi_h n<2> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmnen_fast<3> int<3> en_fast<3> vgnd_io net018<0> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=1.00 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmnen_fast<2> int<2> en_fast<2> vgnd_io net018<1> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=1.00 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmnen_fast<1> int<1> en_fast<1> vgnd_io net018<2> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=1.00 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmnen_fast<0> int<0> en_fast<0> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmpen pu_h_n puen_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.60 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmpin pu_h_n drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=3 w=5.00 l=0.60 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
* .SUBCKT sky130_fd_io__com_pupredrvr_nbias drvhi_h en_h en_h_n nbias pu_h_n puen_h 
* + vcc_io vgnd_io
* *.PININFO drvhi_h:I en_h:I en_h_n:I pu_h_n:I puen_h:I vcc_io:I vgnd_io:I 
* *.PININFO nbias:O
* XICEn<6> n<6> / icecap
* XICEdrvhi_i_h_n drvhi_i_h_n / icecap
* XICEen_h_n en_h_n / icecap
* XICEbias_g bias_g / icecap
* XICEn<2> n<2> / icecap
* XICEn<8> n<8> / icecap
* XICEdrvhi_h drvhi_h / icecap
* XICEen_h en_h / icecap
* XICEnet141 net141 / icecap
* XICEvccio_2vtn vccio_2vtn / icecap
* XICEnbias nbias / icecap
* XICEnet153 net153 / icecap
* XICEpu_h_n pu_h_n / icecap
* XICEnet88 net88 / icecap
* XICEn<7> n<7> / icecap
* XICEn<1> n<1> / icecap
* XICEnet90 net90 / icecap
* XICEpuen_h puen_h / icecap
* XI36 n<2> pu_h_n en_h / sky130_fd_io__tk_opto
* XE5 nbias net88 / sky130_fd_io__tk_em1s
* XE4 n<6> net153 / sky130_fd_io__tk_em1s
* XE7 bias_g net90 / sky130_fd_io__tk_em1s
* XE6 net141 nbias / sky130_fd_io__tk_em1s
* XE1 n<2> n<1> / sky130_fd_io__tk_em1o
* XE2 n<6> nbias / sky130_fd_io__tk_em1o
* mI34 n<1> drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI32 n<1> n<2> n<2> vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI31 bias_g n<1> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI30 bias_g drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI29 bias_g en_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI21 nbias bias_g vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.00 l=0.80 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI12 drvhi_i_h_n drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI47 n<7> bias_g vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI49 net88 bias_g vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.00 l=0.80 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI50 n<1> puen_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI56 vcc_io pu_h_n net90 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=8.00 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI19 n<6> n<6> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=4 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI20 nbias nbias n<6> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=4 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI28 bias_g drvhi_h n<3> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI27 n<3> n<2> n<4> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI26 n<4> en_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI13 drvhi_i_h_n drvhi_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI24 nbias en_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI53 vccio_2vtn drvhi_i_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI25 nbias drvhi_i_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI40 vccio_2vtn vcc_io vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI39 net153 vccio_2vtn vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=4 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI44 n<8> n<8> vccio_2vtn vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI41 n<7> n<7> n<8> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI54 net141 bias_g vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.00 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* .ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pupredrvr_strong drvhi_h pu_h_n<3> pu_h_n<2> 
+ puen_h slow_h_n vcc_io vgnd_io
*.PININFO drvhi_h:I puen_h:I slow_h_n:I vcc_io:I vgnd_io:I pu_h_n<3>:O 
*.PININFO pu_h_n<2>:O
Xnd2b drvhi_h en_fast_h_3<3> en_fast_h_3<2> en_fast_h_3<1> en_fast_h_3<0> 
+ pu_h_n<3> puen_h vcc_io vgnd_io / sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd3
Xnd2a drvhi_h net54 net54 net54 net54 pu_h_n<2> puen_h vcc_io vgnd_io / 
+ sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd2
XI98 en_fast_h_3<0> en_fast_h_3<3> vgnd_io / sky130_fd_io__tk_opti
XI97 en_fast_h_3<1> en_fast_h_3<3> vgnd_io / sky130_fd_io__tk_opti
XI92 en_fast_h_3<3> nbias_out en_fast_h / sky130_fd_io__tk_opto
XI96 en_fast_h_3<2> en_fast_h_3<3> vgnd_io / sky130_fd_io__tk_opto
XI93 net54 nbias_out en_fast_h / sky130_fd_io__tk_opto
Xinv en_fast_h_n en_fast_h vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
Xnbias drvhi_h en_fast_h en_fast_h_n nbias_out pu_h_n<2> puen_h vcc_io vgnd_io 
+ / sky130_fd_io__com_pupredrvr_nbias
Xnand puen_h slow_h_n en_fast_h_n vgnd_io vcc_io / sky130_fd_io__com_nand2_dnw
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_obpredrvr_old drvhi_h drvlo_h_n en_cmos_b nsw_en 
+ pd_h<3> pd_h<2> pd_h<1> pd_h<0> pden_h_n<1> pden_h_n<0> pu_h_n<3> pu_h_n<2> 
+ pu_h_n<1> pu_h_n<0> puen_h<1> puen_h<0> slow_h slow_h_n vcc_io vgnd_io
*.PININFO drvhi_h:I drvlo_h_n:I en_cmos_b:I nsw_en:I pden_h_n<1>:I 
*.PININFO pden_h_n<0>:I puen_h<1>:I puen_h<0>:I slow_h:I slow_h_n:I vcc_io:I 
*.PININFO vgnd_io:I pd_h<3>:O pd_h<2>:O pd_h<1>:O pd_h<0>:O pu_h_n<3>:O 
*.PININFO pu_h_n<2>:O pu_h_n<1>:O pu_h_n<0>:O
XICEpden_h_n<0> pden_h_n<0> / icecap
XICEdrvhi_h drvhi_h / icecap
XICEpd_h<0> pd_h<0> / icecap
XICEpuen_h<1> puen_h<1> / icecap
XICEslow_h slow_h / icecap
XICEpd_h<1> pd_h<1> / icecap
XICEpu_h_n<0> pu_h_n<0> / icecap
XICEslow_h_n slow_h_n / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEen_cmos_b en_cmos_b / icecap
XICEnsw_en nsw_en / icecap
XI23<0> pd_h<3> / icecap
XI23<1> pd_h<2> / icecap
XI22<0> pu_h_n<3> / icecap
XI22<1> pu_h_n<2> / icecap
XICEpuen_h<0> puen_h<0> / icecap
XICEpden_h_n<1> pden_h_n<1> / icecap
XICEpu_h_n<1> pu_h_n<1> / icecap
xI19 vgnd_io vcc_io condiode
Xpu_strong_slow drvhi_h pu_h_n<1> puen_h<1> vcc_io vgnd_io / 
+ sky130_fd_io__com_pupredrvr_strong_slow
Xpu_weak drvhi_h pu_h_n<0> puen_h<0> vcc_io vgnd_io / 
+ sky130_fd_io__com_pupredrvr_weak
XI151 drvlo_h_n pd_h<0> pden_h_n<0> vcc_io vgnd_io / 
+ sky130_fd_io__com_pdpredrvr_weak
Xpd_strong_slow drvlo_h_n pd_h<1> en_cmos_b vcc_io vgnd_io / 
+ sky130_fd_io__com_pdpredrvr_strong_slow
XI150 drvlo_h_n drvlo_h_n en_cmos_b nsw_en pd_h<3> pd_h<2> pden_h_n<1> slow_h 
+ vcc_io vgnd_io / sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_cmos
Xpu_strong drvhi_h pu_h_n<3> pu_h_n<2> puen_h<1> slow_h_n vcc_io vgnd_io / 
+ sky130_fd_io__gpio_ovtv2_pupredrvr_strong
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_obpredrvr_leak_fix drvhi_h drvlo_h_n i2c_mode_h_n 
+ nghs_h oe_i_h_n pad pd_dis_h pd_h<3> pd_h<2> pd_h<1> pd_h<0> pden_h_n<1> 
+ pden_h_n<0> pghs_h pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> puen_h<1> 
+ puen_h<0> pug_h slew_ctl_h<1> slew_ctl_h<0> slew_ctl_h_n<1> slew_ctl_h_n<0> 
+ slow_h slow_h_n vcc_io vgnd_io vpb_drvr vssd
*.PININFO drvhi_h:I drvlo_h_n:I i2c_mode_h_n:I nghs_h:I oe_i_h_n:I pd_dis_h:I 
*.PININFO pden_h_n<1>:I pden_h_n<0>:I pghs_h:I puen_h<1>:I puen_h<0>:I pug_h:I 
*.PININFO slew_ctl_h<1>:I slew_ctl_h<0>:I slew_ctl_h_n<1>:I slew_ctl_h_n<0>:I 
*.PININFO slow_h:I slow_h_n:I vcc_io:I vgnd_io:I vpb_drvr:I vssd:I pd_h<3>:O 
*.PININFO pd_h<2>:O pd_h<1>:O pd_h<0>:O pu_h_n<3>:O pu_h_n<2>:O pu_h_n<1>:O 
*.PININFO pu_h_n<0>:O pad:B
XICEpad pad / icecap
XICEpden_h_n<1> pden_h_n<1> / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEdrvhi_h drvhi_h / icecap
XI375<0> pu_h_n<3> / icecap
XI375<1> pu_h_n<2> / icecap
XI375<2> pu_h_n<1> / icecap
XI375<3> pu_h_n<0> / icecap
XICEvssd vssd / icecap
XI374<0> pd_h<3> / icecap
XI374<1> pd_h<2> / icecap
XI374<2> pd_h<1> / icecap
XI374<3> pd_h<0> / icecap
XICEi2c_mode_h_n i2c_mode_h_n / icecap
XICEpug_h pug_h / icecap
XI376<0> puen_h<1> / icecap
XI376<1> puen_h<0> / icecap
XI377<0> pden_h_n<1> / icecap
XI377<1> pden_h_n<0> / icecap
XICEpd_dis_h pd_dis_h / icecap
XICEnsw_en nsw_en / icecap
XICEslow_h slow_h / icecap
XICEoe_i_h_n oe_i_h_n / icecap
XI380<0> slew_ctl_h_n<1> / icecap
XI380<1> slew_ctl_h_n<0> / icecap
XICEslow_h_n slow_h_n / icecap
XICEvpb_drvr vpb_drvr / icecap
XICEpghs_h pghs_h / icecap
XI379<0> pd_h<3> / icecap
XI379<1> pd_h<2> / icecap
XI378<0> slew_ctl_h<1> / icecap
XI378<1> slew_ctl_h<0> / icecap
XICEen_cmos_b en_cmos_b / icecap
XICEnghs_h nghs_h / icecap
XI192 drvlo_h_n en_cmos_b i2c_mode_h_n nghs_h nsw_en oe_i_h_n pad pd_dis_h 
+ pd_h<3> pd_h<2> pden_h_n<1> pghs_h pug_h slew_ctl_h<1> slew_ctl_h<0> 
+ slew_ctl_h_n<1> slew_ctl_h_n<0> slow_h_n vcc_io vgnd_io vpb_drvr vssd / 
+ sky130_fd_io__gpio_ovtv2_obpredrvr_new_leak_fix
XI191 drvhi_h drvlo_h_n en_cmos_b nsw_en pd_h<3> pd_h<2> pd_h<1> pd_h<0> 
+ pden_h_n<1> pden_h_n<0> pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> puen_h<1> 
+ puen_h<0> slow_h slow_h_n vcc_io vgnd_io / sky130_fd_io__gpio_ovtv2_obpredrvr_old
.ENDS
* .SUBCKT sky130_fd_io__gpio_dat_ls hld_h_n in out_h out_h_n rst_h set_h vcc_io vgnd 
* + vpwr_ka
* *.PININFO hld_h_n:I in:I rst_h:I set_h:I vcc_io:I vgnd:I vpwr_ka:I out_h:O 
* *.PININFO out_h_n:O
* XICEnet107 net107 / icecap
* XICEhld_h_n hld_h_n / icecap
* XICEset_h set_h / icecap
* XICEnet79 net79 / icecap
* XICEnet83 net83 / icecap
* XICEout_h out_h / icecap
* XICErst_h rst_h / icecap
* XICEnet103 net103 / icecap
* XICEin in / icecap
* XICEout_h_n out_h_n / icecap
* XICEin_i in_i / icecap
* XICEfbk fbk / icecap
* XICEin_i_n in_i_n / icecap
* XICEfbk_n fbk_n / icecap
* mI3 fbk fbk_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI4 fbk_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI5 fbk hld_h_n net79 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI6 fbk_n hld_h_n net83 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI7 net107 in_i_n vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=8 w=1.00 l=0.15 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI8 net103 in_i vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=8 w=1.00 l=0.15 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI12 out_h fbk_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI13 out_h_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mmnset fbk_n set_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mmnrst fbk rst_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI34 in_i_n in vgnd vgnd sky130_fd_pr__nfet_01v8 m=2 w=1.00 l=0.25 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI35 in_i in_i_n vgnd vgnd sky130_fd_pr__nfet_01v8 m=2 w=1.00 l=0.25 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI31 net83 vpwr_ka net103 vgnd sky130_fd_pr__nfet_05v0_nvt m=8 w=1.00 l=0.90 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI30 net79 vpwr_ka net107 vgnd sky130_fd_pr__nfet_05v0_nvt m=8 w=1.00 l=0.90 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI1 fbk_n fbk vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI2 fbk fbk_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI33 in_i in_i_n vpwr_ka vpwr_ka sky130_fd_pr__pfet_01v8_hvt m=1 w=3.00 l=0.25 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI11 out_h fbk_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI14 out_h_n fbk vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI32 in_i_n in vpwr_ka vpwr_ka sky130_fd_pr__pfet_01v8_hvt m=1 w=3.00 l=0.25 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__com_cclat_hvnor3 in0 in1 in2 out vcc_io vgnd vnb
* *.PININFO in0:I in1:I in2:I vcc_io:I vgnd:I vnb:I out:O
* XICEin0 in0 / icecap
* XICEin2 in2 / icecap
* XICEout out / icecap
* XICEn<1> n<1> / icecap
* XICEin1 in1 / icecap
* XICEn<0> n<0> / icecap
* mmp0 n<0> in0 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mmp2 out in2 n<1> vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mmp1 n<1> in1 n<0> vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mmn0 out in0 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mmn2 out in2 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mmn1 out in1 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__com_cclat_hvnand3 in0 in1 in2 out vcc_io vgnd vnb
* *.PININFO in0:I in1:I in2:I vcc_io:I vgnd:I vnb:I out:O
* XICEin0 in0 / icecap
* XICEn0 n0 / icecap
* XICEin2 in2 / icecap
* XICEin1 in1 / icecap
* XICEout out / icecap
* XICEn1 n1 / icecap
* mmp0 out in0 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mmp2 out in2 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mmp1 out in1 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mmn2 out in2 n1 vnb sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 sa=265e-3 sb=265e-3 sd=280e-3 
* + topography=normal perim=1.14
* mmn0 n0 in0 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=4 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mmn1 n1 in1 n0 vnb sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 sa=265e-3 sb=265e-3 sd=280e-3 
* + topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__com_cclat_inv_in in out vcc_io vgnd vnb
* *.PININFO in:I vcc_io:I vgnd:I vnb:I out:O
* XICEin in / icecap
* XICEout out / icecap
* mmp1 out in vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mmn1 out in vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__com_cclat_inv_out in out vcc_io vgnd vnb
* *.PININFO in:I vcc_io:I vgnd:I vnb:I out:O
* XICEin in / icecap
* XICEout out / icecap
* mI1 out in vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=6 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI2 out in vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=6 w=3.00 l=0.60 sa=265e-3 sb=265e-3 sd=280e-3 
* + topography=normal perim=1.14
* .ENDS
.SUBCKT sky130_fd_io__com_cclat_i2c_fix drvhi_h drvlo_h_n oe_h pd_dis_h pu_dis_h 
+ vcc_io vgnd
*.PININFO oe_h:I pd_dis_h:I pu_dis_h:I vcc_io:I vgnd:I drvhi_h:O drvlo_h_n:O
XICEpd_dis_h pd_dis_h / icecap
XICEoe_h oe_h / icecap
XICEdrvhi_h drvhi_h / icecap
XICEn0 n0 / icecap
XICEn1 n1 / icecap
XICEoe_i_h_n oe_i_h_n / icecap
XICEpu_dis_h pu_dis_h / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEpu_dis_h_n pu_dis_h_n / icecap
Xnor3 oe_i_h_n drvhi_h pd_dis_h n1 vcc_io vgnd vgnd / sky130_fd_io__com_cclat_hvnor3
Xnand3 oe_h drvlo_h_n pu_dis_h_n n0 vcc_io vgnd vgnd / 
+ sky130_fd_io__com_cclat_hvnand3
Xinv_oe2 oe_h oe_i_h_n vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_in
Xinv_pudis pu_dis_h pu_dis_h_n vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_in
Xinv_out n1 drvlo_h_n vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_out
Xinv_out_1 n0 drvhi_h vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_out
.ENDS
* .SUBCKT sky130_fd_io__hvsbt_inv_x1 in out vgnd vpwr
* *.PININFO in:I vgnd:I vpwr:I out:O
* XICEin in / icecap
* XICEout out / icecap
* mI1 out in vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI2 out in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
.SUBCKT sky130_fd_io__gpio_dat_ls_i2c_fix hld_h_n in out_h_n set_h set_h_n vcc_io 
+ vgnd vpwr_ka
*.PININFO hld_h_n:I in:I set_h:I set_h_n:I vcc_io:I vgnd:I vpwr_ka:I out_h_n:O
XICEnet76 net76 / icecap
XICEin_i_n in_i_n / icecap
XICEset_h set_h / icecap
XICEin in / icecap
XICEnet96 net96 / icecap
XICEout_h_n out_h_n / icecap
XICEhld_h_n hld_h_n / icecap
XICEnet100 net100 / icecap
XICEfbk_n fbk_n / icecap
XICEfbk fbk / icecap
XICEin_i in_i / icecap
XICEnet80 net80 / icecap
XICEset_h_n set_h_n / icecap
mI3 fbk fbk_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI4 fbk_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI5 fbk hld_h_n net76 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI6 fbk_n hld_h_n net80 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI7 net100 in_i_n vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=8 w=1.00 l=0.15 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI8 net96 in_i vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=8 w=1.00 l=0.15 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI13 out_h_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mmnset fbk_n set_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=4 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI34 in_i_n in vgnd vgnd sky130_fd_pr__nfet_01v8 m=2 w=1.00 l=0.25 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI35 in_i in_i_n vgnd vgnd sky130_fd_pr__nfet_01v8 m=2 w=1.00 l=0.25 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI31 net80 vpwr_ka net96 vgnd sky130_fd_pr__nfet_05v0_nvt m=8 w=1.00 l=0.90 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI30 net76 vpwr_ka net100 vgnd sky130_fd_pr__nfet_05v0_nvt m=8 w=1.00 l=0.90 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI1 fbk_n fbk vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI2 fbk fbk_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI33 in_i in_i_n vpwr_ka vpwr_ka sky130_fd_pr__pfet_01v8_hvt m=1 w=3.00 l=0.25 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI14 out_h_n fbk vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI36 fbk set_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI32 in_i_n in vpwr_ka vpwr_ka sky130_fd_pr__pfet_01v8_hvt m=1 w=3.00 l=0.25 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_opath_datoe_i2c_fix drvhi_h drvlo_h_n hld_h_n 
+ hld_i_ovr_h od_i_h_n oe_h oe_n out pd_dis_h vcc_io vgnd vpwr_ka
*.PININFO hld_h_n:I hld_i_ovr_h:I od_i_h_n:I oe_n:I out:I vcc_io:I vgnd:I 
*.PININFO vpwr_ka:I drvhi_h:O drvlo_h_n:O oe_h:O pd_dis_h:O
XICEhld_h_n hld_h_n / icecap
XICEnet56 net56 / icecap
XICEoe_h oe_h / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEout out / icecap
XICEhld_i_ovr_h hld_i_ovr_h / icecap
XICEpu_dis_h pu_dis_h / icecap
XICEpd_dis_h pd_dis_h / icecap
XICEdrvhi_h drvhi_h / icecap
XICEod_i_h_n od_i_h_n / icecap
XICEnet60 net60 / icecap
XICEoe_n oe_n / icecap
Xdat_ls hld_i_ovr_h out pd_dis_h pu_dis_h vgnd net60 vcc_io vgnd vpwr_ka / 
+ sky130_fd_io__gpio_dat_ls
Xcclat drvhi_h drvlo_h_n oe_h pd_dis_h pu_dis_h vcc_io vgnd / 
+ sky130_fd_io__com_cclat_i2c_fix
XI36 od_i_h_n net60 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI37 od_i_h_n net56 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
Xoe_ls hld_i_ovr_h oe_n oe_h net56 od_i_h_n vcc_io vgnd vpwr_ka / 
+ sky130_fd_io__gpio_dat_ls_i2c_fix
.ENDS
* .SUBCKT sky130_fd_io__hvsbt_nor in0 in1 out vgnd vpwr
* *.PININFO in0:I in1:I vgnd:I vpwr:I out:O
* mI3 net16 in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI12 out in1 net16 vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI1 out in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI6 out in1 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__hvsbt_xor in0 in1 out vgnd vpwr
* *.PININFO in0:I in1:I vgnd:I vpwr:I out:O
* XICEin0 in0 / icecap
* XICEin1 in1 / icecap
* XICEout out / icecap
* XICEnet54 net54 / icecap
* XICEnet29 net29 / icecap
* XICEnet70 net70 / icecap
* XICEnet45 net45 / icecap
* mI3 net29 in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI5 out net54 net45 vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI17 net70 in1 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI18 net54 in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI13 net45 in1 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI12 out net70 net29 vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI1 out in1 net58 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI16 net70 in1 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI6 out net70 net62 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI15 net62 net54 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI14 net58 in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI19 net54 in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__hvsbt_inv_x2 in out vgnd vpwr
* *.PININFO in:I vgnd:I vpwr:I out:O
* XICEout out / icecap
* XICEin in / icecap
* mI2 out in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI1 out in vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__com_ctl_ls hld_h_n in out_h out_h_n rst_h set_h vcc_io vgnd 
* + vpwr
* *.PININFO hld_h_n:I in:I rst_h:I set_h:I vcc_io:I vgnd:I vpwr:I out_h:O 
* *.PININFO out_h_n:O
* XICEout_h_n out_h_n / icecap
* XICEset_h set_h / icecap
* XICEfbk_n fbk_n / icecap
* XICErst_h rst_h / icecap
* XICEnet122 net122 / icecap
* XICEnet130 net130 / icecap
* XICEnet94 net94 / icecap
* XICEhld_h_n hld_h_n / icecap
* XICEfbk fbk / icecap
* XICEout_h out_h / icecap
* XICEnet98 net98 / icecap
* XICEin in / icecap
* XICEin_i in_i / icecap
* XICEin_i_n in_i_n / icecap
* mI14 out_h_n fbk vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI34 in_i in_i_n vpwr vpwr sky130_fd_pr__pfet_01v8_hvt m=1 w=1.00 l=0.25 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI29 in_i_n in vpwr vpwr sky130_fd_pr__pfet_01v8_hvt m=1 w=1.00 l=0.25 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI11 out_h fbk_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI2 fbk fbk_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI1 fbk_n fbk vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI13 out_h_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mmnset fbk_n set_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI32 in_i in_i_n vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.25 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI12 out_h fbk_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI58 net130 vpwr net94 vgnd sky130_fd_pr__nfet_05v0_nvt m=4 w=1.00 l=0.90 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmnrst fbk rst_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI59 net122 vpwr net98 vgnd sky130_fd_pr__nfet_05v0_nvt m=4 w=1.00 l=0.90 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI6 fbk_n hld_h_n net122 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI27 in_i_n in vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.25 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI5 fbk hld_h_n net130 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI4 fbk_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI3 fbk fbk_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI8 net98 in_i vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=4 w=1.00 l=0.15 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI7 net94 in_i_n vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=4 w=1.00 l=0.15 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_octl_i2c_fix dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> 
+ dm_h_n<1> dm_h_n<0> hld_i_h_n od_i_h_n pden_h_n<2> pden_h_n<1> pden_h_n<0> 
+ puen_0_h puen_2or1_h puen_h<1> puen_h<0> slow slow_h slow_h_n vcc_io vgnd 
+ vpwr vreg_en_h_n
*.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I 
*.PININFO hld_i_h_n:I od_i_h_n:I slow:I vcc_io:I vgnd:I vpwr:I vreg_en_h_n:I 
*.PININFO pden_h_n<2>:O pden_h_n<1>:O pden_h_n<0>:O puen_0_h:O puen_2or1_h:O 
*.PININFO puen_h<1>:O puen_h<0>:O slow_h:O slow_h_n:O
XI211 n<8> dm_h_n<1> puen_0_h vgnd vcc_io / sky130_fd_io__hvsbt_nor
XI201 dm_h_n<2> dm_h_n<1> n<9> vgnd vcc_io / sky130_fd_io__hvsbt_nor
XI366 dm_h<1> dm_h<0> net87 vgnd vcc_io / sky130_fd_io__hvsbt_nor
XI210 dm_h<2> dm_h<0> n<8> vgnd vcc_io / sky130_fd_io__hvsbt_xor
XI200 dm_h<2> dm_h<1> n<10> vgnd vcc_io / sky130_fd_io__hvsbt_xor
XI185 dm_h_n<0> n<4> net207 vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI186 dm_h_n<2> dm_h_n<1> n<4> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI187 dm_h<1> dm_h<0> n<3> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI208 puen_2or1_h vreg_en_h_n n<5> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI203 n<10> dm_h<0> n<1> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI204 n<9> dm_h_n<0> n<0> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI205 n<1> n<0> puen_2or1_h vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI365 net87 dm_h<2> pden_h_n<2> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI254 puen_h1_n puen_h<1> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
XI256 puen_h0_n puen_h<0> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
XI249 pden_h0 pden_h_n<0> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
XI247 pden_h1 pden_h_n<1> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
XI377 puen_0_h puen_h0_n vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI209 n<5> n<2> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI376 n<2> puen_h1_n vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI374 net207 pden_h1 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI375 n<3> pden_h0 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI381 od_i_h_n n9 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
Xls_slow hld_i_h_n slow slow_h slow_h_n n9 vgnd vcc_io vgnd vpwr / 
+ sky130_fd_io__com_ctl_ls
XICEn<0> n<0> / icecap
XICEn<4> n<4> / icecap
XICEpuen_2or1_h puen_2or1_h / icecap
XICEdm_h<2> dm_h<2> / icecap
XICEpden_h1 pden_h1 / icecap
XICEn<10> n<10> / icecap
XICEslow_h_n slow_h_n / icecap
XICEdm_h_n<1> dm_h_n<1> / icecap
XICEpden_h0 pden_h0 / icecap
XICEdm_h<1> dm_h<1> / icecap
XICEn<8> n<8> / icecap
XICEslow slow / icecap
XICEdm_h<0> dm_h<0> / icecap
XICEpden_h_n<1> pden_h_n<1> / icecap
XICEn<9> n<9> / icecap
XICEpuen_0_h puen_0_h / icecap
XICEpuen_h1_n puen_h1_n / icecap
XICEpuen_h<0> puen_h<0> / icecap
XICEpuen_h0_n puen_h0_n / icecap
XICEdm_h_n<2> dm_h_n<2> / icecap
XICEhld_i_h_n hld_i_h_n / icecap
XICEnet177 net207 / icecap
XICEn<3> n<3> / icecap
XICEvreg_en_h_n vreg_en_h_n / icecap
XICEdm_h_n<0> dm_h_n<0> / icecap
XICEpden_h_n<0> pden_h_n<0> / icecap
XICEn<1> n<1> / icecap
XICEn<2> n<2> / icecap
XICEpuen_h<1> puen_h<1> / icecap
XICEslow_h slow_h / icecap
XICEn<5> n<5> / icecap
XICEnet198 net87 / icecap
.ENDS
.SUBCKT sky130_fd_io__sio_hvsbt_inv_x2 in out vgnd vnb vpb vpwr
*.PININFO in:I vgnd:I vnb:I vpb:I vpwr:I out:O
XICEin in / icecap
XICEout out / icecap
mI1 out in vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.60 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal perim=1.14
mI2 out in vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.60 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_octl_dat_i2c_fix_leak_fix dm_h<2> dm_h<1> dm_h<0> 
+ dm_h_n<2> dm_h_n<1> dm_h_n<0> drvhi_h hld_i_h_n hld_i_ovr_h nghs_h od_i_h_n 
+ oe_hs_h oe_n out pad pd_h<3> pd_h<2> pd_h<1> pd_h<0> pghs_h pu_h_n<3> 
+ pu_h_n<2> pu_h_n<1> pu_h_n<0> pug_h slew_ctl_h<1> slew_ctl_h<0> 
+ slew_ctl_h_n<1> slew_ctl_h_n<0> slow slow_h_n vccd vddio vpb_drvr vpwr_ka 
+ vssd vssio
*.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I 
*.PININFO hld_i_h_n:I hld_i_ovr_h:I nghs_h:I od_i_h_n:I oe_n:I out:I pghs_h:I 
*.PININFO pug_h:I slew_ctl_h<1>:I slew_ctl_h<0>:I slew_ctl_h_n<1>:I 
*.PININFO slew_ctl_h_n<0>:I slow:I vccd:I vddio:I vpb_drvr:I vpwr_ka:I vssd:I 
*.PININFO vssio:I drvhi_h:O oe_hs_h:O pd_h<3>:O pd_h<2>:O pd_h<1>:O pd_h<0>:O 
*.PININFO pu_h_n<3>:O pu_h_n<2>:O pu_h_n<1>:O pu_h_n<0>:O slow_h_n:O pad:B
XI425<0> pd_h<3> / icecap
XI425<1> pd_h<2> / icecap
XI425<2> pd_h<1> / icecap
XI425<3> pd_h<0> / icecap
XICEpden_h_n<2> pden_h_n<2> / icecap
XICEoe_h oe_h / icecap
XICEvpb_drvr vpb_drvr / icecap
XICEod_i_h_n od_i_h_n / icecap
XI431<0> pden_h_n<1> / icecap
XI431<1> pden_h_n<0> / icecap
XICEoe_hs_i_h_n oe_hs_i_h_n / icecap
XICEoe_hs_i_h oe_hs_i_h / icecap
XICEhld_i_ovr_h hld_i_ovr_h / icecap
XICEn<1> n<1> / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEslow_h_n slow_h_n / icecap
XICEnghs_h nghs_h / icecap
XI422<0> pu_h_n<3> / icecap
XI422<1> pu_h_n<2> / icecap
XI422<2> pu_h_n<1> / icecap
XI422<3> pu_h_n<0> / icecap
XI424<0> dm_h<2> / icecap
XI424<1> dm_h<1> / icecap
XI424<2> dm_h<0> / icecap
XI430<0> puen_h<1> / icecap
XI430<1> puen_h<0> / icecap
XI423<0> pd_h<3> / icecap
XI423<1> pd_h<2> / icecap
XI423<2> pd_h<1> / icecap
XI423<3> pd_h<0> / icecap
XICEnet85 net85 / icecap
XICEpad pad / icecap
XI429<0> pu_h_n<3> / icecap
XI429<1> pu_h_n<2> / icecap
XI429<2> pu_h_n<1> / icecap
XI429<3> pu_h_n<0> / icecap
XI432<0> slew_ctl_h_n<1> / icecap
XI432<1> slew_ctl_h_n<0> / icecap
XICEdrvhi_h drvhi_h / icecap
XI426<0> dm_h_n<2> / icecap
XI426<1> dm_h_n<1> / icecap
XI426<2> dm_h_n<0> / icecap
XICEoe_i_h_n oe_i_h_n / icecap
XICEslow_h slow_h / icecap
XICEoe_n oe_n / icecap
XICEpug_h pug_h / icecap
XICEnet86 net86 / icecap
XICEslow slow / icecap
XICEhld_i_h_n hld_i_h_n / icecap
XICEoe_hs_h oe_hs_h / icecap
XICEpghs_h pghs_h / icecap
XICEnet72 net72 / icecap
XI427<0> slew_ctl_h<1> / icecap
XI427<1> slew_ctl_h<0> / icecap
XICEout out / icecap
XI428<0> pden_h_n<2> / icecap
XI428<1> pden_h_n<1> / icecap
XI428<2> pden_h_n<0> / icecap
Xpredrvr drvhi_h drvlo_h_n pden_h_n<2> nghs_h oe_i_h_n pad net72 pd_h<3> 
+ pd_h<2> pd_h<1> pd_h<0> pden_h_n<1> pden_h_n<0> pghs_h pu_h_n<3> pu_h_n<2> 
+ pu_h_n<1> pu_h_n<0> puen_h<1> puen_h<0> pug_h slew_ctl_h<1> slew_ctl_h<0> 
+ slew_ctl_h_n<1> slew_ctl_h_n<0> slow_h slow_h_n vddio vssio vpb_drvr vssd / 
+ sky130_fd_io__gpio_ovtv2_obpredrvr_leak_fix
Xdatoe drvhi_h drvlo_h_n hld_i_h_n hld_i_ovr_h od_i_h_n oe_h oe_n out net72 
+ vddio vssd vpwr_ka / sky130_fd_io__gpio_ovtv2_opath_datoe_i2c_fix
Xctl dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n od_i_h_n 
+ pden_h_n<2> pden_h_n<1> pden_h_n<0> net86 net85 puen_h<1> puen_h<0> slow 
+ slow_h slow_h_n vddio vssd vccd vddio / sky130_fd_io__gpio_ovtv2_octl_i2c_fix
XI354 oe_hs_i_h oe_hs_i_h_n vssd vssd vddio vddio / sky130_fd_io__sio_hvsbt_inv_x1
XI353 oe_h oe_i_h_n vssd vssd vddio vddio / sky130_fd_io__sio_hvsbt_inv_x2
XI355 oe_hs_i_h_n oe_hs_h vssd vssd vddio vddio / sky130_fd_io__sio_hvsbt_inv_x2
XI351 net86 net85 n<1> vssd vssd vddio vddio / sky130_fd_io__sio_hvsbt_nor
XI352 n<1> oe_i_h_n oe_hs_i_h vssd vssd vddio vddio / sky130_fd_io__sio_hvsbt_nor
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_opath_i2c_fix_leak_fix dm_h<2> dm_h<1> dm_h<0> 
+ dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n hld_i_ovr_h nga_pad_vpmp_h 
+ ngb_pad_vpmp_h od_i_h_n oe_n out pad pd_csd_h pghs_h pu_csd_h pug_h<6> 
+ pug_h<5> slew_ctl_h<1> slew_ctl_h<0> slew_ctl_h_n<1> slew_ctl_h_n<0> slow 
+ tie_hi_esd tie_lo_esd vccd vddio vddio_amx vpb_drvr vpwr_ka vssa vssd vssio 
+ vssio_amx
*.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I 
*.PININFO hld_i_h_n:I hld_i_ovr_h:I nga_pad_vpmp_h:I ngb_pad_vpmp_h:I 
*.PININFO od_i_h_n:I oe_n:I out:I pd_csd_h:I pu_csd_h:I slew_ctl_h<1>:I 
*.PININFO slew_ctl_h<0>:I slew_ctl_h_n<1>:I slew_ctl_h_n<0>:I slow:I vccd:I 
*.PININFO vddio:I vpwr_ka:I vssa:I vssd:I vssio:I vssio_amx:I pad:O pghs_h:O 
*.PININFO tie_hi_esd:O tie_lo_esd:O pug_h<6>:B pug_h<5>:B vddio_amx:B 
*.PININFO vpb_drvr:B
Xodrvr tie_lo_esd nga_pad_vpmp_h ngb_pad_vpmp_h nghs_h od_i_h_n oe_hs_h pad 
+ pd_csd_h pd_h<3> pd_h<2> pd_h<1> pd_h<0> pghs_h pu_csd_h pu_h_n<3> pu_h_n<2> 
+ pu_h_n<1> pu_h_n<0> pug_h<7> pug_h<6> pug_h<5> tie_hi_esd tie_lo_esd vddio 
+ vddio_amx vpb_drvr vssa vssd vssio vssio_amx / 
+ sky130_fd_io__gpio_ovtv2_odrvr_i2c_fix_leak_fix
Xopath dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> drvhi_h hld_i_h_n 
+ hld_i_ovr_h nghs_h od_i_h_n oe_hs_h oe_n out pad pd_h<3> pd_h<2> pd_h<1> 
+ pd_h<0> pghs_h pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> pug_h<7> 
+ slew_ctl_h<1> slew_ctl_h<0> slew_ctl_h_n<1> slew_ctl_h_n<0> slow slow_h_n 
+ vccd vddio vpb_drvr vpwr_ka vssd vssio / 
+ sky130_fd_io__gpio_ovtv2_octl_dat_i2c_fix_leak_fix
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_ctl_ls_i2c_fix in in_b out_h rst_h rst_h_n vgnd 
+ vpwr_hv vpwr_lv
*.PININFO in:I in_b:I rst_h:I rst_h_n:I vgnd:I vpwr_hv:I vpwr_lv:I out_h:O
XICEnet70 net70 / icecap
XICEnet75 net75 / icecap
XICErst_h_n rst_h_n / icecap
XICEfbk_n fbk_n / icecap
XICEin in / icecap
XICEnet71 net71 / icecap
XICEin_b in_b / icecap
XICEout_h out_h / icecap
XICErst_h rst_h / icecap
XICEfbk fbk / icecap
mI14 fbk_n rst_h_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=2 w=0.75 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI11 out_h fbk_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=2 w=0.75 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI2 fbk_n fbk vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI1 fbk fbk_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI5 net70 rst_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=4 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI12 out_h fbk_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI58 fbk vpwr_lv net71 vgnd sky130_fd_pr__nfet_05v0_nvt m=4 w=1.00 l=0.90 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mmnrst fbk rst_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.50 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI59 fbk_n vpwr_lv net75 vgnd sky130_fd_pr__nfet_05v0_nvt m=4 w=1.00 l=0.90 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI8 net75 in net70 vgnd sky130_fd_pr__nfet_01v8_lvt m=4 w=1.00 l=0.15 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI7 net71 in_b net70 vgnd sky130_fd_pr__nfet_01v8_lvt m=4 w=1.00 l=0.15 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
* .SUBCKT sky130_fd_io__gpiov2_amux_ls_inv_x1 in out vgnd vpwr
* *.PININFO in:I vgnd:I vpwr:I out:O
* XICEout out / icecap
* XICEin in / icecap
* mI2 out in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI1 out in vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_amux_ctl_lshv2hv in in_b out_h out_h_n rst_h rst_h_n 
* + vgnd vpwr_hv
* *.PININFO in:I in_b:I rst_h:I rst_h_n:I vgnd:I vpwr_hv:I out_h:O out_h_n:O
* XICEnet64 net64 / icecap
* XICEin in / icecap
* XICErst_h_n rst_h_n / icecap
* XICEout_h out_h / icecap
* XICEfbk fbk / icecap
* XICEin_b in_b / icecap
* XICEfbk_n fbk_n / icecap
* XICErst_h rst_h / icecap
* XICEout_h_n out_h_n / icecap
* mI14 out_h_n fbk vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI11 out_h fbk_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI2 fbk fbk_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI1 fbk_n fbk vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI64 net64 rst_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI13 out_h_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI12 out_h fbk_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mmnrst fbk rst_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI8 fbk_n in net64 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI7 fbk in_b net64 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_amux_ctl_inv_1 in out vgnd vpwr
* *.PININFO in:I vgnd:I vpwr:I out:O
* XICEout out / icecap
* XICEin in / icecap
* mI27 out in vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI29 out in vpwr vpwr sky130_fd_pr__pfet_01v8_hvt m=1 w=1.00 l=0.25 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_ls_i2c_fix amux_en_vdda_h amux_en_vdda_h_n 
+ amux_en_vddio_h amux_en_vswitch_h amux_en_vswitch_h_n analog_en 
+ enable_vdda_h enable_vdda_h_n enable_vswitch_h hld_i_h_n vccd vdda vddio_q 
+ vssa vssd vswitch
*.PININFO analog_en:I enable_vdda_h:I enable_vswitch_h:I hld_i_h_n:I vccd:I 
*.PININFO vdda:I vddio_q:I vssa:I vssd:I vswitch:I amux_en_vdda_h:O 
*.PININFO amux_en_vdda_h_n:O amux_en_vddio_h:O amux_en_vswitch_h:O 
*.PININFO amux_en_vswitch_h_n:O enable_vdda_h_n:O
XICEamux_en_vswitch_h amux_en_vswitch_h / icecap
XICEanalog_en analog_en / icecap
XICEnet028 net028 / icecap
XICEhld_i_h_n hld_i_h_n / icecap
XICEamux_en_vdda_h_n amux_en_vdda_h_n / icecap
XICEamux_en_vswitch_h_n amux_en_vswitch_h_n / icecap
XICEnet83 net83 / icecap
XICEana_en_i_n ana_en_i_n / icecap
XICEnet082 net082 / icecap
XICEamux_en_vddio_h amux_en_vddio_h / icecap
XICEenable_vdda_h_n enable_vdda_h_n / icecap
XICEana_en_i ana_en_i / icecap
XICEenable_vswitch_h enable_vswitch_h / icecap
XICEenable_vdda_h enable_vdda_h / icecap
XICEamux_en_vdda_h amux_en_vdda_h / icecap
Xpd_vddio_ls ana_en_i ana_en_i_n amux_en_vddio_h net082 hld_i_h_n vssd vddio_q 
+ vccd / sky130_fd_io__gpiov2_amux_ctl_ls_i2c_fix
XI32 enable_vdda_h enable_vdda_h_n vssa vdda / sky130_fd_io__gpiov2_amux_ls_inv_x1
Xpd_vswitch_ls amux_en_vddio_h net028 amux_en_vswitch_h amux_en_vswitch_h_n 
+ net83 enable_vswitch_h vssa vswitch / sky130_fd_io__gpiov2_amux_ctl_lshv2hv
Xpd_vdda_ls amux_en_vddio_h net028 amux_en_vdda_h amux_en_vdda_h_n 
+ enable_vdda_h_n enable_vdda_h vssa vdda / sky130_fd_io__gpiov2_amux_ctl_lshv2hv
XI15 analog_en ana_en_i_n vssd vccd / sky130_fd_io__gpiov2_amux_ctl_inv_1
XI16 ana_en_i_n ana_en_i vssd vccd / sky130_fd_io__gpiov2_amux_ctl_inv_1
XI18 enable_vswitch_h net83 vssa vswitch / sky130_fd_io__hvsbt_inv_x1
XI36 amux_en_vddio_h net028 vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI35 hld_i_h_n net082 vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3_ver2 in in_b out_h out_h_n 
+ rst2_h rst2_h_n rst_h rst_h_n vgnd vpwr_hv vpwr_lv
*.PININFO in:I in_b:I rst2_h:I rst2_h_n:I rst_h:I rst_h_n:I vgnd:I vpwr_hv:I 
*.PININFO vpwr_lv:I out_h:O out_h_n:O
XICEin_b in_b / icecap
XICEnet76 net76 / icecap
XICEout_h out_h / icecap
XICEnet56 net56 / icecap
XICErst_h rst_h / icecap
XICErst2_h_n rst2_h_n / icecap
XICErst_h_n rst_h_n / icecap
XICEnet52 net52 / icecap
XICEin in / icecap
XICEout_h_n out_h_n / icecap
XICErst2_h rst2_h / icecap
XICEnet72 net72 / icecap
mI11 out_h_n out_h vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI9 out_h out_h_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI29 out_h_n rst2_h_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.50 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI28 out_h_n rst_h_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI21 net56 vpwr_lv net76 vgnd sky130_fd_pr__nfet_05v0_nvt m=2 w=1.00 l=0.90 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI20 net52 vpwr_lv net72 vgnd sky130_fd_pr__nfet_05v0_nvt m=2 w=1.00 l=0.90 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI17 out_h rst_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI6 net76 in vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=2 w=1.00 l=0.15 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI12 net72 in_b vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=2 w=1.00 l=0.15 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI31 out_h rst2_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.50 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI25 out_h rst_h_n net52 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI24 out_h_n rst_h_n net56 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amx_pucsd_buf A Y vda vssa
*.PININFO A:I vda:I vssa:I Y:O
XICEA A / icecap
XICEY Y / icecap
XICEint int / icecap
mI75 int A vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=4 w=0.42 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI6 Y int vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=3 w=0.42 l=0.60 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal perim=1.14
mI74 int A vda vda sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal perim=1.14
mI5 Y int vda vda sky130_fd_pr__pfet_g5v0d10v5 m=5 w=1.00 l=0.60 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3 in in_b out_h out_h_n rst2_h_n 
+ rst_h_n vgnd vpwr_hv vpwr_lv
*.PININFO in:I in_b:I rst2_h_n:I rst_h_n:I vgnd:I vpwr_hv:I vpwr_lv:I out_h:O 
*.PININFO out_h_n:O
XICEout_h_n out_h_n / icecap
XICErst2_h_n rst2_h_n / icecap
XICErst_h_n rst_h_n / icecap
XICEnet074 net074 / icecap
XICEout_h out_h / icecap
XICEnet75 net75 / icecap
XICEnet51 net51 / icecap
XICEnet086 net086 / icecap
XICEin in / icecap
XICEnet55 net55 / icecap
XICEin_b in_b / icecap
XICEnet79 net79 / icecap
XI34 rst_h_n net086 vgnd vpwr_hv / sky130_fd_io__hvsbt_inv_x1
XI33 rst2_h_n net074 vgnd vpwr_hv / sky130_fd_io__hvsbt_inv_x1
mI11 out_h_n out_h vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI9 out_h out_h_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI29 out_h_n rst2_h_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.50 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI28 out_h_n rst_h_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI21 net55 vpwr_lv net79 vgnd sky130_fd_pr__nfet_05v0_nvt m=2 w=1.00 l=0.90 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI20 net51 vpwr_lv net75 vgnd sky130_fd_pr__nfet_05v0_nvt m=2 w=1.00 l=0.90 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI17 out_h net086 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI6 net79 in vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=2 w=1.00 l=0.15 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI12 net75 in_b vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=2 w=1.00 l=0.15 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI31 out_h net074 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.50 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI25 out_h rst_h_n net51 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI24 out_h_n rst_h_n net55 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
* .SUBCKT sky130_fd_io__gpiov2_amux_drvr_lshv2hv in in_b out_h_n rst_h rst_h_n vgnd 
* + vpwr_hv
* *.PININFO in:I in_b:I rst_h:I rst_h_n:I vgnd:I vpwr_hv:I out_h_n:O
* XICErst_h rst_h / icecap
* XICEout_h_n out_h_n / icecap
* XICEin in / icecap
* XICEfbk fbk / icecap
* XICEin_b in_b / icecap
* XICEnet52 net52 / icecap
* XICEfbk_n fbk_n / icecap
* XICErst_h_n rst_h_n / icecap
* mI14 out_h_n fbk vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI2 fbk fbk_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI1 fbk_n fbk vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI64 net52 rst_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI13 out_h_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mmnrst fbk rst_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI8 fbk_n in net52 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI7 fbk in_b net52 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_amx_inv4 A Y vda vssa
* *.PININFO A:I vda:I vssa:I Y:O
* XICEA A / icecap
* XICEY Y / icecap
* mI75 Y A vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=0.42 l=0.60 sa=265e-3 sb=265e-3 sd=280e-3 
* + topography=normal perim=1.14
* mI74 Y A vda vda sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 sa=265e-3 sb=265e-3 sd=280e-3 
* + topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_amx_pdcsd_inv A Y vda vssa
* *.PININFO A:I vda:I vssa:I Y:O
* XICEA A / icecap
* XICEY Y / icecap
* mI414 Y A vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 sa=265e-3 sb=265e-3 sd=280e-3 
* + topography=normal perim=1.14
* mI519 Y vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI517 Y A vda vda sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=2.00 sa=265e-3 sb=265e-3 sd=280e-3 
* + topography=normal perim=1.14
* mI429 Y A vda vda sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=2.00 sa=265e-3 sb=265e-3 sd=280e-3 
* + topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__amx_inv1 A Y vda vssa
* *.PININFO A:I vda:I vssa:I Y:O
* XICEA A / icecap
* XICEY Y / icecap
* mI92 Y A vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 sa=265e-3 sb=265e-3 sd=280e-3 
* + topography=normal perim=1.14
* mI54 Y A vda vda sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 sa=265e-3 sb=265e-3 sd=280e-3 
* + topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_amux_drvr_ls in in_b out_h out_h_n rst_h rst_h_n vgnd 
* + vpwr_hv vpwr_lv
* *.PININFO in:I in_b:I rst_h:I rst_h_n:I vgnd:I vpwr_hv:I vpwr_lv:I out_h:O 
* *.PININFO out_h_n:O
* XICEin_b in_b / icecap
* XICErst_h_n rst_h_n / icecap
* XICEnet42 net42 / icecap
* XICErst_h rst_h / icecap
* XICEnet38 net38 / icecap
* XICEin in / icecap
* XICEnet54 net54 / icecap
* XICEout_h_n out_h_n / icecap
* XICEout_h out_h / icecap
* XICEnet58 net58 / icecap
* mI11 out_h_n out_h vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI9 out_h out_h_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI21 net42 vpwr_lv net58 vgnd sky130_fd_pr__nfet_05v0_nvt m=2 w=1.00 l=0.90 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI20 net38 vpwr_lv net54 vgnd sky130_fd_pr__nfet_05v0_nvt m=2 w=1.00 l=0.90 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI17 out_h rst_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI6 net58 in vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=2 w=1.00 l=0.15 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI12 net54 in_b vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=2 w=1.00 l=0.15 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI25 out_h rst_h_n net38 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI24 out_h_n rst_h_n net42 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* .ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_drvr_i2c_fix amux_en_vdda_h amux_en_vdda_h_n 
+ amux_en_vddio_h amux_en_vswitch_h amux_en_vswitch_h_n amuxbusa_on 
+ amuxbusa_on_n amuxbusb_on amuxbusb_on_n hld_i_h_n nga_amx_vswitch_h 
+ nga_pad_vswitch_h nga_pad_vswitch_h_n ngb_amx_vswitch_h ngb_pad_vswitch_h 
+ ngb_pad_vswitch_h_n nmida_on_n nmida_vccd nmida_vccd_n nmidb_on_n nmidb_vccd 
+ nmidb_vccd_n pd_csd_vswitch_h pd_csd_vswitch_h_n pd_on pd_on_n 
+ pga_amx_vdda_h_n pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n 
+ pu_csd_vddioq_h_n pu_on pu_on_n vccd vdda vddio_q vssa vssd vswitch
*.PININFO amux_en_vdda_h:I amux_en_vdda_h_n:I amux_en_vddio_h:I 
*.PININFO amux_en_vswitch_h:I amux_en_vswitch_h_n:I amuxbusa_on:I 
*.PININFO amuxbusa_on_n:I amuxbusb_on:I amuxbusb_on_n:I hld_i_h_n:I 
*.PININFO nmida_on_n:I nmidb_on_n:I pd_on:I pd_on_n:I pu_on:I pu_on_n:I vccd:I 
*.PININFO vdda:I vddio_q:I vssa:I vssd:I vswitch:I nga_amx_vswitch_h:O 
*.PININFO nga_pad_vswitch_h:O nga_pad_vswitch_h_n:O ngb_amx_vswitch_h:O 
*.PININFO ngb_pad_vswitch_h:O ngb_pad_vswitch_h_n:O nmida_vccd:O 
*.PININFO nmida_vccd_n:O nmidb_vccd:O nmidb_vccd_n:O pd_csd_vswitch_h:O 
*.PININFO pd_csd_vswitch_h_n:O pga_amx_vdda_h_n:O pga_pad_vddioq_h_n:O 
*.PININFO pgb_amx_vdda_h_n:O pgb_pad_vddioq_h_n:O pu_csd_vddioq_h_n:O
XICEhld_i_h_n hld_i_h_n / icecap
XICEnmida_vccd_n nmida_vccd_n / icecap
XICEnmidb_vccd nmidb_vccd / icecap
XICEpu_on_n pu_on_n / icecap
XICEnet295 net295 / icecap
XICEpd_csd_vswitch_h pd_csd_vswitch_h / icecap
XICEnet278 net278 / icecap
XICEnet160 net160 / icecap
XICEnet154 net154 / icecap
XICEhld_i_h hld_i_h / icecap
XICEamuxbusb_on_n amuxbusb_on_n / icecap
XICEnet149 net149 / icecap
XICEpd_on pd_on / icecap
XICEnet284 net284 / icecap
XICEpga_amx_vdda_h_n pga_amx_vdda_h_n / icecap
XICEamuxbusa_on amuxbusa_on / icecap
XICEpga_pad_vddioq_h_n pga_pad_vddioq_h_n / icecap
XICEamux_en_vddio_h amux_en_vddio_h / icecap
XICEpgb_amx_vdda_h_n pgb_amx_vdda_h_n / icecap
XICEamux_en_vswitch_h_n amux_en_vswitch_h_n / icecap
XICEnet296 net296 / icecap
XICEamux_en_vdda_h amux_en_vdda_h / icecap
XICEpd_on_n pd_on_n / icecap
XICEnmidb_vccd_n nmidb_vccd_n / icecap
XICEnet167 net167 / icecap
XICEngb_amx_vswitch_h ngb_amx_vswitch_h / icecap
XICEnet293 net293 / icecap
XICEnet168 net168 / icecap
XICEnga_pad_vswitch_h nga_pad_vswitch_h / icecap
XICEnmida_on_n nmida_on_n / icecap
XICEnga_amx_vswitch_h nga_amx_vswitch_h / icecap
XICEnet287 net287 / icecap
XICEpu_csd_vddioq_h_n pu_csd_vddioq_h_n / icecap
XICEamux_en_vdda_h_n amux_en_vdda_h_n / icecap
XICEamuxbusa_on_n amuxbusa_on_n / icecap
XICEamux_en_vswitch_h amux_en_vswitch_h / icecap
XICEamuxbusb_on amuxbusb_on / icecap
XICEpu_on pu_on / icecap
XICEnet144 net144 / icecap
XICEngb_pad_vswitch_h ngb_pad_vswitch_h / icecap
XICEpgb_pad_vddioq_h_n pgb_pad_vddioq_h_n / icecap
XICEpd_csd_vswitch_h_n pd_csd_vswitch_h_n / icecap
XICEamux_en_vddio_h_n amux_en_vddio_h_n / icecap
XICEngb_pad_vswitch_h_n ngb_pad_vswitch_h_n / icecap
XICEnmida_vccd nmida_vccd / icecap
XICEnmidb_on_n nmidb_on_n / icecap
XICEnga_pad_vswitch_h_n nga_pad_vswitch_h_n / icecap
Xpga_pad_ls amuxbusa_on amuxbusa_on_n net154 net160 hld_i_h hld_i_h_n 
+ amux_en_vddio_h_n amux_en_vddio_h vssd vddio_q vccd / 
+ sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3_ver2
Xpgb_pad_ls amuxbusb_on amuxbusb_on_n net144 net149 hld_i_h hld_i_h_n 
+ amux_en_vddio_h_n amux_en_vddio_h vssd vddio_q vccd / 
+ sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3_ver2
XI38 net168 pu_csd_vddioq_h_n vddio_q vssd / sky130_fd_io__gpiov2_amx_pucsd_buf
Xpu_csd_ls pu_on pu_on_n net167 net168 hld_i_h_n amux_en_vddio_h vssd vddio_q 
+ vccd / sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3
XI111 hld_i_h_n hld_i_h vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI110 amux_en_vddio_h amux_en_vddio_h_n vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI93 nmida_vccd nmida_vccd_n vssd vccd / sky130_fd_io__hvsbt_inv_x1
XI105 nmidb_vccd nmidb_vccd_n vssd vccd / sky130_fd_io__hvsbt_inv_x1
Xpga_amx_ls net154 net160 pga_amx_vdda_h_n amux_en_vdda_h_n amux_en_vdda_h 
+ vssa vdda / sky130_fd_io__gpiov2_amux_drvr_lshv2hv
XI103 net144 net149 pgb_amx_vdda_h_n amux_en_vdda_h_n amux_en_vdda_h vssa vdda 
+ / sky130_fd_io__gpiov2_amux_drvr_lshv2hv
XI45 net295 nga_amx_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_inv4
XI42 net154 pga_pad_vddioq_h_n vddio_q vssd / sky130_fd_io__gpiov2_amx_inv4
XI47 net295 nga_pad_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_inv4
XI62 net144 pgb_pad_vddioq_h_n vddio_q vssd / sky130_fd_io__gpiov2_amx_inv4
XI63 net284 ngb_amx_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_inv4
XI64 net284 ngb_pad_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_inv4
XI53 nmidb_on_n nmidb_vccd vssd vccd / sky130_fd_io__hvsbt_inv_x2
XI89 nmida_on_n nmida_vccd vssd vccd / sky130_fd_io__hvsbt_inv_x2
Xpdcsd_inv net293 pd_csd_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_pdcsd_inv
XI87 nga_pad_vswitch_h nga_pad_vswitch_h_n vswitch vssa / sky130_fd_io__amx_inv1
XI85 ngb_pad_vswitch_h ngb_pad_vswitch_h_n vswitch vssa / sky130_fd_io__amx_inv1
XI90 pd_csd_vswitch_h pd_csd_vswitch_h_n vswitch vssa / sky130_fd_io__amx_inv1
mI76 ngb_amx_vswitch_h amux_en_vdda_h_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI77 ngb_pad_vswitch_h amux_en_vddio_h_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI75 nga_amx_vswitch_h amux_en_vdda_h_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI78 nga_pad_vswitch_h amux_en_vddio_h_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI104 pd_csd_vswitch_h amux_en_vddio_h_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
Xnga_ls amuxbusa_on amuxbusa_on_n net296 net295 amux_en_vswitch_h_n 
+ amux_en_vswitch_h vssa vswitch vccd / sky130_fd_io__gpiov2_amux_drvr_ls
Xpd_csd_ls pd_on pd_on_n net287 net293 amux_en_vswitch_h_n amux_en_vswitch_h 
+ vssa vswitch vccd / sky130_fd_io__gpiov2_amux_drvr_ls
Xngb_ls amuxbusb_on amuxbusb_on_n net278 net284 amux_en_vswitch_h_n 
+ amux_en_vswitch_h vssa vswitch vccd / sky130_fd_io__gpiov2_amux_drvr_ls
.ENDS
* .SUBCKT sky130_fd_io__nor2_1 A B Y vgnd vnb vpb vpwr
* *.PININFO A:I B:I vgnd:I vnb:I vpb:I vpwr:I Y:O
* XICEY Y / icecap
* XICEA A / icecap
* XICEB B / icecap
* mMP0 vpwr A sndPA vpb sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mMP1 sndPA B Y vpb sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mMN0 Y A vgnd vnb sky130_fd_pr__nfet_01v8 m=1 w=740e-3 l=150e-3 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mMN1 Y B vgnd vnb sky130_fd_pr__nfet_01v8 m=1 w=740e-3 l=150e-3 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__nand2_1 A B Y vgnd vnb vpb vpwr
* *.PININFO A:I B:I vgnd:I vnb:I vpb:I vpwr:I Y:O
* XICEA A / icecap
* XICEB B / icecap
* XICEY Y / icecap
* mMP0 Y A vpwr vpb sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mMP1 Y B vpwr vpb sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mMN0 Y A sndA vnb sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mMN1 sndA B vgnd vnb sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_amux_nand5 in0 in1 in2 in3 in4 out vgnd vpwr
* *.PININFO in0:I in1:I in2:I in3:I in4:I vgnd:I vpwr:I out:O
* XICEin4 in4 / icecap
* XICEin3 in3 / icecap
* XICEin1 in1 / icecap
* XICEout out / icecap
* XICEin2 in2 / icecap
* XICEin0 in0 / icecap
* XICEout_n out_n / icecap
* mI3 out in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI20 out out_n vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI21 out_n out vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI1 out in1 net51 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI18 net63 in4 net59 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI6 net59 in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI15 net55 in3 net63 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI14 net51 in2 net55 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI22 out_n out vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI23 vgnd out_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_amux_nand4 in0 in1 in2 in3 out vgnd vpwr
* *.PININFO in0:I in1:I in2:I in3:I vgnd:I vpwr:I out:O
* XICEout_n out_n / icecap
* XICEin1 in1 / icecap
* XICEout out / icecap
* XICEin3 in3 / icecap
* XICEin0 in0 / icecap
* XICEin2 in2 / icecap
* mI3 out in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI19 out_n out vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI20 out out_n vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI1 out in1 net50 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI6 net58 in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI15 net54 in3 net58 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI14 net50 in2 net54 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI18 out_n out vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI21 vgnd out_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__xor2_1 A B X vgnd vpwr
* *.PININFO A:I B:I vgnd:I vpwr:I X:O
* XICEpmid pmid / icecap
* XICEinor inor / icecap
* XICEX X / icecap
* XICEA A / icecap
* XICEB B / icecap
* mMNnor0 inor A vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=840e-3 l=150e-3 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mMNnor1 inor B vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=840e-3 l=150e-3 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mMNaoi10 vgnd A sndNA vgnd sky130_fd_pr__nfet_01v8 m=1 w=840e-3 l=150e-3 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mMNaoi11 sndNA B X vgnd sky130_fd_pr__nfet_01v8 m=1 w=840e-3 l=150e-3 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mMNaoi20 X inor vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=840e-3 l=150e-3 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mMPnor0 vpwr A sndPA vpwr sky130_fd_pr__pfet_01v8_hvt m=1 w=1.26 l=150e-3 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mMPnor1 sndPA B inor vpwr sky130_fd_pr__pfet_01v8_hvt m=1 w=1.26 l=150e-3 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mMPaoi10 pmid A vpwr vpwr sky130_fd_pr__pfet_01v8_hvt m=1 w=1.26 l=150e-3 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mMPaoi11 pmid B vpwr vpwr sky130_fd_pr__pfet_01v8_hvt m=1 w=1.26 l=150e-3 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mMPaoi20 X inor pmid vpwr sky130_fd_pr__pfet_01v8_hvt m=1 w=1.26 l=150e-3 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__inv_1 A Y vgnd vnb vpb vpwr
* *.PININFO A:I vgnd:I vnb:I vpb:I vpwr:I Y:O
* XICEA A / icecap
* XICEY Y / icecap
* mMIN1 Y A vgnd vnb sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mMIP1 Y A vpwr vpb sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_amux_decoder amuxbusa_on amuxbusa_on_n amuxbusb_on 
* + amuxbusb_on_n analog_en analog_pol analog_sel nga_pad_vswitch_h 
* + nga_pad_vswitch_h_n ngb_pad_vswitch_h ngb_pad_vswitch_h_n nmida_on_n 
* + nmida_vccd_n nmidb_on_n nmidb_vccd_n out pd_on pd_on_n pd_vswitch_h_n 
* + pga_amx_vdda_h_n pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n 
* + pu_on pu_on_n pu_vddioq_h_n vccd vssd
* *.PININFO analog_en:I analog_pol:I analog_sel:I nga_pad_vswitch_h:I 
* *.PININFO nga_pad_vswitch_h_n:I ngb_pad_vswitch_h:I ngb_pad_vswitch_h_n:I 
* *.PININFO nmida_vccd_n:I nmidb_vccd_n:I out:I pd_vswitch_h_n:I 
* *.PININFO pga_amx_vdda_h_n:I pga_pad_vddioq_h_n:I pgb_amx_vdda_h_n:I 
* *.PININFO pgb_pad_vddioq_h_n:I pu_vddioq_h_n:I vccd:I vssd:I amuxbusa_on:O 
* *.PININFO amuxbusa_on_n:O amuxbusb_on:O amuxbusb_on_n:O nmida_on_n:O 
* *.PININFO nmidb_on_n:O pd_on:O pd_on_n:O pu_on:O pu_on_n:O
* XICEint_pu_on int_pu_on / icecap
* XICEout_i_n out_i_n / icecap
* XICEpd_vswitch_h_n pd_vswitch_h_n / icecap
* XICEnmida_on_n nmida_on_n / icecap
* XICEnmida_vccd_n nmida_vccd_n / icecap
* XICEnmidb_vccd_n nmidb_vccd_n / icecap
* XICEamuxbusa_on amuxbusa_on / icecap
* XICEnet167 net167 / icecap
* XICEanalog_pol analog_pol / icecap
* XICEnga_pad_vswitch_h_n nga_pad_vswitch_h_n / icecap
* XICEint_pd_on int_pd_on / icecap
* XICEout out / icecap
* XICEana_en_i_n ana_en_i_n / icecap
* XICEpgb_pad_vddioq_h_n pgb_pad_vddioq_h_n / icecap
* XICEint_amuxb_on int_amuxb_on / icecap
* XICEint_pd_on_n int_pd_on_n / icecap
* XICEpu_on pu_on / icecap
* XICEpu_vddioq_h_n pu_vddioq_h_n / icecap
* XICEpga_amx_vdda_h_n pga_amx_vdda_h_n / icecap
* XICEnet212 net212 / icecap
* XICEngb_pad_vswitch_h_n ngb_pad_vswitch_h_n / icecap
* XICEpd_on_n pd_on_n / icecap
* XICEint_amuxa_on int_amuxa_on / icecap
* XICEint_amux_a_on_n int_amux_a_on_n / icecap
* XICEpgb_amx_vdda_h_n pgb_amx_vdda_h_n / icecap
* XICEint_amux_b_on_n int_amux_b_on_n / icecap
* XICEint_fbk_puon_n int_fbk_puon_n / icecap
* XICEnet222 net222 / icecap
* XICEnmidb_on_n nmidb_on_n / icecap
* XICEana_pol_i ana_pol_i / icecap
* XICEamuxbusb_on_n amuxbusb_on_n / icecap
* XICEint_fbk_pdon_n int_fbk_pdon_n / icecap
* XICEnet137 net137 / icecap
* XICEanalog_en analog_en / icecap
* XICEnga_pad_vswitch_h nga_pad_vswitch_h / icecap
* XICEana_sel_i ana_sel_i / icecap
* XICEnet144 net144 / icecap
* XICEpd_on pd_on / icecap
* XICEamuxbusb_on amuxbusb_on / icecap
* XICEanalog_sel analog_sel / icecap
* XICEngb_pad_vswitch_h ngb_pad_vswitch_h / icecap
* XICEpol_xor_out pol_xor_out / icecap
* XICEana_sel_i_n ana_sel_i_n / icecap
* XICEout_i out_i / icecap
* XICEpu_on_n pu_on_n / icecap
* XICEamuxbusa_on_n amuxbusa_on_n / icecap
* XICEint_pu_on_n int_pu_on_n / icecap
* XICEnet172 net172 / icecap
* XICEpga_pad_vddioq_h_n pga_pad_vddioq_h_n / icecap
* XICEana_pol_i_n ana_pol_i_n / icecap
* XI116 ana_en_i_n int_pd_on_n int_pd_on vssd vssd vccd vccd / sky130_fd_io__nor2_1
* XI113 ana_en_i_n net144 int_amuxa_on vssd vssd vccd vccd / sky130_fd_io__nor2_1
* XI115 ana_en_i_n int_pu_on_n int_pu_on vssd vssd vccd vccd / sky130_fd_io__nor2_1
* XI114 ana_en_i_n net137 int_amuxb_on vssd vssd vccd vccd / sky130_fd_io__nor2_1
* XI111 ana_pol_i out_i int_pu_on_n vssd vssd vccd vccd / sky130_fd_io__nand2_1
* XI112 ana_pol_i_n out_i_n int_pd_on_n vssd vssd vccd vccd / sky130_fd_io__nand2_1
* XI109 ana_sel_i_n pol_xor_out net144 vssd vssd vccd vccd / sky130_fd_io__nand2_1
* XI110 pol_xor_out ana_sel_i net137 vssd vssd vccd vccd / sky130_fd_io__nand2_1
* XI106 ngb_pad_vswitch_h net212 net172 vssd vccd / sky130_fd_io__hvsbt_nor
* XI102 nga_pad_vswitch_h net222 net167 vssd vccd / sky130_fd_io__hvsbt_nor
* XI79 int_pu_on pga_pad_vddioq_h_n pgb_pad_vddioq_h_n nga_pad_vswitch_h_n 
* + ngb_pad_vswitch_h_n int_fbk_puon_n vssd vccd / sky130_fd_io__gpiov2_amux_nand5
* XI80 int_pd_on pga_pad_vddioq_h_n pgb_pad_vddioq_h_n nga_pad_vswitch_h_n 
* + ngb_pad_vswitch_h_n int_fbk_pdon_n vssd vccd / sky130_fd_io__gpiov2_amux_nand5
* XI78 int_amuxb_on pu_vddioq_h_n pd_vswitch_h_n nmidb_vccd_n amuxbusb_on_n vssd 
* + vccd / sky130_fd_io__gpiov2_amux_nand4
* XI77 int_amuxa_on pu_vddioq_h_n pd_vswitch_h_n nmida_vccd_n amuxbusa_on_n vssd 
* + vccd / sky130_fd_io__gpiov2_amux_nand4
* XI101 pga_pad_vddioq_h_n pga_amx_vdda_h_n net222 vssd vccd / 
* + sky130_fd_io__hvsbt_nand2
* XI121 int_amux_b_on_n net172 nmidb_on_n vssd vccd / sky130_fd_io__hvsbt_nand2
* XI105 pgb_pad_vddioq_h_n pgb_amx_vdda_h_n net212 vssd vccd / 
* + sky130_fd_io__hvsbt_nand2
* XI120 int_amux_a_on_n net167 nmida_on_n vssd vccd / sky130_fd_io__hvsbt_nand2
* XI45 ana_pol_i out_i pol_xor_out vssd vccd / sky130_fd_io__xor2_1
* XI41 ana_pol_i_n ana_pol_i vssd vssd vccd vccd / sky130_fd_io__inv_1
* XI89 int_amuxa_on int_amux_a_on_n vssd vssd vccd vccd / sky130_fd_io__inv_1
* XI39 analog_sel ana_sel_i_n vssd vssd vccd vccd / sky130_fd_io__inv_1
* XI40 ana_sel_i_n ana_sel_i vssd vssd vccd vccd / sky130_fd_io__inv_1
* XI35 analog_pol ana_pol_i_n vssd vssd vccd vccd / sky130_fd_io__inv_1
* XI74 amuxbusb_on_n amuxbusb_on vssd vssd vccd vccd / sky130_fd_io__inv_1
* XI73 amuxbusa_on_n amuxbusa_on vssd vssd vccd vccd / sky130_fd_io__inv_1
* XI76 int_fbk_pdon_n pd_on vssd vssd vccd vccd / sky130_fd_io__inv_1
* XI58 analog_en ana_en_i_n vssd vssd vccd vccd / sky130_fd_io__inv_1
* XI75 int_fbk_puon_n pu_on vssd vssd vccd vccd / sky130_fd_io__inv_1
* XI43 out out_i_n vssd vssd vccd vccd / sky130_fd_io__inv_1
* XI44 out_i_n out_i vssd vssd vccd vccd / sky130_fd_io__inv_1
* XI91 int_amuxb_on int_amux_b_on_n vssd vssd vccd vccd / sky130_fd_io__inv_1
* XI93 pu_on pu_on_n vssd vssd vccd vccd / sky130_fd_io__inv_1
* XI95 pd_on pd_on_n vssd vssd vccd vccd / sky130_fd_io__inv_1
* .ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_ctl_logic_i2c_fix analog_en analog_pol analog_sel 
+ enable_vdda_h enable_vdda_h_n enable_vswitch_h hld_i_h_n nga_amx_vswitch_h 
+ nga_pad_vswitch_h ngb_amx_vswitch_h ngb_pad_vswitch_h nmida_vccd nmidb_vccd 
+ out pd_csd_vswitch_h pga_amx_vdda_h_n pga_pad_vddioq_h_n pgb_amx_vdda_h_n 
+ pgb_pad_vddioq_h_n pu_csd_vddioq_h_n vccd vdda vddio_q vssa vssd vswitch
*.PININFO analog_en:I analog_pol:I analog_sel:I enable_vdda_h:I 
*.PININFO enable_vswitch_h:I hld_i_h_n:I out:I vccd:I vdda:I vddio_q:I vssa:I 
*.PININFO vssd:I vswitch:I enable_vdda_h_n:O nga_amx_vswitch_h:O 
*.PININFO nga_pad_vswitch_h:O ngb_amx_vswitch_h:O ngb_pad_vswitch_h:O 
*.PININFO nmida_vccd:O nmidb_vccd:O pd_csd_vswitch_h:O pga_amx_vdda_h_n:O 
*.PININFO pga_pad_vddioq_h_n:O pgb_amx_vdda_h_n:O pgb_pad_vddioq_h_n:O 
*.PININFO pu_csd_vddioq_h_n:O
XICEnga_pad_vswitch_h nga_pad_vswitch_h / icecap
XICEngb_pad_vswitch_h ngb_pad_vswitch_h / icecap
XICEpd_csd_vswitch_h pd_csd_vswitch_h / icecap
XICEnmidb_on_n nmidb_on_n / icecap
XICEenable_vswitch_h enable_vswitch_h / icecap
XICEamuxbusb_on_n amuxbusb_on_n / icecap
XICEpu_on pu_on / icecap
XICEpu_csd_vddioq_h_n pu_csd_vddioq_h_n / icecap
XICEnmida_vccd_n nmida_vccd_n / icecap
XICEnga_pad_vswitch_h_n nga_pad_vswitch_h_n / icecap
XICEpd_on pd_on / icecap
XICEamux_en_vswitch_h_n amux_en_vswitch_h_n / icecap
XICEhld_i_h_n hld_i_h_n / icecap
XICEenable_vdda_h_n enable_vdda_h_n / icecap
XICEout out / icecap
XICEpu_on_n pu_on_n / icecap
XICEanalog_en analog_en / icecap
XICEpgb_amx_vdda_h_n pgb_amx_vdda_h_n / icecap
XICEamux_en_vdda_h amux_en_vdda_h / icecap
XICEngb_pad_vswitch_h_n ngb_pad_vswitch_h_n / icecap
XICEpd_on_n pd_on_n / icecap
XICEamux_en_vswitch_h amux_en_vswitch_h / icecap
XICEamux_en_vdda_h_n amux_en_vdda_h_n / icecap
XICEpgb_pad_vddioq_h_n pgb_pad_vddioq_h_n / icecap
XICEnga_amx_vswitch_h nga_amx_vswitch_h / icecap
XICEenable_vdda_h enable_vdda_h / icecap
XICEpd_csd_vswitch_h_n pd_csd_vswitch_h_n / icecap
XICEnmida_vccd nmida_vccd / icecap
XICEamuxbusa_on_n amuxbusa_on_n / icecap
XICEnmidb_vccd nmidb_vccd / icecap
XICEanalog_pol analog_pol / icecap
XICEpga_amx_vdda_h_n pga_amx_vdda_h_n / icecap
XICEamux_en_vddio_h amux_en_vddio_h / icecap
XICEngb_amx_vswitch_h ngb_amx_vswitch_h / icecap
XICEamuxbusa_on amuxbusa_on / icecap
XICEamuxbusb_on amuxbusb_on / icecap
XICEpga_pad_vddioq_h_n pga_pad_vddioq_h_n / icecap
XICEnmida_on_n nmida_on_n / icecap
XICEanalog_sel analog_sel / icecap
XICEnmidb_vccd_n nmidb_vccd_n / icecap
Xamux_ls amux_en_vdda_h amux_en_vdda_h_n amux_en_vddio_h amux_en_vswitch_h 
+ amux_en_vswitch_h_n analog_en enable_vdda_h enable_vdda_h_n enable_vswitch_h 
+ hld_i_h_n vccd vdda vddio_q vssa vssd vswitch / 
+ sky130_fd_io__gpiov2_amux_ls_i2c_fix
Xamux_sw_drvr amux_en_vdda_h amux_en_vdda_h_n amux_en_vddio_h 
+ amux_en_vswitch_h amux_en_vswitch_h_n amuxbusa_on amuxbusa_on_n amuxbusb_on 
+ amuxbusb_on_n hld_i_h_n nga_amx_vswitch_h nga_pad_vswitch_h 
+ nga_pad_vswitch_h_n ngb_amx_vswitch_h ngb_pad_vswitch_h ngb_pad_vswitch_h_n 
+ nmida_on_n nmida_vccd nmida_vccd_n nmidb_on_n nmidb_vccd nmidb_vccd_n 
+ pd_csd_vswitch_h pd_csd_vswitch_h_n pd_on pd_on_n pga_amx_vdda_h_n 
+ pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n pu_csd_vddioq_h_n 
+ pu_on pu_on_n vccd vdda vddio_q vssa vssd vswitch / 
+ sky130_fd_io__gpiov2_amux_drvr_i2c_fix
Xamux_lv_decoder amuxbusa_on amuxbusa_on_n amuxbusb_on amuxbusb_on_n analog_en 
+ analog_pol analog_sel nga_pad_vswitch_h nga_pad_vswitch_h_n 
+ ngb_pad_vswitch_h ngb_pad_vswitch_h_n nmida_on_n nmida_vccd_n nmidb_on_n 
+ nmidb_vccd_n out pd_on pd_on_n pd_csd_vswitch_h_n pga_amx_vdda_h_n 
+ pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n pu_on pu_on_n 
+ pu_csd_vddioq_h_n vccd vssd / sky130_fd_io__gpiov2_amux_decoder
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_amux_switch ag_hv ng_ag_vpmp ng_pad_vpmp nghs_h 
+ nmid_vdda pad_hv_n0 pad_hv_n1 pad_hv_n2 pad_hv_n3 pad_hv_p0 pad_hv_p1 
+ pd_h_vdda pd_h_vddio pg_ag_vdda pg_pad_vddioq pghs_h pug_h vdda vddio 
+ vpb_drvr vssa vssd vssio
*.PININFO ng_ag_vpmp:I ng_pad_vpmp:I nghs_h:I nmid_vdda:I pd_h_vdda:I 
*.PININFO pd_h_vddio:I pg_ag_vdda:I pg_pad_vddioq:I pghs_h:I vdda:I vddio:I 
*.PININFO vssa:I vssd:I vssio:I ag_hv:B pad_hv_n0:B pad_hv_n1:B pad_hv_n2:B 
*.PININFO pad_hv_n3:B pad_hv_p0:B pad_hv_p1:B pug_h:B vpb_drvr:B
XICEnmid_vdda nmid_vdda / icecap
XICEpad_hv_n1 pad_hv_n1 / icecap
XICEpug_h pug_h / icecap
XICEnet85 net85 / icecap
XICEpad_hv_n3 pad_hv_n3 / icecap
XI78<0> mid / icecap
XI78<1> mid1 / icecap
XICEpg_pad_vddioq pg_pad_vddioq / icecap
XICEpd_h_vddio pd_h_vddio / icecap
XICEnghs_h nghs_h / icecap
XICEpg_ag_vdda pg_ag_vdda / icecap
XICEag_hv ag_hv / icecap
XICEvddio vddio / icecap
XICEpad_hv_p1 pad_hv_p1 / icecap
XICEpad_hv_n2 pad_hv_n2 / icecap
XICEmid1 mid1 / icecap
XICEmid mid / icecap
XICEnet83 net83 / icecap
XICEpad_hv_n0 pad_hv_n0 / icecap
XICEpghs_h pghs_h / icecap
XICEpd_h_vdda pd_h_vdda / icecap
XICEng_ag_vpmp ng_ag_vpmp / icecap
XICEng_pad_vpmp ng_pad_vpmp / icecap
XICEpad_hv_p0 pad_hv_p0 / icecap
xI72 vssa vddio condiode
xI71 mid1 vddio condiode
xI70 mid vddio condiode
XI56 vssa net85 / s8_esd_res75only_small
XI12 vssa net83 / s8_esd_res75only_small
mI46 pad_hv_n3 ng_pad_vpmp mid1 mid1 sky130_fd_pr__nfet_g5v0d10v5 m=2 w=10.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI35 mid ng_pad_vpmp pad_hv_n1 mid sky130_fd_pr__nfet_g5v0d10v5 m=2 w=10.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI24 pad_hv_n0 ng_pad_vpmp mid mid sky130_fd_pr__nfet_g5v0d10v5 m=3 w=10.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI45 mid1 ng_pad_vpmp pad_hv_n2 mid1 sky130_fd_pr__nfet_g5v0d10v5 m=3 w=10.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI28 mid ng_ag_vpmp ag_hv mid sky130_fd_pr__nfet_g5v0d10v5 m=5 w=10.0 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI57 mid1 nmid_vdda net85 vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI63 pug_h nghs_h pg_pad_vddioq vssio sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI47 mid1 ng_ag_vpmp ag_hv mid1 sky130_fd_pr__nfet_g5v0d10v5 m=5 w=10.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI75<1> mid pd_h_vdda vssa net050<0> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI75<0> mid1 pd_h_vdda vssa net050<1> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI74<1> mid pd_h_vddio vssa net051<0> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI74<0> mid1 pd_h_vddio vssa net051<1> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI1 mid nmid_vdda net83 vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI22 mid pug_h pad_hv_p1 vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=10.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI36 mid pug_h pad_hv_p0 vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=10.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI62 pg_pad_vddioq pghs_h pug_h vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI26 mid pg_ag_vdda ag_hv vdda sky130_fd_pr__pfet_g5v0d10v5 m=4 w=10.0 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_amux_i2c_fix amuxbus_a amuxbus_b analog_en 
+ analog_pol analog_sel enable_vdda_h enable_vswitch_h hld_i_h_n 
+ nga_pad_vpmp_h ngb_pad_vpmp_h nghs_h out pad pd_csd_h pghs_h pu_csd_h 
+ pug_h<1> pug_h<0> vccd vdda vddio vddio_q vpb_drvr vssa vssd vssio vswitch
*.PININFO analog_en:I analog_pol:I analog_sel:I enable_vdda_h:I 
*.PININFO enable_vswitch_h:I hld_i_h_n:I nghs_h:I out:I pghs_h:I vccd:I vdda:I 
*.PININFO vddio:I vddio_q:I vssa:I vssd:I vssio:I vswitch:I nga_pad_vpmp_h:O 
*.PININFO ngb_pad_vpmp_h:O pd_csd_h:O pu_csd_h:O amuxbus_a:B amuxbus_b:B pad:B 
*.PININFO pug_h<1>:B pug_h<0>:B vpb_drvr:B
XICEpghs_h pghs_h / icecap
XICEnga_pad_vpmp_h nga_pad_vpmp_h / icecap
XICEngb_amx_vpmp_h ngb_amx_vpmp_h / icecap
XICEanalog_pol analog_pol / icecap
XICEvssio vssio / icecap
XICEenable_vdda_h_n enable_vdda_h_n / icecap
XICEpad pad / icecap
XICEnet128 net128 / icecap
XICEenable_vdda_h enable_vdda_h / icecap
XICEnet126 net126 / icecap
XICEpgb_pad_vddioq_h_n pgb_pad_vddioq_h_n / icecap
XICEpug_h<1> pug_h<1> / icecap
XICEamuxbus_a amuxbus_a / icecap
XICEpu_csd_h pu_csd_h / icecap
XICEhld_i_h_n hld_i_h_n / icecap
XICEpga_pad_vddioq_h_n pga_pad_vddioq_h_n / icecap
XICEpgb_amx_vdda_h_n pgb_amx_vdda_h_n / icecap
XICEhld_i_h_amux_sw hld_i_h_amux_sw / icecap
XICEpga_amx_vdda_h_n pga_amx_vdda_h_n / icecap
XICEnet120 net120 / icecap
XICEout out / icecap
XICEnmidb_vccd nmidb_vccd / icecap
XICEnga_amx_vpmp_h nga_amx_vpmp_h / icecap
XICEenable_vswitch_h enable_vswitch_h / icecap
XICEnet142 net142 / icecap
XICEnghs_h nghs_h / icecap
XICEnet139 net139 / icecap
XICEnet124 net124 / icecap
XICEpug_h<0> pug_h<0> / icecap
XICEngb_pad_vpmp_h ngb_pad_vpmp_h / icecap
XICEamuxbus_b amuxbus_b / icecap
XICEnet143 net143 / icecap
XICEanalog_sel analog_sel / icecap
XICEnmida_vccd nmida_vccd / icecap
XICEpd_csd_h pd_csd_h / icecap
XICEnet144 net144 / icecap
XICEanalog_en analog_en / icecap
XI78 hld_i_h_n hld_i_h_amux_sw vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XBBM_logic analog_en analog_pol analog_sel enable_vdda_h enable_vdda_h_n 
+ enable_vswitch_h hld_i_h_n nga_amx_vpmp_h nga_pad_vpmp_h ngb_amx_vpmp_h 
+ ngb_pad_vpmp_h nmida_vccd nmidb_vccd out pd_csd_h pga_amx_vdda_h_n 
+ pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n pu_csd_h vccd vdda 
+ vddio_q vssa vssd vswitch / sky130_fd_io__gpiov2_amux_ctl_logic_i2c_fix
xI77 vssa vdda condiode
XI26 net128 net142 / s8_esd_res75only_small
XI58 net126 net139 / s8_esd_res75only_small
XI28 net124 net144 / s8_esd_res75only_small
XI57 pad net126 / s8_esd_res75only_small
XI27 net120 net143 / s8_esd_res75only_small
XI55 pad net128 / s8_esd_res75only_small
XI54 pad net124 / s8_esd_res75only_small
XI53 pad net120 / s8_esd_res75only_small
Xmux_a amuxbus_a nga_amx_vpmp_h nga_pad_vpmp_h nghs_h nmida_vccd net144 net144 
+ net139 net139 net143 net142 enable_vdda_h_n hld_i_h_amux_sw pga_amx_vdda_h_n 
+ pga_pad_vddioq_h_n pghs_h pug_h<0> vdda vddio vpb_drvr vssa vssd vssio / 
+ sky130_fd_io__gpio_ovtv2_amux_switch
Xmux_b amuxbus_b ngb_amx_vpmp_h ngb_pad_vpmp_h nghs_h nmidb_vccd net144 net144 
+ net139 net139 net143 net142 enable_vdda_h_n hld_i_h_amux_sw pgb_amx_vdda_h_n 
+ pgb_pad_vddioq_h_n pghs_h pug_h<1> vdda vddio vpb_drvr vssa vssd vssio / 
+ sky130_fd_io__gpio_ovtv2_amux_switch
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_ctl_lsbank_i2c_fix dm<2> dm<1> dm<0> dm_h<2> 
+ dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n hyst_trim 
+ hyst_trim_h hyst_trim_h_n ib_mode_sel<1> ib_mode_sel<0> ib_mode_sel_h<1> 
+ ib_mode_sel_h<0> ib_mode_sel_h_n<1> ib_mode_sel_h_n<0> inp_dis inp_dis_h 
+ inp_dis_h_n od_i_h_n slew_ctl<1> slew_ctl<0> slew_ctl_h<1> slew_ctl_h<0> 
+ slew_ctl_h_n<1> slew_ctl_h_n<0> startup_rst_h startup_st_h vcc_io vgnd vpwr 
+ vtrip_sel vtrip_sel_h vtrip_sel_h_n
*.PININFO dm<2>:I dm<1>:I dm<0>:I hld_i_h_n:I hyst_trim:I ib_mode_sel<1>:I 
*.PININFO ib_mode_sel<0>:I inp_dis:I od_i_h_n:I slew_ctl<1>:I slew_ctl<0>:I 
*.PININFO startup_rst_h:I startup_st_h:I vcc_io:I vgnd:I vpwr:I vtrip_sel:I 
*.PININFO dm_h<2>:O dm_h<1>:O dm_h<0>:O dm_h_n<2>:O dm_h_n<1>:O dm_h_n<0>:O 
*.PININFO hyst_trim_h:O hyst_trim_h_n:O ib_mode_sel_h<1>:O ib_mode_sel_h<0>:O 
*.PININFO ib_mode_sel_h_n<1>:O ib_mode_sel_h_n<0>:O inp_dis_h:O inp_dis_h_n:O 
*.PININFO slew_ctl_h<1>:O slew_ctl_h<0>:O slew_ctl_h_n<1>:O slew_ctl_h_n<0>:O 
*.PININFO vtrip_sel_h:O vtrip_sel_h_n:O
XICEdm_h_n<0> dm_h_n<0> / icecap
XI851<0> ib_mode_sel<1> / icecap
XI851<1> ib_mode_sel<0> / icecap
XI837<0> ib_mode_sel_rst_h<1> / icecap
XI837<1> ib_mode_sel_rst_h<0> / icecap
XI843<0> dm_h<2> / icecap
XI843<1> dm_h<1> / icecap
XICEod_i_h od_i_h / icecap
XICEvtrip_sel_h_n vtrip_sel_h_n / icecap
XICEdm_h<0> dm_h<0> / icecap
XICEie_n_st_h ie_n_st_h / icecap
XICEhyst_trim_st_h hyst_trim_st_h / icecap
XICEvtrip_sel vtrip_sel / icecap
XICEinp_dis_h_n inp_dis_h_n / icecap
XICEinp_dis inp_dis / icecap
XICEdm<0> dm<0> / icecap
XICEdm_rst_h<2> dm_rst_h<2> / icecap
XI844<0> slew_ctl<1> / icecap
XI844<1> slew_ctl<0> / icecap
XI846<0> slew_ctl_h<1> / icecap
XI846<1> slew_ctl_h<0> / icecap
XICEhyst_trim_h_n hyst_trim_h_n / icecap
XICEdm_st_h<2> dm_st_h<2> / icecap
XICEhyst_trim_rst_h hyst_trim_rst_h / icecap
XICEdm_rst_h<0> dm_rst_h<0> / icecap
XI845<0> slew_ctl_rst_h<1> / icecap
XI845<1> slew_ctl_rst_h<0> / icecap
XI839<0> dm<2> / icecap
XI839<1> dm<1> / icecap
XICEie_n_rst_h ie_n_rst_h / icecap
XI840<0> dm_h_n<2> / icecap
XI840<1> dm_h_n<1> / icecap
XICEod_i_h_n od_i_h_n / icecap
XICEdm_st_h<0> dm_st_h<0> / icecap
XICEhyst_trim_h hyst_trim_h / icecap
XI838<0> dm_st_h<2> / icecap
XI838<1> dm_st_h<1> / icecap
XICEinp_dis_h inp_dis_h / icecap
XICEdm_rst_h<1> dm_rst_h<1> / icecap
XICEvtrip_sel_h vtrip_sel_h / icecap
XICEstartup_rst_h startup_rst_h / icecap
XICEstartup_st_h startup_st_h / icecap
XICEhyst_trim hyst_trim / icecap
XI841<0> ib_mode_sel_h<1> / icecap
XI841<1> ib_mode_sel_h<0> / icecap
XI848<0> ib_mode_sel_st_h<1> / icecap
XI848<1> ib_mode_sel_st_h<0> / icecap
XICEdm_st_h<1> dm_st_h<1> / icecap
XI847<0> slew_ctl_st_h<1> / icecap
XI847<1> slew_ctl_st_h<0> / icecap
XICEtrip_sel_st_h trip_sel_st_h / icecap
XICEtrip_sel_rst_h trip_sel_rst_h / icecap
XICEhld_i_h_n hld_i_h_n / icecap
XI850<0> slew_ctl_h_n<1> / icecap
XI850<1> slew_ctl_h_n<0> / icecap
XI849<0> ib_mode_sel_h_n<1> / icecap
XI849<1> ib_mode_sel_h_n<0> / icecap
XI842<0> dm_rst_h<2> / icecap
XI842<1> dm_rst_h<1> / icecap
XI836 od_i_h_n od_i_h vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
Xtrip_sel_st trip_sel_st_h od_i_h vgnd / sky130_fd_io__tk_opti
XI803<1> dm_st_h<1> od_i_h vgnd / sky130_fd_io__tk_opti
Xtrip_sel_rst trip_sel_rst_h vgnd od_i_h / sky130_fd_io__tk_opti
XI802<1> dm_st_h<2> od_i_h vgnd / sky130_fd_io__tk_opti
XI804<1> dm_rst_h<2> vgnd od_i_h / sky130_fd_io__tk_opti
XI338<1> dm_rst_h<0> startup_st_h startup_rst_h / sky130_fd_io__tk_opti
XI615 hyst_trim_st_h od_i_h vgnd / sky130_fd_io__tk_opti
XI614 hyst_trim_rst_h vgnd od_i_h / sky130_fd_io__tk_opti
XI598<1> ib_mode_sel_st_h<1> od_i_h vgnd / sky130_fd_io__tk_opti
XI598<0> ib_mode_sel_st_h<0> od_i_h vgnd / sky130_fd_io__tk_opti
XI597<1> ib_mode_sel_rst_h<1> vgnd od_i_h / sky130_fd_io__tk_opti
XI597<0> ib_mode_sel_rst_h<0> vgnd od_i_h / sky130_fd_io__tk_opti
XI337<1> dm_st_h<0> startup_rst_h startup_st_h / sky130_fd_io__tk_opti
XI805<1> dm_rst_h<1> vgnd od_i_h / sky130_fd_io__tk_opti
XI666<1> slew_ctl_st_h<1> od_i_h vgnd / sky130_fd_io__tk_opti
XI666<0> slew_ctl_st_h<0> od_i_h vgnd / sky130_fd_io__tk_opti
XI665<1> slew_ctl_rst_h<1> vgnd od_i_h / sky130_fd_io__tk_opti
XI665<0> slew_ctl_rst_h<0> vgnd od_i_h / sky130_fd_io__tk_opti
XI687 ie_n_st_h startup_st_h startup_rst_h / sky130_fd_io__tk_opti
XI686 ie_n_rst_h startup_rst_h startup_st_h / sky130_fd_io__tk_opti
Xdm_ls_0 hld_i_h_n dm<0> dm_h<0> dm_h_n<0> dm_rst_h<0> dm_st_h<0> vcc_io vgnd 
+ vpwr / sky130_fd_io__com_ctl_ls
Xinp_dis_ls hld_i_h_n inp_dis inp_dis_h inp_dis_h_n ie_n_rst_h ie_n_st_h 
+ vcc_io vgnd vpwr / sky130_fd_io__com_ctl_ls
Xtrip_sel_ls hld_i_h_n vtrip_sel vtrip_sel_h vtrip_sel_h_n trip_sel_rst_h 
+ trip_sel_st_h vcc_io vgnd vpwr / sky130_fd_io__com_ctl_ls
XI616 hld_i_h_n hyst_trim hyst_trim_h hyst_trim_h_n hyst_trim_rst_h 
+ hyst_trim_st_h vcc_io vgnd vpwr / sky130_fd_io__com_ctl_ls
XI595<1> hld_i_h_n ib_mode_sel<1> ib_mode_sel_h<1> ib_mode_sel_h_n<1> 
+ ib_mode_sel_rst_h<1> ib_mode_sel_st_h<1> net58<0> net56<0> net57<0> / 
+ sky130_fd_io__com_ctl_ls
XI595<0> hld_i_h_n ib_mode_sel<0> ib_mode_sel_h<0> ib_mode_sel_h_n<0> 
+ ib_mode_sel_rst_h<0> ib_mode_sel_st_h<0> net58<1> net56<1> net57<1> / 
+ sky130_fd_io__com_ctl_ls
XI667<1> hld_i_h_n slew_ctl<1> slew_ctl_h<1> slew_ctl_h_n<1> slew_ctl_rst_h<1> 
+ slew_ctl_st_h<1> net61<0> net59<0> net60<0> / sky130_fd_io__com_ctl_ls
XI667<0> hld_i_h_n slew_ctl<0> slew_ctl_h<0> slew_ctl_h_n<0> slew_ctl_rst_h<0> 
+ slew_ctl_st_h<0> net61<1> net59<1> net60<1> / sky130_fd_io__com_ctl_ls
Xdm_ls<2> hld_i_h_n dm<2> dm_h<2> dm_h_n<2> dm_rst_h<2> dm_st_h<2> vcc_io vgnd 
+ vpwr / sky130_fd_io__com_ctl_ls
Xdm_ls<1> hld_i_h_n dm<1> dm_h<1> dm_h_n<1> dm_rst_h<1> dm_st_h<1> vcc_io vgnd 
+ vpwr / sky130_fd_io__com_ctl_ls
.ENDS
.SUBCKT sky130_fd_io__enh_nand2_1_sp in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
XICEout out / icecap
XICEin1 in1 / icecap
XICEin0 in0 / icecap
mI3 out in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI5 out in1 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI1 out in1 net25 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI6 net25 in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__enh_nor2_x1 in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
XICEout out / icecap
XICEnet16 net16 / icecap
XICEin0 in0 / icecap
XICEin1 in1 / icecap
mI3 net16 in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI12 out in1 net16 vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI1 out in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI6 out in1 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__enh_nand2_1 in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
XICEout out / icecap
XICEin0 in0 / icecap
XICEin1 in1 / icecap
mI3 out in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI5 out in1 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI1 out in1 net25 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI6 net25 in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__nor2_4_enhpath in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
XICEout out / icecap
XICEnet16 net16 / icecap
XICEin0 in0 / icecap
XICEin1 in1 / icecap
mI3 net16 in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=16 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI12 out in1 net16 vpwr sky130_fd_pr__pfet_g5v0d10v5 m=16 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI1 out in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=8 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI6 out in1 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=8 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__nand2_2_enhpath in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
XICEout out / icecap
XICEin1 in1 / icecap
XICEin0 in0 / icecap
mI3 out in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI5 out in1 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI1 out in1 net25 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI6 net25 in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_ctl_hld_i2c_fix enable_h hld_h_n hld_i_h_n 
+ hld_i_ovr_h hld_ovr od_i_h_n vcc_io vgnd vpwr
*.PININFO enable_h:I hld_h_n:I hld_ovr:I vcc_io:I vgnd:I vpwr:I hld_i_h_n:O 
*.PININFO hld_i_ovr_h:O od_i_h_n:O
Xhld_nand enable_h hld_h_n n1 vgnd vcc_io / sky130_fd_io__enh_nand2_1_sp
XI50 od_i_h_n net45 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI46 n1 n1 n2 vgnd vcc_io / sky130_fd_io__enh_nor2_x1
XI49 od_h od_h od_i_h_n vgnd vcc_io / sky130_fd_io__enh_nor2_x1
XI48 enable_h enable_h od_h vgnd vcc_io / sky130_fd_io__enh_nand2_1
XI155 n3 n3 hld_i_h_n vgnd vcc_io / sky130_fd_io__nor2_4_enhpath
XI154 n2 n2 n3 vgnd vcc_io / sky130_fd_io__nand2_2_enhpath
Xhld_ovr_ls n2 hld_ovr hld_ovr_h net79 od_h vgnd vcc_io vgnd vpwr / 
+ sky130_fd_io__com_ctl_ls
XI30 net45 hld_i_ovr_h_n hld_i_ovr_h vgnd vcc_io / sky130_fd_io__hvsbt_nor
XI26 n2 hld_ovr_h hld_i_ovr_h_n vgnd vcc_io / sky130_fd_io__hvsbt_nor
.ENDS
.SUBCKT sky130_fd_io__gpio_ctlv2_i2c_fix dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> 
+ dm_h_n<2> dm_h_n<1> dm_h_n<0> enable_h enable_inp_h hld_h_n hld_i_h_n 
+ hld_i_ovr_h hld_ovr hyst_trim hyst_trim_h hyst_trim_h_n ib_mode_sel<1> 
+ ib_mode_sel<0> ib_mode_sel_h<1> ib_mode_sel_h<0> ib_mode_sel_h_n<1> 
+ ib_mode_sel_h_n<0> inp_dis inp_dis_h_n od_i_h_n slew_ctl<1> slew_ctl<0> 
+ slew_ctl_h<1> slew_ctl_h<0> slew_ctl_h_n<1> slew_ctl_h_n<0> vccd vddio_q 
+ vssd vtrip_sel vtrip_sel_h
*.PININFO dm<2>:I dm<1>:I dm<0>:I enable_h:I enable_inp_h:I hld_h_n:I 
*.PININFO hld_ovr:I hyst_trim:I ib_mode_sel<1>:I ib_mode_sel<0>:I inp_dis:I 
*.PININFO slew_ctl<1>:I slew_ctl<0>:I vccd:I vddio_q:I vssd:I vtrip_sel:I 
*.PININFO dm_h<2>:O dm_h<1>:O dm_h<0>:O dm_h_n<2>:O dm_h_n<1>:O dm_h_n<0>:O 
*.PININFO hld_i_h_n:O hld_i_ovr_h:O hyst_trim_h:O hyst_trim_h_n:O 
*.PININFO ib_mode_sel_h<1>:O ib_mode_sel_h<0>:O ib_mode_sel_h_n<1>:O 
*.PININFO ib_mode_sel_h_n<0>:O inp_dis_h_n:O od_i_h_n:O slew_ctl_h<1>:O 
*.PININFO slew_ctl_h<0>:O slew_ctl_h_n<1>:O slew_ctl_h_n<0>:O vtrip_sel_h:O
Xls_bank dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
+ dm_h_n<0> hld_i_h_n hyst_trim hyst_trim_h hyst_trim_h_n ib_mode_sel<1> 
+ ib_mode_sel<0> ib_mode_sel_h<1> ib_mode_sel_h<0> ib_mode_sel_h_n<1> 
+ ib_mode_sel_h_n<0> inp_dis net83 inp_dis_h_n od_i_h_n slew_ctl<1> 
+ slew_ctl<0> slew_ctl_h<1> slew_ctl_h<0> slew_ctl_h_n<1> slew_ctl_h_n<0> 
+ startup_rst_h inp_startup_en_h vddio_q vssd vccd vtrip_sel vtrip_sel_h net77 
+ / sky130_fd_io__gpio_ovtv2_ctl_lsbank_i2c_fix
Xhld_dis_blk enable_h hld_h_n hld_i_h_n hld_i_ovr_h hld_ovr od_i_h_n vddio_q 
+ vssd vccd / sky130_fd_io__gpio_ovtv2_ctl_hld_i2c_fix
XI75 enable_inp_h enable_h startup_rst_h vssd vddio_q / sky130_fd_io__hvsbt_nor
XI56 net109 enable_inp_h net108 vssd vddio_q / sky130_fd_io__hvsbt_nand2
XI77 od_i_h_n net109 vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI57 net108 inp_startup_en_h vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_ipath_lvls enable_vddio_lv in out out_b vcchib vssd
*.PININFO enable_vddio_lv:I in:I vcchib:I vssd:I out:O out_b:O
XICEin in / icecap
XICEenable_vddio_lv enable_vddio_lv / icecap
XICEout out / icecap
XICEfbk fbk / icecap
XICEout_b out_b / icecap
XICEfbk_n fbk_n / icecap
mI248 fbk_n in vcchib vcchib sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI271 out out_b vcchib vcchib sky130_fd_pr__pfet_01v8_hvt m=2 w=5.00 l=0.25 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI281 fbk_n enable_vddio_lv vcchib vcchib sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI272 out_b fbk vcchib vcchib sky130_fd_pr__pfet_01v8_hvt m=1 w=5.00 l=0.25 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI277 fbk fbk_n vcchib vcchib sky130_fd_pr__pfet_01v8_hvt m=1 w=5.00 l=0.25 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI273 out out_b vssd vssd sky130_fd_pr__nfet_01v8 m=2 w=3.00 l=0.25 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI278 fbk fbk_n vssd vssd sky130_fd_pr__nfet_01v8 m=1 w=3.00 l=0.25 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI305 out_b fbk vssd vssd sky130_fd_pr__nfet_01v8 m=1 w=3.00 l=0.25 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI535 fbk_n in vssd_1 vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI279 vssd_1 enable_vddio_lv vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_ipath_hvls en_h_n in inb out out_b vddio_q vssd
*.PININFO en_h_n:I in:I inb:I vddio_q:I vssd:I out:O out_b:O
XICEfbk_b fbk_b / icecap
XICEout out / icecap
XICEinb inb / icecap
XICEout_b out_b / icecap
XICEen_h_n en_h_n / icecap
XICEfbk fbk / icecap
XICEin in / icecap
mI250 fbk fbk_b vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI253 out out_b vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=5 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI249 fbk_b fbk vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI248 out_b fbk vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI247 out_b fbk vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI252 out out_b vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI304 fbk inb vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI262 fbk en_h_n vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI246 fbk_b in vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_in_buf en_h en_h_n enable_vddio_lv in_h in_vt 
+ mode_normal_n mode_ref_3v_n mode_ref_n mode_vccd_n out out_n vcchib vddio_q 
+ vrefin vssd vtrip_sel_h vtrip_sel_h_n
*.PININFO en_h:I en_h_n:I enable_vddio_lv:I in_h:I in_vt:I mode_normal_n:I 
*.PININFO mode_ref_3v_n:I mode_ref_n:I mode_vccd_n:I vcchib:I vddio_q:I 
*.PININFO vrefin:I vssd:I vtrip_sel_h:I vtrip_sel_h_n:I out:O out_n:O
XICEmode_ref_3v_n mode_ref_3v_n / icecap
XICEvirt_pwr virt_pwr / icecap
XICEvddio_ref vddio_ref / icecap
XICEvcchib_int1 vcchib_int1 / icecap
XICEvddio_ref1 vddio_ref1 / icecap
XICEenable_vddio_lv enable_vddio_lv / icecap
XICEvtrip_sel_h vtrip_sel_h / icecap
XICEfbk fbk / icecap
XICEin_h in_h / icecap
XICEen_h en_h / icecap
XICEen_h_n en_h_n / icecap
XICEout out / icecap
XICEmode_vccd_n mode_vccd_n / icecap
XICEvrefin vrefin / icecap
XICEvtrip_sel_h_n vtrip_sel_h_n / icecap
XICEvcchib_int vcchib_int / icecap
XICEmode_ref_n mode_ref_n / icecap
XICEvirt_pwr2 virt_pwr2 / icecap
XICEin_b in_b / icecap
XICEmode_normal_cmos_h mode_normal_cmos_h / icecap
XICEout_n out_n / icecap
XICEenable_vddio_lv_n enable_vddio_lv_n / icecap
XICEmode_normal_cmos_h_n mode_normal_cmos_h_n / icecap
XICEmode_normal_n mode_normal_n / icecap
XICEvirt_pwr1 virt_pwr1 / icecap
XICEin_vt in_vt / icecap
XICEfbk1 fbk1 / icecap
XICEfbk2 fbk2 / icecap
XI35 enable_vddio_lv en_h enable_vddio_lv_n vssd vcchib / sky130_fd_io__hvsbt_nand2
xI405 virt_pwr1 vddio_q condiode
xI404 virt_pwr vddio_q condiode
XI488 vtrip_sel_h mode_normal_n mode_normal_cmos_h vssd vddio_q / 
+ sky130_fd_io__hvsbt_nor
XI43 mode_normal_cmos_h mode_normal_cmos_h_n vssd vddio_q / 
+ sky130_fd_io__hvsbt_inv_x1
mI630 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.00 l=0.80 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI105 fbk1 in_b fbk vssd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.80 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI620 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.00 l=0.80 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI441 in_vt vtrip_sel_h_n vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI417 out en_h_n vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI419 out_n en_h_n vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI394 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.00 l=0.80 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI494 fbk in_h vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=6 w=5.00 l=0.80 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI12 fbk2 in_b fbk vssd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.00 l=0.80 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI26 out in_b vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI49 vddio_ref vrefin virt_pwr virt_pwr sky130_fd_pr__nfet_05v0_nvt m=3 w=10.0 l=0.90 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI451 fbk in_vt vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=12 w=5.00 l=0.80 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI453 in_b in_h fbk vssd sky130_fd_pr__nfet_g5v0d10v5 m=6 w=5.00 l=0.80 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI111 vddio_ref1 vrefin virt_pwr1 virt_pwr1 sky130_fd_pr__nfet_05v0_nvt m=3 w=10.0 l=0.90 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI446 out_n out vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI389 virt_pwr vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.80 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI450 in_b in_vt fbk vssd sky130_fd_pr__nfet_g5v0d10v5 m=6 w=5.00 l=0.80 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI274 fbk1 mode_ref_n virt_pwr1 virt_pwr1 sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI116 virt_pwr mode_normal_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI109 in_b in_h virt_pwr virt_pwr sky130_fd_pr__pfet_g5v0d10v5 m=3 w=5.00 l=0.80 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI25 out in_b virt_pwr1 virt_pwr1 sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI13 fbk2 mode_normal_cmos_h_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI611 fbk1 mode_normal_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI396 vddio_ref1 mode_ref_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI115 virt_pwr mode_vccd_n vcchib_int virt_pwr sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI478 vcchib_int1 enable_vddio_lv_n vcchib vcchib sky130_fd_pr__pfet_01v8 m=8 w=5.00 l=0.25 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI373 vddio_ref mode_ref_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI403 out in_b virt_pwr2 virt_pwr2 sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI376 fbk2 mode_ref_3v_n virt_pwr1 virt_pwr1 sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI477 vcchib_int enable_vddio_lv_n vcchib vcchib sky130_fd_pr__pfet_01v8 m=8 w=5.00 l=0.25 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI401 in_b in_h virt_pwr2 virt_pwr2 sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.80 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI457 out_n out virt_pwr1 virt_pwr1 sky130_fd_pr__pfet_g5v0d10v5 m=5 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI486 fbk1 mode_vccd_n vcchib_int virt_pwr1 sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI400 virt_pwr2 mode_vccd_n vcchib_int virt_pwr2 sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI381 virt_pwr1 mode_vccd_n vcchib_int1 virt_pwr1 sky130_fd_pr__pfet_g5v0d10v5 m=6 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI380 virt_pwr1 mode_normal_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_ibuf_se en_h en_h_n enable_vddio_lv ibufmux_out 
+ ibufmux_out_h in_h in_vt mode_normal_n mode_ref_3v_n mode_ref_n mode_vccd_n 
+ vcchib vddio_q vrefin vssd vtrip_sel_h vtrip_sel_h_n
*.PININFO en_h:I en_h_n:I enable_vddio_lv:I in_h:I in_vt:I mode_normal_n:I 
*.PININFO mode_ref_3v_n:I mode_ref_n:I mode_vccd_n:I vcchib:I vddio_q:I 
*.PININFO vrefin:I vssd:I vtrip_sel_h:I vtrip_sel_h_n:I ibufmux_out:O 
*.PININFO ibufmux_out_h:O
XICEnet43 net43 / icecap
XICEin_h in_h / icecap
XICEout_n out_n / icecap
XICEmode_vccd_n mode_vccd_n / icecap
XICEin_vt in_vt / icecap
XICEvrefin vrefin / icecap
XICEvtrip_sel_h vtrip_sel_h / icecap
XICEen_h_n en_h_n / icecap
XICEibufmux_out_h ibufmux_out_h / icecap
XICEibufmux_out ibufmux_out / icecap
XICEen_h en_h / icecap
XICEout out / icecap
XICEmode_normal_n mode_normal_n / icecap
XICEmode_ref_3v_n mode_ref_3v_n / icecap
XICEmode_ref_n mode_ref_n / icecap
XICEenable_vddio_lv enable_vddio_lv / icecap
XICEnet49 net49 / icecap
XICEvtrip_sel_h_n vtrip_sel_h_n / icecap
Xlvls enable_vddio_lv out ibufmux_out net43 vcchib vssd / 
+ sky130_fd_io__gpio_ovtv2_ipath_lvls
Xhvls en_h_n out out_n ibufmux_out_h net49 vddio_q vssd / 
+ sky130_fd_io__gpio_ovtv2_ipath_hvls
Xbuf en_h en_h_n enable_vddio_lv in_h in_vt mode_normal_n mode_ref_3v_n 
+ mode_ref_n mode_vccd_n out out_n vcchib vddio_q vrefin vssd vtrip_sel_h 
+ vtrip_sel_h_n / sky130_fd_io__gpio_ovtv2_in_buf
.ENDS
* .SUBCKT s8_esd_res250only_small pad rout
* *.PININFO pad:B rout:B
* rI175 net12 net16 sky130_fd_pr__res_generic_po m=1 w=2 l=10.07
* rI229 net16 rout sky130_fd_pr__res_generic_po m=1 w=2 l=0.17
* rI228 pad net12 sky130_fd_pr__res_generic_po m=1 w=2 l=0.17
* rI237<1> net16 rout short
* rI237<2> net16 rout short
* rI234<1> pad net12 short
* rI234<2> pad net12 short
* .ENDS
* .SUBCKT sky130_fd_io__gpio_ovtv2_buf_localesd in_h out_h out_vt vddio_q vssd 
* + vtrip_sel_h
* *.PININFO in_h:I vtrip_sel_h:I out_h:O out_vt:O vddio_q:B vssd:B
* XICEvtrip_sel_h vtrip_sel_h / icecap
* XICEin_h in_h / icecap
* XICEout_vt out_vt / icecap
* XICEout_h out_h / icecap
* mhv_passgate out_h vtrip_sel_h out_vt vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* Xesd_res in_h out_h / s8_esd_res250only_small
* Xggnfet6 vssd vddio_q vssd vddio_q out_h / s8_esd_signal_5_sym_hv_local_5term
* Xggnfet1 vssd out_h vssd vddio_q vssd / s8_esd_signal_5_sym_hv_local_5term
* .ENDS
* .SUBCKT sky130_fd_io__gpio_ovtv2_ictl_logic dm_h_n<2> dm_h_n<1> dm_h_n<0> hys_trim 
* + ibuf_mode_sel<0> ibuf_mode_sel<1> inp_dis_h_n inp_dis_i_h inp_dis_i_h_n 
* + mode_normal_n mode_ref_3v_n mode_ref_n mode_vccd_n tripsel_i_h tripsel_i_h_n 
* + vddio_q vssd vtrip_sel_h
* *.PININFO dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I hys_trim:I ibuf_mode_sel<0>:I 
* *.PININFO ibuf_mode_sel<1>:I inp_dis_h_n:I vddio_q:I vssd:I vtrip_sel_h:I 
* *.PININFO inp_dis_i_h:O inp_dis_i_h_n:O mode_normal_n:O mode_ref_3v_n:O 
* *.PININFO mode_ref_n:O mode_vccd_n:O tripsel_i_h:O tripsel_i_h_n:O
* XICEtripsel_i_h_n tripsel_i_h_n / icecap
* XICEmode_vccd_n mode_vccd_n / icecap
* XICEmode_ref_n mode_ref_n / icecap
* XICEibuf_mode_sel<1> ibuf_mode_sel<1> / icecap
* XICEinp_dis_i_h_n inp_dis_i_h_n / icecap
* XICEnet55 net55 / icecap
* XICEinp_dis_h_n inp_dis_h_n / icecap
* XICEinp_dis_i_h inp_dis_i_h / icecap
* XICEibuf_mode_sel<0> ibuf_mode_sel<0> / icecap
* XICEmode_ref_3v_n mode_ref_3v_n / icecap
* XICEtripsel_i_h tripsel_i_h / icecap
* XICEnand_dm01 nand_dm01 / icecap
* XICEmode_normal_n mode_normal_n / icecap
* XICEdm_h_n<0> dm_h_n<0> / icecap
* XICEand_dm01 and_dm01 / icecap
* XICEnet60 net60 / icecap
* XICEnet66 net66 / icecap
* XICEdm_buf_dis dm_buf_dis / icecap
* XICEdm_h_n<1> dm_h_n<1> / icecap
* XICEvtrip_sel_h vtrip_sel_h / icecap
* XICEmode_ref mode_ref / icecap
* XICEnet70 net70 / icecap
* XICEhys_trim hys_trim / icecap
* XICEdm_h_n<2> dm_h_n<2> / icecap
* XI41 net66 mode_normal_n tripsel_i_h vssd vddio_q / sky130_fd_io__hvsbt_nor
* XI34 ibuf_mode_sel<1> net70 net60 vssd vddio_q / sky130_fd_io__hvsbt_nor
* XI33 ibuf_mode_sel<1> ibuf_mode_sel<0> net55 vssd vddio_q / sky130_fd_io__hvsbt_nor
* Xdm10nand_inv nand_dm01 and_dm01 vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
* XI68 inp_dis_i_h inp_dis_i_h_n vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
* XI43 tripsel_i_h tripsel_i_h_n vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
* XI50 mode_ref_n mode_ref vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
* XI39 ibuf_mode_sel<0> net70 vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
* XI61 vtrip_sel_h net66 vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
* Xinpdis dm_buf_dis inp_dis_h_n inp_dis_i_h vssd vddio_q / sky130_fd_io__hvsbt_nand2
* Xdm210 dm_h_n<2> and_dm01 dm_buf_dis vssd vddio_q / sky130_fd_io__hvsbt_nand2
* Xdm10 dm_h_n<1> dm_h_n<0> nand_dm01 vssd vddio_q / sky130_fd_io__hvsbt_nand2
* XI40 inp_dis_i_h_n ibuf_mode_sel<1> mode_ref_n vssd vddio_q / 
* + sky130_fd_io__hvsbt_nand2
* XI36 inp_dis_i_h_n net60 mode_vccd_n vssd vddio_q / sky130_fd_io__hvsbt_nand2
* XI35 inp_dis_i_h_n net55 mode_normal_n vssd vddio_q / sky130_fd_io__hvsbt_nand2
* XI52 mode_ref hys_trim mode_ref_3v_n vssd vddio_q / sky130_fd_io__hvsbt_nand2
* .ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_ipath dm_h_n<2> dm_h_n<1> dm_h_n<0> 
+ enable_vddio_lv hys_trim_h ib_mode_sel_h<1> ib_mode_sel_h<0> inp_dis_h_n out 
+ out_h pad vcchib vddio_q vinref vssd vtrip_sel_h
*.PININFO dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I enable_vddio_lv:I hys_trim_h:I 
*.PININFO ib_mode_sel_h<1>:I ib_mode_sel_h<0>:I inp_dis_h_n:I vcchib:I 
*.PININFO vddio_q:I vssd:I vtrip_sel_h:I out:O out_h:O pad:B vinref:B
XICEib_mode_sel_h<0> ib_mode_sel_h<0> / icecap
XICEmode_ref_n mode_ref_n / icecap
XICEvtrip_sel_h vtrip_sel_h / icecap
XICEhys_trim_h hys_trim_h / icecap
XICEib_mode_sel_h<1> ib_mode_sel_h<1> / icecap
XICEinp_dis_h_n inp_dis_h_n / icecap
XI111<0> dm_h_n<2> / icecap
XI111<1> dm_h_n<1> / icecap
XI111<2> dm_h_n<0> / icecap
XICEin_vt in_vt / icecap
XICEen_h_n en_h_n / icecap
XICEmode_normal_n mode_normal_n / icecap
XICEpad pad / icecap
XICEtripsel_i_h_n tripsel_i_h_n / icecap
XICEout out / icecap
XICEenable_vddio_lv enable_vddio_lv / icecap
XICEen_h en_h / icecap
XICEvinref vinref / icecap
XICEmode_ref_3v_n mode_ref_3v_n / icecap
XICEmode_vccd_n mode_vccd_n / icecap
XICEtripsel_i_h tripsel_i_h / icecap
XICEin_h in_h / icecap
XICEout_h out_h / icecap
Xibuf_se en_h en_h_n enable_vddio_lv out out_h in_h in_vt mode_normal_n 
+ mode_ref_3v_n mode_ref_n mode_vccd_n vcchib vddio_q vinref vssd tripsel_i_h 
+ tripsel_i_h_n / sky130_fd_io__gpio_ovtv2_ibuf_se
Xesd pad in_h in_vt vddio_q vssd tripsel_i_h / sky130_fd_io__gpio_ovtv2_buf_localesd
Xlogic dm_h_n<2> dm_h_n<1> dm_h_n<0> hys_trim_h ib_mode_sel_h<0> 
+ ib_mode_sel_h<1> inp_dis_h_n en_h_n en_h mode_normal_n mode_ref_3v_n 
+ mode_ref_n mode_vccd_n tripsel_i_h tripsel_i_h_n vddio_q vssd vtrip_sel_h / 
+ sky130_fd_io__gpio_ovtv2_ictl_logic
.ENDS
.SUBCKT sky130_fd_io__top_gpio_ovtv2 amuxbus_a amuxbus_b analog_en analog_pol 
+ analog_sel dm<2> dm<1> dm<0> enable_h enable_inp_h enable_vdda_h 
+ enable_vddio enable_vswitch_h hld_h_n hld_ovr hys_trim ib_mode_sel<1> 
+ ib_mode_sel<0> in in_h inp_dis oe_n out pad pad_a_esd_0_h pad_a_esd_1_h 
+ pad_a_noesd_h slew_ctl<1> slew_ctl<0> slow tie_hi_esd tie_lo_esd vccd vcchib 
+ vdda vddio vddio_q vinref vssa vssd vssio vssio_q vswitch vtrip_sel
*.PININFO analog_en:I analog_pol:I analog_sel:I dm<2>:I dm<1>:I dm<0>:I 
*.PININFO enable_h:I enable_inp_h:I enable_vdda_h:I enable_vddio:I 
*.PININFO enable_vswitch_h:I hld_h_n:I hld_ovr:I hys_trim:I ib_mode_sel<1>:I 
*.PININFO ib_mode_sel<0>:I inp_dis:I oe_n:I out:I slew_ctl<1>:I slew_ctl<0>:I 
*.PININFO slow:I vinref:I vtrip_sel:I in:O in_h:O tie_hi_esd:O tie_lo_esd:O 
*.PININFO amuxbus_a:B amuxbus_b:B pad:B pad_a_esd_0_h:B pad_a_esd_1_h:B 
*.PININFO pad_a_noesd_h:B vccd:B vcchib:B vdda:B vddio:B vddio_q:B vssa:B 
*.PININFO vssd:B vssio:B vssio_q:B vswitch:B
Xopath dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n 
+ hld_i_ovr_h nga_pad_vpmp_h ngb_pad_vpmp_h od_i_h_n oe_n out pad pd_csd_h 
+ pghs_h pu_csd_h pug_h<6> pug_h<5> slew_ctl_h<1> slew_ctl_h<0> 
+ slew_ctl_h_n<1> slew_ctl_h_n<0> slow tie_hi_esd tie_lo_esd vccd vddio 
+ vddio_q vpb_drvr vcchib vssa vssd vssio vssio_q / 
+ sky130_fd_io__gpio_ovtv2_opath_i2c_fix_leak_fix
Xovt_amux amuxbus_a amuxbus_b analog_en analog_pol analog_sel enable_vdda_h 
+ enable_vswitch_h hld_i_h_n nga_pad_vpmp_h ngb_pad_vpmp_h tie_hi_esd out pad 
+ pd_csd_h pghs_h pu_csd_h pug_h<6> pug_h<5> vccd vdda vddio vddio_q vpb_drvr 
+ vssa vssd vssio vswitch / sky130_fd_io__gpio_ovtv2_amux_i2c_fix
Xctrl dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> 
+ enable_h enable_inp_h hld_h_n hld_i_h_n hld_i_ovr_h hld_ovr hys_trim 
+ hyst_trim_h net164 ib_mode_sel<1> ib_mode_sel<0> ib_mode_sel_h<1> 
+ ib_mode_sel_h<0> net166<0> net166<1> inp_dis inp_dis_h_n od_i_h_n 
+ slew_ctl<1> slew_ctl<0> slew_ctl_h<1> slew_ctl_h<0> slew_ctl_h_n<1> 
+ slew_ctl_h_n<0> vccd vddio_q vssd vtrip_sel vtrip_sel_h / 
+ sky130_fd_io__gpio_ctlv2_i2c_fix
XI336 net193 pad_a_esd_1_h / s8_esd_res75only_small
XI335 pad net193 / s8_esd_res75only_small
XI334 net189 pad_a_esd_0_h / s8_esd_res75only_small
Xresd4 pad net189 / s8_esd_res75only_small
rS0 pad pad_a_noesd_h short
Xipath dm_h_n<2> dm_h_n<1> dm_h_n<0> enable_vddio hyst_trim_h ib_mode_sel_h<1> 
+ ib_mode_sel_h<0> inp_dis_h_n in in_h pad vcchib vddio_q vinref vssd 
+ vtrip_sel_h / sky130_fd_io__gpio_ovtv2_ipath
.ENDS
* .SUBCKT sky130_fd_io__gpiov2_amux_switch amuxbus_hv ng_amx_vpmp_h ng_pad_vpmp_h 
* + nmid_vccd pad_hv_n0 pad_hv_n1 pad_hv_n2 pad_hv_n3 pad_hv_p0 pad_hv_p1 
* + pd_h_vdda pd_h_vddio pg_amx_vdda_h_n pg_pad_vddioq_h_n vdda vddio vssa vssd
* *.PININFO ng_amx_vpmp_h:I ng_pad_vpmp_h:I nmid_vccd:I pd_h_vdda:I pd_h_vddio:I 
* *.PININFO pg_amx_vdda_h_n:I pg_pad_vddioq_h_n:I vdda:I vddio:I vssa:I vssd:I 
* *.PININFO amuxbus_hv:B pad_hv_n0:B pad_hv_n1:B pad_hv_n2:B pad_hv_n3:B 
* *.PININFO pad_hv_p0:B pad_hv_p1:B
* XICEnet79 net79 / icecap
* XICEpad_hv_n1 pad_hv_n1 / icecap
* XICEpad_hv_n3 pad_hv_n3 / icecap
* XICEpd_h_vdda pd_h_vdda / icecap
* XICEng_pad_vpmp_h ng_pad_vpmp_h / icecap
* XICEpg_pad_vddioq_h_n pg_pad_vddioq_h_n / icecap
* XICEpg_amx_vdda_h_n pg_amx_vdda_h_n / icecap
* XICEpad_hv_n0 pad_hv_n0 / icecap
* XICEpad_hv_n2 pad_hv_n2 / icecap
* XICEng_amx_vpmp_h ng_amx_vpmp_h / icecap
* XICEnet77 net77 / icecap
* XICEpad_hv_p0 pad_hv_p0 / icecap
* XI85<0> mid / icecap
* XI85<1> mid1 / icecap
* XICEpad_hv_p1 pad_hv_p1 / icecap
* XICEamuxbus_hv amuxbus_hv / icecap
* XICEmid1 mid1 / icecap
* XICEpd_h_vddio pd_h_vddio / icecap
* XICEmid mid / icecap
* XICEnmid_vccd nmid_vccd / icecap
* xI72 vssa vdda condiode
* xI71 mid1 vdda condiode
* xI70 mid vdda condiode
* XI56 vssa net79 / s8_esd_res75only_small
* XI12 vssa net77 / s8_esd_res75only_small
* mI46 pad_hv_n3 ng_pad_vpmp_h mid1 mid1 sky130_fd_pr__nfet_g5v0d10v5 m=4 w=7.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI35 mid ng_pad_vpmp_h pad_hv_n1 mid sky130_fd_pr__nfet_g5v0d10v5 m=4 w=7.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI24 pad_hv_n0 ng_pad_vpmp_h mid mid sky130_fd_pr__nfet_g5v0d10v5 m=3 w=7.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI45 mid1 ng_pad_vpmp_h pad_hv_n2 mid1 sky130_fd_pr__nfet_g5v0d10v5 m=4 w=7.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI28 mid ng_amx_vpmp_h amuxbus_hv mid sky130_fd_pr__nfet_g5v0d10v5 m=7 w=7.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI57 mid1 nmid_vccd net79 vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI47 mid1 ng_amx_vpmp_h amuxbus_hv mid1 sky130_fd_pr__nfet_g5v0d10v5 m=7 w=7.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI78<1> mid pd_h_vdda vssa net043<0> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI78<0> mid1 pd_h_vdda vssa net043<1> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI77<1> mid pd_h_vddio vssa net044<0> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI77<0> mid1 pd_h_vddio vssa net044<1> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI1 mid nmid_vccd net77 vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI26 mid pg_amx_vdda_h_n amuxbus_hv vdda sky130_fd_pr__pfet_g5v0d10v5 m=5 w=7.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI22 mid pg_pad_vddioq_h_n pad_hv_p1 vddio sky130_fd_pr__pfet_g5v0d10v5 m=3 w=7.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI36 mid pg_pad_vddioq_h_n pad_hv_p0 vddio sky130_fd_pr__pfet_g5v0d10v5 m=3 w=7.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_amx_pucsd_inv A Y vda vssa
* *.PININFO A:I vda:I vssa:I Y:O
* XICEA A / icecap
* XICEY Y / icecap
* mI75 Y A vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=7 w=0.42 l=0.60 sa=265e-3 sb=265e-3 sd=280e-3 
* + topography=normal perim=1.14
* mI74 Y A vda vda sky130_fd_pr__pfet_g5v0d10v5 m=7 w=1.00 l=0.60 sa=265e-3 sb=265e-3 sd=280e-3 
* + topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_amux_drvr amux_en_vdda_h amux_en_vdda_h_n 
* + amux_en_vddio_h amux_en_vddio_h_n amux_en_vswitch_h amux_en_vswitch_h_n 
* + amuxbusa_on amuxbusa_on_n amuxbusb_on amuxbusb_on_n nga_amx_vswitch_h 
* + nga_pad_vswitch_h nga_pad_vswitch_h_n ngb_amx_vswitch_h ngb_pad_vswitch_h 
* + ngb_pad_vswitch_h_n nmida_on_n nmida_vccd nmida_vccd_n nmidb_on_n nmidb_vccd 
* + nmidb_vccd_n pd_csd_vswitch_h pd_csd_vswitch_h_n pd_on pd_on_n 
* + pga_amx_vdda_h_n pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n 
* + pu_csd_vddioq_h_n pu_on pu_on_n vccd vdda vddio_q vssa vssd vswitch
* *.PININFO amux_en_vdda_h:I amux_en_vdda_h_n:I amux_en_vddio_h:I 
* *.PININFO amux_en_vddio_h_n:I amux_en_vswitch_h:I amux_en_vswitch_h_n:I 
* *.PININFO amuxbusa_on:I amuxbusa_on_n:I amuxbusb_on:I amuxbusb_on_n:I 
* *.PININFO nmida_on_n:I nmidb_on_n:I pd_on:I pd_on_n:I pu_on:I pu_on_n:I vccd:I 
* *.PININFO vdda:I vddio_q:I vssa:I vssd:I vswitch:I nga_amx_vswitch_h:O 
* *.PININFO nga_pad_vswitch_h:O nga_pad_vswitch_h_n:O ngb_amx_vswitch_h:O 
* *.PININFO ngb_pad_vswitch_h:O ngb_pad_vswitch_h_n:O nmida_vccd:O 
* *.PININFO nmida_vccd_n:O nmidb_vccd:O nmidb_vccd_n:O pd_csd_vswitch_h:O 
* *.PININFO pd_csd_vswitch_h_n:O pga_amx_vdda_h_n:O pga_pad_vddioq_h_n:O 
* *.PININFO pgb_amx_vdda_h_n:O pgb_pad_vddioq_h_n:O pu_csd_vddioq_h_n:O
* XICEnmidb_vccd nmidb_vccd / icecap
* XICEamux_en_vddio_h amux_en_vddio_h / icecap
* XICEnga_pad_vswitch_h nga_pad_vswitch_h / icecap
* XICEnmidb_vccd_n nmidb_vccd_n / icecap
* XICEpu_on_n pu_on_n / icecap
* XICEnet272 net272 / icecap
* XICEamux_en_vswitch_h_n amux_en_vswitch_h_n / icecap
* XICEpd_on_n pd_on_n / icecap
* XICEnet236 net236 / icecap
* XICEngb_pad_vswitch_h ngb_pad_vswitch_h / icecap
* XICEamux_en_vdda_h_n amux_en_vdda_h_n / icecap
* XICEamux_en_vdda_h amux_en_vdda_h / icecap
* XICEpgb_amx_vdda_h_n pgb_amx_vdda_h_n / icecap
* XICEamux_en_vddio_h_n amux_en_vddio_h_n / icecap
* XICEnga_amx_vswitch_h nga_amx_vswitch_h / icecap
* XICEnet239 net239 / icecap
* XICEnet256 net256 / icecap
* XICEpgb_pad_vddioq_h_n pgb_pad_vddioq_h_n / icecap
* XICEamuxbusa_on amuxbusa_on / icecap
* XICEamux_en_vswitch_h amux_en_vswitch_h / icecap
* XICEpu_on pu_on / icecap
* XICEnet265 net265 / icecap
* XICEnmidb_on_n nmidb_on_n / icecap
* XICEnet274 net274 / icecap
* XICEnmida_vccd_n nmida_vccd_n / icecap
* XICEngb_pad_vswitch_h_n ngb_pad_vswitch_h_n / icecap
* XICEnet254 net254 / icecap
* XICEpga_pad_vddioq_h_n pga_pad_vddioq_h_n / icecap
* XICEngb_amx_vswitch_h ngb_amx_vswitch_h / icecap
* XICEnet275 net275 / icecap
* XICEpd_csd_vswitch_h_n pd_csd_vswitch_h_n / icecap
* XICEnmida_on_n nmida_on_n / icecap
* XICEnet248 net248 / icecap
* XICEnet257 net257 / icecap
* XICEpd_on pd_on / icecap
* XICEpd_csd_vswitch_h pd_csd_vswitch_h / icecap
* XICEpu_csd_vddioq_h_n pu_csd_vddioq_h_n / icecap
* XICEnet230 net230 / icecap
* XICEnga_pad_vswitch_h_n nga_pad_vswitch_h_n / icecap
* XICEamuxbusb_on_n amuxbusb_on_n / icecap
* XICEamuxbusb_on amuxbusb_on / icecap
* XICEnet245 net245 / icecap
* XICEnmida_vccd nmida_vccd / icecap
* XICEamuxbusa_on_n amuxbusa_on_n / icecap
* XICEpga_amx_vdda_h_n pga_amx_vdda_h_n / icecap
* XI93 nmida_vccd nmida_vccd_n vssd vccd / sky130_fd_io__hvsbt_inv_x1
* XI105 nmidb_vccd nmidb_vccd_n vssd vccd / sky130_fd_io__hvsbt_inv_x1
* XI38 net274 pu_csd_vddioq_h_n vddio_q vssd / sky130_fd_io__gpiov2_amx_pucsd_inv
* Xpga_amx_ls net265 net272 pga_amx_vdda_h_n amux_en_vdda_h_n amux_en_vdda_h 
* + vssa vdda / sky130_fd_io__gpiov2_amux_drvr_lshv2hv
* XI103 net239 net245 pgb_amx_vdda_h_n amux_en_vdda_h_n amux_en_vdda_h vssa vdda 
* + / sky130_fd_io__gpiov2_amux_drvr_lshv2hv
* XI45 net256 nga_amx_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_inv4
* XI42 net265 pga_pad_vddioq_h_n vddio_q vssd / sky130_fd_io__gpiov2_amx_inv4
* XI47 net256 nga_pad_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_inv4
* XI62 net239 pgb_pad_vddioq_h_n vddio_q vssd / sky130_fd_io__gpiov2_amx_inv4
* XI63 net236 ngb_amx_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_inv4
* XI64 net236 ngb_pad_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_inv4
* XI53 nmidb_on_n nmidb_vccd vssd vccd / sky130_fd_io__hvsbt_inv_x2
* XI89 nmida_on_n nmida_vccd vssd vccd / sky130_fd_io__hvsbt_inv_x2
* Xpdcsd_inv net254 pd_csd_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_pdcsd_inv
* XI90 pd_csd_vswitch_h pd_csd_vswitch_h_n vswitch vssa / sky130_fd_io__amx_inv1
* XI85 ngb_pad_vswitch_h ngb_pad_vswitch_h_n vswitch vssa / sky130_fd_io__amx_inv1
* XI87 nga_pad_vswitch_h nga_pad_vswitch_h_n vswitch vssa / sky130_fd_io__amx_inv1
* mI76 ngb_amx_vswitch_h amux_en_vdda_h_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI77 ngb_pad_vswitch_h amux_en_vddio_h_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI75 nga_amx_vswitch_h amux_en_vdda_h_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI78 nga_pad_vswitch_h amux_en_vddio_h_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI104 pd_csd_vswitch_h amux_en_vddio_h_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* Xpu_csd_ls pu_on pu_on_n net274 net275 amux_en_vddio_h_n amux_en_vddio_h vssd 
* + vddio_q vccd / sky130_fd_io__gpiov2_amux_drvr_ls
* Xpga_pad_ls amuxbusa_on amuxbusa_on_n net265 net272 amux_en_vddio_h_n 
* + amux_en_vddio_h vssd vddio_q vccd / sky130_fd_io__gpiov2_amux_drvr_ls
* Xnga_ls amuxbusa_on amuxbusa_on_n net257 net256 amux_en_vswitch_h_n 
* + amux_en_vswitch_h vssa vswitch vccd / sky130_fd_io__gpiov2_amux_drvr_ls
* Xpd_csd_ls pd_on pd_on_n net248 net254 amux_en_vswitch_h_n amux_en_vswitch_h 
* + vssa vswitch vccd / sky130_fd_io__gpiov2_amux_drvr_ls
* Xpgb_pad_ls amuxbusb_on amuxbusb_on_n net239 net245 amux_en_vddio_h_n 
* + amux_en_vddio_h vssd vddio_q vccd / sky130_fd_io__gpiov2_amux_drvr_ls
* Xngb_ls amuxbusb_on amuxbusb_on_n net230 net236 amux_en_vswitch_h_n 
* + amux_en_vswitch_h vssa vswitch vccd / sky130_fd_io__gpiov2_amux_drvr_ls
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_amux_ctl_ls in in_b out_h out_h_n rst_h rst_h_n vgnd 
* + vpwr_hv vpwr_lv
* *.PININFO in:I in_b:I rst_h:I rst_h_n:I vgnd:I vpwr_hv:I vpwr_lv:I out_h:O 
* *.PININFO out_h_n:O
* XICEout_h out_h / icecap
* XICEout_h_n out_h_n / icecap
* XICEnet61 net61 / icecap
* XICEfbk_n fbk_n / icecap
* XICEfbk fbk / icecap
* XICEin_b in_b / icecap
* XICErst_h rst_h / icecap
* XICEnet66 net66 / icecap
* XICEnet62 net62 / icecap
* XICEin in / icecap
* XICErst_h_n rst_h_n / icecap
* mI14 out_h fbk_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI11 out_h_n fbk vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI2 fbk_n fbk vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI1 fbk fbk_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI5 net61 rst_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=4 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI13 out_h fbk_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI12 out_h_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI58 fbk vpwr_lv net62 vgnd sky130_fd_pr__nfet_05v0_nvt m=4 w=1.00 l=0.90 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmnrst fbk rst_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI59 fbk_n vpwr_lv net66 vgnd sky130_fd_pr__nfet_05v0_nvt m=4 w=1.00 l=0.90 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI8 net66 in net61 vgnd sky130_fd_pr__nfet_01v8_lvt m=4 w=1.00 l=0.15 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI7 net62 in_b net61 vgnd sky130_fd_pr__nfet_01v8_lvt m=4 w=1.00 l=0.15 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_amux_ls amux_en_vdda_h amux_en_vdda_h_n 
* + amux_en_vddio_h amux_en_vddio_h_n amux_en_vswitch_h amux_en_vswitch_h_n 
* + analog_en enable_vdda_h enable_vdda_h_n enable_vswitch_h hld_i_h hld_i_h_n 
* + vccd vdda vddio_q vssa vssd vswitch
* *.PININFO analog_en:I enable_vdda_h:I enable_vswitch_h:I hld_i_h:I hld_i_h_n:I 
* *.PININFO vccd:I vdda:I vddio_q:I vssa:I vssd:I vswitch:I amux_en_vdda_h:O 
* *.PININFO amux_en_vdda_h_n:O amux_en_vddio_h:O amux_en_vddio_h_n:O 
* *.PININFO amux_en_vswitch_h:O amux_en_vswitch_h_n:O enable_vdda_h_n:O
* XICEanalog_en analog_en / icecap
* XICEenable_vswitch_h enable_vswitch_h / icecap
* XICEamux_en_vswitch_h amux_en_vswitch_h / icecap
* XICEhld_i_h_n hld_i_h_n / icecap
* XICEamux_en_vswitch_h_n amux_en_vswitch_h_n / icecap
* XICEenable_vdda_h_n enable_vdda_h_n / icecap
* XICEana_en_i_n ana_en_i_n / icecap
* XICEamux_en_vdda_h amux_en_vdda_h / icecap
* XICEhld_i_h hld_i_h / icecap
* XICEamux_en_vddio_h amux_en_vddio_h / icecap
* XICEana_en_i ana_en_i / icecap
* XICEenable_vdda_h enable_vdda_h / icecap
* XICEamux_en_vddio_h_n amux_en_vddio_h_n / icecap
* XICEnet74 net74 / icecap
* XICEamux_en_vdda_h_n amux_en_vdda_h_n / icecap
* XI32 enable_vdda_h enable_vdda_h_n vssa vdda / sky130_fd_io__gpiov2_amux_ls_inv_x1
* Xpd_vswitch_ls amux_en_vddio_h amux_en_vddio_h_n amux_en_vswitch_h 
* + amux_en_vswitch_h_n net74 enable_vswitch_h vssa vswitch / 
* + sky130_fd_io__gpiov2_amux_ctl_lshv2hv
* Xpd_vdda_ls amux_en_vddio_h amux_en_vddio_h_n amux_en_vdda_h amux_en_vdda_h_n 
* + enable_vdda_h_n enable_vdda_h vssa vdda / sky130_fd_io__gpiov2_amux_ctl_lshv2hv
* XI15 analog_en ana_en_i_n vssd vccd / sky130_fd_io__gpiov2_amux_ctl_inv_1
* XI16 ana_en_i_n ana_en_i vssd vccd / sky130_fd_io__gpiov2_amux_ctl_inv_1
* XI18 enable_vswitch_h net74 vssa vswitch / sky130_fd_io__hvsbt_inv_x1
* Xpd_vddio_ls ana_en_i ana_en_i_n amux_en_vddio_h amux_en_vddio_h_n hld_i_h 
* + hld_i_h_n vssd vddio_q vccd / sky130_fd_io__gpiov2_amux_ctl_ls
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_amux_ctl_logic analog_en analog_pol analog_sel 
* + enable_vdda_h enable_vdda_h_n enable_vswitch_h hld_i_h hld_i_h_n 
* + nga_amx_vswitch_h nga_pad_vswitch_h ngb_amx_vswitch_h ngb_pad_vswitch_h 
* + nmida_vccd nmidb_vccd out pd_csd_vswitch_h pga_amx_vdda_h_n 
* + pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n pu_csd_vddioq_h_n 
* + vccd vdda vddio_q vssa vssd vswitch
* *.PININFO analog_en:I analog_pol:I analog_sel:I enable_vdda_h:I 
* *.PININFO enable_vswitch_h:I hld_i_h:I hld_i_h_n:I out:I vccd:I vdda:I 
* *.PININFO vddio_q:I vssa:I vssd:I vswitch:I enable_vdda_h_n:O 
* *.PININFO nga_amx_vswitch_h:O nga_pad_vswitch_h:O ngb_amx_vswitch_h:O 
* *.PININFO ngb_pad_vswitch_h:O nmida_vccd:O nmidb_vccd:O pd_csd_vswitch_h:O 
* *.PININFO pga_amx_vdda_h_n:O pga_pad_vddioq_h_n:O pgb_amx_vdda_h_n:O 
* *.PININFO pgb_pad_vddioq_h_n:O pu_csd_vddioq_h_n:O
* XICEngb_pad_vswitch_h_n ngb_pad_vswitch_h_n / icecap
* XICEnga_pad_vswitch_h nga_pad_vswitch_h / icecap
* XICEnmida_vccd_n nmida_vccd_n / icecap
* XICEanalog_pol analog_pol / icecap
* XICEamux_en_vswitch_h_n amux_en_vswitch_h_n / icecap
* XICEnga_pad_vswitch_h_n nga_pad_vswitch_h_n / icecap
* XICEamux_en_vddio_h amux_en_vddio_h / icecap
* XICEngb_pad_vswitch_h ngb_pad_vswitch_h / icecap
* XICEenable_vdda_h_n enable_vdda_h_n / icecap
* XICEpga_pad_vddioq_h_n pga_pad_vddioq_h_n / icecap
* XICEamuxbusa_on_n amuxbusa_on_n / icecap
* XICEnmidb_vccd nmidb_vccd / icecap
* XICEpd_on_n pd_on_n / icecap
* XICEanalog_en analog_en / icecap
* XICEngb_amx_vswitch_h ngb_amx_vswitch_h / icecap
* XICEpgb_pad_vddioq_h_n pgb_pad_vddioq_h_n / icecap
* XICEamuxbusb_on_n amuxbusb_on_n / icecap
* XICEpd_csd_vswitch_h pd_csd_vswitch_h / icecap
* XICEpu_csd_vddioq_h_n pu_csd_vddioq_h_n / icecap
* XICEamux_en_vswitch_h amux_en_vswitch_h / icecap
* XICEhld_i_h hld_i_h / icecap
* XICEnmida_on_n nmida_on_n / icecap
* XICEamuxbusa_on amuxbusa_on / icecap
* XICEout out / icecap
* XICEnga_amx_vswitch_h nga_amx_vswitch_h / icecap
* XICEpd_csd_vswitch_h_n pd_csd_vswitch_h_n / icecap
* XICEpu_on_n pu_on_n / icecap
* XICEnmidb_on_n nmidb_on_n / icecap
* XICEpga_amx_vdda_h_n pga_amx_vdda_h_n / icecap
* XICEenable_vdda_h enable_vdda_h / icecap
* XICEenable_vswitch_h enable_vswitch_h / icecap
* XICEpd_on pd_on / icecap
* XICEhld_i_h_n hld_i_h_n / icecap
* XICEnmidb_vccd_n nmidb_vccd_n / icecap
* XICEnmida_vccd nmida_vccd / icecap
* XICEamux_en_vddio_h_n amux_en_vddio_h_n / icecap
* XICEamuxbusb_on amuxbusb_on / icecap
* XICEpu_on pu_on / icecap
* XICEpgb_amx_vdda_h_n pgb_amx_vdda_h_n / icecap
* XICEamux_en_vdda_h_n amux_en_vdda_h_n / icecap
* XICEamux_en_vdda_h amux_en_vdda_h / icecap
* XICEanalog_sel analog_sel / icecap
* Xamux_sw_drvr amux_en_vdda_h amux_en_vdda_h_n amux_en_vddio_h 
* + amux_en_vddio_h_n amux_en_vswitch_h amux_en_vswitch_h_n amuxbusa_on 
* + amuxbusa_on_n amuxbusb_on amuxbusb_on_n nga_amx_vswitch_h nga_pad_vswitch_h 
* + nga_pad_vswitch_h_n ngb_amx_vswitch_h ngb_pad_vswitch_h ngb_pad_vswitch_h_n 
* + nmida_on_n nmida_vccd nmida_vccd_n nmidb_on_n nmidb_vccd nmidb_vccd_n 
* + pd_csd_vswitch_h pd_csd_vswitch_h_n pd_on pd_on_n pga_amx_vdda_h_n 
* + pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n pu_csd_vddioq_h_n 
* + pu_on pu_on_n vccd vdda vddio_q vssa vssd vswitch / sky130_fd_io__gpiov2_amux_drvr
* Xamux_lv_decoder amuxbusa_on amuxbusa_on_n amuxbusb_on amuxbusb_on_n analog_en 
* + analog_pol analog_sel nga_pad_vswitch_h nga_pad_vswitch_h_n 
* + ngb_pad_vswitch_h ngb_pad_vswitch_h_n nmida_on_n nmida_vccd_n nmidb_on_n 
* + nmidb_vccd_n out pd_on pd_on_n pd_csd_vswitch_h_n pga_amx_vdda_h_n 
* + pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n pu_on pu_on_n 
* + pu_csd_vddioq_h_n vccd vssd / sky130_fd_io__gpiov2_amux_decoder
* Xamux_ls amux_en_vdda_h amux_en_vdda_h_n amux_en_vddio_h amux_en_vddio_h_n 
* + amux_en_vswitch_h amux_en_vswitch_h_n analog_en enable_vdda_h 
* + enable_vdda_h_n enable_vswitch_h hld_i_h hld_i_h_n vccd vdda vddio_q vssa 
* + vssd vswitch / sky130_fd_io__gpiov2_amux_ls
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_amux amuxbus_a amuxbus_b analog_en analog_pol 
* + analog_sel enable_vdda_h enable_vswitch_h hld_i_h hld_i_h_n out pad vccd 
* + vdda vddio_q vssa vssd vssio_q vswitch
* *.PININFO analog_en:I analog_pol:I analog_sel:I enable_vdda_h:I 
* *.PININFO enable_vswitch_h:I hld_i_h:I hld_i_h_n:I out:I vccd:I vdda:I 
* *.PININFO vddio_q:I vssa:I vssd:I vssio_q:I vswitch:I amuxbus_a:B amuxbus_b:B 
* *.PININFO pad:B
* XICEnet168 net168 / icecap
* XICEhld_i_h_n hld_i_h_n / icecap
* XICEamuxbus_a amuxbus_a / icecap
* XICEnet101 net101 / icecap
* XICEpga_pad_vddioq_h_n pga_pad_vddioq_h_n / icecap
* XICEanalog_pol analog_pol / icecap
* XICEpgb_pad_vddioq_h_n pgb_pad_vddioq_h_n / icecap
* XICEnet0127 net0127 / icecap
* XICEnet166 net166 / icecap
* XICEnmidb_vccd nmidb_vccd / icecap
* XICEanalog_en analog_en / icecap
* XICEnet99 net99 / icecap
* XICEenable_vdda_h enable_vdda_h / icecap
* XICEnet85 net85 / icecap
* XICEpgb_amx_vdda_h_n pgb_amx_vdda_h_n / icecap
* XICEpga_amx_vdda_h_n pga_amx_vdda_h_n / icecap
* XICEenable_vswitch_h enable_vswitch_h / icecap
* XICEpad pad / icecap
* XICEanalog_sel analog_sel / icecap
* XICEnet97 net97 / icecap
* XICEamuxbus_b amuxbus_b / icecap
* XICEnga_amx_vpmp_h nga_amx_vpmp_h / icecap
* XICEnet81 net81 / icecap
* XICEpd_csd_vswitch_h pd_csd_vswitch_h / icecap
* XICEout out / icecap
* XICEnet100 net100 / icecap
* XICEpu_csd_vddioq_h_n pu_csd_vddioq_h_n / icecap
* XICEnga_pad_vpmp_h nga_pad_vpmp_h / icecap
* XICEnmida_vccd nmida_vccd / icecap
* XICEngb_pad_vpmp_h ngb_pad_vpmp_h / icecap
* XICEhld_i_h hld_i_h / icecap
* XICEngb_amx_vpmp_h ngb_amx_vpmp_h / icecap
* xI43 vssio_q vdda condiode
* xI78 vssa vswitch condiode
* mI52 net81 pu_csd_vddioq_h_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=3 w=15.0 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mMP_PU net85 pu_csd_vddioq_h_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=4 w=15.0 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI49 net81 pd_csd_vswitch_h vssio_q vssio_q sky130_fd_pr__nfet_g5v0d10v5 m=6 w=5.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mMN_PD net85 pd_csd_vswitch_h vssio_q vssio_q sky130_fd_pr__nfet_g5v0d10v5 m=8 w=5.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* Xmux_a amuxbus_a nga_amx_vpmp_h nga_pad_vpmp_h nmida_vccd net101 net101 net97 
* + net97 net100 net99 net0127 hld_i_h pga_amx_vdda_h_n pga_pad_vddioq_h_n vdda 
* + vddio_q vssa vssd / sky130_fd_io__gpiov2_amux_switch
* Xmux_b amuxbus_b ngb_amx_vpmp_h ngb_pad_vpmp_h nmidb_vccd net101 net101 net97 
* + net97 net100 net99 net0127 hld_i_h pgb_amx_vdda_h_n pgb_pad_vddioq_h_n vdda 
* + vddio_q vssa vssd / sky130_fd_io__gpiov2_amux_switch
* XBBM_logic analog_en analog_pol analog_sel enable_vdda_h net0127 
* + enable_vswitch_h hld_i_h hld_i_h_n nga_amx_vpmp_h nga_pad_vpmp_h 
* + ngb_amx_vpmp_h ngb_pad_vpmp_h nmida_vccd nmidb_vccd out pd_csd_vswitch_h 
* + pga_amx_vdda_h_n pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n 
* + pu_csd_vddioq_h_n vccd vdda vddio_q vssa vssd vswitch / 
* + sky130_fd_io__gpiov2_amux_ctl_logic
* XI26 pad net99 / s8_esd_res75only_small
* XI58 net168 net97 / s8_esd_res75only_small
* XI28 net166 net101 / s8_esd_res75only_small
* XI57 pad net168 / s8_esd_res75only_small
* XI27 pad net100 / s8_esd_res75only_small
* XI55 pad pad / s8_esd_res75only_small
* XI54 pad net166 / s8_esd_res75only_small
* XI53 pad pad / s8_esd_res75only_small
* XI39 pad net81 / s8_esd_res75only_small
* XI40 pad net85 / s8_esd_res75only_small
* .ENDS
* .SUBCKT sky130_fd_io__com_pddrvr_unit_2_5 nd ngin ns
* *.PININFO ngin:I nd:B ns:B
* XICEngin ngin / icecap
* XICEnet10 ngin / icecap
* XICEnd nd / icecap
* mndrv nd ngin ns ns sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.60 sa=265e-3 sb=265e-3 sd=280e-3 
* + topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_pddrvr_strong pad pd_h<3> pd_h<2> pd_h_i2c tie_lo_esd 
* + vcc_io vgnd_io
* *.PININFO pd_h<3>:I pd_h<2>:I pd_h_i2c:I vcc_io:I vgnd_io:I pad:O tie_lo_esd:O
* XICEpd_h<2> pd_h<2> / icecap
* XICEpad pad / icecap
* XICEpd_h<3> pd_h<3> / icecap
* XICEnet78 net78 / icecap
* XICEnet80 net80 / icecap
* XICEpd_h_i2c pd_h_i2c / icecap
* XICEtie_lo_esd tie_lo_esd / icecap
* XICEnet66 net66 / icecap
* XICEnet76 net76 / icecap
* XICEnet68 net68 / icecap
* XICEnet72 net72 / icecap
* XICEnet46 net46 / icecap
* XI97 pd_h<3> net80 / sky130_fd_io__tk_em2s
* XI108 pd_h<3> net78 / sky130_fd_io__tk_em2s
* XI109 tie_lo_esd net76 / sky130_fd_io__tk_em2s
* XI102 pd_h<3> net72 / sky130_fd_io__tk_em2s
* XI104 pd_h<3> net68 / sky130_fd_io__tk_em2s
* XI96 pd_h<3> net66 / sky130_fd_io__tk_em2s
* XI113 pd_h<2> net46 / sky130_fd_io__tk_em2s
* XI99 tie_lo_esd net80 / sky130_fd_io__tk_em2o
* XI98 pd_h<2> net80 / sky130_fd_io__tk_em2o
* XI106 pd_h<2> net78 / sky130_fd_io__tk_em2o
* XI107 tie_lo_esd net78 / sky130_fd_io__tk_em2o
* XI110 pd_h<3> net76 / sky130_fd_io__tk_em2o
* XI111 pd_h<2> net76 / sky130_fd_io__tk_em2o
* XI100 tie_lo_esd net72 / sky130_fd_io__tk_em2o
* XI101 pd_h<2> net72 / sky130_fd_io__tk_em2o
* XI103 tie_lo_esd net68 / sky130_fd_io__tk_em2o
* XI105 pd_h<2> net68 / sky130_fd_io__tk_em2o
* XI95 pd_h<2> net66 / sky130_fd_io__tk_em2o
* XI94 tie_lo_esd net66 / sky130_fd_io__tk_em2o
* XI88 pd_h<3> net46 / sky130_fd_io__tk_em2o
* XI87 tie_lo_esd net46 / sky130_fd_io__tk_em2o
* XI49 vgnd_io tie_lo_esd / sky130_fd_io__tk_tie_r_out_esd
* Xn24<2> pad net80 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn24<1> pad net80 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn24<0> pad net80 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn23<2> pad net66 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn23<1> pad net66 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn23<0> pad net66 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn22<2> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn22<1> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn22<0> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn21<2> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn21<1> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn21<0> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn12 pad pd_h_i2c vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn32<2> pad net68 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn32<1> pad net68 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn32<0> pad net68 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn33<2> pad net78 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn33<1> pad net78 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn33<0> pad net78 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn34<3> pad net76 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn34<2> pad net76 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn34<1> pad net76 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn34<0> pad net76 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn11<2> pad pd_h<2> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn11<1> pad pd_h<2> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn11<0> pad pd_h<2> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn13 pad net46 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* Xn31 pad net72 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
* xI72 vgnd_io vcc_io condiode
* .ENDS
* .SUBCKT sky130_fd_io__gpio_pudrvr_unit_2_5 pd pgin ps
* *.PININFO pgin:I pd:B ps:B
* XICEnet10 pgin / icecap
* XICEpgin pgin / icecap
* XICEpd pd / icecap
* mpdrv pd pgin ps ps sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.60 sa=265e-3 sb=265e-3 sd=280e-3 
* + topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpio_pudrvr_strong pad pu_h_n<3> pu_h_n<2> tie_hi_esd vcc_io 
* + vnb
* *.PININFO pu_h_n<3>:I pu_h_n<2>:I vcc_io:I vnb:I pad:O tie_hi_esd:O
* XI112 pu_h_n<2> net43 / sky130_fd_io__tk_em2s
* XI108 tie_hi_esd net59 / sky130_fd_io__tk_em2s
* XI109 tie_hi_esd net53 / sky130_fd_io__tk_em2s
* XI104 pu_h_n<3> net49 / sky130_fd_io__tk_em2s
* XI125 pu_h_n<3> net45 / sky130_fd_io__tk_em2s
* XI83 pu_h_n<3> net43 / sky130_fd_io__tk_em2o
* XI82 tie_hi_esd net43 / sky130_fd_io__tk_em2o
* XI106 pu_h_n<2> net59 / sky130_fd_io__tk_em2o
* XI107 pu_h_n<3> net59 / sky130_fd_io__tk_em2o
* XI110 pu_h_n<3> net53 / sky130_fd_io__tk_em2o
* XI111 pu_h_n<2> net53 / sky130_fd_io__tk_em2o
* XI103 tie_hi_esd net49 / sky130_fd_io__tk_em2o
* XI105 pu_h_n<2> net49 / sky130_fd_io__tk_em2o
* XI124 tie_hi_esd net45 / sky130_fd_io__tk_em2o
* XI123 pu_h_n<2> net45 / sky130_fd_io__tk_em2o
* XI49 vcc_io tie_hi_esd / sky130_fd_io__tk_tie_r_out_esd
* Xn24<2> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn24<1> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn24<0> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn23<2> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn23<1> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn23<0> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn22 pad net45 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn21 pad pu_h_n<2> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn12<2> pad net43 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn12<1> pad net43 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn12<0> pad net43 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn32<2> pad net49 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn32<1> pad net49 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn32<0> pad net49 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn33<1> pad net59 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn33<0> pad net59 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn34<2> pad net53 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn34<1> pad net53 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn34<0> pad net53 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn11<2> pad pu_h_n<2> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn11<1> pad pu_h_n<2> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn11<0> pad pu_h_n<2> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn13<2> pad pu_h_n<2> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn13<1> pad pu_h_n<2> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn13<0> pad pu_h_n<2> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn31<2> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn31<1> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* Xn31<0> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
* .ENDS
* .SUBCKT sky130_fd_io__com_pudrvr_weak pad pu_h_n vcc_io vgnd_io vpb_drvr
* *.PININFO pu_h_n:I vcc_io:I vgnd_io:I vpb_drvr:I pad:O
* XICEpad pad / icecap
* XICEpu_h_n pu_h_n / icecap
* mpdrv pad pu_h_n vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=4 w=7.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI29 pad pu_h_n vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__com_pudrvr_strong_slow pad pu_h_n vcc_io vgnd_io vpb_drvr
* *.PININFO pu_h_n:I vcc_io:I vgnd_io:I vpb_drvr:I pad:O
* XICEpu_h_n pu_h_n / icecap
* XICEpad pad / icecap
* mpdrv pad pu_h_n vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=8 w=7.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_odrvr_sub force_hi_h_n pad pd_h<3> pd_h<2> pd_h<1> 
* + pd_h<0> pd_h_i2c pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> tie_hi_esd 
* + tie_lo_esd vcc_io vgnd vgnd_io
* *.PININFO force_hi_h_n:I pd_h<3>:I pd_h<2>:I pd_h<1>:I pd_h<0>:I pd_h_i2c:I 
* *.PININFO pu_h_n<3>:I pu_h_n<2>:I pu_h_n<1>:I pu_h_n<0>:I vcc_io:I vgnd:I 
* *.PININFO vgnd_io:I pad:O tie_hi_esd:B tie_lo_esd:B
* XICEpad pad / icecap
* XICEpu_h_n<0> pu_h_n<0> / icecap
* XICEpad_r250 pad_r250 / icecap
* XICEtie_hi_esd tie_hi_esd / icecap
* XICEweak_pad weak_pad / icecap
* XI75<0> pu_h_n<3> / icecap
* XI75<1> pu_h_n<2> / icecap
* XICEvgnd vgnd / icecap
* XI74<0> pd_h<3> / icecap
* XI74<1> pd_h<2> / icecap
* XICEpu_h_n<1> pu_h_n<1> / icecap
* XICEpd_h<1> pd_h<1> / icecap
* XICEpd_h_i2c pd_h_i2c / icecap
* XICEforce_hi_h_n force_hi_h_n / icecap
* XICEtie_lo_esd tie_lo_esd / icecap
* XICEstrong_slow_pad strong_slow_pad / icecap
* XICEpd_h<0> pd_h<0> / icecap
* Xpddrvr_strong pad pd_h<3> pd_h<2> pd_h_i2c tie_lo_esd vcc_io vgnd_io / 
* + sky130_fd_io__gpiov2_pddrvr_strong
* Xpudrvr_strong pad pu_h_n<3> pu_h_n<2> tie_hi_esd vcc_io vgnd / 
* + sky130_fd_io__gpio_pudrvr_strong
* Xpudrvr_weak weak_pad pu_h_n<0> vcc_io vgnd vcc_io / sky130_fd_io__com_pudrvr_weak
* Xpddrvr_weak weak_pad pd_h<0> vcc_io vgnd_io / sky130_fd_io__gpio_pddrvr_weak
* Xstrong_slow_pddrvr strong_slow_pad pd_h<1> vcc_io vgnd_io / 
* + sky130_fd_io__gpio_pddrvr_strong_slow
* Xstrong_slow_pudrvr strong_slow_pad pu_h_n<1> vcc_io vgnd vcc_io / 
* + sky130_fd_io__com_pudrvr_strong_slow
* Xres strong_slow_pad pad_r250 vgnd_io / sky130_fd_io__com_res_strong_slow
* Xres_weak weak_pad pad_r250 vgnd_io / sky130_fd_io__com_res_weak
* Xresd pad pad_r250 / s8_esd_res250only_small
* xI60 vgnd_io vcc_io condiode
* xI59 vgnd_io vcc_io condiode
* xI58 vgnd_io vcc_io condiode
* xI72 vgnd_io vcc_io condiode
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_odrvr force_hi_h_n pad pd_h<3> pd_h<2> pd_h<1> pd_h<0> 
* + pd_h_i2c pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> tie_hi_esd tie_lo_esd 
* + vcc_io vgnd vgnd_io
* *.PININFO force_hi_h_n:I pd_h<3>:I pd_h<2>:I pd_h<1>:I pd_h<0>:I pd_h_i2c:I 
* *.PININFO pu_h_n<3>:I pu_h_n<2>:I pu_h_n<1>:I pu_h_n<0>:I vcc_io:I vgnd:I 
* *.PININFO vgnd_io:I pad:O tie_hi_esd:O tie_lo_esd:O
* Xodrvr force_hi_h_n pad pd_h<3> pd_h<2> pd_h<1> pd_h<0> pd_h_i2c pu_h_n<3> 
* + pu_h_n<2> pu_h_n<1> pu_h_n<0> tie_hi_esd tie_lo_esd vcc_io vgnd vgnd_io / 
* + sky130_fd_io__gpiov2_odrvr_sub
* Xbondpad pad vgnd_io / sky130_fd_io__com_pad
* .ENDS
* .SUBCKT sky130_fd_io__com_cclat drvhi_h drvlo_h_n oe_h_n pd_dis_h pu_dis_h vcc_io 
* + vgnd
* *.PININFO oe_h_n:I pd_dis_h:I pu_dis_h:I vcc_io:I vgnd:I drvhi_h:O drvlo_h_n:O
* XICEpu_dis_h_n pu_dis_h_n / icecap
* XICEn0 n0 / icecap
* XICEn1 n1 / icecap
* XICEoe_i_h_n oe_i_h_n / icecap
* XICEpu_dis_h pu_dis_h / icecap
* XICEoe_h_n oe_h_n / icecap
* XICEdrvlo_h_n drvlo_h_n / icecap
* XICEoe_i_h oe_i_h / icecap
* XICEpd_dis_h pd_dis_h / icecap
* XICEdrvhi_h drvhi_h / icecap
* Xnor3 oe_i_h_n drvhi_h pd_dis_h n1 vcc_io vgnd vgnd / sky130_fd_io__com_cclat_hvnor3
* Xnand3 oe_i_h drvlo_h_n pu_dis_h_n n0 vcc_io vgnd vgnd / 
* + sky130_fd_io__com_cclat_hvnand3
* Xinv_oe1 oe_h_n oe_i_h vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_in
* Xinv_oe2 oe_i_h oe_i_h_n vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_in
* Xinv_pudis pu_dis_h pu_dis_h_n vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_in
* Xinv_out n1 drvlo_h_n vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_out
* Xinv_out_1 n0 drvhi_h vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_out
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_opath_datoe drvhi_h drvlo_h_n hld_h_n hld_i_ovr_h od_h 
* + oe_h oe_n out vcc_io vgnd vpwr_ka
* *.PININFO hld_h_n:I hld_i_ovr_h:I od_h:I oe_n:I out:I vcc_io:I vgnd:I 
* *.PININFO vpwr_ka:I drvhi_h:O drvlo_h_n:O oe_h:O
* XICEhld_h_n hld_h_n / icecap
* XICEdrvhi_h drvhi_h / icecap
* XICEout out / icecap
* XICEod_h od_h / icecap
* XICEoe_n oe_n / icecap
* XICEoe_h oe_h / icecap
* XICEoe_h_n oe_h_n / icecap
* XICEpd_dis_h pd_dis_h / icecap
* XICEpu_dis_h pu_dis_h / icecap
* XICEhld_i_ovr_h hld_i_ovr_h / icecap
* XICEdrvlo_h_n drvlo_h_n / icecap
* Xdat_ls hld_i_ovr_h out pd_dis_h pu_dis_h vgnd od_h vcc_io vgnd vpwr_ka / 
* + sky130_fd_io__gpio_dat_ls
* Xoe_ls hld_i_ovr_h oe_n oe_h_n oe_h vgnd od_h vcc_io vgnd vpwr_ka / 
* + sky130_fd_io__gpio_dat_ls
* Xcclat drvhi_h drvlo_h_n oe_h_n pd_dis_h pu_dis_h vcc_io vgnd / 
* + sky130_fd_io__com_cclat
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_octl dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
* + dm_h_n<0> hld_i_h_n od_h pden_h_n<2> pden_h_n<1> pden_h_n<0> puen_0_h 
* + puen_2or1_h puen_h<1> puen_h<0> slow slow_h slow_h_n vcc_io vgnd vpwr 
* + vreg_en_h_n
* *.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I 
* *.PININFO hld_i_h_n:I od_h:I slow:I vcc_io:I vgnd:I vpwr:I vreg_en_h_n:I 
* *.PININFO pden_h_n<2>:O pden_h_n<1>:O pden_h_n<0>:O puen_0_h:O puen_2or1_h:O 
* *.PININFO puen_h<1>:O puen_h<0>:O slow_h:O slow_h_n:O
* XICEn<5> n<5> / icecap
* XICEpuen_h<1> puen_h<1> / icecap
* XICEod_h od_h / icecap
* XICEvreg_en_h_n vreg_en_h_n / icecap
* XICEn<4> n<4> / icecap
* XICEpden_h0 pden_h0 / icecap
* XICEn<1> n<1> / icecap
* XICEn<2> n<2> / icecap
* XICEdm_h_n<0> dm_h_n<0> / icecap
* XICEpuen_h1_n puen_h1_n / icecap
* XICEn<3> n<3> / icecap
* XICEdm_h_n<2> dm_h_n<2> / icecap
* XICEnet70 net70 / icecap
* XICEpden_h_n<0> pden_h_n<0> / icecap
* XICEslow_h slow_h / icecap
* XICEslow slow / icecap
* XICEpuen_h0_n puen_h0_n / icecap
* XICEslow_h_n slow_h_n / icecap
* XICEn<9> n<9> / icecap
* XICEpuen_0_h puen_0_h / icecap
* XICEpuen_2or1_h puen_2or1_h / icecap
* XICEn<0> n<0> / icecap
* XICEn<8> n<8> / icecap
* XICEdm_h_n<1> dm_h_n<1> / icecap
* XICEdm_h<1> dm_h<1> / icecap
* XICEdm_h<2> dm_h<2> / icecap
* XICEpden_h_n<2> pden_h_n<2> / icecap
* XICEdm_h<0> dm_h<0> / icecap
* XICEpuen_h<0> puen_h<0> / icecap
* XICEnet130 net130 / icecap
* XICEpden_h_n<1> pden_h_n<1> / icecap
* XICEhld_i_h_n hld_i_h_n / icecap
* XICEn<10> n<10> / icecap
* XICEpden_h1 pden_h1 / icecap
* XI211 n<8> dm_h_n<1> puen_0_h vgnd vcc_io / sky130_fd_io__hvsbt_nor
* XI201 dm_h_n<2> dm_h_n<1> n<9> vgnd vcc_io / sky130_fd_io__hvsbt_nor
* XI381 dm_h<1> dm_h<0> net70 vgnd vcc_io / sky130_fd_io__hvsbt_nor
* XI210 dm_h<2> dm_h<0> n<8> vgnd vcc_io / sky130_fd_io__hvsbt_xor
* XI200 dm_h<2> dm_h<1> n<10> vgnd vcc_io / sky130_fd_io__hvsbt_xor
* XI185 dm_h_n<0> n<4> net130 vgnd vcc_io / sky130_fd_io__hvsbt_nand2
* XI186 dm_h_n<2> dm_h_n<1> n<4> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
* XI187 dm_h<1> dm_h<0> n<3> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
* XI208 puen_2or1_h vreg_en_h_n n<5> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
* XI203 n<10> dm_h<0> n<1> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
* XI204 n<9> dm_h_n<0> n<0> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
* XI205 n<1> n<0> puen_2or1_h vgnd vcc_io / sky130_fd_io__hvsbt_nand2
* XI382 dm_h<2> net70 pden_h_n<2> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
* XI254 puen_h1_n puen_h<1> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
* XI256 puen_h0_n puen_h<0> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
* XI249 pden_h0 pden_h_n<0> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
* XI247 pden_h1 pden_h_n<1> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
* XI377 puen_0_h puen_h0_n vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
* XI209 n<5> n<2> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
* XI376 n<2> puen_h1_n vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
* XI374 net130 pden_h1 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
* XI375 n<3> pden_h0 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
* Xls_slow hld_i_h_n slow slow_h slow_h_n od_h vgnd vcc_io vgnd vpwr / 
* + sky130_fd_io__com_ctl_ls
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_pupredrvr_strong_nd2 drvhi_h en_fast<3> en_fast<2> 
* + en_fast<1> en_fast<0> pu_h_n puen_h vcc_io vgnd_io
* *.PININFO drvhi_h:I en_fast<3>:I en_fast<2>:I en_fast<1>:I en_fast<0>:I 
* *.PININFO puen_h:I vcc_io:I vgnd_io:I pu_h_n:O
* XICEpuen_h puen_h / icecap
* XICEpu_h_n pu_h_n / icecap
* XI134<0> en_fast<3> / icecap
* XI134<1> en_fast<2> / icecap
* XI134<2> en_fast<1> / icecap
* XI134<3> en_fast<0> / icecap
* XICEint_res int_res / icecap
* XICEnet24 net24 / icecap
* XICEdrvhi_h drvhi_h / icecap
* XE1 net24 pu_h_n / sky130_fd_io__tk_em1s
* rrespu1 int_res net24 sky130_fd_pr__res_generic_po m=1 w=0.33 l=11
* rrespu2 pu_h_n int_res sky130_fd_pr__res_generic_po m=1 w=0.33 l=4
* mmnin_fast<3> net24 drvhi_h int<3> net013<0> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmnin_fast<2> net24 drvhi_h int<2> net013<1> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmnin_fast<1> net24 drvhi_h int<1> net013<2> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmnin_fast<0> net24 drvhi_h int<0> net013<3> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmnen_slow1 n<2> puen_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.00 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmnin_slow pu_h_n drvhi_h n<2> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.00 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmnen_fast<3> int<3> en_fast<3> vgnd_io net014<0> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=1.00 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmnen_fast<2> int<2> en_fast<2> vgnd_io net014<1> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=1.00 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmnen_fast<1> int<1> en_fast<1> vgnd_io net014<2> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=1.00 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmnen_fast<0> int<0> en_fast<0> vgnd_io net014<3> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=1.00 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmpen pu_h_n puen_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmpin pu_h_n drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=3 w=5.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_pupredrvr_strong drvhi_h pu_h_n<3> pu_h_n<2> puen_h 
* + slow_h_n vcc_io vgnd_io
* *.PININFO drvhi_h:I puen_h:I slow_h_n:I vcc_io:I vgnd_io:I pu_h_n<3>:O 
* *.PININFO pu_h_n<2>:O
* Xnd2b drvhi_h en_fast_h_3<3> en_fast_h_3<2> en_fast_h_3<1> en_fast_h_3<0> 
* + pu_h_n<3> puen_h vcc_io vgnd_io / sky130_fd_io__gpiov2_pupredrvr_strong_nd2
* Xnd2a drvhi_h net54 net54 net54 net54 pu_h_n<2> puen_h vcc_io vgnd_io / 
* + sky130_fd_io__gpiov2_pupredrvr_strong_nd2
* XI98 en_fast_h_3<0> en_fast_h_3<3> vgnd_io / sky130_fd_io__tk_opti
* XI97 en_fast_h_3<1> en_fast_h_3<3> vgnd_io / sky130_fd_io__tk_opti
* XI92 en_fast_h_3<3> nbias_out en_fast_h / sky130_fd_io__tk_opto
* XI96 en_fast_h_3<2> en_fast_h_3<3> vgnd_io / sky130_fd_io__tk_opto
* XI93 net54 nbias_out en_fast_h / sky130_fd_io__tk_opto
* Xinv en_fast_h_n en_fast_h vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
* Xnbias drvhi_h en_fast_h en_fast_h_n nbias_out pu_h_n<2> puen_h vcc_io vgnd_io 
* + / sky130_fd_io__com_pupredrvr_nbias
* Xnand puen_h slow_h_n en_fast_h_n vgnd_io vcc_io / sky130_fd_io__com_nand2_dnw
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_octl_mux a_h b_h sel_h sel_h_n vccio vssio y_h
* *.PININFO a_h:I b_h:I sel_h:I sel_h_n:I vccio:I vssio:I y_h:O
* XICEsel_h sel_h / icecap
* XICEy_h y_h / icecap
* XICEa_h a_h / icecap
* XICEsel_h_n sel_h_n / icecap
* XICEb_h b_h / icecap
* mI2 y_h sel_h b_h vccio sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI3 y_h sel_h_n a_h vccio sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI1 b_h sel_h_n y_h vssio sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI4 a_h sel_h y_h vssio sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_pdpredrvr_strong_nr2 drvlo_h_n en_fast_n<1> 
* + en_fast_n<0> i2c_mode_h pd_h pd_i2c_h pden_h_n vcc_io vgnd_io
* *.PININFO drvlo_h_n:I en_fast_n<1>:I en_fast_n<0>:I i2c_mode_h:I pden_h_n:I 
* *.PININFO vcc_io:I vgnd_io:I pd_h:O pd_i2c_h:O
* XICEpden_h_n pden_h_n / icecap
* XI105<0> net53<0> / icecap
* XI105<1> net53<1> / icecap
* XICEnet62 net62 / icecap
* XICEpd_i2c_h pd_i2c_h / icecap
* XICEi2c_mode_h i2c_mode_h / icecap
* XICEpd_h pd_h / icecap
* XI104<0> en_fast_n<1> / icecap
* XI104<1> en_fast_n<0> / icecap
* XICEen_fast_n<1> en_fast_n<1> / icecap
* XICEdrvlo_h_n drvlo_h_n / icecap
* XICEnet42 net42 / icecap
* mmpin_slow pd_i2c_h drvlo_h_n int_slow vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.00 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmpen_slow int_slow pden_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.00 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmpin_fast<1> pd_i2c_h drvlo_h_n net62 net030<0> sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmpin_fast<0> pd_i2c_h drvlo_h_n net62 net030<1> sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmpen_fast1 net62 en_fast_n<1> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI72<1> net53<0> en_fast_n<1> net42 net031<0> sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI72<0> net53<1> en_fast_n<0> net42 net031<1> sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI74<1> pd_h drvlo_h_n net53<0> net032<0> sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI74<0> pd_h drvlo_h_n net53<1> net032<1> sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI75 net039 pden_h_n net42 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.00 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI76 pd_h drvlo_h_n net45 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.00 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI73 net42 i2c_mode_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=3 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI101 net45 pden_h_n net039 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.00 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI94 pd_h i2c_mode_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmnin pd_i2c_h drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmnen pd_i2c_h pden_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI78 pd_h pden_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI77 pd_h drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_pdpredrvr_strong_nr3 drvlo_h_n en_fast_n<1> 
* + en_fast_n<0> i2c_mode_h pd_h pden_h_n vcc_io vgnd_io
* *.PININFO drvlo_h_n:I en_fast_n<1>:I en_fast_n<0>:I i2c_mode_h:I pden_h_n:I 
* *.PININFO vcc_io:I vgnd_io:I pd_h:O
* XI110<0> en_fast_n<1> / icecap
* XI110<1> en_fast_n<0> / icecap
* XICEint1 int1 / icecap
* XICEpden_h_n pden_h_n / icecap
* XICEpd_h pd_h / icecap
* XICEi2c_mode_h i2c_mode_h / icecap
* XICEint2 int2 / icecap
* XICEdrvlo_h_n drvlo_h_n / icecap
* mI85 int1 i2c_mode_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmpin_slow pd_h drvlo_h_n int_slow vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=2.00 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmpen_slow int_slow pden_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.00 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmpin_fast<1> pd_h drvlo_h_n int_nor<1> vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmpin_fast<0> pd_h drvlo_h_n int_nor<0> vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmpen_fast<1> int_nor<1> en_fast_n<1> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmpen_fast<0> int_nor<0> en_fast_n<0> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI90 pd_h drvlo_h_n net43 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=2.00 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI56 net43 pden_h_n int1 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=2.00 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI87<1> pd_h drvlo_h_n int2 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI87<0> pd_h drvlo_h_n int2 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI86<1> int2 en_fast_n<1> int1 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI86<0> int2 en_fast_n<0> int1 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmnin pd_h drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=5 w=3.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mmnen pd_h pden_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__com_pdpredrvr_pbias drvlo_h_n en_h en_h_n pbias pd_h pden_h_n 
* + vcc_io vgnd_io
* *.PININFO drvlo_h_n:I en_h:I en_h_n:I pd_h:I pden_h_n:I vcc_io:I vgnd_io:I 
* *.PININFO pbias:O
* XICEpbias pbias / icecap
* XICEpden_h_n pden_h_n / icecap
* XICEbias_g bias_g / icecap
* XICEnet157 net157 / icecap
* XICEnet108 net108 / icecap
* XICEn<101> n<101> / icecap
* XICEdrvlo_h_n drvlo_h_n / icecap
* XICEdrvlo_i_h drvlo_i_h / icecap
* XICEen_h en_h / icecap
* XICEpbias1 pbias1 / icecap
* XICEnet84 net84 / icecap
* XICEn<0> n<0> / icecap
* XICEn<1> n<1> / icecap
* XICE2vtp N0 / icecap
* XICEen_h_n en_h_n / icecap
* XICEpd_h pd_h / icecap
* XICEnet88 net88 / icecap
* XICEnet161 net161 / icecap
* XI27 n<0> pd_h en_h_n / sky130_fd_io__tk_opto
* XE1 n<1> n<0> / sky130_fd_io__tk_em1o
* XE2 pbias pbias1 / sky130_fd_io__tk_em1o
* XE3 pbias1 net88 / sky130_fd_io__tk_em1s
* XE4 net108 pbias / sky130_fd_io__tk_em1s
* XE6 pbias net84 / sky130_fd_io__tk_em1s
* XE5 n<101> bias_g / sky130_fd_io__tk_em1s
* mI47 pbias bias_g vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=1.00 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI24 n<1> drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI18 bias_g drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI23 n<0> n<0> n<1> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI13 drvlo_i_h drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI20 bias_g n<1> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI19 bias_g en_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI34 net157 bias_g vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI36 net108 bias_g vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=1.00 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI38 n<1> pden_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI48 n<100> pd_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.00 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI41 n<101> pd_h n<100> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.00 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI44 pbias pbias pbias1 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI45 pbias1 pbias1 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI15 net183 en_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI16 net171 n<0> net183 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI6 pbias en_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI12 drvlo_i_h drvlo_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI17 bias_g drvlo_h_n net171 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI14 pbias drvlo_i_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI33 N0 vgnd_io vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=8.00 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI32 net161 net161 N0 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI31 net157 net157 net161 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI30 net88 N0 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI43 net84 bias_g vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.00 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI40 N0 drvlo_i_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_pdpredrvr_strong drvlo_h_n i2c_mode_h_n pd_h<4> 
* + pd_h<3> pd_h<2> pden_h_n slow_h tie_hi_esd vcc_io vgnd vgnd_io
* *.PININFO drvlo_h_n:I i2c_mode_h_n:I pden_h_n:I slow_h:I tie_hi_esd:I vcc_io:I 
* *.PININFO vgnd:I vgnd_io:I pd_h<4>:O pd_h<3>:O pd_h<2>:O
* XICEpd_h<2> pd_h<2> / icecap
* XI162<0> en_fast2_n<1> / icecap
* XI162<1> en_fast2_n<0> / icecap
* XICEpden_h_n pden_h_n / icecap
* XICEmod_drvlo_h_n mod_drvlo_h_n / icecap
* XICEtie_hi_esd tie_hi_esd / icecap
* XICEnet142 net142 / icecap
* XICEen_fast2_n<0> en_fast2_n<0> / icecap
* XICEpd_h<3> pd_h<3> / icecap
* XICEmod_slow_h mod_slow_h / icecap
* XICEi2c_mode_h i2c_mode_h / icecap
* XICEnet75 net75 / icecap
* XICEen_fast_h_n en_fast_h_n / icecap
* XICEen_fast2_n<1> en_fast2_n<1> / icecap
* XICEdrvlo_h_n drvlo_h_n / icecap
* XICEslow_h slow_h / icecap
* XICEen_fast_h en_fast_h / icecap
* XI163<0> pbias_out / icecap
* XI163<1> pbias_out / icecap
* XICEint_slow1 int_slow1 / icecap
* XICEpbias_out pbias_out / icecap
* XICEi2c_mode_h_n i2c_mode_h_n / icecap
* XICEpd_h<4> pd_h<4> / icecap
* XICEmod_drvlo_h_n_i2c mod_drvlo_h_n_i2c / icecap
* XICEnet118 net118 / icecap
* mI87 mod_drvlo_h_n_i2c pd_h<4> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI88 mod_drvlo_h_n_i2c pd_h<4> vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* XI160 i2c_mode_h_n slow_h net75 vgnd vcc_io / sky130_fd_io__hvsbt_nand2
* XI98 i2c_mode_h slow_h int_slow1 vgnd vcc_io / sky130_fd_io__hvsbt_nand2
* XI161 net75 net142 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
* XI97 int_slow1 mod_slow_h vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
* XI93 i2c_mode_h_n i2c_mode_h vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
* Xmux mod_drvlo_h_n_i2c drvlo_h_n i2c_mode_h i2c_mode_h_n vcc_io vgnd_io 
* + mod_drvlo_h_n / sky130_fd_io__gpiov2_octl_mux
* Xnr3 drvlo_h_n pbias_out pbias_out mod_slow_h pd_h<2> pd_h<4> pden_h_n vcc_io 
* + vgnd_io / sky130_fd_io__gpiov2_pdpredrvr_strong_nr2
* Xnr2 mod_drvlo_h_n en_fast2_n<1> en_fast2_n<0> mod_slow_h pd_h<3> pden_h_n 
* + vcc_io vgnd_io / sky130_fd_io__gpiov2_pdpredrvr_strong_nr3
* XI77 en_fast2_n<1> pbias_out en_fast_h_n / sky130_fd_io__tk_opto
* XI76 net118 pbias_out en_fast_h_n / sky130_fd_io__tk_opto
* XI79 en_fast2_n<0> en_fast2_n<1> vcc_io / sky130_fd_io__tk_opti
* Xinv en_fast_h en_fast_h_n vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
* Xbias drvlo_h_n en_fast_h en_fast_h_n pbias_out pd_h<4> pden_h_n vcc_io 
* + vgnd_io / sky130_fd_io__com_pdpredrvr_pbias
* Xnor net142 pden_h_n en_fast_h vgnd_io vcc_io / sky130_fd_io__com_nor2_dnw
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_obpredrvr drvhi_h drvlo_h_n i2c_mode_h_n pd_h<4> 
* + pd_h<3> pd_h<2> pd_h<1> pd_h<0> pden_h_n<1> pden_h_n<0> pu_h_n<3> pu_h_n<2> 
* + pu_h_n<1> pu_h_n<0> puen_h<1> puen_h<0> slow_h slow_h_n tie_hi_esd vcc_io 
* + vgnd vgnd_io
* *.PININFO drvhi_h:I drvlo_h_n:I i2c_mode_h_n:I pden_h_n<1>:I pden_h_n<0>:I 
* *.PININFO puen_h<1>:I puen_h<0>:I slow_h:I slow_h_n:I tie_hi_esd:I vcc_io:I 
* *.PININFO vgnd:I vgnd_io:I pd_h<4>:O pd_h<3>:O pd_h<2>:O pd_h<1>:O pd_h<0>:O 
* *.PININFO pu_h_n<3>:O pu_h_n<2>:O pu_h_n<1>:O pu_h_n<0>:O
* XICEtie_hi_esd tie_hi_esd / icecap
* XICEpden_h_n<1> pden_h_n<1> / icecap
* XICEpu_h_n<0> pu_h_n<0> / icecap
* XICEpuen_h<1> puen_h<1> / icecap
* XICEslow_h slow_h / icecap
* XICEslow_h_n slow_h_n / icecap
* XICEpden_h_n<0> pden_h_n<0> / icecap
* XI125<0> pu_h_n<3> / icecap
* XI125<1> pu_h_n<2> / icecap
* XI126<0> pd_h<4> / icecap
* XI126<1> pd_h<3> / icecap
* XI126<2> pd_h<2> / icecap
* XICEi2c_mode_h_n i2c_mode_h_n / icecap
* XICEdrvhi_h drvhi_h / icecap
* XICEdrvlo_h_n drvlo_h_n / icecap
* XICEpu_h_n<1> pu_h_n<1> / icecap
* XICEpd_h<1> pd_h<1> / icecap
* XICEpuen_h<0> puen_h<0> / icecap
* XICEpd_h<0> pd_h<0> / icecap
* Xpu_strong drvhi_h pu_h_n<3> pu_h_n<2> puen_h<1> slow_h_n vcc_io vgnd_io / 
* + sky130_fd_io__gpiov2_pupredrvr_strong
* Xpd_strong drvlo_h_n i2c_mode_h_n pd_h<4> pd_h<3> pd_h<2> pden_h_n<1> slow_h 
* + tie_hi_esd vcc_io vgnd vgnd_io / sky130_fd_io__gpiov2_pdpredrvr_strong
* Xpu_weak drvhi_h pu_h_n<0> puen_h<0> vcc_io vgnd_io / 
* + sky130_fd_io__com_pupredrvr_weak
* Xpd_weak drvlo_h_n pd_h<0> pden_h_n<0> vcc_io vgnd_io / 
* + sky130_fd_io__com_pdpredrvr_weak
* Xpu_strong_slow drvhi_h pu_h_n<1> puen_h<1> vcc_io vgnd_io / 
* + sky130_fd_io__com_pupredrvr_strong_slow
* Xpd_strong_slow drvlo_h_n pd_h<1> pden_h_n<1> vcc_io vgnd_io / 
* + sky130_fd_io__com_pdpredrvr_strong_slow
* xI15 vgnd_io vcc_io condiode
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_octl_dat dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
* + dm_h_n<0> drvhi_h hld_i_h_n hld_i_ovr_h od_h oe_n out pd_h<4> pd_h<3> 
* + pd_h<2> pd_h<1> pd_h<0> pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> slow 
* + slow_h_n tie_hi_esd vcc_io vgnd vgnd_io vpwr vpwr_ka
* *.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I 
* *.PININFO hld_i_h_n:I hld_i_ovr_h:I od_h:I oe_n:I out:I slow:I tie_hi_esd:I 
* *.PININFO vcc_io:I vgnd:I vgnd_io:I vpwr:I vpwr_ka:I drvhi_h:O pd_h<4>:O 
* *.PININFO pd_h<3>:O pd_h<2>:O pd_h<1>:O pd_h<0>:O pu_h_n<3>:O pu_h_n<2>:O 
* *.PININFO pu_h_n<1>:O pu_h_n<0>:O slow_h_n:O
* XICEhld_i_h_n hld_i_h_n / icecap
* XI204<0> pden_h_n<2> / icecap
* XI204<1> pden_h_n<1> / icecap
* XI204<2> pden_h_n<0> / icecap
* XICEtie_hi_esd tie_hi_esd / icecap
* XI202<0> pd_h<4> / icecap
* XI202<1> pd_h<3> / icecap
* XI202<2> pd_h<2> / icecap
* XI202<3> pd_h<1> / icecap
* XI202<4> pd_h<0> / icecap
* XICEdrvlo_h_n drvlo_h_n / icecap
* XI200<0> pu_h_n<3> / icecap
* XI200<1> pu_h_n<2> / icecap
* XI200<2> pu_h_n<1> / icecap
* XI200<3> pu_h_n<0> / icecap
* XI203<0> pd_h<4> / icecap
* XI203<1> pd_h<3> / icecap
* XI203<2> pd_h<2> / icecap
* XI203<3> pd_h<1> / icecap
* XI203<4> pd_h<0> / icecap
* XI205<0> pu_h_n<3> / icecap
* XI205<1> pu_h_n<2> / icecap
* XI205<2> pu_h_n<1> / icecap
* XI205<3> pu_h_n<0> / icecap
* XICEpuen_0_h puen_0_h / icecap
* XI207<0> pden_h_n<1> / icecap
* XI207<1> pden_h_n<0> / icecap
* XICEhld_i_ovr_h hld_i_ovr_h / icecap
* XI201<0> dm_h_n<2> / icecap
* XI201<1> dm_h_n<1> / icecap
* XI201<2> dm_h_n<0> / icecap
* XICEod_h od_h / icecap
* XI206<0> puen_h<1> / icecap
* XI206<1> puen_h<0> / icecap
* XICEoe_n oe_n / icecap
* XICEout out / icecap
* XI199<0> dm_h<2> / icecap
* XI199<1> dm_h<1> / icecap
* XI199<2> dm_h<0> / icecap
* XICEpden_h_n<2> pden_h_n<2> / icecap
* XICEslow_h_n slow_h_n / icecap
* XICEpuen_2or1_h puen_2or1_h / icecap
* XICEslow_h slow_h / icecap
* XICEdrvhi_h drvhi_h / icecap
* XICEslow slow / icecap
* XICEoe_h oe_h / icecap
* Xdatoe drvhi_h drvlo_h_n hld_i_h_n hld_i_ovr_h od_h oe_h oe_n out vcc_io vgnd 
* + vpwr_ka / sky130_fd_io__gpiov2_opath_datoe
* Xctl dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n od_h 
* + pden_h_n<2> pden_h_n<1> pden_h_n<0> puen_0_h puen_2or1_h puen_h<1> puen_h<0> 
* + slow slow_h slow_h_n vcc_io vgnd vpwr vcc_io / sky130_fd_io__gpiov2_octl
* Xpredrvr drvhi_h drvlo_h_n pden_h_n<2> pd_h<4> pd_h<3> pd_h<2> pd_h<1> pd_h<0> 
* + pden_h_n<1> pden_h_n<0> pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> puen_h<1> 
* + puen_h<0> slow_h slow_h_n tie_hi_esd vcc_io vgnd vgnd_io / 
* + sky130_fd_io__gpiov2_obpredrvr
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_opath dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
* + dm_h_n<0> hld_i_h_n hld_i_ovr_h od_h oe_n out pad slow tie_hi_esd tie_lo_esd 
* + vcc_io vgnd vgnd_io vpwr vpwr_ka
* *.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I 
* *.PININFO hld_i_h_n:I hld_i_ovr_h:I od_h:I oe_n:I out:I slow:I vcc_io:I vgnd:I 
* *.PININFO vgnd_io:I vpwr:I vpwr_ka:I pad:O tie_hi_esd:O tie_lo_esd:O
* Xodrvr net70 pad pd_h<3> pd_h<2> pd_h<1> pd_h<0> pd_h<4> pu_h_n<3> pu_h_n<2> 
* + pu_h_n<1> pu_h_n<0> tie_hi_esd tie_lo_esd vcc_io vgnd vgnd_io / 
* + sky130_fd_io__gpiov2_odrvr
* Xopath dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> drvhi_h hld_i_h_n 
* + hld_i_ovr_h od_h oe_n out pd_h<4> pd_h<3> pd_h<2> pd_h<1> pd_h<0> pu_h_n<3> 
* + pu_h_n<2> pu_h_n<1> pu_h_n<0> slow slow_h_n tie_hi_esd vcc_io vgnd vgnd_io 
* + vpwr vpwr_ka / sky130_fd_io__gpiov2_octl_dat
* .ENDS
* .SUBCKT sky130_fd_io__hvsbt_inv_x4 in out vgnd vpwr
* *.PININFO in:I vgnd:I vpwr:I out:O
* XICEin in / icecap
* XICEout out / icecap
* mI1 out in vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=8 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI2 out in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=4 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__hvsbt_inv_x8 in out vgnd vpwr
* *.PININFO in:I vgnd:I vpwr:I out:O
* XICEout out / icecap
* XICEin in / icecap
* mI2 out in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=8 w=0.70 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI1 out in vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=16 w=1.00 l=0.60 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_ctl_hld enable_h hld_h_n hld_i_h hld_i_h_n hld_i_ovr_h 
* + hld_ovr od_i_h vcc_io vgnd vpwr
* *.PININFO enable_h:I hld_h_n:I hld_ovr:I vcc_io:I vgnd:I vpwr:I hld_i_h:O 
* *.PININFO hld_i_h_n:O hld_i_ovr_h:O od_i_h:O
* XICEenable_vdda_h_n enable_vdda_h_n / icecap
* XICEhld_ovr hld_ovr / icecap
* XICEod_i_h od_i_h / icecap
* XICEhld_h_n hld_h_n / icecap
* XICEod_h od_h / icecap
* XICEhld_ovr_h hld_ovr_h / icecap
* XICEod_i_h_n od_i_h_n / icecap
* XICEnet37 net37 / icecap
* XICEhld_i_ovr_h_n hld_i_ovr_h_n / icecap
* XICEnet65 net65 / icecap
* XICEenable_h enable_h / icecap
* XICEnet64 net64 / icecap
* XICEhld_i_ovr_h hld_i_ovr_h / icecap
* Xhld_ovr_ls net65 hld_ovr hld_ovr_h net37 od_h vgnd vcc_io vgnd vpwr / 
* + sky130_fd_io__com_ctl_ls
* XI30 od_i_h hld_i_ovr_h_n hld_i_ovr_h vgnd vcc_io / sky130_fd_io__hvsbt_nor
* XI26 net65 hld_ovr_h hld_i_ovr_h_n vgnd vcc_io / sky130_fd_io__hvsbt_nor
* Xhld_i_h_inv4 net65 enable_vdda_h_n vgnd vcc_io / sky130_fd_io__hvsbt_inv_x4
* XI31 od_i_h_n od_i_h vgnd vcc_io / sky130_fd_io__hvsbt_inv_x4
* Xhld_nand enable_h hld_h_n net64 vgnd vcc_io / sky130_fd_io__hvsbt_nand2
* Xod_h_inv enable_h od_h vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
* Xhld_i_h_inv1 net64 net65 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
* XI32 od_h od_i_h_n vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
* Xhld_i_h_inv8<1> enable_vdda_h_n hld_i_h_n_net<1> net019<0> net018<0> / 
* + sky130_fd_io__hvsbt_inv_x8
* Xhld_i_h_inv8<0> enable_vdda_h_n hld_i_h_n_net<0> net019<1> net018<1> / 
* + sky130_fd_io__hvsbt_inv_x8
* rshort<1> hld_i_h_n_net<1> hld_i_h_n short
* rshort<0> hld_i_h_n_net<0> hld_i_h_n short
* rshort_hld_i_h enable_vdda_h_n hld_i_h short
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_ctl_lsbank dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> 
* + dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n ib_mode_sel ib_mode_sel_h 
* + ib_mode_sel_h_n inp_dis inp_dis_h inp_dis_h_n od_i_h startup_rst_h 
* + startup_st_h vcc_io vgnd vpwr vtrip_sel vtrip_sel_h vtrip_sel_h_n
* *.PININFO dm<2>:I dm<1>:I dm<0>:I hld_i_h_n:I ib_mode_sel:I inp_dis:I od_i_h:I 
* *.PININFO startup_rst_h:I startup_st_h:I vcc_io:I vgnd:I vpwr:I vtrip_sel:I 
* *.PININFO dm_h<2>:O dm_h<1>:O dm_h<0>:O dm_h_n<2>:O dm_h_n<1>:O dm_h_n<0>:O 
* *.PININFO ib_mode_sel_h:O ib_mode_sel_h_n:O inp_dis_h:O inp_dis_h_n:O 
* *.PININFO vtrip_sel_h:O vtrip_sel_h_n:O
* XICEdm_h_n<0> dm_h_n<0> / icecap
* XICEie_n_rst_h ie_n_rst_h / icecap
* XICEdm_st_h<2> dm_st_h<2> / icecap
* XI660<0> dm_h_n<2> / icecap
* XI660<1> dm_h_n<1> / icecap
* XICEvtrip_sel_h vtrip_sel_h / icecap
* XICEinp_dis inp_dis / icecap
* XICEhld_i_h_n hld_i_h_n / icecap
* XICEib_mode_sel_h_n ib_mode_sel_h_n / icecap
* XICEdm_rst_h<2> dm_rst_h<2> / icecap
* XICEinp_dis_h inp_dis_h / icecap
* XICEtrip_sel_rst_h trip_sel_rst_h / icecap
* XICEvtrip_sel_h_n vtrip_sel_h_n / icecap
* XICEstartup_rst_h startup_rst_h / icecap
* XI659<0> dm_st_h<2> / icecap
* XI659<1> dm_st_h<1> / icecap
* XICEib_mode_sel_rst_h ib_mode_sel_rst_h / icecap
* XI663<0> dm_h<2> / icecap
* XI663<1> dm_h<1> / icecap
* XI662<0> dm_rst_h<2> / icecap
* XI662<1> dm_rst_h<1> / icecap
* XICEdm_st_h<1> dm_st_h<1> / icecap
* XICEvtrip_sel vtrip_sel / icecap
* XICEdm<0> dm<0> / icecap
* XICEib_mode_sel ib_mode_sel / icecap
* XICEdm_rst_h<1> dm_rst_h<1> / icecap
* XICEstartup_st_h startup_st_h / icecap
* XICEdm_h<0> dm_h<0> / icecap
* XICEdm_rst_h<0> dm_rst_h<0> / icecap
* XICEod_i_h od_i_h / icecap
* XICEib_mode_sel_h ib_mode_sel_h / icecap
* XICEinp_dis_h_n inp_dis_h_n / icecap
* XICEib_mode_sel_st_h ib_mode_sel_st_h / icecap
* XICEie_n_st_h ie_n_st_h / icecap
* XI661<0> dm<2> / icecap
* XI661<1> dm<1> / icecap
* XICEdm_st_h<0> dm_st_h<0> / icecap
* XICEtrip_sel_st_h trip_sel_st_h / icecap
* Xtrip_sel_st trip_sel_st_h od_i_h vgnd / sky130_fd_io__tk_opti
* Xtrip_sel_rst trip_sel_rst_h vgnd od_i_h / sky130_fd_io__tk_opti
* Xie_n_rst ie_n_rst_h startup_rst_h startup_st_h / sky130_fd_io__tk_opti
* Xie_n_st ie_n_st_h startup_st_h startup_rst_h / sky130_fd_io__tk_opti
* XI338<1> dm_rst_h<0> startup_st_h startup_rst_h / sky130_fd_io__tk_opti
* XI803<1> dm_st_h<1> od_i_h vgnd / sky130_fd_io__tk_opti
* XI802<1> dm_st_h<2> od_i_h vgnd / sky130_fd_io__tk_opti
* XI804<1> dm_rst_h<2> vgnd od_i_h / sky130_fd_io__tk_opti
* XI805<1> dm_rst_h<1> vgnd od_i_h / sky130_fd_io__tk_opti
* XI598 ib_mode_sel_st_h od_i_h vgnd / sky130_fd_io__tk_opti
* XI597 ib_mode_sel_rst_h vgnd od_i_h / sky130_fd_io__tk_opti
* XI337<1> dm_st_h<0> startup_rst_h startup_st_h / sky130_fd_io__tk_opti
* Xdm_ls<0> hld_i_h_n dm<0> dm_h<0> dm_h_n<0> dm_rst_h<0> dm_st_h<0> vcc_io vgnd 
* + vpwr / sky130_fd_io__com_ctl_ls
* Xinp_dis_ls hld_i_h_n inp_dis inp_dis_h inp_dis_h_n ie_n_rst_h ie_n_st_h 
* + vcc_io vgnd vpwr / sky130_fd_io__com_ctl_ls
* Xtrip_sel_ls hld_i_h_n vtrip_sel vtrip_sel_h vtrip_sel_h_n trip_sel_rst_h 
* + trip_sel_st_h vcc_io vgnd vpwr / sky130_fd_io__com_ctl_ls
* Xdm_ls<2> hld_i_h_n dm<2> dm_h<2> dm_h_n<2> dm_rst_h<2> dm_st_h<2> vcc_io vgnd 
* + vpwr / sky130_fd_io__com_ctl_ls
* Xdm_ls<1> hld_i_h_n dm<1> dm_h<1> dm_h_n<1> dm_rst_h<1> dm_st_h<1> vcc_io vgnd 
* + vpwr / sky130_fd_io__com_ctl_ls
* XI595 hld_i_h_n ib_mode_sel ib_mode_sel_h ib_mode_sel_h_n ib_mode_sel_rst_h 
* + ib_mode_sel_st_h vcc_io vgnd vpwr / sky130_fd_io__com_ctl_ls
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_ctl dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> 
* + dm_h_n<2> dm_h_n<1> dm_h_n<0> enable_h enable_inp_h hld_h_n hld_i_h 
* + hld_i_h_n hld_i_ovr_h hld_ovr ib_mode_sel ib_mode_sel_h ib_mode_sel_h_n 
* + inp_dis inp_dis_h_n od_i_h vcc_io vgnd vpwr vtrip_sel vtrip_sel_h 
* + vtrip_sel_h_n
* *.PININFO dm<2>:I dm<1>:I dm<0>:I enable_h:I enable_inp_h:I hld_h_n:I 
* *.PININFO hld_ovr:I ib_mode_sel:I inp_dis:I vcc_io:I vgnd:I vpwr:I vtrip_sel:I 
* *.PININFO dm_h<2>:O dm_h<1>:O dm_h<0>:O dm_h_n<2>:O dm_h_n<1>:O dm_h_n<0>:O 
* *.PININFO hld_i_h:O hld_i_h_n:O hld_i_ovr_h:O ib_mode_sel_h:O 
* *.PININFO ib_mode_sel_h_n:O inp_dis_h_n:O od_i_h:O vtrip_sel_h:O 
* *.PININFO vtrip_sel_h_n:O
* XICEnet92 net92 / icecap
* XICEvtrip_sel_h_n vtrip_sel_h_n / icecap
* XICEvtrip_sel vtrip_sel / icecap
* XICEstartup_rst_h startup_rst_h / icecap
* XICEinp_startup_en_h inp_startup_en_h / icecap
* XICEhld_i_h_n hld_i_h_n / icecap
* XICEib_mode_sel_h ib_mode_sel_h / icecap
* XI78<0> dm_h_n<2> / icecap
* XI78<1> dm_h_n<1> / icecap
* XI78<2> dm_h_n<0> / icecap
* XICEenable_h enable_h / icecap
* XICEib_mode_sel_h_n ib_mode_sel_h_n / icecap
* XICEib_mode_sel ib_mode_sel / icecap
* XICEhld_ovr hld_ovr / icecap
* XI76<0> dm_h<2> / icecap
* XI76<1> dm_h<1> / icecap
* XI76<2> dm_h<0> / icecap
* XICEinp_dis inp_dis / icecap
* XICEvtrip_sel_h vtrip_sel_h / icecap
* XICEnet80 net80 / icecap
* XICEhld_i_h hld_i_h / icecap
* XICEenable_inp_h enable_inp_h / icecap
* XICEhld_i_ovr_h hld_i_ovr_h / icecap
* XI77<0> dm<2> / icecap
* XI77<1> dm<1> / icecap
* XI77<2> dm<0> / icecap
* XICEod_i_h od_i_h / icecap
* XICEhld_h_n hld_h_n / icecap
* XICEinp_dis_h_n inp_dis_h_n / icecap
* XI75 enable_inp_h enable_h startup_rst_h vgnd vcc_io / sky130_fd_io__hvsbt_nor
* Xhld_dis_blk enable_h hld_h_n hld_i_h hld_i_h_n hld_i_ovr_h hld_ovr od_i_h 
* + vcc_io vgnd vpwr / sky130_fd_io__gpiov2_ctl_hld
* Xls_bank dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
* + dm_h_n<0> hld_i_h_n ib_mode_sel ib_mode_sel_h ib_mode_sel_h_n inp_dis net80 
* + inp_dis_h_n od_i_h startup_rst_h inp_startup_en_h vcc_io vgnd vpwr vtrip_sel 
* + vtrip_sel_h vtrip_sel_h_n / sky130_fd_io__gpiov2_ctl_lsbank
* XI56 od_i_h enable_inp_h net92 vgnd vcc_io / sky130_fd_io__hvsbt_nand2
* XI57 net92 inp_startup_en_h vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_inbuf_lvinv_x1 in out vgnd vnb vpb vpwr
* *.PININFO in:I vgnd:I vnb:I vpb:I vpwr:I out:O
* XICEout out / icecap
* XICEin in / icecap
* mI2 out in vgnd vnb sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.25 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI1 out in vpwr vpb sky130_fd_pr__pfet_01v8_hvt m=1 w=3.00 l=0.25 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_ipath_lvls in_vcchib in_vddio mode_normal_lv 
* + mode_normal_lv_n mode_vcchib_lv mode_vcchib_lv_n out out_b vcchib vssd
* *.PININFO in_vcchib:I in_vddio:I mode_normal_lv:I mode_normal_lv_n:I 
* *.PININFO mode_vcchib_lv:I mode_vcchib_lv_n:I vcchib:I vssd:I out:O out_b:O
* XICEin_vcchib in_vcchib / icecap
* XICEout out / icecap
* XICEmode_normal_lv mode_normal_lv / icecap
* XICEfbk_n fbk_n / icecap
* XICEmode_vcchib_lv mode_vcchib_lv / icecap
* XICEnet50 net50 / icecap
* XICEnet78 net78 / icecap
* XICEfbk fbk / icecap
* XICEmode_normal_lv_n mode_normal_lv_n / icecap
* XICEin_vddio in_vddio / icecap
* XICEnet95 net95 / icecap
* XICEmode_vcchib_lv_n mode_vcchib_lv_n / icecap
* XICEnet115 net115 / icecap
* XICEnet111 net111 / icecap
* XICEout_b out_b / icecap
* mI345 fbk_n in_vddio vcchib vcchib sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI344 net70 mode_vcchib_lv vcchib vcchib sky130_fd_pr__pfet_01v8 m=1 w=3.00 l=0.25 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI343 out_b fbk net78 vcchib sky130_fd_pr__pfet_01v8 m=2 w=3.00 l=0.25 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI342 net78 mode_normal_lv_n vcchib vcchib sky130_fd_pr__pfet_01v8 m=2 w=3.00 l=0.25 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI341 out_b mode_normal_lv net70 vcchib sky130_fd_pr__pfet_01v8 m=1 w=3.00 l=0.25 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI340 net50 mode_vcchib_lv_n vcchib vcchib sky130_fd_pr__pfet_01v8 m=2 w=3.00 l=0.25 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI339 fbk_n mode_normal_lv vcchib vcchib sky130_fd_pr__pfet_01v8 m=1 w=5.00 l=0.25 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI338 fbk fbk_n vcchib vcchib sky130_fd_pr__pfet_01v8 m=1 w=5.00 l=0.25 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI337 out out_b vcchib vcchib sky130_fd_pr__pfet_01v8 m=4 w=3.00 l=0.25 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI336 out_b in_vcchib net50 vcchib sky130_fd_pr__pfet_01v8 m=2 w=3.00 l=0.25 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI351 net111 mode_normal_lv vssd vssd sky130_fd_pr__nfet_01v8 m=2 w=3.00 l=0.25 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI350 out_b fbk net111 vssd sky130_fd_pr__nfet_01v8 m=2 w=3.00 l=0.25 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI349 out out_b vssd vssd sky130_fd_pr__nfet_01v8 m=2 w=3.00 l=0.25 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI348 fbk fbk_n vssd vssd sky130_fd_pr__nfet_01v8 m=1 w=3.00 l=0.25 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI347 net95 mode_vcchib_lv vssd vssd sky130_fd_pr__nfet_01v8 m=2 w=3.00 l=0.25 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI346 out_b in_vcchib net95 vssd sky130_fd_pr__nfet_01v8 m=2 w=3.00 l=0.25 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI353 fbk_n in_vddio net115 vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI352 net115 mode_normal_lv vssd vssd sky130_fd_pr__nfet_01v8 m=1 w=3.00 l=0.25 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_ipath_hvls in_vcchib in_vddio inb_vcchib mode_normal 
* + mode_normal_n mode_vcchib mode_vcchib_n out out_b vddio_q vssd
* *.PININFO in_vcchib:I in_vddio:I inb_vcchib:I mode_normal:I mode_normal_n:I 
* *.PININFO mode_vcchib:I mode_vcchib_n:I vddio_q:I vssd:I out:O out_b:O
* XICEinb_vcchib inb_vcchib / icecap
* XICEin_vcchib in_vcchib / icecap
* XICEnet75 net75 / icecap
* XICEin_vddio in_vddio / icecap
* XICEnet84 net84 / icecap
* XICEout out / icecap
* XICEout_b out_b / icecap
* XICEmode_vcchib_n mode_vcchib_n / icecap
* XICEnet92 net92 / icecap
* XICEfbk fbk / icecap
* XICEmode_normal mode_normal / icecap
* XICEfbk_b fbk_b / icecap
* XICEnet116 net116 / icecap
* XICEmode_normal_n mode_normal_n / icecap
* XICEnet55 net55 / icecap
* XICEmode_vcchib mode_vcchib / icecap
* mI325 fbk fbk_b vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI324 fbk_b fbk vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI323 net63 mode_normal vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI322 out_b in_vddio net75 vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI321 net75 mode_normal_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI320 out out_b vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=5 w=5.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI319 out_b mode_vcchib net63 vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI318 net55 mode_vcchib_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI317 out_b net84 net55 vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI336 net84 fbk_b vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI335 out_b net84 net88 vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI334 fbk inb_vcchib net116 vssd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI333 net116 mode_vcchib vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI332 net112 mode_normal vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI331 out out_b vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI330 out_b in_vddio net112 vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI329 fbk_b in_vcchib net92 vssd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI328 fbk mode_vcchib_n vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI327 net92 mode_vcchib vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI326 net88 mode_vcchib vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI337 net84 fbk_b vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_vcchib_in_buf in_h mode_vcchib_lv_n out out_n vcchib 
* + vssd
* *.PININFO in_h:I mode_vcchib_lv_n:I vcchib:I vssd:I out:O out_n:O
* XICEnet57 net57 / icecap
* XICEnet81 net81 / icecap
* XICEnet112 net112 / icecap
* XICEmode_vcchib_lv_n mode_vcchib_lv_n / icecap
* XICEout out / icecap
* XICEout_n out_n / icecap
* XICEnet108 net108 / icecap
* XICEin_b in_b / icecap
* XICEfbk fbk / icecap
* XICEin_h in_h / icecap
* mI420 net57 in_b fbk vssd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.00 l=0.80 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI552 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.80 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI544 fbk in_h vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.80 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI551 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.80 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI424 net81 in_b vssd vssd sky130_fd_pr__nfet_01v8 m=2 w=1.00 l=0.25 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI423 out_n net81 vssd vssd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.25 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI545 in_b in_h fbk vssd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.80 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI487 out out_n vssd vssd sky130_fd_pr__nfet_01v8 m=3 w=1.00 l=0.25 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI541 net81 mode_vcchib_lv_n vssd vssd sky130_fd_pr__nfet_01v8 m=2 w=1.00 l=0.25 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI549 net57 mode_vcchib_lv_n vcchib vcchib sky130_fd_pr__pfet_01v8 m=1 w=5.00 l=0.25 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI436 net81 in_b net112 vcchib sky130_fd_pr__pfet_01v8 m=2 w=1.00 l=0.25 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI543 in_b in_h net108 vcchib sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.80 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI429 out_n net81 vcchib vcchib sky130_fd_pr__pfet_01v8 m=1 w=5.00 l=0.25 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI538 net112 mode_vcchib_lv_n vcchib vcchib sky130_fd_pr__pfet_01v8 m=1 w=3.00 l=0.25 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI489 out out_n vcchib vcchib sky130_fd_pr__pfet_01v8 m=1 w=5.00 l=0.25 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI547 net108 mode_vcchib_lv_n vcchib vcchib sky130_fd_pr__pfet_01v8 m=3 w=5.00 l=0.25 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_in_buf in_h in_vt mode_normal_n out out_n vddio_q vssd 
* + vtrip_sel_h vtrip_sel_h_n
* *.PININFO in_h:I in_vt:I mode_normal_n:I vddio_q:I vssd:I vtrip_sel_h:I 
* *.PININFO vtrip_sel_h_n:I out:O out_n:O
* XICEmode_normal_n mode_normal_n / icecap
* XICEvtrip_sel_h vtrip_sel_h / icecap
* XICEnet122 net122 / icecap
* XICEin_h in_h / icecap
* XICEin_vt in_vt / icecap
* XICEnet158 net158 / icecap
* XICEnet103 net103 / icecap
* XICEmode_normal_cmos_h_n mode_normal_cmos_h_n / icecap
* XICEnet138 net138 / icecap
* XICEmode_normal_cmos_h mode_normal_cmos_h / icecap
* XICEnet91 net91 / icecap
* XICEvtrip_sel_h_n vtrip_sel_h_n / icecap
* XICEout out / icecap
* XICEfbk fbk / icecap
* XICEfbk2 fbk2 / icecap
* XICEout_n out_n / icecap
* XICEin_b in_b / icecap
* XI43 mode_normal_cmos_h mode_normal_cmos_h_n vssd vddio_q / 
* + sky130_fd_io__hvsbt_inv_x1
* XI488 vtrip_sel_h mode_normal_n mode_normal_cmos_h vssd vddio_q / 
* + sky130_fd_io__hvsbt_nor
* mI583 in_vt vtrip_sel_h_n vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI644 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.80 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI646 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.80 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI593 net91 mode_normal_n vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI592 net103 in_b fbk vssd sky130_fd_pr__nfet_g5v0d10v5 m=4 w=1.00 l=0.80 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI591 fbk in_h vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=6 w=5.00 l=0.80 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI590 fbk2 in_b fbk vssd sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.00 l=0.80 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI589 net91 in_b vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI588 fbk in_vt vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.80 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI587 in_b in_h fbk vssd sky130_fd_pr__nfet_g5v0d10v5 m=5 w=5.00 l=0.80 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI586 out_n net91 vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI642 out out_n vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
* + sd=280e-3 topography=normal perim=1.14
* mI629 in_b in_h net158 vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.80 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI636 net158 mode_normal_cmos_h_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI632 net122 mode_normal_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI647 vddio_q vddio_q vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.80 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI600 net103 mode_normal_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI598 net91 in_b net138 vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI597 fbk2 mode_normal_cmos_h_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI596 out_n net91 vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI595 net138 mode_normal_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 
* + sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI631 in_b in_h net122 vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.80 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* mI643 out out_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
* + sb=265e-3 sd=280e-3 topography=normal perim=1.14
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_ibuf_se enable_vddio_lv ibufmux_out ibufmux_out_h in_h 
* + in_vt mode_normal_n mode_vcchib_n vcchib vddio_q vssd vtrip_sel_h 
* + vtrip_sel_h_n
* *.PININFO enable_vddio_lv:I in_h:I in_vt:I mode_normal_n:I mode_vcchib_n:I 
* *.PININFO vcchib:I vddio_q:I vssd:I vtrip_sel_h:I vtrip_sel_h_n:I 
* *.PININFO ibufmux_out:O ibufmux_out_h:O
* XICEvtrip_sel_h vtrip_sel_h / icecap
* XICEout_n_vddio out_n_vddio / icecap
* XICEmode_vcchib mode_vcchib / icecap
* XICEmode_vcchib_lv_n mode_vcchib_lv_n / icecap
* XICEout_n_vcchib out_n_vcchib / icecap
* XICEmode_normal_lv_n mode_normal_lv_n / icecap
* XICEmode_normal mode_normal / icecap
* XICEin_h in_h / icecap
* XICEvtrip_sel_h_n vtrip_sel_h_n / icecap
* XICEout_vcchib out_vcchib / icecap
* XICEnet57 net57 / icecap
* XICEibufmux_out ibufmux_out / icecap
* XICEmode_vcchib_n mode_vcchib_n / icecap
* XICEibufmux_out_h ibufmux_out_h / icecap
* XICEmode_normal_lv mode_normal_lv / icecap
* XICEnet68 net68 / icecap
* XICEmode_normal_n mode_normal_n / icecap
* XICEout_vddio out_vddio / icecap
* XICEmode_vcchib_lv mode_vcchib_lv / icecap
* XICEin_vt in_vt / icecap
* XICEenable_vddio_lv enable_vddio_lv / icecap
* XI148 enable_vddio_lv mode_vcchib mode_vcchib_lv_n vssd vcchib / 
* + sky130_fd_io__hvsbt_nand2
* XI149 enable_vddio_lv mode_normal mode_normal_lv_n vssd vcchib / 
* + sky130_fd_io__hvsbt_nand2
* XI112 mode_normal_lv_n mode_normal_lv vssd vssd vcchib vcchib / 
* + sky130_fd_io__gpiov2_inbuf_lvinv_x1
* XI111 mode_vcchib_lv_n mode_vcchib_lv vssd vssd vcchib vcchib / 
* + sky130_fd_io__gpiov2_inbuf_lvinv_x1
* Xlvls out_vcchib out_vddio mode_normal_lv mode_normal_lv_n mode_vcchib_lv 
* + mode_vcchib_lv_n ibufmux_out net57 vcchib vssd / sky130_fd_io__gpiov2_ipath_lvls
* Xhvls out_vcchib out_vddio out_n_vcchib mode_normal mode_normal_n mode_vcchib 
* + mode_vcchib_n ibufmux_out_h net68 vddio_q vssd / sky130_fd_io__gpiov2_ipath_hvls
* XI88 in_h mode_vcchib_lv_n out_vcchib out_n_vcchib vcchib vssd / 
* + sky130_fd_io__gpiov2_vcchib_in_buf
* Xbuf in_h in_vt mode_normal_n out_vddio out_n_vddio vddio_q vssd vtrip_sel_h 
* + vtrip_sel_h_n / sky130_fd_io__gpiov2_in_buf
* XI491 mode_normal_n mode_normal vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
* XI105 mode_vcchib_n mode_vcchib vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_ictl_logic dm_h_n<2> dm_h_n<1> dm_h_n<0> ib_mode_sel_h 
* + ib_mode_sel_h_n inp_dis_h_n inp_dis_i_h inp_dis_i_h_n mode_normal_n 
* + mode_vcchib_n tripsel_i_h tripsel_i_h_n vddio_q vssd vtrip_sel_h_n
* *.PININFO dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I ib_mode_sel_h:I 
* *.PININFO ib_mode_sel_h_n:I inp_dis_h_n:I vddio_q:I vssd:I vtrip_sel_h_n:I 
* *.PININFO inp_dis_i_h:O inp_dis_i_h_n:O mode_normal_n:O mode_vcchib_n:O 
* *.PININFO tripsel_i_h:O tripsel_i_h_n:O
* XICEdm_buf_dis_n dm_buf_dis_n / icecap
* XICEvtrip_sel_h_n vtrip_sel_h_n / icecap
* XICEand_dm01 and_dm01 / icecap
* XICEdm_h_n<1> dm_h_n<1> / icecap
* XICEib_mode_sel_h_n ib_mode_sel_h_n / icecap
* XICEinp_dis_i_h inp_dis_i_h / icecap
* XICEnand_dm01 nand_dm01 / icecap
* XICEtripsel_i_h_n tripsel_i_h_n / icecap
* XICEinp_dis_h_n inp_dis_h_n / icecap
* XICEinp_dis_i_h_n inp_dis_i_h_n / icecap
* XICEtripsel_i_h tripsel_i_h / icecap
* XICEdm_h_n<2> dm_h_n<2> / icecap
* XICEmode_normal_n mode_normal_n / icecap
* XICEmode_vcchib_n mode_vcchib_n / icecap
* XICEdm_h_n<0> dm_h_n<0> / icecap
* XICEib_mode_sel_h ib_mode_sel_h / icecap
* XI71 vtrip_sel_h_n mode_normal_n tripsel_i_h vssd vddio_q / sky130_fd_io__hvsbt_nor
* XI80 dm_buf_dis_n inp_dis_h_n inp_dis_i_h vssd vddio_q / sky130_fd_io__hvsbt_nand2
* XI79 dm_h_n<2> and_dm01 dm_buf_dis_n vssd vddio_q / sky130_fd_io__hvsbt_nand2
* XI78 dm_h_n<1> dm_h_n<0> nand_dm01 vssd vddio_q / sky130_fd_io__hvsbt_nand2
* XI36 inp_dis_i_h_n ib_mode_sel_h mode_vcchib_n vssd vddio_q / 
* + sky130_fd_io__hvsbt_nand2
* XI35 inp_dis_i_h_n ib_mode_sel_h_n mode_normal_n vssd vddio_q / 
* + sky130_fd_io__hvsbt_nand2
* XI111 inp_dis_i_h inp_dis_i_h_n vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
* XI75 nand_dm01 and_dm01 vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
* XI74 tripsel_i_h tripsel_i_h_n vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
* .ENDS
* .SUBCKT sky130_fd_io__gpiov2_ipath dm_h_n<2> dm_h_n<1> dm_h_n<0> enable_vddio_lv 
* + ib_mode_sel_h ib_mode_sel_h_n inp_dis_h_n out out_h pad vcchib vddio_q vssd 
* + vtrip_sel_h_n
* *.PININFO dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I enable_vddio_lv:I 
* *.PININFO ib_mode_sel_h:I ib_mode_sel_h_n:I inp_dis_h_n:I vcchib:I vddio_q:I 
* *.PININFO vssd:I vtrip_sel_h_n:I out:O out_h:O pad:B
* XICEinp_dis_h_n inp_dis_h_n / icecap
* XICEin_h in_h / icecap
* XICEmode_normal_n mode_normal_n / icecap
* XICEen_h_n en_h_n / icecap
* XICEpad pad / icecap
* XICEen_h en_h / icecap
* XICEout_h out_h / icecap
* XICEin_vt in_vt / icecap
* XICEvtrip_sel_h_n vtrip_sel_h_n / icecap
* XICEenable_vddio_lv enable_vddio_lv / icecap
* XICEtripsel_i_h tripsel_i_h / icecap
* XICEib_mode_sel_h_n ib_mode_sel_h_n / icecap
* XI152<0> dm_h_n<2> / icecap
* XI152<1> dm_h_n<1> / icecap
* XI152<2> dm_h_n<0> / icecap
* XICEtripsel_i_h_n tripsel_i_h_n / icecap
* XICEib_mode_sel_h ib_mode_sel_h / icecap
* XICEmode_vcchib_n mode_vcchib_n / icecap
* XICEout out / icecap
* XI106 enable_vddio_lv out out_h in_h in_vt mode_normal_n mode_vcchib_n vcchib 
* + vddio_q vssd tripsel_i_h tripsel_i_h_n / sky130_fd_io__gpiov2_ibuf_se
* XI107 dm_h_n<2> dm_h_n<1> dm_h_n<0> ib_mode_sel_h ib_mode_sel_h_n inp_dis_h_n 
* + en_h_n en_h mode_normal_n mode_vcchib_n tripsel_i_h tripsel_i_h_n vddio_q 
* + vssd vtrip_sel_h_n / sky130_fd_io__gpiov2_ictl_logic
* XI120 pad in_h in_vt vddio_q vssd tripsel_i_h / 
* + sky130_fd_io__gpio_ovtv2_buf_localesd
* .ENDS
* .SUBCKT sky130_fd_io__top_gpiov2 amuxbus_a amuxbus_b analog_en analog_pol 
* + analog_sel dm<2> dm<1> dm<0> enable_h enable_inp_h enable_vdda_h 
* + enable_vddio enable_vswitch_h hld_h_n hld_ovr ib_mode_sel in in_h inp_dis 
* + oe_n out pad pad_a_esd_0_h pad_a_esd_1_h pad_a_noesd_h slow tie_hi_esd 
* + tie_lo_esd vccd vcchib vdda vddio vddio_q vssa vssd vssio vssio_q vswitch 
* + vtrip_sel
* *.PININFO analog_en:I analog_pol:I analog_sel:I dm<2>:I dm<1>:I dm<0>:I 
* *.PININFO enable_h:I enable_inp_h:I enable_vdda_h:I enable_vddio:I 
* *.PININFO enable_vswitch_h:I hld_h_n:I hld_ovr:I ib_mode_sel:I inp_dis:I 
* *.PININFO oe_n:I out:I slow:I vtrip_sel:I in:O in_h:O tie_hi_esd:O 
* *.PININFO tie_lo_esd:O amuxbus_a:B amuxbus_b:B pad:B pad_a_esd_0_h:B 
* *.PININFO pad_a_esd_1_h:B pad_a_noesd_h:B vccd:B vcchib:B vdda:B vddio:B 
* *.PININFO vddio_q:B vssa:B vssd:B vssio:B vssio_q:B vswitch:B
* Xamux amuxbus_a amuxbus_b analog_en analog_pol analog_sel enable_vdda_h 
* + enable_vswitch_h hld_i_h hld_i_h_n out pad vccd vdda vddio_q vssa vssd 
* + vssio_q vswitch / sky130_fd_io__gpiov2_amux
* Xopath dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n 
* + hld_i_ovr_h od_i_h oe_n out pad slow tie_hi_esd tie_lo_esd vddio vssd vssio 
* + vccd vcchib / sky130_fd_io__gpiov2_opath
* Xctrl dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> 
* + enable_h enable_inp_h hld_h_n hld_i_h hld_i_h_n hld_i_ovr_h hld_ovr 
* + ib_mode_sel ib_mode_sel_h ib_mode_sel_h_n inp_dis inp_dis_h_n od_i_h vddio_q 
* + vssd vccd vtrip_sel vtrip_sel_h vtrip_sel_h_n / sky130_fd_io__gpiov2_ctl
* Xipath dm_h_n<2> dm_h_n<1> dm_h_n<0> enable_vddio ib_mode_sel_h 
* + ib_mode_sel_h_n inp_dis_h_n in in_h pad vcchib vddio_q vssd vtrip_sel_h_n / 
* + sky130_fd_io__gpiov2_ipath
* Xresd3 pad_a_esd_1_h net210 / s8_esd_res75only_small
* Xresd1 net204 pad / s8_esd_res75only_small
* Xresd4 net210 pad / s8_esd_res75only_small
* Xresd2 pad_a_esd_0_h net204 / s8_esd_res75only_small
* XICEoe_n oe_n / icecap
* XICEhld_h_n hld_h_n / icecap
* XICEslow slow / icecap
* XICEpad pad / icecap
* XICEtie_hi_esd tie_hi_esd / icecap
* XI259<0> dm_h_n<2> / icecap
* XI259<1> dm_h_n<1> / icecap
* XI259<2> dm_h_n<0> / icecap
* XI257<0> dm_h<2> / icecap
* XI257<1> dm_h<1> / icecap
* XI257<2> dm_h<0> / icecap
* XICEhld_i_h_n hld_i_h_n / icecap
* XICEtie_lo_esd tie_lo_esd / icecap
* XI258<0> dm<2> / icecap
* XI258<1> dm<1> / icecap
* XI258<2> dm<0> / icecap
* XICEinp_dis inp_dis / icecap
* XICEhld_i_ovr_h hld_i_ovr_h / icecap
* XICEhld_ovr hld_ovr / icecap
* XICEout out / icecap
* XICEvtrip_sel vtrip_sel / icecap
* XICEod_h od_i_h / icecap
* rS0<2> pad pad_a_noesd_h short
* rS0<1> pad pad_a_noesd_h short
* rS0<0> pad pad_a_noesd_h short
* .ENDS

.SUBCKT s8_esd_gnd2gnd_120x2_lv_isosub vssi vssn vsub
*.PININFO vssi:B vssn:B vsub:B
dI9 vssn vssi sky130_fd_pr__diode_pd2nw_05v5 m=4 pj=33
dI10 vssi vssn sky130_fd_pr__diode_pd2nw_05v5 m=4 pj=33
.ENDS

.SUBCKT sky130_fd_io__top_power_lvc_wpad amuxbus_a amuxbus_b bdy2_b2b drn_lvc1 
+ drn_lvc2 ogc_lvc p_core p_pad src_bdy_lvc1 src_bdy_lvc2 vccd vcchib vdda 
+ vddio vddio_q vssa vssd vssio vssio_q vswitch
*.PININFO amuxbus_a:B amuxbus_b:B bdy2_b2b:B drn_lvc1:B drn_lvc2:B ogc_lvc:B 
*.PININFO p_core:B p_pad:B src_bdy_lvc1:B src_bdy_lvc2:B vccd:B vcchib:B 
*.PININFO vdda:B vddio:B vddio_q:B vssa:B vssd:B vssio:B vssio_q:B vswitch:B
Xesd bdy2_b2b src_bdy_lvc1 vssd / s8_esd_gnd2gnd_120x2_lv_isosub
xI54 src_bdy_lvc2 vddio condiode
xI50 src_bdy_lvc1 vddio condiode
rI21 p_pad p_core short
mpre_p1 g_nclamp_lvc1 g_pdpre_lvc1 drn_lvc1 drn_lvc1 sky130_fd_pr__pfet_01v8 m=20 w=7.00 l=0.18 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI40 g_nclamp_lvc2 g_pdpre_lvc2 drn_lvc2 drn_lvc2 sky130_fd_pr__pfet_01v8 m=20 w=7.00 l=0.18 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mclamp_xtor drn_lvc1 g_nclamp_lvc1 src_bdy_lvc1 src_bdy_lvc1 sky130_fd_pr__nfet_01v8 m=166 
+ w=7.00 l=0.18 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ perim=1.14
mI42 drn_lvc2 g_nclamp_lvc2 src_bdy_lvc2 src_bdy_lvc2 sky130_fd_pr__nfet_01v8 m=152 w=7.00 
+ l=0.18 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ perim=1.14
mI61 drn_lvc2 g_nclamp_lvc2 src_bdy_lvc2 src_bdy_lvc2 sky130_fd_pr__nfet_01v8 m=38 w=5.00 
+ l=0.18 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ perim=1.14
mI62 drn_lvc1 g_nclamp_lvc1 src_bdy_lvc1 src_bdy_lvc1 sky130_fd_pr__nfet_01v8 m=20 w=5.00 
+ l=0.18 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ perim=1.14
mncap src_bdy_lvc1 g_pdpre_lvc1 src_bdy_lvc1 src_bdy_lvc1 sky130_fd_pr__nfet_01v8 m=15 w=7.00 
+ l=8.00 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ perim=1.14
mpre_n1 g_nclamp_lvc1 g_pdpre_lvc1 src_bdy_lvc1 src_bdy_lvc1 sky130_fd_pr__nfet_01v8 m=3 w=7.00 
+ l=0.18 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ perim=1.14
mI43 g_nclamp_lvc2 g_pdpre_lvc2 src_bdy_lvc2 src_bdy_lvc2 sky130_fd_pr__nfet_01v8 m=2 w=7.00 
+ l=0.18 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ perim=1.14
mI58 src_bdy_lvc2 g_pdpre_lvc2 src_bdy_lvc2 src_bdy_lvc2 sky130_fd_pr__nfet_01v8 m=6 w=5.00 
+ l=8.00 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ perim=1.14
mI60 src_bdy_lvc2 g_pdpre_lvc2 src_bdy_lvc2 src_bdy_lvc2 sky130_fd_pr__nfet_01v8 m=1 w=5.00 
+ l=4.00 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ perim=1.14
mI59 src_bdy_lvc2 g_pdpre_lvc2 src_bdy_lvc2 src_bdy_lvc2 sky130_fd_pr__nfet_01v8 m=10 w=7.00 
+ l=8.00 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ perim=1.14
rrc_res g_pdpre_lvc1 drn_lvc1 sky130_fd_pr__res_generic_po m=1 w=0.33 l=1950
rI44 drn_lvc2 net161 sky130_fd_pr__res_generic_po m=1 w=0.33 l=900
rI47 net161 net155 sky130_fd_pr__res_generic_po m=1 w=0.33 l=300
rI46 g_pdpre_lvc2 net157 sky130_fd_pr__res_generic_po m=1 w=0.33 l=200
rI45 net157 net155 sky130_fd_pr__res_generic_po m=1 w=0.33 l=720
.ENDS

.SUBCKT sky130_fd_io__top_ground_lvc_wpad amuxbus_a amuxbus_b bdy2_b2b drn_lvc1 
+ drn_lvc2 g_core g_pad ogc_lvc src_bdy_lvc1 src_bdy_lvc2 vccd vcchib vdda 
+ vddio vddio_q vssa vssd vssio vssio_q vswitch
*.PININFO amuxbus_a:B amuxbus_b:B bdy2_b2b:B drn_lvc1:B drn_lvc2:B g_core:B 
*.PININFO g_pad:B ogc_lvc:B src_bdy_lvc1:B src_bdy_lvc2:B vccd:B vcchib:B 
*.PININFO vdda:B vddio:B vddio_q:B vssa:B vssd:B vssio:B vssio_q:B vswitch:B
Xesd bdy2_b2b src_bdy_lvc1 vssd / s8_esd_gnd2gnd_120x2_lv_isosub
xI54 src_bdy_lvc2 vddio condiode
xI50 src_bdy_lvc1 vddio condiode
rI21 g_pad g_core short
mpre_p1 g_nclamp_lvc1 g_pdpre_lvc1 drn_lvc1 drn_lvc1 sky130_fd_pr__pfet_01v8 m=20 w=7.00 l=0.18 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI40 g_nclamp_lvc2 g_pdpre_lvc2 drn_lvc2 drn_lvc2 sky130_fd_pr__pfet_01v8 m=20 w=7.00 l=0.18 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mclamp_xtor drn_lvc1 g_nclamp_lvc1 src_bdy_lvc1 src_bdy_lvc1 sky130_fd_pr__nfet_01v8 m=166 
+ w=7.00 l=0.18 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ perim=1.14
mI42 drn_lvc2 g_nclamp_lvc2 src_bdy_lvc2 src_bdy_lvc2 sky130_fd_pr__nfet_01v8 m=152 w=7.00 
+ l=0.18 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ perim=1.14
mI61 drn_lvc2 g_nclamp_lvc2 src_bdy_lvc2 src_bdy_lvc2 sky130_fd_pr__nfet_01v8 m=38 w=5.00 
+ l=0.18 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ perim=1.14
mI62 drn_lvc1 g_nclamp_lvc1 src_bdy_lvc1 src_bdy_lvc1 sky130_fd_pr__nfet_01v8 m=20 w=5.00 
+ l=0.18 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ perim=1.14
mncap src_bdy_lvc1 g_pdpre_lvc1 src_bdy_lvc1 src_bdy_lvc1 sky130_fd_pr__nfet_01v8 m=15 w=7.00 
+ l=8.00 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ perim=1.14
mpre_n1 g_nclamp_lvc1 g_pdpre_lvc1 src_bdy_lvc1 src_bdy_lvc1 sky130_fd_pr__nfet_01v8 m=3 w=7.00 
+ l=0.18 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ perim=1.14
mI43 g_nclamp_lvc2 g_pdpre_lvc2 src_bdy_lvc2 src_bdy_lvc2 sky130_fd_pr__nfet_01v8 m=2 w=7.00 
+ l=0.18 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ perim=1.14
mI58 src_bdy_lvc2 g_pdpre_lvc2 src_bdy_lvc2 src_bdy_lvc2 sky130_fd_pr__nfet_01v8 m=6 w=5.00 
+ l=8.00 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ perim=1.14
mI60 src_bdy_lvc2 g_pdpre_lvc2 src_bdy_lvc2 src_bdy_lvc2 sky130_fd_pr__nfet_01v8 m=1 w=5.00 
+ l=4.00 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ perim=1.14
mI59 src_bdy_lvc2 g_pdpre_lvc2 src_bdy_lvc2 src_bdy_lvc2 sky130_fd_pr__nfet_01v8 m=10 w=7.00 
+ l=8.00 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ perim=1.14
rrc_res g_pdpre_lvc1 drn_lvc1 sky130_fd_pr__res_generic_po m=1 w=0.33 l=1950
rI44 drn_lvc2 net161 sky130_fd_pr__res_generic_po m=1 w=0.33 l=900
rI47 net161 net155 sky130_fd_pr__res_generic_po m=1 w=0.33 l=300
rI46 g_pdpre_lvc2 net157 sky130_fd_pr__res_generic_po m=1 w=0.33 l=200
rI45 net157 net155 sky130_fd_pr__res_generic_po m=1 w=0.33 l=720
.ENDS

.SUBCKT sky130_fd_io__top_ground_hvc_wpad amuxbus_a amuxbus_b drn_hvc g_core g_pad 
+ ogc_hvc src_bdy_hvc vccd vcchib vdda vddio vddio_q vssa vssd vssio vssio_q 
+ vswitch
*.PININFO amuxbus_a:B amuxbus_b:B drn_hvc:B g_core:B g_pad:B ogc_hvc:B 
*.PININFO src_bdy_hvc:B vccd:B vcchib:B vdda:B vddio:B vddio_q:B vssa:B vssd:B 
*.PININFO vssio:B vssio_q:B vswitch:B
mcxtor2 drn_hvc g_nclamp src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=22 w=10.0 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mnc2 src_bdy_hvc g_pdpre src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=5 w=5.00 l=4.00 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mnc1 src_bdy_hvc g_pdpre src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=15 w=5.00 l=8.00 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mpre_n1 g_nclamp g_pdpre src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=15 w=7.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mclamp_xtor drn_hvc g_nclamp src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=120 w=20.0 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
rrc_res g_pdpre net94 sky130_fd_pr__res_generic_po m=1 w=0.33 l=470
rI38 net90 drn_hvc sky130_fd_pr__res_generic_po m=1 w=0.33 l=700
rI37 net94 net90 sky130_fd_pr__res_generic_po m=1 w=0.33 l=1550
mpre_p1 g_nclamp g_pdpre drn_hvc drn_hvc sky130_fd_pr__pfet_g5v0d10v5 m=50 w=7.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
xI39 src_bdy_hvc vddio condiode
rI13 g_pad g_core short
.ENDS
.SUBCKT sky130_fd_io__top_hvclamp_wopadv2 drn_hvc ogc_hvc src_bdy_hvc vssd
*.PININFO drn_hvc:B ogc_hvc:B src_bdy_hvc:B vssd:B
xI39 src_bdy_hvc ogc_hvc condiode
mpre_p1 g_nclamp g_pdpre drn_hvc drn_hvc sky130_fd_pr__pfet_g5v0d10v5 m=50 w=7.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
rrc_res g_pdpre net41 sky130_fd_pr__res_generic_po m=1 w=0.33 l=470
rI38 net37 drn_hvc sky130_fd_pr__res_generic_po m=1 w=0.33 l=700
rI37 net41 net37 sky130_fd_pr__res_generic_po m=1 w=0.33 l=1550
mclamp_xtor drn_hvc g_nclamp src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=120 w=20.0 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mpre_n1 g_nclamp g_pdpre src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=15 w=7.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mnc1 src_bdy_hvc g_pdpre src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=15 w=5.00 l=8.00 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mnc2 src_bdy_hvc g_pdpre src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=5 w=5.00 l=4.00 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mcxtor2 drn_hvc g_nclamp src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=22 w=10.0 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__top_power_hvc_wpadv2 amuxbus_a amuxbus_b drn_hvc ogc_hvc 
+ p_core p_pad src_bdy_hvc vccd vcchib vdda vddio vddio_q vssa vssd vssio 
+ vssio_q vswitch
*.PININFO amuxbus_a:B amuxbus_b:B drn_hvc:B ogc_hvc:B p_core:B p_pad:B 
*.PININFO src_bdy_hvc:B vccd:B vcchib:B vdda:B vddio:B vddio_q:B vssa:B vssd:B 
*.PININFO vssio:B vssio_q:B vswitch:B
xI39 src_bdy_hvc vddio condiode
mpre_p1 g_nclamp g_pdpre drn_hvc drn_hvc sky130_fd_pr__pfet_g5v0d10v5 m=50 w=7.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
rrc_res g_pdpre net67 sky130_fd_pr__res_generic_po m=1 w=0.33 l=470
rI38 net63 drn_hvc sky130_fd_pr__res_generic_po m=1 w=0.33 l=700
rI37 net67 net63 sky130_fd_pr__res_generic_po m=1 w=0.33 l=1550
mclamp_xtor drn_hvc g_nclamp src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=120 w=20.0 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mpre_n1 g_nclamp g_pdpre src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=15 w=7.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mnc1 src_bdy_hvc g_pdpre src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=15 w=5.00 l=8.00 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mnc2 src_bdy_hvc g_pdpre src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=5 w=5.00 l=4.00 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mcxtor2 drn_hvc g_nclamp src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=22 w=10.0 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
rI13 p_pad p_core short
.ENDS
.SUBCKT sky130_fd_io__top_vrefcapv2 amuxbus_a amuxbus_b cneg cpos vccd vcchib vdda 
+ vddio vddio_q vssa vssd vssio vssio_q vswitch
*.PININFO amuxbus_a:B amuxbus_b:B cneg:B cpos:B vccd:B vcchib:B vdda:B vddio:B 
*.PININFO vddio_q:B vssa:B vssd:B vssio:B vssio_q:B vswitch:B
xI271 cneg vddio_q condiode
mI334 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt m=180 w=10.0 l=0.90 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__xres4v2_in_buf enable_hv enable_vddio_lv in_h in_h_n pad 
+ vcchib vddio vgnd vnormal vnormal_b
*.PININFO enable_hv:I enable_vddio_lv:I pad:I vcchib:I vddio:I vgnd:I 
*.PININFO vnormal:I vnormal_b:I in_h:O in_h_n:O
XICEnet152 net152 / icecap
XICEnet193 net193 / icecap
XICEenable_vddio_lv_n enable_vddio_lv_n / icecap
XICEnet110 net110 / icecap
XICEpad_inv pad_inv / icecap
XICEvnormal_b vnormal_b / icecap
XICEpad1 pad1 / icecap
XICEvcchib_int vcchib_int / icecap
XICEnet116 net116 / icecap
XICEnet124 net124 / icecap
XICEenable_vddio_lv enable_vddio_lv / icecap
XICEnet106 net106 / icecap
XICEmode_vcchib mode_vcchib / icecap
XICEnet235 net235 / icecap
XICEin_h in_h / icecap
XICEin_h_n in_h_n / icecap
XICEenable_hv_b enable_hv_b / icecap
XICEpad pad / icecap
XICEnet140 net140 / icecap
XICEnet112 net112 / icecap
XICEvcchib vcchib / icecap
XICEnet207 net207 / icecap
XICEnet206 net206 / icecap
XICEvnormal vnormal / icecap
XICEenable_hv enable_hv / icecap
XICEfbk fbk / icecap
XICEnet120 net120 / icecap
XICEnet108 net108 / icecap
XI165 enable_vddio_lv enable_vddio_lv_n vgnd vgnd vcchib vcchib / 
+ sky130_fd_io__inv_1
XI61 net106 mode_vcchib vgnd vddio / sky130_fd_io__hvsbt_inv_x1
XI35 vnormal_b enable_hv net106 vgnd vddio / sky130_fd_io__hvsbt_nand2
rI132 net207 net110 sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=1077.19
rI159 net235 net108 sky130_fd_pr__res_generic_po m=1 w=0.4 l=713.695
mI8 net193 pad1 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI86 pad1 pad_inv vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI85 pad_inv pad net140 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.80 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI114 net152 pad_inv net140 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.00 l=0.80 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI145 enable_hv_b enable_hv vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI251 in_h in_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI83 net140 pad vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.80 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI7 fbk pad_inv vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI213 in_h_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI152 vgnd vgnd vgnd vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI113 net124 pad net152 vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=1.00 l=0.90 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI154 net120 mode_vcchib net206 vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=1.00 l=0.90 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI151 net116 mode_vcchib vcchib_int vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI150 net112 pad_inv net140 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.80 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI116 pad1 pad_inv net235 vddio sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI143 net124 vnormal vddio vddio sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI156 net116 enable_vddio_lv_n vcchib vcchib sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI252 in_h in_h_n vddio vddio sky130_fd_pr__pfet_g5v0d10v5 m=3 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI107 net108 mode_vcchib vddio vddio sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI146 enable_hv_b enable_hv vddio vddio sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI88 pad_inv pad vcchib_int vcchib_int sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.80 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI89 pad_inv pad net207 vddio sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI90 pad1 pad_inv net206 net206 sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI133 net110 mode_vcchib vddio vddio sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI2 net193 fbk vddio vddio sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI219 fbk net193 vddio vddio sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI14 in_h_n fbk vddio vddio sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI158 net120 enable_vddio_lv_n vcchib vcchib sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI139 net207 vnormal_b net110 vddio sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI136 net112 vnormal_b vddio vddio sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI153 vcchib_int vcchib_int vcchib_int vcchib_int sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.80 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI160 net235 vnormal_b net108 vddio sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_buf_localesd in_h out_h out_vt vcc_io vgnd vtrip_sel_h
*.PININFO in_h:I vtrip_sel_h:I out_h:O out_vt:O vcc_io:B vgnd:B
XICEout_vt out_vt / icecap
XICEin_h in_h / icecap
XICEout_h out_h / icecap
XICEvtrip_sel_h vtrip_sel_h / icecap
mhv_passgate out_h vtrip_sel_h out_vt vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
Xesd_res in_h out_h / s8_esd_res250only_small
Xggnfet2 vgnd out_vt vgnd vcc_io vgnd / s8_esd_signal_5_sym_hv_local_5term
Xggnfet6 vgnd vcc_io vgnd vcc_io out_h / s8_esd_signal_5_sym_hv_local_5term
Xggnfet5 vgnd vcc_io vgnd vcc_io out_vt / s8_esd_signal_5_sym_hv_local_5term
Xggnfet1 vgnd out_h vgnd vcc_io vgnd / s8_esd_signal_5_sym_hv_local_5term
.ENDS
.SUBCKT sky130_fd_io__gpio_pddrvr_strong force_lo_h force_lovol_h pad pd_h<3> 
+ pd_h<2> tie_lo_esd vcc_io vgnd_io vssio_amx
*.PININFO force_lo_h:I force_lovol_h:I pd_h<3>:I pd_h<2>:I vcc_io:I vgnd_io:I 
*.PININFO vssio_amx:I pad:O tie_lo_esd:O
XI112 pd_h<2> net61 / sky130_fd_io__tk_em2s
XI113 pd_h<2> net59 / sky130_fd_io__tk_em2s
XI97 pd_h<3> net85 / sky130_fd_io__tk_em2s
XI108 tie_lo_esd net83 / sky130_fd_io__tk_em2s
XI109 tie_lo_esd net77 / sky130_fd_io__tk_em2s
XI102 pd_h<3> net73 / sky130_fd_io__tk_em2s
XI104 pd_h<3> net69 / sky130_fd_io__tk_em2s
XI96 pd_h<3> net67 / sky130_fd_io__tk_em2s
XI87 tie_lo_esd net59 / sky130_fd_io__tk_em2o
XI83 pd_h<3> net61 / sky130_fd_io__tk_em2o
XI99 tie_lo_esd net85 / sky130_fd_io__tk_em2o
XI82 tie_lo_esd net61 / sky130_fd_io__tk_em2o
XI98 pd_h<2> net85 / sky130_fd_io__tk_em2o
XI106 pd_h<2> net83 / sky130_fd_io__tk_em2o
XI107 pd_h<3> net83 / sky130_fd_io__tk_em2o
XI110 pd_h<3> net77 / sky130_fd_io__tk_em2o
XI111 pd_h<2> net77 / sky130_fd_io__tk_em2o
XI100 tie_lo_esd net73 / sky130_fd_io__tk_em2o
XI101 pd_h<2> net73 / sky130_fd_io__tk_em2o
XI103 tie_lo_esd net69 / sky130_fd_io__tk_em2o
XI105 pd_h<2> net69 / sky130_fd_io__tk_em2o
XI95 pd_h<2> net67 / sky130_fd_io__tk_em2o
XI94 tie_lo_esd net67 / sky130_fd_io__tk_em2o
XI88 pd_h<3> net59 / sky130_fd_io__tk_em2o
XI49 vgnd_io tie_lo_esd / sky130_fd_io__tk_tie_r_out_esd
Xn24<2> pad net85 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn24<1> pad net85 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn24<0> pad net85 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn23<2> pad net67 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn23<1> pad net67 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn23<0> pad net67 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn22<2> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn22<1> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn22<0> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn21<2> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn21<1> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn21<0> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn12 pad net61 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn32<2> pad net69 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn32<1> pad net69 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn32<0> pad net69 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn33<2> pad net83 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn33<1> pad net83 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn33<0> pad net83 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn34<3> pad net77 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn34<2> pad net77 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn34<1> pad net77 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn34<0> pad net77 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn11<2> pad pd_h<2> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn11<1> pad pd_h<2> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn11<0> pad pd_h<2> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn13 pad net59 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn31 pad net73 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
xI72 vgnd_io vcc_io condiode
.ENDS
.SUBCKT sky130_fd_io__xres_esd out_h out_vt pad vddio vssd vssio
*.PININFO out_h:B out_vt:B pad:B vddio:B vssd:B vssio:B
Xesd pad out_h out_vt vddio vssd vssd / sky130_fd_io__gpio_buf_localesd
Xpddrvr_strong tie_lo_esd tie_lo_esd pad tie_lo_esd tie_lo_esd tie_lo_esd 
+ vddio vssio vssio / sky130_fd_io__gpio_pddrvr_strong
Xpudrvr_strong pad tie_hi_esd tie_hi_esd tie_hi_esd vddio vssd / 
+ sky130_fd_io__gpio_pudrvr_strong
xI271 vssio vddio condiode
.ENDS
.SUBCKT sky130_fd_io__xres_wpu pad vddio vssd
*.PININFO pad:B vddio:B vssd:B
Xesdr pad net15 / s8_esd_res250only_small
X5kres vddio net15 vssd / sky130_fd_io__com_res_weak
.ENDS
.SUBCKT sky130_fd_io__com_xres_weak_pu ra rb vgnd_io
*.PININFO vgnd_io:I ra:B rb:B
XICEn<3> n<3> / icecap
XICEn<2> n<2> / icecap
XICErb rb / icecap
XICEn<0> n<0> / icecap
XICEn<4> n<4> / icecap
XICEra ra / icecap
XICEnet64 net64 / icecap
XICEn<1> n<1> / icecap
XICEn<5> n<5> / icecap
Xe9 n<0> n<1> / sky130_fd_io__tk_em1s
Xe11 n<2> n<3> / sky130_fd_io__tk_em1s
Xe10 n<1> n<2> / sky130_fd_io__tk_em1s
Xe12 n<3> rb / sky130_fd_io__tk_em1s
Xe13 n<4> n<0> / sky130_fd_io__tk_em1s
Xe14 n<5> n<4> / sky130_fd_io__tk_em1o
rI84 n<0> n<1> sky130_fd_pr__res_generic_po m=1 w=0.8 l=1.5
rI62 n<3> rb sky130_fd_pr__res_generic_po m=1 w=0.8 l=1.5
rI82 n<2> n<3> sky130_fd_pr__res_generic_po m=1 w=0.8 l=1.5
rI85 ra net64 sky130_fd_pr__res_generic_po m=1 w=0.8 l=50
rI83 n<1> n<2> sky130_fd_pr__res_generic_po m=1 w=0.8 l=1.5
rI116 net64 n<5> sky130_fd_pr__res_generic_po m=1 w=0.8 l=12
rI104 n<4> n<0> sky130_fd_pr__res_generic_po m=1 w=0.8 l=6
rI134 n<5> n<4> sky130_fd_pr__res_generic_po m=1 w=0.8 l=6
.ENDS
.SUBCKT sky130_fd_io__xres_tk_emlo a b
*.PININFO a:B b:B
rI2 b net8 short
rI1 a net3 short
.ENDS
.SUBCKT sky130_fd_io__xres_tk_emlc a
*.PININFO a:B
rI2 a net7 short
rI1 a net2 short
.ENDS
.SUBCKT sky130_fd_io__xres_rcfilter_lpf_res_sub in out vgnd
*.PININFO in:I out:O vgnd:B
Xe1 in / sky130_fd_io__xres_tk_emlc
Xe2 out net30 / sky130_fd_io__xres_tk_emlo
rropti out net30 sky130_fd_pr__res_generic_nd m=1 w=0.5 l=14 isHV=FALSE
rr1 net30 in sky130_fd_pr__res_generic_nd m=1 w=0.5 l=47 isHV=FALSE
rropto in in sky130_fd_pr__res_generic_nd m=1 w=0.5 l=14 isHV=FALSE
.ENDS
.SUBCKT sky130_fd_io__xres_rcfilter_lpf_rcunit in out vgnd vnb vpwr
*.PININFO in:I out:O vgnd:B vnb:B vpwr:B
Xr1b net14 out vnb / sky130_fd_io__xres_rcfilter_lpf_res_sub
Xr1a in net14 vnb / sky130_fd_io__xres_rcfilter_lpf_res_sub
mI242 vgnd out vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=7.00 l=4.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI244 vpwr out vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=7.00 l=4.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__xres_rcfilter_lpf in out vcc_io vssd
*.PININFO in:I out:O vcc_io:B vssd:B
Xe5 net65 net40 / sky130_fd_io__xres_tk_emlo
Xe1 net135 net67 / sky130_fd_io__xres_tk_emlo
Xe4 net43 net65 / sky130_fd_io__xres_tk_emlo
XI200 net59 out / sky130_fd_io__xres_tk_emlo
XI199 net62 out / sky130_fd_io__xres_tk_emlo
XI198 vssd net59 / sky130_fd_io__xres_tk_emlo
XI197 vssd net57 / sky130_fd_io__xres_tk_emlo
XI194 net57 out / sky130_fd_io__xres_tk_emlo
XI193 net45 out / sky130_fd_io__xres_tk_emlo
XI191 net42 out / sky130_fd_io__xres_tk_emlo
XI190 net40 out / sky130_fd_io__xres_tk_emlo
XI187 vssd out / sky130_fd_io__xres_tk_emlo
XI186 vssd net45 / sky130_fd_io__xres_tk_emlo
Xe2 net67 net43 / sky130_fd_io__xres_tk_emlo
XI183 net42 vssd / sky130_fd_io__xres_tk_emlo
XI181 net40 vssd / sky130_fd_io__xres_tk_emlo
XI202 vssd / sky130_fd_io__xres_tk_emlc
XI201 vssd / sky130_fd_io__xres_tk_emlc
XI192 out / sky130_fd_io__xres_tk_emlc
XI189 vssd / sky130_fd_io__xres_tk_emlc
XI188 vssd / sky130_fd_io__xres_tk_emlc
XI180 net40 / sky130_fd_io__xres_tk_emlc
XI182 net42 / sky130_fd_io__xres_tk_emlc
Xe3 net43 / sky130_fd_io__xres_tk_emlc
XI172 in net135 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI184 vssd net57 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI185 vssd net45 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI196 vssd net62 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI195 vssd net59 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI179 net43 net65 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI178 net65 net40 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI177 net40 net42 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI176 net42 out vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI175 net67 net43 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI174 net43 net43 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI173 net135 net67 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
.ENDS
.SUBCKT sky130_fd_io__xres_inv_hys in_h out_h vcc_io vssd
*.PININFO in_h:I vcc_io:I vssd:I out_h:O
XICEpmid1 pmid1 / icecap
XICEout_h_n out_h_n / icecap
XICEout_h out_h / icecap
XICEin_h in_h / icecap
XICEnmid1 nmid1 / icecap
mI7 pmid1 in_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI8 out_h_n in_h pmid1 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI9 out_h out_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI10 pmid1 out_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI4 out_h_n in_h nmid1 vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=1.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI5 nmid1 in_h vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=1.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI6 out_h out_h_n vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
mI11 nmid1 out_h vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.00 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal perim=1.14
.ENDS
.SUBCKT sky130_fd_io__top_xres4v2 amuxbus_a amuxbus_b disable_pullup_h 
+ en_vddio_sig_h enable_h enable_vddio filt_in_h inp_sel_h pad pad_a_esd_h 
+ pullup_h tie_hi_esd tie_lo_esd tie_weak_hi_h vccd vcchib vdda vddio vddio_q 
+ vssa vssd vssio vssio_q vswitch xres_h_n
*.PININFO disable_pullup_h:I en_vddio_sig_h:I enable_h:I enable_vddio:I 
*.PININFO filt_in_h:I inp_sel_h:I vccd:I vcchib:I vdda:I vddio:I vddio_q:I 
*.PININFO vssa:I vssd:I vssio:I vssio_q:I vswitch:I tie_hi_esd:O tie_lo_esd:O 
*.PININFO xres_h_n:O amuxbus_a:B amuxbus_b:B pad:B pad_a_esd_h:B pullup_h:B 
*.PININFO tie_weak_hi_h:B
XI326 vssio tie_lo_esd / sky130_fd_io__tk_tie_r_out_esd
XI49 vddio tie_hi_esd / sky130_fd_io__tk_tie_r_out_esd
Xgpio_inbuf enable_h enable_vddio net79 net83 in_h vcchib vddio_q vssd 
+ en_vddio_sig_h en_vddio_sig_h_n / sky130_fd_io__xres4v2_in_buf
Xxresesd in_h net86 pad vddio vssd vssio / sky130_fd_io__xres_esd
Xweakpullup tie_weak_hi_h vddio vssd / sky130_fd_io__xres_wpu
Xesd_res pad pad_a_esd_h / s8_esd_res250only_small
XI335 net97 pullup_h vssd / sky130_fd_io__com_xres_weak_pu
XI363 inp_sel_h inp_sel_h_n vssd vddio_q / sky130_fd_io__hvsbt_inv_x2
XI334 net103 net107 vssd vddio / sky130_fd_io__hvsbt_inv_x2
XI333 disable_pullup_h net103 vssd vddio / sky130_fd_io__hvsbt_inv_x2
XI374 en_vddio_sig_h en_vddio_sig_h_n vssd vddio_q / sky130_fd_io__hvsbt_inv_x2
mI361 net124 inp_sel_h_n filt_in_h vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI358 net124 inp_sel_h net79 vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI332 net97 net107 vddio vddio sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI360 net124 inp_sel_h filt_in_h vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
mI357 net124 inp_sel_h_n net79 vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal perim=1.14
XI368 net124 out_rcfilt_h vddio_q vssd / sky130_fd_io__xres_rcfilter_lpf
XI367 out_rcfilt_h out_hysbuf_h vddio_q vssd / sky130_fd_io__xres_inv_hys
XI365 out_hysbuf_h out_h_n vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI364<1> out_h_n xres_h_n vssd vddio_q / sky130_fd_io__hvsbt_inv_x4
XI364<0> out_h_n xres_h_n vssd vddio_q / sky130_fd_io__hvsbt_inv_x4
.ENDS

* .SUBCKT condiode pin0 pin1
* .ENDS condiode
*********************************************************
* Copyright (c) 2017 by Cypress Semiconductor
* Cypress Confidential Information
*********************************************************

*.BIPOLAR
*.RESI=1
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.LDD
*.SCALE MICRON
*.MEGA
*.PARAM
*.OPTION SCALE=1E-6

************************************************************************
* auCdl Netlist:
*
* Library Name: s8iom0s8
* Top Cell Name: sky130_fd_io__top_gpiov2
* View Name: schematic
* Netlisted on: ... XX XX:XX:XX 2...
************************************************************************




************************************************************************
* Library Name: s8_esd
* Cell Name: s8_esd_res75only_small
* View Name: schematic
************************************************************************

.SUBCKT s8_esd_res75only_small pad rout
*.PININFO pad:B rout:B
RI175 pad rout sky130_fd_pr__res_generic_po l=3.15 m=1 w=2
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_amux_switch
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_amux_switch amuxbus_hv ng_amx_vpmp_h ng_pad_vpmp_h nmid_vccd pad_hv_n0
+ pad_hv_n1 pad_hv_n2 pad_hv_n3 pad_hv_p0 pad_hv_p1 pd_h_vdda pd_h_vddio pg_amx_vdda_h_n
+ pg_pad_vddioq_h_n vdda vddio vssa vssd
*.PININFO ng_amx_vpmp_h:I ng_pad_vpmp_h:I nmid_vccd:I pd_h_vdda:I pd_h_vddio:I
*.PININFO pg_amx_vdda_h_n:I pg_pad_vddioq_h_n:I vdda:I vddio:I vssa:I vssd:I
*.PININFO amuxbus_hv:B pad_hv_n0:B pad_hv_n1:B pad_hv_n2:B pad_hv_n3:B
*.PININFO pad_hv_p0:B pad_hv_p1:B
XI70 mid vdda condiode
XI71 mid1 vdda condiode
XI72 vssa vdda condiode
XI12 vssa net77 / s8_esd_res75only_small
XI56 vssa net79 / s8_esd_res75only_small
XMI45 mid1 ng_pad_vpmp_h pad_hv_n2 mid1 sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(7.00)*(0.50) l=0.50 m=4*1 p=2*(7.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=7.00
XMI24 pad_hv_n0 ng_pad_vpmp_h mid mid sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(7.00)*(0.50) l=0.50 m=3*1 p=2*(7.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=7.00
XMI35 mid ng_pad_vpmp_h pad_hv_n1 mid sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(7.00)*(0.50) l=0.50 m=4*1 p=2*(7.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=7.00
XMI46 pad_hv_n3 ng_pad_vpmp_h mid1 mid1 sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(7.00)*(0.50) l=0.50 m=4*1 p=2*(7.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=7.00
XMI1 mid nmid_vccd net77 vssa sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI77<1> mid pd_h_vddio vssa vssa sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(0.50) l=0.50 m=1*1 p=2*(0.42)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI77<0> mid1 pd_h_vddio vssa vssa sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(0.50) l=0.50 m=1*1 p=2*(0.42)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI78<1> mid pd_h_vdda vssa vssa sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(0.50) l=0.50 m=1*1 p=2*(0.42)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI78<0> mid1 pd_h_vdda vssa vssa sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(0.50) l=0.50 m=1*1 p=2*(0.42)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI47 mid1 ng_amx_vpmp_h amuxbus_hv mid1 sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(7.00)*(0.50) l=0.50 m=7*1 p=2*(7.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=7.00
XMI57 mid1 nmid_vccd net79 vssa sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI28 mid ng_amx_vpmp_h amuxbus_hv mid sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(7.00)*(0.50) l=0.50 m=7*1 p=2*(7.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=7.00
XMI26 mid pg_amx_vdda_h_n amuxbus_hv vdda sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(7.00)*(0.50) l=0.50 m=5*1 p=2*(7.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=7.00
XMI36 mid pg_pad_vddioq_h_n pad_hv_p0 vddio sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(7.00)*(0.50) l=0.50 m=3*1 p=2*(7.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=7.00
XMI22 mid pg_pad_vddioq_h_n pad_hv_p1 vddio sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(7.00)*(0.50) l=0.50 m=3*1 p=2*(7.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=7.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__hvsbt_inv_x1
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__hvsbt_inv_x1 in out vgnd vpwr
*.PININFO in:I vgnd:I vpwr:I out:O
XMI1 out in vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=2*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI2 out in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.70)*(0.60) l=0.60 m=1*1 p=2*(0.70)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.70
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_amx_pucsd_inv
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_amx_pucsd_inv A Y vda vssa
*.PININFO A:I vda:I vssa:I Y:O
XMI75 Y A vssa vssa sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(0.60) l=0.60 m=7*1 p=2*(0.42)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI74 Y A vda vda sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=7*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_amux_drvr_lshv2hv
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_amux_drvr_lshv2hv in in_b out_h_n rst_h rst_h_n vgnd vpwr_hv
*.PININFO in:I in_b:I rst_h:I rst_h_n:I vgnd:I vpwr_hv:I out_h_n:O
XMI1 fbk_n fbk vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(1.00) l=1.00 m=1*1 p=2*(0.42)+2*(1.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI2 fbk fbk_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(1.00) l=1.00 m=1*1 p=2*(0.42)+2*(1.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI14 out_h_n fbk vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=2*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI64 net52 rst_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI7 fbk in_b net52 vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=3*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI8 fbk_n in net52 vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=3*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMmnrst fbk rst_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=1*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI13 out_h_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=1*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_amx_inv4
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_amx_inv4 A Y vda vssa
*.PININFO A:I vda:I vssa:I Y:O
XMI75 Y A vssa vssa sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(0.60) l=0.60 m=2*1 p=2*(0.42)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI74 Y A vda vda sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=2*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__hvsbt_inv_x2
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__hvsbt_inv_x2 in out vgnd vpwr
*.PININFO in:I vgnd:I vpwr:I out:O
XMI2 out in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.70)*(0.60) l=0.60 m=2*1 p=2*(0.70)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.70
XMI1 out in vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=4*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_amx_pdcsd_inv
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_amx_pdcsd_inv A Y vda vssa
*.PININFO A:I vda:I vssa:I Y:O
XMI519 Y vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMI414 Y A vssa vssa sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMI429 Y A vda vda sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.75)*(2.00) l=2.00 m=1*1 p=2*(0.75)+2*(2.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.75
XMI517 Y A vda vda sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.75)*(2.00) l=2.00 m=1*1 p=2*(0.75)+2*(2.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.75
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__amx_inv1
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__amx_inv1 A Y vda vssa
*.PININFO A:I vda:I vssa:I Y:O
XMI92 Y A vssa vssa sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.75)*(0.50) l=0.50 m=1*1 p=2*(0.75)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.75
XMI54 Y A vda vda sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_amux_drvr_ls
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_amux_drvr_ls in in_b out_h out_h_n rst_h rst_h_n vgnd vpwr_hv
+ vpwr_lv
*.PININFO in:I in_b:I rst_h:I rst_h_n:I vgnd:I vpwr_hv:I vpwr_lv:I out_h:O
*.PININFO out_h_n:O
XMI9 out_h out_h_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.70)*(0.60) l=0.60 m=1*1 p=2*(0.70)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.70
XMI11 out_h_n out_h vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.70)*(0.60) l=0.60 m=1*1 p=2*(0.70)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.70
XMI20 net38 vpwr_lv net54 vgnd sky130_fd_pr__nfet_05v0_nvt AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.90) l=0.90 m=2*1 p=2*(1.00)+2*(0.90) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI21 net42 vpwr_lv net58 vgnd sky130_fd_pr__nfet_05v0_nvt AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.90) l=0.90 m=2*1 p=2*(1.00)+2*(0.90) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI24 out_h_n rst_h_n net42 vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=2*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMI25 out_h rst_h_n net38 vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=2*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMI12 net54 in_b vgnd vgnd sky130_fd_pr__nfet_01v8_lvt AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.15) l=0.15 m=2*1 p=2*(1.00)+2*(0.15) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI6 net58 in vgnd vgnd sky130_fd_pr__nfet_01v8_lvt AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.15) l=0.15 m=2*1 p=2*(1.00)+2*(0.15) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI17 out_h rst_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=2*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_amux_drvr
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_amux_drvr amux_en_vdda_h amux_en_vdda_h_n amux_en_vddio_h amux_en_vddio_h_n
+ amux_en_vswitch_h amux_en_vswitch_h_n amuxbusa_on amuxbusa_on_n amuxbusb_on amuxbusb_on_n
+ nga_amx_vswitch_h nga_pad_vswitch_h nga_pad_vswitch_h_n ngb_amx_vswitch_h ngb_pad_vswitch_h
+ ngb_pad_vswitch_h_n nmida_on_n nmida_vccd nmida_vccd_n nmidb_on_n nmidb_vccd nmidb_vccd_n
+ pd_csd_vswitch_h pd_csd_vswitch_h_n pd_on pd_on_n pga_amx_vdda_h_n pga_pad_vddioq_h_n
+ pgb_amx_vdda_h_n pgb_pad_vddioq_h_n pu_csd_vddioq_h_n pu_on pu_on_n vccd vdda vddio_q vssa vssd
+ vswitch
*.PININFO amux_en_vdda_h:I amux_en_vdda_h_n:I amux_en_vddio_h:I
*.PININFO amux_en_vddio_h_n:I amux_en_vswitch_h:I amux_en_vswitch_h_n:I
*.PININFO amuxbusa_on:I amuxbusa_on_n:I amuxbusb_on:I amuxbusb_on_n:I
*.PININFO nmida_on_n:I nmidb_on_n:I pd_on:I pd_on_n:I pu_on:I pu_on_n:I vccd:I
*.PININFO vdda:I vddio_q:I vssa:I vssd:I vswitch:I nga_amx_vswitch_h:O
*.PININFO nga_pad_vswitch_h:O nga_pad_vswitch_h_n:O ngb_amx_vswitch_h:O
*.PININFO ngb_pad_vswitch_h:O ngb_pad_vswitch_h_n:O nmida_vccd:O
*.PININFO nmida_vccd_n:O nmidb_vccd:O nmidb_vccd_n:O pd_csd_vswitch_h:O
*.PININFO pd_csd_vswitch_h_n:O pga_amx_vdda_h_n:O pga_pad_vddioq_h_n:O
*.PININFO pgb_amx_vdda_h_n:O pgb_pad_vddioq_h_n:O pu_csd_vddioq_h_n:O
XI105 nmidb_vccd nmidb_vccd_n vssd vccd / sky130_fd_io__hvsbt_inv_x1
XI93 nmida_vccd nmida_vccd_n vssd vccd / sky130_fd_io__hvsbt_inv_x1
XI38 net274 pu_csd_vddioq_h_n vddio_q vssd / sky130_fd_io__gpiov2_amx_pucsd_inv
XI103 net239 net245 pgb_amx_vdda_h_n amux_en_vdda_h_n amux_en_vdda_h vssa vdda /
+ sky130_fd_io__gpiov2_amux_drvr_lshv2hv
Xpga_amx_ls net265 net272 pga_amx_vdda_h_n amux_en_vdda_h_n amux_en_vdda_h vssa vdda /
+ sky130_fd_io__gpiov2_amux_drvr_lshv2hv
XI64 net236 ngb_pad_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_inv4
XI63 net236 ngb_amx_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_inv4
XI62 net239 pgb_pad_vddioq_h_n vddio_q vssd / sky130_fd_io__gpiov2_amx_inv4
XI47 net256 nga_pad_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_inv4
XI42 net265 pga_pad_vddioq_h_n vddio_q vssd / sky130_fd_io__gpiov2_amx_inv4
XI45 net256 nga_amx_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_inv4
XI89 nmida_on_n nmida_vccd vssd vccd / sky130_fd_io__hvsbt_inv_x2
XI53 nmidb_on_n nmidb_vccd vssd vccd / sky130_fd_io__hvsbt_inv_x2
Xpdcsd_inv net254 pd_csd_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_pdcsd_inv
XI90 pd_csd_vswitch_h pd_csd_vswitch_h_n vswitch vssa / sky130_fd_io__amx_inv1
XI85 ngb_pad_vswitch_h ngb_pad_vswitch_h_n vswitch vssa / sky130_fd_io__amx_inv1
XI87 nga_pad_vswitch_h nga_pad_vswitch_h_n vswitch vssa / sky130_fd_io__amx_inv1
XMI104 pd_csd_vswitch_h amux_en_vddio_h_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=1*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI78 nga_pad_vswitch_h amux_en_vddio_h_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=1*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI75 nga_amx_vswitch_h amux_en_vdda_h_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=1*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI77 ngb_pad_vswitch_h amux_en_vddio_h_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=1*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI76 ngb_amx_vswitch_h amux_en_vdda_h_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=1*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
Xngb_ls amuxbusb_on amuxbusb_on_n net230 net236 amux_en_vswitch_h_n amux_en_vswitch_h vssa vswitch
+ vccd / sky130_fd_io__gpiov2_amux_drvr_ls
Xpgb_pad_ls amuxbusb_on amuxbusb_on_n net239 net245 amux_en_vddio_h_n amux_en_vddio_h vssd vddio_q
+ vccd / sky130_fd_io__gpiov2_amux_drvr_ls
Xpd_csd_ls pd_on pd_on_n net248 net254 amux_en_vswitch_h_n amux_en_vswitch_h vssa vswitch vccd
+ / sky130_fd_io__gpiov2_amux_drvr_ls
Xnga_ls amuxbusa_on amuxbusa_on_n net257 net256 amux_en_vswitch_h_n amux_en_vswitch_h vssa vswitch
+ vccd / sky130_fd_io__gpiov2_amux_drvr_ls
Xpga_pad_ls amuxbusa_on amuxbusa_on_n net265 net272 amux_en_vddio_h_n amux_en_vddio_h vssd vddio_q
+ vccd / sky130_fd_io__gpiov2_amux_drvr_ls
Xpu_csd_ls pu_on pu_on_n net274 net275 amux_en_vddio_h_n amux_en_vddio_h vssd vddio_q vccd
+ / sky130_fd_io__gpiov2_amux_drvr_ls
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__nor2_1
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__nor2_1 A B Y vgnd vnb vpb vpwr
*.PININFO A:I B:I vgnd:I vnb:I vpb:I vpwr:I Y:O
XMMP1 sndPA B Y vpb sky130_fd_pr__pfet_01v8_hvt AD=0 AS=0 PD=0 PS=0
+ a=(1.12)*(0.15) l=0.15 m=1*1 p=2*(1.12)+2*(0.15) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.12
XMMP0 vpwr A sndPA vpb sky130_fd_pr__pfet_01v8_hvt AD=0 AS=0 PD=0 PS=0
+ a=(1.12)*(0.15) l=0.15 m=1*1 p=2*(1.12)+2*(0.15) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.12
XMMN1 Y B vgnd vnb sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(740e-3)*(150e-3) l=150e-3 m=1*1 p=2*(740e-3)+2*(150e-3) sa=265e-3
+ sb=265e-3 sd=280e-3 w=740e-3
XMMN0 Y A vgnd vnb sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(740e-3)*(150e-3) l=150e-3 m=1*1 p=2*(740e-3)+2*(150e-3) sa=265e-3
+ sb=265e-3 sd=280e-3 w=740e-3
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__nand2_1
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__nand2_1 A B Y vgnd vnb vpb vpwr
*.PININFO A:I B:I vgnd:I vnb:I vpb:I vpwr:I Y:O
XMMP1 Y B vpwr vpb sky130_fd_pr__pfet_01v8_hvt AD=0 AS=0 PD=0 PS=0
+ a=(1.12)*(0.15) l=0.15 m=1*1 p=2*(1.12)+2*(0.15) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.12
XMMP0 Y A vpwr vpb sky130_fd_pr__pfet_01v8_hvt AD=0 AS=0 PD=0 PS=0
+ a=(1.12)*(0.15) l=0.15 m=1*1 p=2*(1.12)+2*(0.15) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.12
XMMN1 sndA B vgnd vnb sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(0.74)*(0.15) l=0.15 m=1*1 p=2*(0.74)+2*(0.15) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.74
XMMN0 Y A sndA vnb sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(0.74)*(0.15) l=0.15 m=1*1 p=2*(0.74)+2*(0.15) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.74
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__hvsbt_nor
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__hvsbt_nor in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
XMI12 out in1 net16 vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=1*2 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI3 net16 in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=1*2 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI6 out in1 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.70)*(0.60) l=0.60 m=1*1 p=2*(0.70)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.70
XMI1 out in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.70)*(0.60) l=0.60 m=1*1 p=2*(0.70)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.70
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_amux_nand5
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_amux_nand5 in0 in1 in2 in3 in4 out vgnd vpwr
*.PININFO in0:I in1:I in2:I in3:I in4:I vgnd:I vpwr:I out:O
XMI21 out_n out vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=2*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI20 out out_n vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(0.50) l=0.50 m=1*1 p=2*(0.42)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI3 out in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=2*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI23 vgnd out_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(0.50) l=0.50 m=1*1 p=2*(0.42)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI22 out_n out vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(0.50) l=0.50 m=1*1 p=2*(0.42)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI14 net51 in2 net55 vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI15 net55 in3 net63 vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI6 net59 in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI18 net63 in4 net59 vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI1 out in1 net51 vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_amux_nand4
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_amux_nand4 in0 in1 in2 in3 out vgnd vpwr
*.PININFO in0:I in1:I in2:I in3:I vgnd:I vpwr:I out:O
XMI20 out out_n vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(0.50) l=0.50 m=1*1 p=2*(0.42)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI19 out_n out vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=2*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI3 out in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=2*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI21 vgnd out_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(0.50) l=0.50 m=1*1 p=2*(0.42)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI18 out_n out vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(0.50) l=0.50 m=1*1 p=2*(0.42)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI14 net50 in2 net54 vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI15 net54 in3 net58 vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI6 net58 in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI1 out in1 net50 vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__hvsbt_nand2
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__hvsbt_nand2 in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
XMI5 out in1 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=2*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI3 out in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=2*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI6 net25 in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.70)*(0.60) l=0.60 m=1*1 p=2*(0.70)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.70
XMI1 out in1 net25 vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.70)*(0.60) l=0.60 m=1*1 p=2*(0.70)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.70
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__xor2_1
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__xor2_1 A B X vgnd vpwr
*.PININFO A:I B:I vgnd:I vpwr:I X:O
XMMNaoi20 X inor vgnd vgnd sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(840e-3)*(150e-3) l=150e-3 m=1*1 p=2*(840e-3)+2*(150e-3) sa=265e-3
+ sb=265e-3 sd=280e-3 w=840e-3
XMMNaoi11 sndNA B X vgnd sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(840e-3)*(150e-3) l=150e-3 m=1*1 p=2*(840e-3)+2*(150e-3) sa=265e-3
+ sb=265e-3 sd=280e-3 w=840e-3
XMMNaoi10 vgnd A sndNA vgnd sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(840e-3)*(150e-3) l=150e-3 m=1*1 p=2*(840e-3)+2*(150e-3) sa=265e-3
+ sb=265e-3 sd=280e-3 w=840e-3
XMMNnor1 inor B vgnd vgnd sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(840e-3)*(150e-3) l=150e-3 m=1*1 p=2*(840e-3)+2*(150e-3) sa=265e-3
+ sb=265e-3 sd=280e-3 w=840e-3
XMMNnor0 inor A vgnd vgnd sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(840e-3)*(150e-3) l=150e-3 m=1*1 p=2*(840e-3)+2*(150e-3) sa=265e-3
+ sb=265e-3 sd=280e-3 w=840e-3
XMMPaoi20 X inor pmid vpwr sky130_fd_pr__pfet_01v8_hvt AD=0 AS=0 PD=0 PS=0
+ a=(1.26)*(150e-3) l=150e-3 m=1*1 p=2*(1.26)+2*(150e-3) sa=265e-3
+ sb=265e-3 sd=280e-3 w=1.26
XMMPaoi11 pmid B vpwr vpwr sky130_fd_pr__pfet_01v8_hvt AD=0 AS=0 PD=0 PS=0
+ a=(1.26)*(150e-3) l=150e-3 m=1*1 p=2*(1.26)+2*(150e-3) sa=265e-3
+ sb=265e-3 sd=280e-3 w=1.26
XMMPaoi10 pmid A vpwr vpwr sky130_fd_pr__pfet_01v8_hvt AD=0 AS=0 PD=0 PS=0
+ a=(1.26)*(150e-3) l=150e-3 m=1*1 p=2*(1.26)+2*(150e-3) sa=265e-3
+ sb=265e-3 sd=280e-3 w=1.26
XMMPnor1 sndPA B inor vpwr sky130_fd_pr__pfet_01v8_hvt AD=0 AS=0 PD=0 PS=0
+ a=(1.26)*(150e-3) l=150e-3 m=1*1 p=2*(1.26)+2*(150e-3) sa=265e-3
+ sb=265e-3 sd=280e-3 w=1.26
XMMPnor0 vpwr A sndPA vpwr sky130_fd_pr__pfet_01v8_hvt AD=0 AS=0 PD=0 PS=0
+ a=(1.26)*(150e-3) l=150e-3 m=1*1 p=2*(1.26)+2*(150e-3) sa=265e-3
+ sb=265e-3 sd=280e-3 w=1.26
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__inv_1
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__inv_1 A Y vgnd vnb vpb vpwr
*.PININFO A:I vgnd:I vnb:I vpb:I vpwr:I Y:O
XMMIN1 Y A vgnd vnb sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(0.74)*(0.15) l=0.15 m=1*1 p=2*(0.74)+2*(0.15) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.74
XMMIP1 Y A vpwr vpb sky130_fd_pr__pfet_01v8_hvt AD=0 AS=0 PD=0 PS=0
+ a=(1.12)*(0.15) l=0.15 m=1*1 p=2*(1.12)+2*(0.15) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.12
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_amux_decoder
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_amux_decoder amuxbusa_on amuxbusa_on_n amuxbusb_on amuxbusb_on_n analog_en
+ analog_pol analog_sel nga_pad_vswitch_h nga_pad_vswitch_h_n ngb_pad_vswitch_h ngb_pad_vswitch_h_n
+ nmida_on_n nmida_vccd_n nmidb_on_n nmidb_vccd_n out pd_on pd_on_n pd_vswitch_h_n pga_amx_vdda_h_n
+ pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n pu_on pu_on_n pu_vddioq_h_n vccd vssd
*.PININFO analog_en:I analog_pol:I analog_sel:I nga_pad_vswitch_h:I
*.PININFO nga_pad_vswitch_h_n:I ngb_pad_vswitch_h:I ngb_pad_vswitch_h_n:I
*.PININFO nmida_vccd_n:I nmidb_vccd_n:I out:I pd_vswitch_h_n:I
*.PININFO pga_amx_vdda_h_n:I pga_pad_vddioq_h_n:I pgb_amx_vdda_h_n:I
*.PININFO pgb_pad_vddioq_h_n:I pu_vddioq_h_n:I vccd:I vssd:I amuxbusa_on:O
*.PININFO amuxbusa_on_n:O amuxbusb_on:O amuxbusb_on_n:O nmida_on_n:O
*.PININFO nmidb_on_n:O pd_on:O pd_on_n:O pu_on:O pu_on_n:O
XI114 ana_en_i_n net137 int_amuxb_on vssd vssd vccd vccd / sky130_fd_io__nor2_1
XI115 ana_en_i_n int_pu_on_n int_pu_on vssd vssd vccd vccd / sky130_fd_io__nor2_1
XI113 ana_en_i_n net144 int_amuxa_on vssd vssd vccd vccd / sky130_fd_io__nor2_1
XI116 ana_en_i_n int_pd_on_n int_pd_on vssd vssd vccd vccd / sky130_fd_io__nor2_1
XI110 pol_xor_out ana_sel_i net137 vssd vssd vccd vccd / sky130_fd_io__nand2_1
XI109 ana_sel_i_n pol_xor_out net144 vssd vssd vccd vccd / sky130_fd_io__nand2_1
XI112 ana_pol_i_n out_i_n int_pd_on_n vssd vssd vccd vccd / sky130_fd_io__nand2_1
XI111 ana_pol_i out_i int_pu_on_n vssd vssd vccd vccd / sky130_fd_io__nand2_1
XI102 nga_pad_vswitch_h net222 net167 vssd vccd / sky130_fd_io__hvsbt_nor
XI106 ngb_pad_vswitch_h net212 net172 vssd vccd / sky130_fd_io__hvsbt_nor
XI80 int_pd_on pga_pad_vddioq_h_n pgb_pad_vddioq_h_n nga_pad_vswitch_h_n ngb_pad_vswitch_h_n
+ int_fbk_pdon_n vssd vccd / sky130_fd_io__gpiov2_amux_nand5
XI79 int_pu_on pga_pad_vddioq_h_n pgb_pad_vddioq_h_n nga_pad_vswitch_h_n ngb_pad_vswitch_h_n
+ int_fbk_puon_n vssd vccd / sky130_fd_io__gpiov2_amux_nand5
XI77 int_amuxa_on pu_vddioq_h_n pd_vswitch_h_n nmida_vccd_n amuxbusa_on_n vssd vccd /
+ sky130_fd_io__gpiov2_amux_nand4
XI78 int_amuxb_on pu_vddioq_h_n pd_vswitch_h_n nmidb_vccd_n amuxbusb_on_n vssd vccd /
+ sky130_fd_io__gpiov2_amux_nand4
XI120 int_amux_a_on_n net167 nmida_on_n vssd vccd / sky130_fd_io__hvsbt_nand2
XI105 pgb_pad_vddioq_h_n pgb_amx_vdda_h_n net212 vssd vccd / sky130_fd_io__hvsbt_nand2
XI121 int_amux_b_on_n net172 nmidb_on_n vssd vccd / sky130_fd_io__hvsbt_nand2
XI101 pga_pad_vddioq_h_n pga_amx_vdda_h_n net222 vssd vccd / sky130_fd_io__hvsbt_nand2
XI45 ana_pol_i out_i pol_xor_out vssd vccd / sky130_fd_io__xor2_1
XI95 pd_on pd_on_n vssd vssd vccd vccd / sky130_fd_io__inv_1
XI93 pu_on pu_on_n vssd vssd vccd vccd / sky130_fd_io__inv_1
XI91 int_amuxb_on int_amux_b_on_n vssd vssd vccd vccd / sky130_fd_io__inv_1
XI44 out_i_n out_i vssd vssd vccd vccd / sky130_fd_io__inv_1
XI43 out out_i_n vssd vssd vccd vccd / sky130_fd_io__inv_1
XI75 int_fbk_puon_n pu_on vssd vssd vccd vccd / sky130_fd_io__inv_1
XI58 analog_en ana_en_i_n vssd vssd vccd vccd / sky130_fd_io__inv_1
XI76 int_fbk_pdon_n pd_on vssd vssd vccd vccd / sky130_fd_io__inv_1
XI73 amuxbusa_on_n amuxbusa_on vssd vssd vccd vccd / sky130_fd_io__inv_1
XI74 amuxbusb_on_n amuxbusb_on vssd vssd vccd vccd / sky130_fd_io__inv_1
XI35 analog_pol ana_pol_i_n vssd vssd vccd vccd / sky130_fd_io__inv_1
XI40 ana_sel_i_n ana_sel_i vssd vssd vccd vccd / sky130_fd_io__inv_1
XI39 analog_sel ana_sel_i_n vssd vssd vccd vccd / sky130_fd_io__inv_1
XI89 int_amuxa_on int_amux_a_on_n vssd vssd vccd vccd / sky130_fd_io__inv_1
XI41 ana_pol_i_n ana_pol_i vssd vssd vccd vccd / sky130_fd_io__inv_1
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_amux_ls_inv_x1
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_amux_ls_inv_x1 in out vgnd vpwr
*.PININFO in:I vgnd:I vpwr:I out:O
XMI2 out in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=1*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI1 out in vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=2*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_amux_ctl_lshv2hv
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_amux_ctl_lshv2hv in in_b out_h out_h_n rst_h rst_h_n vgnd vpwr_hv
*.PININFO in:I in_b:I rst_h:I rst_h_n:I vgnd:I vpwr_hv:I out_h:O out_h_n:O
XMI1 fbk_n fbk vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(1.00) l=1.00 m=1*1 p=2*(0.42)+2*(1.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI2 fbk fbk_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(1.00) l=1.00 m=1*1 p=2*(0.42)+2*(1.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI11 out_h fbk_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMI14 out_h_n fbk vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMI64 net64 rst_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI7 fbk in_b net64 vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=3*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI8 fbk_n in net64 vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=3*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMmnrst fbk rst_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=1*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI12 out_h fbk_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=1*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI13 out_h_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=1*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_amux_ctl_inv_1
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_amux_ctl_inv_1 in out vgnd vpwr
*.PININFO in:I vgnd:I vpwr:I out:O
XMI27 out in vgnd vgnd sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(0.74)*(0.15) l=0.15 m=1*1 p=2*(0.74)+2*(0.15) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.74
XMI29 out in vpwr vpwr sky130_fd_pr__pfet_01v8_hvt AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.25) l=0.25 m=1*1 p=2*(1.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_amux_ctl_ls
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_amux_ctl_ls in in_b out_h out_h_n rst_h rst_h_n vgnd vpwr_hv
+ vpwr_lv
*.PININFO in:I in_b:I rst_h:I rst_h_n:I vgnd:I vpwr_hv:I vpwr_lv:I out_h:O
*.PININFO out_h_n:O
XMI1 fbk fbk_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.75)*(0.50) l=0.50 m=1*1 p=2*(0.75)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.75
XMI2 fbk_n fbk vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.75)*(0.50) l=0.50 m=1*1 p=2*(0.75)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.75
XMI11 out_h_n fbk vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMI14 out_h fbk_n vpwr_hv vpwr_hv sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMI5 net61 rst_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=4*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI7 net62 in_b net61 vgnd sky130_fd_pr__nfet_01v8_lvt AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.15) l=0.15 m=4*1 p=2*(1.00)+2*(0.15) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI8 net66 in net61 vgnd sky130_fd_pr__nfet_01v8_lvt AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.15) l=0.15 m=4*1 p=2*(1.00)+2*(0.15) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI59 fbk_n vpwr_lv net66 vgnd sky130_fd_pr__nfet_05v0_nvt AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.90) l=0.90 m=4*1 p=2*(1.00)+2*(0.90) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMmnrst fbk rst_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=1*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI58 fbk vpwr_lv net62 vgnd sky130_fd_pr__nfet_05v0_nvt AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.90) l=0.90 m=4*1 p=2*(1.00)+2*(0.90) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI12 out_h_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=1*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI13 out_h fbk_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=1*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_amux_ls
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_amux_ls amux_en_vdda_h amux_en_vdda_h_n amux_en_vddio_h amux_en_vddio_h_n
+ amux_en_vswitch_h amux_en_vswitch_h_n analog_en enable_vdda_h enable_vdda_h_n enable_vswitch_h
+ hld_i_h hld_i_h_n vccd vdda vddio_q vssa vssd vswitch
*.PININFO analog_en:I enable_vdda_h:I enable_vswitch_h:I hld_i_h:I hld_i_h_n:I
*.PININFO vccd:I vdda:I vddio_q:I vssa:I vssd:I vswitch:I amux_en_vdda_h:O
*.PININFO amux_en_vdda_h_n:O amux_en_vddio_h:O amux_en_vddio_h_n:O
*.PININFO amux_en_vswitch_h:O amux_en_vswitch_h_n:O enable_vdda_h_n:O
XI32 enable_vdda_h enable_vdda_h_n vssa vdda / sky130_fd_io__gpiov2_amux_ls_inv_x1
Xpd_vdda_ls amux_en_vddio_h amux_en_vddio_h_n amux_en_vdda_h amux_en_vdda_h_n enable_vdda_h_n
+ enable_vdda_h vssa vdda / sky130_fd_io__gpiov2_amux_ctl_lshv2hv
Xpd_vswitch_ls amux_en_vddio_h amux_en_vddio_h_n amux_en_vswitch_h amux_en_vswitch_h_n net74
+ enable_vswitch_h vssa vswitch / sky130_fd_io__gpiov2_amux_ctl_lshv2hv
XI16 ana_en_i_n ana_en_i vssd vccd / sky130_fd_io__gpiov2_amux_ctl_inv_1
XI15 analog_en ana_en_i_n vssd vccd / sky130_fd_io__gpiov2_amux_ctl_inv_1
XI18 enable_vswitch_h net74 vssa vswitch / sky130_fd_io__hvsbt_inv_x1
Xpd_vddio_ls ana_en_i ana_en_i_n amux_en_vddio_h amux_en_vddio_h_n hld_i_h hld_i_h_n vssd vddio_q
+ vccd / sky130_fd_io__gpiov2_amux_ctl_ls
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_amux_ctl_logic
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_amux_ctl_logic analog_en analog_pol analog_sel enable_vdda_h enable_vdda_h_n
+ enable_vswitch_h hld_i_h hld_i_h_n nga_amx_vswitch_h nga_pad_vswitch_h ngb_amx_vswitch_h
+ ngb_pad_vswitch_h nmida_vccd nmidb_vccd out pd_csd_vswitch_h pga_amx_vdda_h_n pga_pad_vddioq_h_n
+ pgb_amx_vdda_h_n pgb_pad_vddioq_h_n pu_csd_vddioq_h_n vccd vdda vddio_q vssa vssd vswitch
*.PININFO analog_en:I analog_pol:I analog_sel:I enable_vdda_h:I
*.PININFO enable_vswitch_h:I hld_i_h:I hld_i_h_n:I out:I vccd:I vdda:I
*.PININFO vddio_q:I vssa:I vssd:I vswitch:I enable_vdda_h_n:O
*.PININFO nga_amx_vswitch_h:O nga_pad_vswitch_h:O ngb_amx_vswitch_h:O
*.PININFO ngb_pad_vswitch_h:O nmida_vccd:O nmidb_vccd:O pd_csd_vswitch_h:O
*.PININFO pga_amx_vdda_h_n:O pga_pad_vddioq_h_n:O pgb_amx_vdda_h_n:O
*.PININFO pgb_pad_vddioq_h_n:O pu_csd_vddioq_h_n:O
Xamux_sw_drvr amux_en_vdda_h amux_en_vdda_h_n amux_en_vddio_h amux_en_vddio_h_n amux_en_vswitch_h
+ amux_en_vswitch_h_n amuxbusa_on amuxbusa_on_n amuxbusb_on amuxbusb_on_n nga_amx_vswitch_h
+ nga_pad_vswitch_h nga_pad_vswitch_h_n ngb_amx_vswitch_h ngb_pad_vswitch_h ngb_pad_vswitch_h_n
+ nmida_on_n nmida_vccd nmida_vccd_n nmidb_on_n nmidb_vccd nmidb_vccd_n pd_csd_vswitch_h
+ pd_csd_vswitch_h_n pd_on pd_on_n pga_amx_vdda_h_n pga_pad_vddioq_h_n pgb_amx_vdda_h_n
+ pgb_pad_vddioq_h_n pu_csd_vddioq_h_n pu_on pu_on_n vccd vdda vddio_q vssa vssd vswitch /
+ sky130_fd_io__gpiov2_amux_drvr
Xamux_lv_decoder amuxbusa_on amuxbusa_on_n amuxbusb_on amuxbusb_on_n analog_en analog_pol analog_sel
+ nga_pad_vswitch_h nga_pad_vswitch_h_n ngb_pad_vswitch_h ngb_pad_vswitch_h_n nmida_on_n
+ nmida_vccd_n nmidb_on_n nmidb_vccd_n out pd_on pd_on_n pd_csd_vswitch_h_n pga_amx_vdda_h_n
+ pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n pu_on pu_on_n pu_csd_vddioq_h_n vccd vssd
+ / sky130_fd_io__gpiov2_amux_decoder
Xamux_ls amux_en_vdda_h amux_en_vdda_h_n amux_en_vddio_h amux_en_vddio_h_n amux_en_vswitch_h
+ amux_en_vswitch_h_n analog_en enable_vdda_h enable_vdda_h_n enable_vswitch_h hld_i_h hld_i_h_n
+ vccd vdda vddio_q vssa vssd vswitch / sky130_fd_io__gpiov2_amux_ls
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_amux
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_amux amuxbus_a amuxbus_b analog_en analog_pol analog_sel enable_vdda_h
+ enable_vswitch_h hld_i_h hld_i_h_n out pad vccd vdda vddio_q vssa vssd vssio_q
+ vswitch
*.PININFO analog_en:I analog_pol:I analog_sel:I enable_vdda_h:I
*.PININFO enable_vswitch_h:I hld_i_h:I hld_i_h_n:I out:I vccd:I vdda:I
*.PININFO vddio_q:I vssa:I vssd:I vssio_q:I vswitch:I amuxbus_a:B amuxbus_b:B
*.PININFO pad:B
XI78 vssa vswitch condiode
XI43 vssio_q vdda condiode
XMMP_PU net85 pu_csd_vddioq_h_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(15.0)*(0.50) l=0.50 m=4*1 p=2*(15.0)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=15.0
XMI52 net81 pu_csd_vddioq_h_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(15.0)*(0.50) l=0.50 m=3*1 p=2*(15.0)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=15.0
XMI49 net81 pd_csd_vswitch_h vssio_q vssio_q sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=6*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMMN_PD net85 pd_csd_vswitch_h vssio_q vssio_q sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=8*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
Xmux_b amuxbus_b ngb_amx_vpmp_h ngb_pad_vpmp_h nmidb_vccd net101 net101 net97 net97 net100
+ net99 net0127 hld_i_h pgb_amx_vdda_h_n pgb_pad_vddioq_h_n vdda vddio_q vssa vssd /
+ sky130_fd_io__gpiov2_amux_switch
Xmux_a amuxbus_a nga_amx_vpmp_h nga_pad_vpmp_h nmida_vccd net101 net101 net97 net97 net100
+ net99 net0127 hld_i_h pga_amx_vdda_h_n pga_pad_vddioq_h_n vdda vddio_q vssa vssd /
+ sky130_fd_io__gpiov2_amux_switch
XBBM_logic analog_en analog_pol analog_sel enable_vdda_h net0127 enable_vswitch_h hld_i_h hld_i_h_n
+ nga_amx_vpmp_h nga_pad_vpmp_h ngb_amx_vpmp_h ngb_pad_vpmp_h nmida_vccd nmidb_vccd out
+ pd_csd_vswitch_h pga_amx_vdda_h_n pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n
+ pu_csd_vddioq_h_n vccd vdda vddio_q vssa vssd vswitch / sky130_fd_io__gpiov2_amux_ctl_logic
XI40 pad net85 / s8_esd_res75only_small
XI39 pad net81 / s8_esd_res75only_small
XI53 pad pad / s8_esd_res75only_small
XI54 pad net166 / s8_esd_res75only_small
XI55 pad pad / s8_esd_res75only_small
XI27 pad net100 / s8_esd_res75only_small
XI57 pad net168 / s8_esd_res75only_small
XI28 net166 net101 / s8_esd_res75only_small
XI58 net168 net97 / s8_esd_res75only_small
XI26 pad net99 / s8_esd_res75only_small
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__tk_em2s
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__tk_em2s a b
*.PININFO a:B b:B
RI2 b net8 short m=1
RI1 a net8 short m=1
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__tk_em2o
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__tk_em2o a b
*.PININFO a:B b:B
RI2 b net7 short m=1
RI1 a net11 short m=1
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__tk_tie_r_out_esd
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__tk_tie_r_out_esd a b
*.PININFO a:B b:B
Resd_r a b sky130_fd_pr__res_generic_po l=10.2 m=1 w=0.5
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__com_pddrvr_unit_2_5
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__com_pddrvr_unit_2_5 nd ngin ns
*.PININFO ngin:I nd:B ns:B
XMndrv nd ngin ns ns sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.60) l=0.60 m=2*1 p=2*(5.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_pddrvr_strong
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_pddrvr_strong pad pd_h<3> pd_h<2> pd_h_i2c tie_lo_esd vcc_io vgnd_io
*.PININFO pd_h<3>:I pd_h<2>:I pd_h_i2c:I vcc_io:I vgnd_io:I pad:O tie_lo_esd:O
XI113 pd_h<2> net46 / sky130_fd_io__tk_em2s
XI96 pd_h<3> net66 / sky130_fd_io__tk_em2s
XI104 pd_h<3> net68 / sky130_fd_io__tk_em2s
XI102 pd_h<3> net72 / sky130_fd_io__tk_em2s
XI109 tie_lo_esd net76 / sky130_fd_io__tk_em2s
XI108 pd_h<3> net78 / sky130_fd_io__tk_em2s
XI97 pd_h<3> net80 / sky130_fd_io__tk_em2s
XI87 tie_lo_esd net46 / sky130_fd_io__tk_em2o
XI88 pd_h<3> net46 / sky130_fd_io__tk_em2o
XI94 tie_lo_esd net66 / sky130_fd_io__tk_em2o
XI95 pd_h<2> net66 / sky130_fd_io__tk_em2o
XI105 pd_h<2> net68 / sky130_fd_io__tk_em2o
XI103 tie_lo_esd net68 / sky130_fd_io__tk_em2o
XI101 pd_h<2> net72 / sky130_fd_io__tk_em2o
XI100 tie_lo_esd net72 / sky130_fd_io__tk_em2o
XI111 pd_h<2> net76 / sky130_fd_io__tk_em2o
XI110 pd_h<3> net76 / sky130_fd_io__tk_em2o
XI107 tie_lo_esd net78 / sky130_fd_io__tk_em2o
XI106 pd_h<2> net78 / sky130_fd_io__tk_em2o
XI98 pd_h<2> net80 / sky130_fd_io__tk_em2o
XI99 tie_lo_esd net80 / sky130_fd_io__tk_em2o
XI49 vgnd_io tie_lo_esd / sky130_fd_io__tk_tie_r_out_esd
Xn31 pad net72 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn13 pad net46 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn11<2> pad pd_h<2> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn11<1> pad pd_h<2> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn11<0> pad pd_h<2> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn34<3> pad net76 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn34<2> pad net76 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn34<1> pad net76 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn34<0> pad net76 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn33<2> pad net78 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn33<1> pad net78 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn33<0> pad net78 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn32<2> pad net68 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn32<1> pad net68 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn32<0> pad net68 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn12 pad pd_h_i2c vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn21<2> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn21<1> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn21<0> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn22<2> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn22<1> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn22<0> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn23<2> pad net66 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn23<1> pad net66 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn23<0> pad net66 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn24<2> pad net80 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn24<1> pad net80 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn24<0> pad net80 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
XI72 vgnd_io vcc_io condiode
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpio_pudrvr_unit_2_5
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpio_pudrvr_unit_2_5 pd pgin ps
*.PININFO pgin:I pd:B ps:B
XMpdrv pd pgin ps ps sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.60) l=0.60 m=2*1 p=2*(5.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpio_pudrvr_strong
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpio_pudrvr_strong pad pu_h_n<3> pu_h_n<2> tie_hi_esd vcc_io vnb
*.PININFO pu_h_n<3>:I pu_h_n<2>:I vcc_io:I vnb:I pad:O tie_hi_esd:O
XI125 pu_h_n<3> net45 / sky130_fd_io__tk_em2s
XI104 pu_h_n<3> net49 / sky130_fd_io__tk_em2s
XI109 tie_hi_esd net53 / sky130_fd_io__tk_em2s
XI108 tie_hi_esd net59 / sky130_fd_io__tk_em2s
XI112 pu_h_n<2> net43 / sky130_fd_io__tk_em2s
XI123 pu_h_n<2> net45 / sky130_fd_io__tk_em2o
XI124 tie_hi_esd net45 / sky130_fd_io__tk_em2o
XI105 pu_h_n<2> net49 / sky130_fd_io__tk_em2o
XI103 tie_hi_esd net49 / sky130_fd_io__tk_em2o
XI111 pu_h_n<2> net53 / sky130_fd_io__tk_em2o
XI110 pu_h_n<3> net53 / sky130_fd_io__tk_em2o
XI107 pu_h_n<3> net59 / sky130_fd_io__tk_em2o
XI106 pu_h_n<2> net59 / sky130_fd_io__tk_em2o
XI82 tie_hi_esd net43 / sky130_fd_io__tk_em2o
XI83 pu_h_n<3> net43 / sky130_fd_io__tk_em2o
XI49 vcc_io tie_hi_esd / sky130_fd_io__tk_tie_r_out_esd
Xn31<2> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn31<1> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn31<0> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn13<2> pad pu_h_n<2> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn13<1> pad pu_h_n<2> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn13<0> pad pu_h_n<2> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn11<2> pad pu_h_n<2> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn11<1> pad pu_h_n<2> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn11<0> pad pu_h_n<2> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn34<2> pad net53 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn34<1> pad net53 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn34<0> pad net53 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn33<1> pad net59 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn33<0> pad net59 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn32<2> pad net49 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn32<1> pad net49 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn32<0> pad net49 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn12<2> pad net43 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn12<1> pad net43 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn12<0> pad net43 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn21 pad pu_h_n<2> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn22 pad net45 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn23<2> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn23<1> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn23<0> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn24<2> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn24<1> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn24<0> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__com_pudrvr_weak
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__com_pudrvr_weak pad pu_h_n vcc_io vgnd_io vpb_drvr
*.PININFO pu_h_n:I vcc_io:I vgnd_io:I vpb_drvr:I pad:O
XMI29 pad pu_h_n vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=4*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMpdrv pad pu_h_n vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(7.00)*(0.50) l=0.50 m=4*1 p=2*(7.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=7.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpio_pddrvr_weak
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpio_pddrvr_weak pad pd_h vcc_io vgnd_io
*.PININFO pd_h:I vcc_io:I vgnd_io:I pad:O
XMndrv1 pad pd_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.60) l=0.60 m=6*1 p=2*(5.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpio_pddrvr_strong_slow
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpio_pddrvr_strong_slow pad pd_h vcc_io vgnd_io
*.PININFO pd_h:I vcc_io:I vgnd_io:I pad:O
XMndrv pad pd_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.60) l=0.60 m=4*1 p=2*(5.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__com_pudrvr_strong_slow
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__com_pudrvr_strong_slow pad pu_h_n vcc_io vgnd_io vpb_drvr
*.PININFO pu_h_n:I vcc_io:I vgnd_io:I vpb_drvr:I pad:O
XMpdrv pad pu_h_n vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(7.00)*(0.50) l=0.50 m=8*1 p=2*(7.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=7.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__tk_em1s
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__tk_em1s a b
*.PININFO a:B b:B
RI2 b net8 short m=1
RI1 a net8 short m=1
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__com_res_strong_slow
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__com_res_strong_slow ra rb vgnd_io
*.PININFO vgnd_io:I ra:B rb:B
XI28 net34 net30 / sky130_fd_io__tk_em1s
Rr1 net34 ra sky130_fd_pr__res_generic_po l=5 m=1 w=2
RI29 net30 net34 sky130_fd_pr__res_generic_po l=3 m=1 w=2
RI32 rb net30 sky130_fd_pr__res_generic_po l=2 m=1 w=2
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__tk_em1o
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__tk_em1o a b
*.PININFO a:B b:B
RI2 b net7 short m=1
RI1 a net11 short m=1
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__com_res_weak
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__com_res_weak ra rb vgnd_io
*.PININFO vgnd_io:I ra:B rb:B
Xe13 n<4> n<0> / sky130_fd_io__tk_em1s
Xe12 n<3> rb / sky130_fd_io__tk_em1s
Xe10 n<1> n<2> / sky130_fd_io__tk_em1s
Xe11 n<2> n<3> / sky130_fd_io__tk_em1s
Xe9 n<0> n<1> / sky130_fd_io__tk_em1s
Xe14 n<5> n<4> / sky130_fd_io__tk_em1o
RI134 n<5> n<4> sky130_fd_pr__res_generic_po l=6 m=1 w=0.8
RI104 n<4> n<0> sky130_fd_pr__res_generic_po l=6 m=1 w=0.8
RI116 net64 n<5> sky130_fd_pr__res_generic_po l=12 m=1 w=0.8
RI83 n<1> n<2> sky130_fd_pr__res_generic_po l=1.5 m=1 w=0.8
RI85 ra net64 sky130_fd_pr__res_generic_po l=50 m=1 w=0.8
RI82 n<2> n<3> sky130_fd_pr__res_generic_po l=1.5 m=1 w=0.8
RI62 n<3> rb sky130_fd_pr__res_generic_po l=1.5 m=1 w=0.8
RI84 n<0> n<1> sky130_fd_pr__res_generic_po l=1.5 m=1 w=0.8
.ENDS

************************************************************************
* Library Name: s8_esd
* Cell Name: s8_esd_res250only_small
* View Name: schematic
************************************************************************

.SUBCKT s8_esd_res250only_small pad rout
*.PININFO pad:B rout:B
RI228 pad net12 sky130_fd_pr__res_generic_po l=0.17 m=1 w=2
RI229 net16 rout sky130_fd_pr__res_generic_po l=0.17 m=1 w=2
RI175 net12 net16 sky130_fd_pr__res_generic_po l=10.07 m=1 w=2
RI234<1> pad net12 short m=1
RI234<2> pad net12 short m=1
RI237<1> net16 rout short m=1
RI237<2> net16 rout short m=1
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_odrvr_sub
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_odrvr_sub force_hi_h_n pad pd_h<3> pd_h<2> pd_h<1> pd_h<0> pd_h_i2c
+ pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> tie_hi_esd tie_lo_esd vcc_io vgnd vgnd_io
*.PININFO force_hi_h_n:I pd_h<3>:I pd_h<2>:I pd_h<1>:I pd_h<0>:I pd_h_i2c:I
*.PININFO pu_h_n<3>:I pu_h_n<2>:I pu_h_n<1>:I pu_h_n<0>:I vcc_io:I vgnd:I
*.PININFO vgnd_io:I pad:O tie_hi_esd:B tie_lo_esd:B
Xpddrvr_strong pad pd_h<3> pd_h<2> pd_h_i2c tie_lo_esd vcc_io vgnd_io /
+ sky130_fd_io__gpiov2_pddrvr_strong
Xpudrvr_strong pad pu_h_n<3> pu_h_n<2> tie_hi_esd vcc_io vgnd / sky130_fd_io__gpio_pudrvr_strong
Xpudrvr_weak weak_pad pu_h_n<0> vcc_io vgnd vcc_io / sky130_fd_io__com_pudrvr_weak
Xpddrvr_weak weak_pad pd_h<0> vcc_io vgnd_io / sky130_fd_io__gpio_pddrvr_weak
Xstrong_slow_pddrvr strong_slow_pad pd_h<1> vcc_io vgnd_io / sky130_fd_io__gpio_pddrvr_strong_slow
Xstrong_slow_pudrvr strong_slow_pad pu_h_n<1> vcc_io vgnd vcc_io / sky130_fd_io__com_pudrvr_strong_slow
Xres strong_slow_pad pad_r250 vgnd_io / sky130_fd_io__com_res_strong_slow
Xres_weak weak_pad pad_r250 vgnd_io / sky130_fd_io__com_res_weak
Xresd pad pad_r250 / s8_esd_res250only_small
XI72 vgnd_io vcc_io condiode
XI58 vgnd_io vcc_io condiode
XI59 vgnd_io vcc_io condiode
XI60 vgnd_io vcc_io condiode
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__com_pad
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__com_pad pad vgnd_io
*.PININFO pad:B vgnd_io:B
XDummyInstance is a cad_dummy_open_device
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_odrvr
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_odrvr force_hi_h_n pad pd_h<3> pd_h<2> pd_h<1> pd_h<0> pd_h_i2c pu_h_n<3>
+ pu_h_n<2> pu_h_n<1> pu_h_n<0> tie_hi_esd tie_lo_esd vcc_io vgnd vgnd_io
*.PININFO force_hi_h_n:I pd_h<3>:I pd_h<2>:I pd_h<1>:I pd_h<0>:I pd_h_i2c:I
*.PININFO pu_h_n<3>:I pu_h_n<2>:I pu_h_n<1>:I pu_h_n<0>:I vcc_io:I vgnd:I
*.PININFO vgnd_io:I pad:O tie_hi_esd:O tie_lo_esd:O
Xodrvr force_hi_h_n pad pd_h<3> pd_h<2> pd_h<1> pd_h<0> pd_h_i2c pu_h_n<3> pu_h_n<2>
+ pu_h_n<1> pu_h_n<0> tie_hi_esd tie_lo_esd vcc_io vgnd vgnd_io / sky130_fd_io__gpiov2_odrvr_sub
Xbondpad pad vgnd_io / sky130_fd_io__com_pad
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpio_dat_ls
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpio_dat_ls hld_h_n in out_h out_h_n rst_h set_h vcc_io vgnd
+ vpwr_ka
*.PININFO hld_h_n:I in:I rst_h:I set_h:I vcc_io:I vgnd:I vpwr_ka:I out_h:O
*.PININFO out_h_n:O
XMI30 net79 vpwr_ka net107 vgnd sky130_fd_pr__nfet_05v0_nvt AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.90) l=0.90 m=8*1 p=2*(1.00)+2*(0.90) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI31 net83 vpwr_ka net103 vgnd sky130_fd_pr__nfet_05v0_nvt AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.90) l=0.90 m=8*1 p=2*(1.00)+2*(0.90) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI35 in_i in_i_n vgnd vgnd sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.25) l=0.25 m=2*1 p=2*(1.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI34 in_i_n in vgnd vgnd sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.25) l=0.25 m=2*1 p=2*(1.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMmnrst fbk rst_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMmnset fbk_n set_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI13 out_h_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=1*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI12 out_h fbk_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=1*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI8 net103 in_i vgnd vgnd sky130_fd_pr__nfet_01v8_lvt AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.15) l=0.15 m=8*1 p=2*(1.00)+2*(0.15) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI7 net107 in_i_n vgnd vgnd sky130_fd_pr__nfet_01v8_lvt AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.15) l=0.15 m=8*1 p=2*(1.00)+2*(0.15) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI6 fbk_n hld_h_n net83 vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI5 fbk hld_h_n net79 vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI4 fbk_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.70)*(0.60) l=0.60 m=1*1 p=2*(0.70)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.70
XMI3 fbk fbk_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.70)*(0.60) l=0.60 m=1*1 p=2*(0.70)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.70
XMI32 in_i_n in vpwr_ka vpwr_ka sky130_fd_pr__pfet_01v8_hvt AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.25) l=0.25 m=1*1 p=2*(3.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI14 out_h_n fbk vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI11 out_h fbk_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI33 in_i in_i_n vpwr_ka vpwr_ka sky130_fd_pr__pfet_01v8_hvt AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.25) l=0.25 m=1*1 p=2*(3.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI2 fbk fbk_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=1*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI1 fbk_n fbk vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=1*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__com_cclat_hvnor3
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__com_cclat_hvnor3 in0 in1 in2 out vcc_io vgnd vnb
*.PININFO in0:I in1:I in2:I vcc_io:I vgnd:I vnb:I out:O
XMmp1 n<1> in1 n<0> vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=4*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMmp2 out in2 n<1> vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=4*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMmp0 n<0> in0 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.60) l=0.60 m=8*1 p=2*(5.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMmn1 out in1 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=2*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMmn2 out in2 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=2*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMmn0 out in0 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=2*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__com_cclat_hvnand3
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__com_cclat_hvnand3 in0 in1 in2 out vcc_io vgnd vnb
*.PININFO in0:I in1:I in2:I vcc_io:I vgnd:I vnb:I out:O
XMmp1 out in1 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMmp2 out in2 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMmp0 out in0 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMmn1 n1 in1 n0 vnb sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=2*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMmn0 n0 in0 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=4*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMmn2 out in2 n1 vnb sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=2*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__com_cclat_inv_in
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__com_cclat_inv_in in out vcc_io vgnd vnb
*.PININFO in:I vcc_io:I vgnd:I vnb:I out:O
XMmp1 out in vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMmn1 out in vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__com_cclat_inv_out
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__com_cclat_inv_out in out vcc_io vgnd vnb
*.PININFO in:I vcc_io:I vgnd:I vnb:I out:O
XMI1 out in vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=6*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI2 out in vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=6*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__com_cclat
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__com_cclat drvhi_h drvlo_h_n oe_h_n pd_dis_h pu_dis_h vcc_io vgnd
*.PININFO oe_h_n:I pd_dis_h:I pu_dis_h:I vcc_io:I vgnd:I drvhi_h:O drvlo_h_n:O
Xnor3 oe_i_h_n drvhi_h pd_dis_h n1 vcc_io vgnd vgnd / sky130_fd_io__com_cclat_hvnor3
Xnand3 oe_i_h drvlo_h_n pu_dis_h_n n0 vcc_io vgnd vgnd / sky130_fd_io__com_cclat_hvnand3
Xinv_pudis pu_dis_h pu_dis_h_n vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_in
Xinv_oe2 oe_i_h oe_i_h_n vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_in
Xinv_oe1 oe_h_n oe_i_h vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_in
Xinv_out_1 n0 drvhi_h vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_out
Xinv_out n1 drvlo_h_n vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_out
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_opath_datoe
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_opath_datoe drvhi_h drvlo_h_n hld_h_n hld_i_ovr_h od_h oe_h oe_n out
+ vcc_io vgnd vpwr_ka
*.PININFO hld_h_n:I hld_i_ovr_h:I od_h:I oe_n:I out:I vcc_io:I vgnd:I
*.PININFO vpwr_ka:I drvhi_h:O drvlo_h_n:O oe_h:O
Xoe_ls hld_i_ovr_h oe_n oe_h_n oe_h vgnd od_h vcc_io vgnd vpwr_ka
+ / sky130_fd_io__gpio_dat_ls
Xdat_ls hld_i_ovr_h out pd_dis_h pu_dis_h vgnd od_h vcc_io vgnd vpwr_ka
+ / sky130_fd_io__gpio_dat_ls
Xcclat drvhi_h drvlo_h_n oe_h_n pd_dis_h pu_dis_h vcc_io vgnd / sky130_fd_io__com_cclat
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__hvsbt_xor
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__hvsbt_xor in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
XMI12 out net70 net29 vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=2*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI13 net45 in1 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=2*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI18 net54 in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=2*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI17 net70 in1 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=2*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI5 out net54 net45 vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=2*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI3 net29 in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=2*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI19 net54 in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.70)*(0.60) l=0.60 m=1*1 p=2*(0.70)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.70
XMI14 net58 in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.70)*(0.60) l=0.60 m=1*1 p=2*(0.70)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.70
XMI15 net62 net54 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.70)*(0.60) l=0.60 m=1*1 p=2*(0.70)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.70
XMI6 out net70 net62 vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.70)*(0.60) l=0.60 m=1*1 p=2*(0.70)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.70
XMI16 net70 in1 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.70)*(0.60) l=0.60 m=1*1 p=2*(0.70)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.70
XMI1 out in1 net58 vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.70)*(0.60) l=0.60 m=1*1 p=2*(0.70)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.70
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__com_ctl_ls
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__com_ctl_ls hld_h_n in out_h out_h_n rst_h set_h vcc_io vgnd
+ vpwr
*.PININFO hld_h_n:I in:I rst_h:I set_h:I vcc_io:I vgnd:I vpwr:I out_h:O
*.PININFO out_h_n:O
XMI1 fbk_n fbk vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.75)*(0.50) l=0.50 m=1*1 p=2*(0.75)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.75
XMI2 fbk fbk_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.75)*(0.50) l=0.50 m=1*1 p=2*(0.75)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.75
XMI11 out_h fbk_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI29 in_i_n in vpwr vpwr sky130_fd_pr__pfet_01v8_hvt AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.25) l=0.25 m=1*1 p=2*(1.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI34 in_i in_i_n vpwr vpwr sky130_fd_pr__pfet_01v8_hvt AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.25) l=0.25 m=1*1 p=2*(1.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI14 out_h_n fbk vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI7 net94 in_i_n vgnd vgnd sky130_fd_pr__nfet_01v8_lvt AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.15) l=0.15 m=4*1 p=2*(1.00)+2*(0.15) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI8 net98 in_i vgnd vgnd sky130_fd_pr__nfet_01v8_lvt AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.15) l=0.15 m=4*1 p=2*(1.00)+2*(0.15) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI3 fbk fbk_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.75)*(1.00) l=1.00 m=1*1 p=2*(0.75)+2*(1.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.75
XMI4 fbk_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.75)*(1.00) l=1.00 m=1*1 p=2*(0.75)+2*(1.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.75
XMI5 fbk hld_h_n net130 vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI27 in_i_n in vgnd vgnd sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.25) l=0.25 m=1*1 p=2*(1.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI6 fbk_n hld_h_n net122 vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI59 net122 vpwr net98 vgnd sky130_fd_pr__nfet_05v0_nvt AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.90) l=0.90 m=4*1 p=2*(1.00)+2*(0.90) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMmnrst fbk rst_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI58 net130 vpwr net94 vgnd sky130_fd_pr__nfet_05v0_nvt AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.90) l=0.90 m=4*1 p=2*(1.00)+2*(0.90) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI12 out_h fbk_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=1*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI32 in_i in_i_n vgnd vgnd sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.25) l=0.25 m=1*1 p=2*(1.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMmnset fbk_n set_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI13 out_h_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=1*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_octl
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_octl dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n od_h
+ pden_h_n<2> pden_h_n<1> pden_h_n<0> puen_0_h puen_2or1_h puen_h<1> puen_h<0> slow slow_h slow_h_n
+ vcc_io vgnd vpwr vreg_en_h_n
*.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I
*.PININFO hld_i_h_n:I od_h:I slow:I vcc_io:I vgnd:I vpwr:I vreg_en_h_n:I
*.PININFO pden_h_n<2>:O pden_h_n<1>:O pden_h_n<0>:O puen_0_h:O puen_2or1_h:O
*.PININFO puen_h<1>:O puen_h<0>:O slow_h:O slow_h_n:O
XI381 dm_h<1> dm_h<0> net70 vgnd vcc_io / sky130_fd_io__hvsbt_nor
XI201 dm_h_n<2> dm_h_n<1> n<9> vgnd vcc_io / sky130_fd_io__hvsbt_nor
XI211 n<8> dm_h_n<1> puen_0_h vgnd vcc_io / sky130_fd_io__hvsbt_nor
XI200 dm_h<2> dm_h<1> n<10> vgnd vcc_io / sky130_fd_io__hvsbt_xor
XI210 dm_h<2> dm_h<0> n<8> vgnd vcc_io / sky130_fd_io__hvsbt_xor
XI382 dm_h<2> net70 pden_h_n<2> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI205 n<1> n<0> puen_2or1_h vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI204 n<9> dm_h_n<0> n<0> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI203 n<10> dm_h<0> n<1> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI208 puen_2or1_h vreg_en_h_n n<5> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI187 dm_h<1> dm_h<0> n<3> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI186 dm_h_n<2> dm_h_n<1> n<4> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI185 dm_h_n<0> n<4> net130 vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI247 pden_h1 pden_h_n<1> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
XI249 pden_h0 pden_h_n<0> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
XI256 puen_h0_n puen_h<0> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
XI254 puen_h1_n puen_h<1> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
XI375 n<3> pden_h0 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI374 net130 pden_h1 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI376 n<2> puen_h1_n vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI209 n<5> n<2> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI377 puen_0_h puen_h0_n vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
Xls_slow hld_i_h_n slow slow_h slow_h_n od_h vgnd vcc_io vgnd vpwr
+ / sky130_fd_io__com_ctl_ls
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_pupredrvr_strong_nd2
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_pupredrvr_strong_nd2 drvhi_h en_fast<3> en_fast<2> en_fast<1> en_fast<0>
+ pu_h_n puen_h vcc_io vgnd_io
*.PININFO drvhi_h:I en_fast<3>:I en_fast<2>:I en_fast<1>:I en_fast<0>:I
*.PININFO puen_h:I vcc_io:I vgnd_io:I pu_h_n:O
XE1 net24 pu_h_n / sky130_fd_io__tk_em1s
Rrespu2 pu_h_n int_res sky130_fd_pr__res_generic_po l=4 m=1 w=0.33
Rrespu1 int_res net24 sky130_fd_pr__res_generic_po l=11 m=1 w=0.33
XMmnen_fast<3> int<3> en_fast<3> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(1.00) l=1.00 m=1*1 p=2*(1.50)+2*(1.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMmnen_fast<2> int<2> en_fast<2> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(1.00) l=1.00 m=1*1 p=2*(1.50)+2*(1.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMmnen_fast<1> int<1> en_fast<1> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(1.00) l=1.00 m=1*1 p=2*(1.50)+2*(1.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMmnen_fast<0> int<0> en_fast<0> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(1.00) l=1.00 m=1*1 p=2*(1.50)+2*(1.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMmnin_slow pu_h_n drvhi_h n<2> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(4.00) l=4.00 m=1*1 p=2*(0.42)+2*(4.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMmnen_slow1 n<2> puen_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(4.00) l=4.00 m=1*1 p=2*(0.42)+2*(4.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMmnin_fast<3> net24 drvhi_h int<3> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMmnin_fast<2> net24 drvhi_h int<2> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMmnin_fast<1> net24 drvhi_h int<1> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMmnin_fast<0> net24 drvhi_h int<0> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMmpin pu_h_n drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.60) l=0.60 m=3*1 p=2*(5.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMmpen pu_h_n puen_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.60) l=0.60 m=1*1 p=2*(5.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__tk_opti
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__tk_opti out spd spu
*.PININFO out:B spd:B spu:B
Xe2 spd out / sky130_fd_io__tk_em1o
Xe1 out spu / sky130_fd_io__tk_em1s
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__tk_opto
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__tk_opto out spd spu
*.PININFO out:B spd:B spu:B
Xe1 spu out / sky130_fd_io__tk_em1o
Xe2 out spd / sky130_fd_io__tk_em1s
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__com_inv_x1_dnw
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__com_inv_x1_dnw in out vgnd vpwr
*.PININFO in:I vgnd:I vpwr:I out:O
XMI1 out in vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI2 out in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=1*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__com_pupredrvr_nbias
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__com_pupredrvr_nbias drvhi_h en_h en_h_n nbias pu_h_n puen_h vcc_io vgnd_io
*.PININFO drvhi_h:I en_h:I en_h_n:I pu_h_n:I puen_h:I vcc_io:I vgnd_io:I
*.PININFO nbias:O
XI36 n<2> pu_h_n en_h / sky130_fd_io__tk_opto
XE6 net141 nbias / sky130_fd_io__tk_em1s
XE7 bias_g net90 / sky130_fd_io__tk_em1s
XE4 n<6> net153 / sky130_fd_io__tk_em1s
XE5 nbias net88 / sky130_fd_io__tk_em1s
XE2 n<6> nbias / sky130_fd_io__tk_em1o
XE1 n<2> n<1> / sky130_fd_io__tk_em1o
XMI56 vcc_io pu_h_n net90 vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(8.00) l=8.00 m=1*1 p=2*(0.42)+2*(8.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI50 n<1> puen_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=1*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI49 net88 bias_g vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.80) l=0.80 m=4*1 p=2*(1.00)+2*(0.80) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI47 n<7> bias_g vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=2*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI12 drvhi_i_h_n drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=2*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI21 nbias bias_g vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.80) l=0.80 m=4*1 p=2*(1.00)+2*(0.80) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI29 bias_g en_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=1*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI30 bias_g drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=1*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI31 bias_g n<1> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=4*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI32 n<1> n<2> n<2> vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI34 n<1> drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=1*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI54 net141 bias_g vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(4.00) l=4.00 m=1*1 p=2*(0.42)+2*(4.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI41 n<7> n<7> n<8> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=2*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI44 n<8> n<8> vccio_2vtn vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=2*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI39 net153 vccio_2vtn vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=4*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI40 vccio_2vtn vcc_io vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(8.00) l=8.00 m=1*1 p=2*(0.42)+2*(8.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI25 nbias drvhi_i_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI53 vccio_2vtn drvhi_i_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI24 nbias en_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI13 drvhi_i_h_n drvhi_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=1*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI26 n<4> en_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMI27 n<3> n<2> n<4> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMI28 bias_g drvhi_h n<3> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMI20 nbias nbias n<6> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=4*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI19 n<6> n<6> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=4*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__com_nand2_dnw
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__com_nand2_dnw in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
XMI5 out in1 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI3 out in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI6 net25 in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=1*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI1 out in1 net25 vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=1*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_pupredrvr_strong
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_pupredrvr_strong drvhi_h pu_h_n<3> pu_h_n<2> puen_h slow_h_n vcc_io vgnd_io
*.PININFO drvhi_h:I puen_h:I slow_h_n:I vcc_io:I vgnd_io:I pu_h_n<3>:O
*.PININFO pu_h_n<2>:O
Xnd2a drvhi_h net54 net54 net54 net54 pu_h_n<2> puen_h vcc_io vgnd_io
+ / sky130_fd_io__gpiov2_pupredrvr_strong_nd2
Xnd2b drvhi_h en_fast_h_3<3> en_fast_h_3<2> en_fast_h_3<1> en_fast_h_3<0> pu_h_n<3> puen_h vcc_io
+ vgnd_io / sky130_fd_io__gpiov2_pupredrvr_strong_nd2
XI97 en_fast_h_3<1> en_fast_h_3<3> vgnd_io / sky130_fd_io__tk_opti
XI98 en_fast_h_3<0> en_fast_h_3<3> vgnd_io / sky130_fd_io__tk_opti
XI93 net54 nbias_out en_fast_h / sky130_fd_io__tk_opto
XI96 en_fast_h_3<2> en_fast_h_3<3> vgnd_io / sky130_fd_io__tk_opto
XI92 en_fast_h_3<3> nbias_out en_fast_h / sky130_fd_io__tk_opto
Xinv en_fast_h_n en_fast_h vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
Xnbias drvhi_h en_fast_h en_fast_h_n nbias_out pu_h_n<2> puen_h vcc_io vgnd_io /
+ sky130_fd_io__com_pupredrvr_nbias
Xnand puen_h slow_h_n en_fast_h_n vgnd_io vcc_io / sky130_fd_io__com_nand2_dnw
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_octl_mux
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_octl_mux a_h b_h sel_h sel_h_n vccio vssio y_h
*.PININFO a_h:I b_h:I sel_h:I sel_h_n:I vccio:I vssio:I y_h:O
XMI3 y_h sel_h_n a_h vccio sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI2 y_h sel_h b_h vccio sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI4 a_h sel_h y_h vssio sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI1 b_h sel_h_n y_h vssio sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_pdpredrvr_strong_nr2
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_pdpredrvr_strong_nr2 drvlo_h_n en_fast_n<1> en_fast_n<0> i2c_mode_h pd_h
+ pd_i2c_h pden_h_n vcc_io vgnd_io
*.PININFO drvlo_h_n:I en_fast_n<1>:I en_fast_n<0>:I i2c_mode_h:I pden_h_n:I
*.PININFO vcc_io:I vgnd_io:I pd_h:O pd_i2c_h:O
XMI101 net45 pden_h_n net039 vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(4.00) l=4.00 m=1*1 p=2*(0.42)+2*(4.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI73 net42 i2c_mode_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=3*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI76 pd_h drvlo_h_n net45 vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(4.00) l=4.00 m=1*1 p=2*(0.42)+2*(4.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI75 net039 pden_h_n net42 vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(4.00) l=4.00 m=1*1 p=2*(0.42)+2*(4.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI74<1> pd_h drvlo_h_n net53<0> vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=2*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI74<0> pd_h drvlo_h_n net53<1> vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=2*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI72<1> net53<0> en_fast_n<1> net42 vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI72<0> net53<1> en_fast_n<0> net42 vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMmpen_fast1 net62 en_fast_n<1> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(1.00) l=1.00 m=1*1 p=2*(0.42)+2*(1.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMmpin_fast<1> pd_i2c_h drvlo_h_n net62 vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(1.00) l=1.00 m=1*1 p=2*(0.42)+2*(1.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMmpin_fast<0> pd_i2c_h drvlo_h_n net62 vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(1.00) l=1.00 m=1*1 p=2*(0.42)+2*(1.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMmpen_slow int_slow pden_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(4.00) l=4.00 m=1*1 p=2*(0.42)+2*(4.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMmpin_slow pd_i2c_h drvlo_h_n int_slow vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(4.00) l=4.00 m=1*1 p=2*(0.42)+2*(4.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI77 pd_h drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=2*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI78 pd_h pden_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMmnen pd_i2c_h pden_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMmnin pd_i2c_h drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=2*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI94 pd_h i2c_mode_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_pdpredrvr_strong_nr3
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_pdpredrvr_strong_nr3 drvlo_h_n en_fast_n<1> en_fast_n<0> i2c_mode_h pd_h
+ pden_h_n vcc_io vgnd_io
*.PININFO drvlo_h_n:I en_fast_n<1>:I en_fast_n<0>:I i2c_mode_h:I pden_h_n:I
*.PININFO vcc_io:I vgnd_io:I pd_h:O
XMI85 int1 i2c_mode_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=2*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI86<1> int2 en_fast_n<1> int1 vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(0.50) l=0.50 m=1*1 p=2*(0.42)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI86<0> int2 en_fast_n<0> int1 vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(0.50) l=0.50 m=1*1 p=2*(0.42)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI87<1> pd_h drvlo_h_n int2 vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(0.50) l=0.50 m=1*1 p=2*(0.42)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI87<0> pd_h drvlo_h_n int2 vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(0.50) l=0.50 m=1*1 p=2*(0.42)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI56 net43 pden_h_n int1 vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(2.00) l=2.00 m=1*1 p=2*(0.42)+2*(2.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI90 pd_h drvlo_h_n net43 vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(2.00) l=2.00 m=1*1 p=2*(0.42)+2*(2.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMmpen_fast<1> int_nor<1> en_fast_n<1> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMmpen_fast<0> int_nor<0> en_fast_n<0> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMmpin_fast<1> pd_h drvlo_h_n int_nor<1> vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMmpin_fast<0> pd_h drvlo_h_n int_nor<0> vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMmpen_slow int_slow pden_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(4.00) l=4.00 m=1*1 p=2*(0.42)+2*(4.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMmpin_slow pd_h drvlo_h_n int_slow vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(2.00) l=2.00 m=1*1 p=2*(0.42)+2*(2.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMmnen pd_h pden_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=2*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMmnin pd_h drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=5*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__com_pdpredrvr_pbias
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__com_pdpredrvr_pbias drvlo_h_n en_h en_h_n pbias pd_h pden_h_n vcc_io vgnd_io
*.PININFO drvlo_h_n:I en_h:I en_h_n:I pd_h:I pden_h_n:I vcc_io:I vgnd_io:I
*.PININFO pbias:O
XI27 n<0> pd_h en_h_n / sky130_fd_io__tk_opto
XE2 pbias pbias1 / sky130_fd_io__tk_em1o
XE1 n<1> n<0> / sky130_fd_io__tk_em1o
XE5 n<101> bias_g / sky130_fd_io__tk_em1s
XE6 pbias net84 / sky130_fd_io__tk_em1s
XE4 net108 pbias / sky130_fd_io__tk_em1s
XE3 pbias1 net88 / sky130_fd_io__tk_em1s
XMI41 n<101> pd_h n<100> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(4.00) l=4.00 m=1*1 p=2*(0.42)+2*(4.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI48 n<100> pd_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(4.00) l=4.00 m=1*1 p=2*(0.42)+2*(4.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI38 n<1> pden_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=1*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI36 net108 bias_g vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(1.00) l=1.00 m=2*1 p=2*(1.00)+2*(1.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI34 net157 bias_g vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.60) l=0.60 m=1*1 p=2*(5.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI19 bias_g en_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=1*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI20 bias_g n<1> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.60) l=0.60 m=1*1 p=2*(5.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI13 drvlo_i_h drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=1*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI23 n<0> n<0> n<1> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI18 bias_g drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=1*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI24 n<1> drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=1*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI47 pbias bias_g vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(1.00) l=1.00 m=2*1 p=2*(1.00)+2*(1.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI40 2vtp drvlo_i_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI43 net84 bias_g vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(4.00) l=4.00 m=1*1 p=2*(0.42)+2*(4.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI30 net88 2vtp vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=8*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI31 net157 net157 net161 vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=4*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI32 net161 net161 2vtp vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=4*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI33 2vtp vgnd_io vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(8.00) l=8.00 m=1*1 p=2*(0.42)+2*(8.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XMI14 pbias drvlo_i_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI17 bias_g drvlo_h_n net171 vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI12 drvlo_i_h drvlo_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.50) l=0.50 m=2*1 p=2*(1.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI6 pbias en_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI16 net171 n<0> net183 vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI15 net183 en_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI45 pbias1 pbias1 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=8*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI44 pbias pbias pbias1 vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=8*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__com_nor2_dnw
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__com_nor2_dnw in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
XMI12 out in1 net17 vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI3 net17 in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI6 out in1 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=1*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI1 out in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=1*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_pdpredrvr_strong
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_pdpredrvr_strong drvlo_h_n i2c_mode_h_n pd_h<4> pd_h<3> pd_h<2> pden_h_n
+ slow_h tie_hi_esd vcc_io vgnd vgnd_io
*.PININFO drvlo_h_n:I i2c_mode_h_n:I pden_h_n:I slow_h:I tie_hi_esd:I vcc_io:I
*.PININFO vgnd:I vgnd_io:I pd_h<4>:O pd_h<3>:O pd_h<2>:O
XMI87 mod_drvlo_h_n_i2c pd_h<4> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI88 mod_drvlo_h_n_i2c pd_h<4> vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.42)*(0.50) l=0.50 m=1*1 p=2*(0.42)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.42
XI98 i2c_mode_h slow_h int_slow1 vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI160 i2c_mode_h_n slow_h net75 vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI93 i2c_mode_h_n i2c_mode_h vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI97 int_slow1 mod_slow_h vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI161 net75 net142 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
Xmux mod_drvlo_h_n_i2c drvlo_h_n i2c_mode_h i2c_mode_h_n vcc_io vgnd_io mod_drvlo_h_n /
+ sky130_fd_io__gpiov2_octl_mux
Xnr3 drvlo_h_n pbias_out pbias_out mod_slow_h pd_h<2> pd_h<4> pden_h_n vcc_io vgnd_io
+ / sky130_fd_io__gpiov2_pdpredrvr_strong_nr2
Xnr2 mod_drvlo_h_n en_fast2_n<1> en_fast2_n<0> mod_slow_h pd_h<3> pden_h_n vcc_io vgnd_io /
+ sky130_fd_io__gpiov2_pdpredrvr_strong_nr3
XI76 net118 pbias_out en_fast_h_n / sky130_fd_io__tk_opto
XI77 en_fast2_n<1> pbias_out en_fast_h_n / sky130_fd_io__tk_opto
XI79 en_fast2_n<0> en_fast2_n<1> vcc_io / sky130_fd_io__tk_opti
Xinv en_fast_h en_fast_h_n vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
Xbias drvlo_h_n en_fast_h en_fast_h_n pbias_out pd_h<4> pden_h_n vcc_io vgnd_io /
+ sky130_fd_io__com_pdpredrvr_pbias
Xnor net142 pden_h_n en_fast_h vgnd_io vcc_io / sky130_fd_io__com_nor2_dnw
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__com_pupredrvr_weak
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__com_pupredrvr_weak drvhi_h pu_h_n puen_h vcc_io vgnd_io
*.PININFO drvhi_h:I puen_h:I vcc_io:I vgnd_io:I pu_h_n:O
XMI39 net21 puen_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI3 pu_h_n drvhi_h net21 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI37 pu_h_n drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.60) l=0.60 m=2*1 p=2*(5.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI38 pu_h_n puen_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.60) l=0.60 m=1*1 p=2*(5.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__com_pdpredrvr_weak
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__com_pdpredrvr_weak drvlo_h_n pd_h pden_h_n vcc_io vgnd_io
*.PININFO drvlo_h_n:I pden_h_n:I vcc_io:I vgnd_io:I pd_h:O
XMI25 pd_h drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI26 pd_h pden_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI23 pd_h drvlo_h_n net25 vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI24 net25 pden_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=2*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__com_pupredrvr_strong_slow
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__com_pupredrvr_strong_slow drvhi_h pu_h_n puen_h vcc_io vgnd_io
*.PININFO drvhi_h:I puen_h:I vcc_io:I vgnd_io:I pu_h_n:O
XMI39 net17 puen_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=2*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI3 pu_h_n drvhi_h net17 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=2*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI37 pu_h_n drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=3*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI38 pu_h_n puen_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__com_pdpredrvr_strong_slow
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__com_pdpredrvr_strong_slow drvlo_h_n pd_h pden_h_n vcc_io vgnd_io
*.PININFO drvlo_h_n:I pden_h_n:I vcc_io:I vgnd_io:I pd_h:O
XMI25 pd_h drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI26 pd_h pden_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.60) l=0.60 m=1*1 p=2*(3.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI23 pd_h drvlo_h_n net25 vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=2*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI24 net25 pden_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=2*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_obpredrvr
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_obpredrvr drvhi_h drvlo_h_n i2c_mode_h_n pd_h<4> pd_h<3> pd_h<2> pd_h<1>
+ pd_h<0> pden_h_n<1> pden_h_n<0> pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> puen_h<1> puen_h<0>
+ slow_h slow_h_n tie_hi_esd vcc_io vgnd vgnd_io
*.PININFO drvhi_h:I drvlo_h_n:I i2c_mode_h_n:I pden_h_n<1>:I pden_h_n<0>:I
*.PININFO puen_h<1>:I puen_h<0>:I slow_h:I slow_h_n:I tie_hi_esd:I vcc_io:I
*.PININFO vgnd:I vgnd_io:I pd_h<4>:O pd_h<3>:O pd_h<2>:O pd_h<1>:O pd_h<0>:O
*.PININFO pu_h_n<3>:O pu_h_n<2>:O pu_h_n<1>:O pu_h_n<0>:O
Xpu_strong drvhi_h pu_h_n<3> pu_h_n<2> puen_h<1> slow_h_n vcc_io vgnd_io /
+ sky130_fd_io__gpiov2_pupredrvr_strong
Xpd_strong drvlo_h_n i2c_mode_h_n pd_h<4> pd_h<3> pd_h<2> pden_h_n<1> slow_h tie_hi_esd vcc_io
+ vgnd vgnd_io / sky130_fd_io__gpiov2_pdpredrvr_strong
Xpu_weak drvhi_h pu_h_n<0> puen_h<0> vcc_io vgnd_io / sky130_fd_io__com_pupredrvr_weak
Xpd_weak drvlo_h_n pd_h<0> pden_h_n<0> vcc_io vgnd_io / sky130_fd_io__com_pdpredrvr_weak
Xpu_strong_slow drvhi_h pu_h_n<1> puen_h<1> vcc_io vgnd_io / sky130_fd_io__com_pupredrvr_strong_slow
Xpd_strong_slow drvlo_h_n pd_h<1> pden_h_n<1> vcc_io vgnd_io / sky130_fd_io__com_pdpredrvr_strong_slow
XI15 vgnd_io vcc_io condiode
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_octl_dat
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_octl_dat dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> drvhi_h
+ hld_i_h_n hld_i_ovr_h od_h oe_n out pd_h<4> pd_h<3> pd_h<2> pd_h<1> pd_h<0> pu_h_n<3>
+ pu_h_n<2> pu_h_n<1> pu_h_n<0> slow slow_h_n tie_hi_esd vcc_io vgnd vgnd_io vpwr vpwr_ka
*.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I
*.PININFO hld_i_h_n:I hld_i_ovr_h:I od_h:I oe_n:I out:I slow:I tie_hi_esd:I
*.PININFO vcc_io:I vgnd:I vgnd_io:I vpwr:I vpwr_ka:I drvhi_h:O pd_h<4>:O
*.PININFO pd_h<3>:O pd_h<2>:O pd_h<1>:O pd_h<0>:O pu_h_n<3>:O pu_h_n<2>:O
*.PININFO pu_h_n<1>:O pu_h_n<0>:O slow_h_n:O
Xdatoe drvhi_h drvlo_h_n hld_i_h_n hld_i_ovr_h od_h oe_h oe_n out vcc_io
+ vgnd vpwr_ka / sky130_fd_io__gpiov2_opath_datoe
Xctl dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n od_h pden_h_n<2>
+ pden_h_n<1> pden_h_n<0> puen_0_h puen_2or1_h puen_h<1> puen_h<0> slow slow_h slow_h_n vcc_io vgnd
+ vpwr vcc_io / sky130_fd_io__gpiov2_octl
Xpredrvr drvhi_h drvlo_h_n pden_h_n<2> pd_h<4> pd_h<3> pd_h<2> pd_h<1> pd_h<0> pden_h_n<1>
+ pden_h_n<0> pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> puen_h<1> puen_h<0> slow_h slow_h_n
+ tie_hi_esd vcc_io vgnd vgnd_io / sky130_fd_io__gpiov2_obpredrvr
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_opath
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_opath dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n
+ hld_i_ovr_h od_h oe_n out pad slow tie_hi_esd tie_lo_esd vcc_io vgnd vgnd_io
+ vpwr vpwr_ka
*.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I
*.PININFO hld_i_h_n:I hld_i_ovr_h:I od_h:I oe_n:I out:I slow:I vcc_io:I vgnd:I
*.PININFO vgnd_io:I vpwr:I vpwr_ka:I pad:O tie_hi_esd:O tie_lo_esd:O
Xodrvr net70 pad pd_h<3> pd_h<2> pd_h<1> pd_h<0> pd_h<4> pu_h_n<3> pu_h_n<2>
+ pu_h_n<1> pu_h_n<0> tie_hi_esd tie_lo_esd vcc_io vgnd vgnd_io / sky130_fd_io__gpiov2_odrvr
Xopath dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> drvhi_h hld_i_h_n hld_i_ovr_h
+ od_h oe_n out pd_h<4> pd_h<3> pd_h<2> pd_h<1> pd_h<0> pu_h_n<3> pu_h_n<2> pu_h_n<1>
+ pu_h_n<0> slow slow_h_n tie_hi_esd vcc_io vgnd vgnd_io vpwr vpwr_ka / sky130_fd_io__gpiov2_octl_dat
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__hvsbt_inv_x4
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__hvsbt_inv_x4 in out vgnd vpwr
*.PININFO in:I vgnd:I vpwr:I out:O
XMI1 out in vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=8*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI2 out in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.70)*(0.60) l=0.60 m=4*1 p=2*(0.70)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.70
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__hvsbt_inv_x8
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__hvsbt_inv_x8 in out vgnd vpwr
*.PININFO in:I vgnd:I vpwr:I out:O
XMI2 out in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(0.70)*(0.60) l=0.60 m=8*1 p=2*(0.70)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=0.70
XMI1 out in vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.60) l=0.60 m=16*1 p=2*(1.00)+2*(0.60) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_ctl_hld
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_ctl_hld enable_h hld_h_n hld_i_h hld_i_h_n hld_i_ovr_h hld_ovr od_i_h vcc_io
+ vgnd vpwr
*.PININFO enable_h:I hld_h_n:I hld_ovr:I vcc_io:I vgnd:I vpwr:I hld_i_h:O
*.PININFO hld_i_h_n:O hld_i_ovr_h:O od_i_h:O
Xhld_ovr_ls net65 hld_ovr hld_ovr_h net37 od_h vgnd vcc_io vgnd vpwr
+ / sky130_fd_io__com_ctl_ls
XI26 net65 hld_ovr_h hld_i_ovr_h_n vgnd vcc_io / sky130_fd_io__hvsbt_nor
XI30 od_i_h hld_i_ovr_h_n hld_i_ovr_h vgnd vcc_io / sky130_fd_io__hvsbt_nor
XI31 od_i_h_n od_i_h vgnd vcc_io / sky130_fd_io__hvsbt_inv_x4
Xhld_i_h_inv4 net65 enable_vdda_h_n vgnd vcc_io / sky130_fd_io__hvsbt_inv_x4
Xhld_nand enable_h hld_h_n net64 vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI32 od_h od_i_h_n vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
Xhld_i_h_inv1 net64 net65 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
Xod_h_inv enable_h od_h vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
Xhld_i_h_inv8<1> enable_vdda_h_n hld_i_h_n_net<1> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x8
Xhld_i_h_inv8<0> enable_vdda_h_n hld_i_h_n_net<0> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x8
Rshort_hld_i_h enable_vdda_h_n hld_i_h short m=1
Rshort<1> hld_i_h_n_net<1> hld_i_h_n short m=1
Rshort<0> hld_i_h_n_net<0> hld_i_h_n short m=1
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_ctl_lsbank
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_ctl_lsbank dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1>
+ dm_h_n<0> hld_i_h_n ib_mode_sel ib_mode_sel_h ib_mode_sel_h_n inp_dis inp_dis_h inp_dis_h_n
+ od_i_h startup_rst_h startup_st_h vcc_io vgnd vpwr vtrip_sel vtrip_sel_h vtrip_sel_h_n
*.PININFO dm<2>:I dm<1>:I dm<0>:I hld_i_h_n:I ib_mode_sel:I inp_dis:I od_i_h:I
*.PININFO startup_rst_h:I startup_st_h:I vcc_io:I vgnd:I vpwr:I vtrip_sel:I
*.PININFO dm_h<2>:O dm_h<1>:O dm_h<0>:O dm_h_n<2>:O dm_h_n<1>:O dm_h_n<0>:O
*.PININFO ib_mode_sel_h:O ib_mode_sel_h_n:O inp_dis_h:O inp_dis_h_n:O
*.PININFO vtrip_sel_h:O vtrip_sel_h_n:O
XI337<1> dm_st_h<0> startup_rst_h startup_st_h / sky130_fd_io__tk_opti
XI597 ib_mode_sel_rst_h vgnd od_i_h / sky130_fd_io__tk_opti
XI598 ib_mode_sel_st_h od_i_h vgnd / sky130_fd_io__tk_opti
XI805<1> dm_rst_h<1> vgnd od_i_h / sky130_fd_io__tk_opti
XI804<1> dm_rst_h<2> vgnd od_i_h / sky130_fd_io__tk_opti
XI802<1> dm_st_h<2> od_i_h vgnd / sky130_fd_io__tk_opti
XI803<1> dm_st_h<1> od_i_h vgnd / sky130_fd_io__tk_opti
XI338<1> dm_rst_h<0> startup_st_h startup_rst_h / sky130_fd_io__tk_opti
Xie_n_st ie_n_st_h startup_st_h startup_rst_h / sky130_fd_io__tk_opti
Xie_n_rst ie_n_rst_h startup_rst_h startup_st_h / sky130_fd_io__tk_opti
Xtrip_sel_rst trip_sel_rst_h vgnd od_i_h / sky130_fd_io__tk_opti
Xtrip_sel_st trip_sel_st_h od_i_h vgnd / sky130_fd_io__tk_opti
XI595 hld_i_h_n ib_mode_sel ib_mode_sel_h ib_mode_sel_h_n ib_mode_sel_rst_h ib_mode_sel_st_h vcc_io
+ vgnd vpwr / sky130_fd_io__com_ctl_ls
Xdm_ls<2> hld_i_h_n dm<2> dm_h<2> dm_h_n<2> dm_rst_h<2> dm_st_h<2> vcc_io vgnd vpwr
+ / sky130_fd_io__com_ctl_ls
Xdm_ls<1> hld_i_h_n dm<1> dm_h<1> dm_h_n<1> dm_rst_h<1> dm_st_h<1> vcc_io vgnd vpwr
+ / sky130_fd_io__com_ctl_ls
Xtrip_sel_ls hld_i_h_n vtrip_sel vtrip_sel_h vtrip_sel_h_n trip_sel_rst_h trip_sel_st_h vcc_io vgnd
+ vpwr / sky130_fd_io__com_ctl_ls
Xinp_dis_ls hld_i_h_n inp_dis inp_dis_h inp_dis_h_n ie_n_rst_h ie_n_st_h vcc_io vgnd vpwr
+ / sky130_fd_io__com_ctl_ls
Xdm_ls<0> hld_i_h_n dm<0> dm_h<0> dm_h_n<0> dm_rst_h<0> dm_st_h<0> vcc_io vgnd vpwr
+ / sky130_fd_io__com_ctl_ls
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_ctl
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_ctl dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1>
+ dm_h_n<0> enable_h enable_inp_h hld_h_n hld_i_h hld_i_h_n hld_i_ovr_h hld_ovr ib_mode_sel
+ ib_mode_sel_h ib_mode_sel_h_n inp_dis inp_dis_h_n od_i_h vcc_io vgnd vpwr vtrip_sel vtrip_sel_h
+ vtrip_sel_h_n
*.PININFO dm<2>:I dm<1>:I dm<0>:I enable_h:I enable_inp_h:I hld_h_n:I
*.PININFO hld_ovr:I ib_mode_sel:I inp_dis:I vcc_io:I vgnd:I vpwr:I vtrip_sel:I
*.PININFO dm_h<2>:O dm_h<1>:O dm_h<0>:O dm_h_n<2>:O dm_h_n<1>:O dm_h_n<0>:O
*.PININFO hld_i_h:O hld_i_h_n:O hld_i_ovr_h:O ib_mode_sel_h:O
*.PININFO ib_mode_sel_h_n:O inp_dis_h_n:O od_i_h:O vtrip_sel_h:O
*.PININFO vtrip_sel_h_n:O
XI75 enable_inp_h enable_h startup_rst_h vgnd vcc_io / sky130_fd_io__hvsbt_nor
Xhld_dis_blk enable_h hld_h_n hld_i_h hld_i_h_n hld_i_ovr_h hld_ovr od_i_h vcc_io vgnd
+ vpwr / sky130_fd_io__gpiov2_ctl_hld
Xls_bank dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0>
+ hld_i_h_n ib_mode_sel ib_mode_sel_h ib_mode_sel_h_n inp_dis net80 inp_dis_h_n od_i_h
+ startup_rst_h inp_startup_en_h vcc_io vgnd vpwr vtrip_sel vtrip_sel_h vtrip_sel_h_n /
+ sky130_fd_io__gpiov2_ctl_lsbank
XI56 od_i_h enable_inp_h net92 vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI57 net92 inp_startup_en_h vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_inbuf_lvinv_x1
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_inbuf_lvinv_x1 in out vgnd vnb vpb vpwr
*.PININFO in:I vgnd:I vnb:I vpb:I vpwr:I out:O
XMI2 out in vgnd vnb sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.25) l=0.25 m=1*1 p=2*(1.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI1 out in vpwr vpb sky130_fd_pr__pfet_01v8_hvt AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.25) l=0.25 m=1*1 p=2*(3.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_ipath_lvls
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_ipath_lvls in_vcchib in_vddio mode_normal_lv mode_normal_lv_n mode_vcchib_lv
+ mode_vcchib_lv_n out out_b vcchib vssd
*.PININFO in_vcchib:I in_vddio:I mode_normal_lv:I mode_normal_lv_n:I
*.PININFO mode_vcchib_lv:I mode_vcchib_lv_n:I vcchib:I vssd:I out:O out_b:O
XMI336 out_b in_vcchib net50 vcchib sky130_fd_pr__pfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.25) l=0.25 m=2*1 p=2*(3.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI337 out out_b vcchib vcchib sky130_fd_pr__pfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.25) l=0.25 m=4*1 p=2*(3.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI338 fbk fbk_n vcchib vcchib sky130_fd_pr__pfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.25) l=0.25 m=1*1 p=2*(5.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI339 fbk_n mode_normal_lv vcchib vcchib sky130_fd_pr__pfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.25) l=0.25 m=1*1 p=2*(5.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI340 net50 mode_vcchib_lv_n vcchib vcchib sky130_fd_pr__pfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.25) l=0.25 m=2*1 p=2*(3.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI341 out_b mode_normal_lv net70 vcchib sky130_fd_pr__pfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.25) l=0.25 m=1*1 p=2*(3.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI342 net78 mode_normal_lv_n vcchib vcchib sky130_fd_pr__pfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.25) l=0.25 m=2*1 p=2*(3.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI343 out_b fbk net78 vcchib sky130_fd_pr__pfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.25) l=0.25 m=2*1 p=2*(3.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI344 net70 mode_vcchib_lv vcchib vcchib sky130_fd_pr__pfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.25) l=0.25 m=1*1 p=2*(3.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI345 fbk_n in_vddio vcchib vcchib sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=2*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI346 out_b in_vcchib net95 vssd sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.25) l=0.25 m=2*1 p=2*(3.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI347 net95 mode_vcchib_lv vssd vssd sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.25) l=0.25 m=2*1 p=2*(3.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI348 fbk fbk_n vssd vssd sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.25) l=0.25 m=1*1 p=2*(3.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI349 out out_b vssd vssd sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.25) l=0.25 m=2*1 p=2*(3.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI350 out_b fbk net111 vssd sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.25) l=0.25 m=2*1 p=2*(3.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI351 net111 mode_normal_lv vssd vssd sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.25) l=0.25 m=2*1 p=2*(3.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI352 net115 mode_normal_lv vssd vssd sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.25) l=0.25 m=1*1 p=2*(3.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI353 fbk_n in_vddio net115 vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_ipath_hvls
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_ipath_hvls in_vcchib in_vddio inb_vcchib mode_normal mode_normal_n
+ mode_vcchib mode_vcchib_n out out_b vddio_q vssd
*.PININFO in_vcchib:I in_vddio:I inb_vcchib:I mode_normal:I mode_normal_n:I
*.PININFO mode_vcchib:I mode_vcchib_n:I vddio_q:I vssd:I out:O out_b:O
XMI336 net84 fbk_b vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMI317 out_b net84 net55 vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=2*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI318 net55 mode_vcchib_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=2*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI319 out_b mode_vcchib net63 vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI320 out out_b vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=5*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI321 net75 mode_normal_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=2*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI322 out_b in_vddio net75 vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=2*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI323 net63 mode_normal vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI324 fbk_b fbk vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMI325 fbk fbk_b vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMI337 net84 fbk_b vssd vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.50)*(0.50) l=0.50 m=1*1 p=2*(1.50)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.50
XMI326 net88 mode_vcchib vssd vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI327 net92 mode_vcchib vssd vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=4*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI328 fbk mode_vcchib_n vssd vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI329 fbk_b in_vcchib net92 vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=3*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI330 out_b in_vddio net112 vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI331 out out_b vssd vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=3*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI332 net112 mode_normal vssd vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI333 net116 mode_vcchib vssd vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=4*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI334 fbk inb_vcchib net116 vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=3*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI335 out_b net84 net88 vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_vcchib_in_buf
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_vcchib_in_buf in_h mode_vcchib_lv_n out out_n vcchib vssd
*.PININFO in_h:I mode_vcchib_lv_n:I vcchib:I vssd:I out:O out_n:O
XMI552 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.80) l=0.80 m=1*1 p=2*(1.00)+2*(0.80) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI420 net57 in_b fbk vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.80) l=0.80 m=3*1 p=2*(1.00)+2*(0.80) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI541 net81 mode_vcchib_lv_n vssd vssd sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.25) l=0.25 m=2*1 p=2*(1.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI487 out out_n vssd vssd sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.25) l=0.25 m=3*1 p=2*(1.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI545 in_b in_h fbk vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.80) l=0.80 m=2*1 p=2*(5.00)+2*(0.80) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI423 out_n net81 vssd vssd sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.25) l=0.25 m=1*1 p=2*(1.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI424 net81 in_b vssd vssd sky130_fd_pr__nfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.25) l=0.25 m=2*1 p=2*(1.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI551 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.80) l=0.80 m=1*1 p=2*(5.00)+2*(0.80) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI544 fbk in_h vssd vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.80) l=0.80 m=2*1 p=2*(5.00)+2*(0.80) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI547 net108 mode_vcchib_lv_n vcchib vcchib sky130_fd_pr__pfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.25) l=0.25 m=3*1 p=2*(5.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI489 out out_n vcchib vcchib sky130_fd_pr__pfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.25) l=0.25 m=1*1 p=2*(5.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI538 net112 mode_vcchib_lv_n vcchib vcchib sky130_fd_pr__pfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.25) l=0.25 m=1*1 p=2*(3.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI429 out_n net81 vcchib vcchib sky130_fd_pr__pfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.25) l=0.25 m=1*1 p=2*(5.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI543 in_b in_h net108 vcchib sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.80) l=0.80 m=2*1 p=2*(5.00)+2*(0.80) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI436 net81 in_b net112 vcchib sky130_fd_pr__pfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.25) l=0.25 m=2*1 p=2*(1.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI549 net57 mode_vcchib_lv_n vcchib vcchib sky130_fd_pr__pfet_01v8 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.25) l=0.25 m=1*1 p=2*(5.00)+2*(0.25) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_in_buf
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_in_buf in_h in_vt mode_normal_n out out_n vddio_q vssd vtrip_sel_h
+ vtrip_sel_h_n
*.PININFO in_h:I in_vt:I mode_normal_n:I vddio_q:I vssd:I vtrip_sel_h:I
*.PININFO vtrip_sel_h_n:I out:O out_n:O
XI43 mode_normal_cmos_h mode_normal_cmos_h_n vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI488 vtrip_sel_h mode_normal_n mode_normal_cmos_h vssd vddio_q / sky130_fd_io__hvsbt_nor
XMI583 in_vt vtrip_sel_h_n vssd vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(1.00) l=1.00 m=1*1 p=2*(3.00)+2*(1.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI642 out out_n vssd vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI586 out_n net91 vssd vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI587 in_b in_h fbk vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.80) l=0.80 m=5*1 p=2*(5.00)+2*(0.80) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI588 fbk in_vt vssd vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.80) l=0.80 m=1*1 p=2*(5.00)+2*(0.80) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI589 net91 in_b vssd vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=2*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI590 fbk2 in_b fbk vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.80) l=0.80 m=4*1 p=2*(5.00)+2*(0.80) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI591 fbk in_h vssd vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.80) l=0.80 m=6*1 p=2*(5.00)+2*(0.80) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI592 net103 in_b fbk vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(1.00)*(0.80) l=0.80 m=4*1 p=2*(1.00)+2*(0.80) sa=265e-3 sb=265e-3
+ sd=280e-3 w=1.00
XMI593 net91 mode_normal_n vssd vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=2*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI646 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.80) l=0.80 m=1*1 p=2*(5.00)+2*(0.80) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI644 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.80) l=0.80 m=1*1 p=2*(5.00)+2*(0.80) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI643 out out_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI631 in_b in_h net122 vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.80) l=0.80 m=1*1 p=2*(5.00)+2*(0.80) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI595 net138 mode_normal_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI596 out_n net91 vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=1*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI597 fbk2 mode_normal_cmos_h_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=2*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI598 net91 in_b net138 vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(0.50) l=0.50 m=1*1 p=2*(3.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
XMI600 net103 mode_normal_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=2*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI647 vddio_q vddio_q vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.80) l=0.80 m=1*1 p=2*(5.00)+2*(0.80) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI632 net122 mode_normal_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=2*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI636 net158 mode_normal_cmos_h_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.50) l=0.50 m=2*1 p=2*(5.00)+2*(0.50) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
XMI629 in_b in_h net158 vddio_q sky130_fd_pr__pfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.00)*(0.80) l=0.80 m=1*1 p=2*(5.00)+2*(0.80) sa=265e-3 sb=265e-3
+ sd=280e-3 w=5.00
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_ibuf_se
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_ibuf_se enable_vddio_lv ibufmux_out ibufmux_out_h in_h in_vt mode_normal_n
+ mode_vcchib_n vcchib vddio_q vssd vtrip_sel_h vtrip_sel_h_n
*.PININFO enable_vddio_lv:I in_h:I in_vt:I mode_normal_n:I mode_vcchib_n:I
*.PININFO vcchib:I vddio_q:I vssd:I vtrip_sel_h:I vtrip_sel_h_n:I
*.PININFO ibufmux_out:O ibufmux_out_h:O
XI149 enable_vddio_lv mode_normal mode_normal_lv_n vssd vcchib / sky130_fd_io__hvsbt_nand2
XI148 enable_vddio_lv mode_vcchib mode_vcchib_lv_n vssd vcchib / sky130_fd_io__hvsbt_nand2
XI111 mode_vcchib_lv_n mode_vcchib_lv vssd vssd vcchib vcchib / sky130_fd_io__gpiov2_inbuf_lvinv_x1
XI112 mode_normal_lv_n mode_normal_lv vssd vssd vcchib vcchib / sky130_fd_io__gpiov2_inbuf_lvinv_x1
Xlvls out_vcchib out_vddio mode_normal_lv mode_normal_lv_n mode_vcchib_lv mode_vcchib_lv_n
+ ibufmux_out net57 vcchib vssd / sky130_fd_io__gpiov2_ipath_lvls
Xhvls out_vcchib out_vddio out_n_vcchib mode_normal mode_normal_n mode_vcchib mode_vcchib_n
+ ibufmux_out_h net68 vddio_q vssd / sky130_fd_io__gpiov2_ipath_hvls
XI88 in_h mode_vcchib_lv_n out_vcchib out_n_vcchib vcchib vssd / sky130_fd_io__gpiov2_vcchib_in_buf
Xbuf in_h in_vt mode_normal_n out_vddio out_n_vddio vddio_q vssd vtrip_sel_h vtrip_sel_h_n
+ / sky130_fd_io__gpiov2_in_buf
XI105 mode_vcchib_n mode_vcchib vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI491 mode_normal_n mode_normal vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_ictl_logic
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_ictl_logic dm_h_n<2> dm_h_n<1> dm_h_n<0> ib_mode_sel_h ib_mode_sel_h_n
+ inp_dis_h_n inp_dis_i_h inp_dis_i_h_n mode_normal_n mode_vcchib_n tripsel_i_h tripsel_i_h_n
+ vddio_q vssd vtrip_sel_h_n
*.PININFO dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I ib_mode_sel_h:I
*.PININFO ib_mode_sel_h_n:I inp_dis_h_n:I vddio_q:I vssd:I vtrip_sel_h_n:I
*.PININFO inp_dis_i_h:O inp_dis_i_h_n:O mode_normal_n:O mode_vcchib_n:O
*.PININFO tripsel_i_h:O tripsel_i_h_n:O
XI71 vtrip_sel_h_n mode_normal_n tripsel_i_h vssd vddio_q / sky130_fd_io__hvsbt_nor
XI35 inp_dis_i_h_n ib_mode_sel_h_n mode_normal_n vssd vddio_q / sky130_fd_io__hvsbt_nand2
XI36 inp_dis_i_h_n ib_mode_sel_h mode_vcchib_n vssd vddio_q / sky130_fd_io__hvsbt_nand2
XI78 dm_h_n<1> dm_h_n<0> nand_dm01 vssd vddio_q / sky130_fd_io__hvsbt_nand2
XI79 dm_h_n<2> and_dm01 dm_buf_dis_n vssd vddio_q / sky130_fd_io__hvsbt_nand2
XI80 dm_buf_dis_n inp_dis_h_n inp_dis_i_h vssd vddio_q / sky130_fd_io__hvsbt_nand2
XI74 tripsel_i_h tripsel_i_h_n vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI75 nand_dm01 and_dm01 vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI111 inp_dis_i_h inp_dis_i_h_n vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
.ENDS

************************************************************************
* Library Name: s8_esd
* Cell Name: s8_esd_signal_5_sym_hv_local_5term
* View Name: schematic
************************************************************************

.SUBCKT s8_esd_signal_5_sym_hv_local_5term gate in nbody nwellRing vgnd
*.PININFO gate:I in:B nbody:B nwellRing:B vgnd:B
XMI1 in gate vgnd nbody sky130_fd_pr__esd_nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(5.40)*(0.60) l=0.60 m=1*1 p=2*(5.40)+2*(0.60) sa=0.0 sb=0.0 sd=0.0
+ w=5.40
RI8 net16 nwellRing short m=1
RI9 net18 nbody short m=1
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpio_ovtv2_buf_localesd
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpio_ovtv2_buf_localesd in_h out_h out_vt vddio_q vssd vtrip_sel_h
*.PININFO in_h:I vtrip_sel_h:I out_h:O out_vt:O vddio_q:B vssd:B
XMhv_passgate out_h vtrip_sel_h out_vt vssd sky130_fd_pr__nfet_g5v0d10v5 AD=0 AS=0 PD=0 PS=0
+ a=(3.00)*(1.00) l=1.00 m=1*1 p=2*(3.00)+2*(1.00) sa=265e-3 sb=265e-3
+ sd=280e-3 w=3.00
Xesd_res in_h out_h / s8_esd_res250only_small
Xggnfet1 vssd out_h vssd vddio_q vssd / s8_esd_signal_5_sym_hv_local_5term
Xggnfet6 vssd vddio_q vssd vddio_q out_h / s8_esd_signal_5_sym_hv_local_5term
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__gpiov2_ipath
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__gpiov2_ipath dm_h_n<2> dm_h_n<1> dm_h_n<0> enable_vddio_lv ib_mode_sel_h
+ ib_mode_sel_h_n inp_dis_h_n out out_h pad vcchib vddio_q vssd vtrip_sel_h_n
*.PININFO dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I enable_vddio_lv:I
*.PININFO ib_mode_sel_h:I ib_mode_sel_h_n:I inp_dis_h_n:I vcchib:I vddio_q:I
*.PININFO vssd:I vtrip_sel_h_n:I out:O out_h:O pad:B
XI106 enable_vddio_lv out out_h in_h in_vt mode_normal_n mode_vcchib_n vcchib vddio_q
+ vssd tripsel_i_h tripsel_i_h_n / sky130_fd_io__gpiov2_ibuf_se
XI107 dm_h_n<2> dm_h_n<1> dm_h_n<0> ib_mode_sel_h ib_mode_sel_h_n inp_dis_h_n en_h_n en_h
+ mode_normal_n mode_vcchib_n tripsel_i_h tripsel_i_h_n vddio_q vssd vtrip_sel_h_n /
+ sky130_fd_io__gpiov2_ictl_logic
XI120 pad in_h in_vt vddio_q vssd tripsel_i_h / sky130_fd_io__gpio_ovtv2_buf_localesd
.ENDS

************************************************************************
* Library Name: s8iom0s8
* Cell Name: sky130_fd_io__top_gpiov2
* View Name: schematic
************************************************************************

.SUBCKT sky130_fd_io__top_gpiov2 amuxbus_a amuxbus_b analog_en analog_pol analog_sel dm[2] dm[1] dm[0]
+ enable_h enable_inp_h enable_vdda_h enable_vddio enable_vswitch_h hld_h_n hld_ovr ib_mode_sel in
+ in_h inp_dis oe_n out pad pad_a_esd_0_h pad_a_esd_1_h pad_a_noesd_h slow tie_hi_esd tie_lo_esd
+ vccd vcchib vdda vddio vddio_q vssa vssd vssio vssio_q vswitch vtrip_sel
*.PININFO analog_en:I analog_pol:I analog_sel:I dm[2]:I dm[1]:I dm[0]:I
*.PININFO enable_h:I enable_inp_h:I enable_vdda_h:I enable_vddio:I
*.PININFO enable_vswitch_h:I hld_h_n:I hld_ovr:I ib_mode_sel:I inp_dis:I
*.PININFO oe_n:I out:I slow:I vtrip_sel:I in:O in_h:O tie_hi_esd:O
*.PININFO tie_lo_esd:O amuxbus_a:B amuxbus_b:B pad:B pad_a_esd_0_h:B
*.PININFO pad_a_esd_1_h:B pad_a_noesd_h:B vccd:B vcchib:B vdda:B vddio:B
*.PININFO vddio_q:B vssa:B vssd:B vssio:B vssio_q:B vswitch:B
Xamux amuxbus_a amuxbus_b analog_en analog_pol analog_sel enable_vdda_h enable_vswitch_h hld_i_h
+ hld_i_h_n out pad vccd vdda vddio_q vssa vssd vssio_q vswitch /
+ sky130_fd_io__gpiov2_amux
Xopath dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n hld_i_ovr_h od_i_h
+ oe_n out pad slow tie_hi_esd tie_lo_esd vddio vssd vssio vccd vcchib
+ / sky130_fd_io__gpiov2_opath
Xctrl dm[2] dm[1] dm[0] dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0>
+ enable_h enable_inp_h hld_h_n hld_i_h hld_i_h_n hld_i_ovr_h hld_ovr ib_mode_sel ib_mode_sel_h
+ ib_mode_sel_h_n inp_dis inp_dis_h_n od_i_h vddio_q vssd vccd vtrip_sel vtrip_sel_h vtrip_sel_h_n
+ / sky130_fd_io__gpiov2_ctl
Xipath dm_h_n<2> dm_h_n<1> dm_h_n<0> enable_vddio ib_mode_sel_h ib_mode_sel_h_n inp_dis_h_n in in_h
+ pad vcchib vddio_q vssd vtrip_sel_h_n / sky130_fd_io__gpiov2_ipath
Xresd2 pad_a_esd_0_h net204 / s8_esd_res75only_small
Xresd4 net210 pad / s8_esd_res75only_small
Xresd1 net204 pad / s8_esd_res75only_small
Xresd3 pad_a_esd_1_h net210 / s8_esd_res75only_small
RS0<2> pad pad_a_noesd_h short m=1
RS0<1> pad pad_a_noesd_h short m=1
RS0<0> pad pad_a_noesd_h short m=1
.ENDS

.SUBCKT cad_dummy_open_device pin0 pin1
.ENDS cad_dummy_open_device
.SUBCKT condiode pin0 pin1
.ENDS condiode
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_02p4x04p6_m1m2_noshield C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB sky130_fd_pr__cap_vpp_02p4x04p6_m1m2_noshield
.ENDS sky130_fd_pr__cap_vpp_02p4x04p6_m1m2_noshield


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_02p7x06p1_m1m2m3m4_shieldl1_fingercap C0 C1 SUB Name= Formula= 2= 3= 4= 5= techLibCellName=-1
*.PININFO C0:? C1:? SUB:?
X1
.ENDS sky130_fd_pr__cap_vpp_02p7x06p1_m1m2m3m4_shieldl1_fingercap


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_02p7x11p1_m1m2m3m4_shieldl1_fingercap C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB
+ sky130_fd_pr__cap_vpp_02p7x11p1_m1m2m3m4_shieldl1_fingercap
.ENDS sky130_fd_pr__cap_vpp_02p7x11p1_m1m2m3m4_shieldl1_fingercap


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_02p7x21p1_m1m2m3m4_shieldl1_fingercap C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB
+ sky130_fd_pr__cap_vpp_02p7x21p1_m1m2m3m4_shieldl1_fingercap
.ENDS sky130_fd_pr__cap_vpp_02p7x21p1_m1m2m3m4_shieldl1_fingercap


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_02p7x41p1_m1m2m3m4_shieldl1_fingercap C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB
+ sky130_fd_pr__cap_vpp_02p7x41p1_m1m2m3m4_shieldl1_fingercap
.ENDS sky130_fd_pr__cap_vpp_02p7x41p1_m1m2m3m4_shieldl1_fingercap


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_02p9x06p1_m1m2m3m4_shieldl1_fingercap2 C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB
+ sky130_fd_pr__cap_vpp_02p9x06p1_m1m2m3m4_shieldl1_fingercap2
.ENDS sky130_fd_pr__cap_vpp_02p9x06p1_m1m2m3m4_shieldl1_fingercap2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_03p9x03p9_m1m2_shieldl1_floatm3 C0 C1 SUB MET3
*.PININFO C0:? C1:? SUB:? MET3:?
X1 C0 C1 SUB MET3
+ sky130_fd_pr__cap_vpp_03p9x03p9_m1m2_shieldl1_floatm3
.ENDS sky130_fd_pr__cap_vpp_03p9x03p9_m1m2_shieldl1_floatm3


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield
.ENDS sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield_o1 C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield_o1
.ENDS sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield_o1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_shieldpo_floatm3 C0 C1 SUB MET3
*.PININFO C0:? C1:? SUB:? MET3:?
X1 C0 C1 SUB MET3
+ sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_shieldpo_floatm3
.ENDS sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_shieldpo_floatm3


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield
.ENDS sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield_o2 C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield_o2
.ENDS sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield_o2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_shieldl1 C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_shieldl1
.ENDS sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_shieldl1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_04p4x04p6_m1m2m3_shieldl1 C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB sky130_fd_pr__cap_vpp_04p4x04p6_m1m2m3_shieldl1
.ENDS sky130_fd_pr__cap_vpp_04p4x04p6_m1m2m3_shieldl1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_04p4x04p6_m1m2m3_shieldl1m5_floatm4 C0 C1 MET5 SUB
*.PININFO C0:? C1:? MET5:? SUB:?
X1 C0 C1 SUB MET5
+ sky130_fd_pr__cap_vpp_04p4x04p6_m1m2m3_shieldl1m5_floatm4
.ENDS sky130_fd_pr__cap_vpp_04p4x04p6_m1m2m3_shieldl1m5_floatm4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_05p9x05p9_m1m2m3m4_shieldl1_wafflecap C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB
+ sky130_fd_pr__cap_vpp_05p9x05p9_m1m2m3m4_shieldl1_wafflecap
.ENDS sky130_fd_pr__cap_vpp_05p9x05p9_m1m2m3m4_shieldl1_wafflecap


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2m3_shieldpom4 C0 C1 MET4 SUB
*.PININFO C0:? C1:? MET4:? SUB:?
X1 C0 C1 SUB MET4 sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2m3_shieldpom4
.ENDS sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2m3_shieldpom4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_06p8x06p1_m1m2m3_shieldl1m4 C0 C1 MET4 SUB
*.PININFO C0:? C1:? MET4:? SUB:?
X1 C0 C1 SUB MET4 sky130_fd_pr__cap_vpp_06p8x06p1_m1m2m3_shieldl1m4
.ENDS sky130_fd_pr__cap_vpp_06p8x06p1_m1m2m3_shieldl1m4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield C0 C1 SUB MET3
*.PININFO C0:? C1:? SUB:? MET3:?
X1 C0 C1 SUB MET3 sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield
.ENDS sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield_o1 C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield_o1
.ENDS sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield_o1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3 C0 C1 SUB MET3
*.PININFO C0:? C1:? SUB:? MET3:?
X1 C0 C1 SUB MET3
+ sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3
.ENDS sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_noshield C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_noshield
.ENDS sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_noshield


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_shieldl1 C0 C1 SUB MET3
*.PININFO C0:? C1:? SUB:? MET3:?
X1 C0 C1 SUB MET3 sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_shieldl1
.ENDS sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_shieldl1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1 C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1
.ENDS sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1m5_floatm4 C0 C1 MET5 SUB
*.PININFO C0:? C1:? MET5:? SUB:?
X1 C0 C1 SUB MET5
+ sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1m5_floatm4
.ENDS sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1m5_floatm4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_11p3x11p3_m1m2m3m4_shieldl1_wafflecap C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB
+ sky130_fd_pr__cap_vpp_11p3x11p3_m1m2m3m4_shieldl1_wafflecap
.ENDS sky130_fd_pr__cap_vpp_11p3x11p3_m1m2m3m4_shieldl1_wafflecap


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_11p3x11p8_l1m1m2m3m4_shieldm5_nhv C0 C1 MET5
*.PININFO C0:? C1:? MET5:?
X1 C0 C1 C1 MET5
+ sky130_fd_pr__cap_vpp_11p3x11p8_l1m1m2m3m4_shieldm5_nhv
.ENDS sky130_fd_pr__cap_vpp_11p3x11p8_l1m1m2m3m4_shieldm5_nhv


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_noshield C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_noshield
.ENDS sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_noshield


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_shieldpom3 C0 C1 SUB MET3
*.PININFO C0:? C1:? SUB:? MET3:?
X1 C0 C1 SUB MET3 sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_shieldpom3
.ENDS sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_shieldpom3


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldm4 C0 C1 MET4 SUB
*.PININFO C0:? C1:? MET4:? SUB:?
X1 C0 C1 SUB MET4 sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldm4
.ENDS sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldm4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldpom4 C0 C1 MET4 SUB
*.PININFO C0:? C1:? MET4:? SUB:?
X1 C0 C1 SUB MET4 sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldpom4
.ENDS sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldpom4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldm5 C0 C1 MET5 SUB
*.PININFO C0:? C1:? MET5:? SUB:?
X1 C0 C1 SUB MET5 sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldm5
.ENDS sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldm5


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5 C0 C1 MET5 SUB
*.PININFO C0:? C1:? MET5:? SUB:?
X1 C0 C1 SUB MET5
+ sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5
.ENDS sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5_x C0 C1 MET5 SUB
*.PININFO C0:? C1:? MET5:? SUB:?
X1 C0 C1 SUB MET5
+ sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5_x
.ENDS sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5_x


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_noshield C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_noshield
.ENDS sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_noshield


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_shieldl1 C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_shieldl1
.ENDS sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_shieldl1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1 C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1
.ENDS sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1m5_floatm4 C0 C1 MET5 SUB
*.PININFO C0:? C1:? MET5:? SUB:?
X1 C0 C1 SUB MET5
+ sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1m5_floatm4
.ENDS sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1m5_floatm4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5 C0 C1 MET5 SUB
*.PININFO C0:? C1:? MET5:? SUB:?
X1 C0 C1 SUB MET5 sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5
.ENDS sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldm5 C0 C1 MET5 SUB
*.PININFO C0:? C1:? MET5:? SUB:?
X1 C0 C1 SUB MET5 sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldm5
.ENDS sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldm5


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_m1m4_noshield C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB sky130_fd_pr__cap_vpp_11p5x11p7_m1m4_noshield
.ENDS sky130_fd_pr__cap_vpp_11p5x11p7_m1m4_noshield


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__cap_vpp_44p7x23p1_pol1m1m2m3m4m5_noshield C0 C1 SUB
*.PININFO C0:? C1:? SUB:?
X1 C0 C1 SUB sky130_fd_pr__cap_vpp_44p7x23p1_pol1m1m2m3m4m5_noshield
.ENDS sky130_fd_pr__cap_vpp_44p7x23p1_pol1m1m2m3m4m5_noshield


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_aM02W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
.ENDS sky130_fd_pr__nfet_01v8_aM02W1p65L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_aM02W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
.ENDS sky130_fd_pr__nfet_01v8_aM02W1p65L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_aM02W1p65L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
.ENDS sky130_fd_pr__nfet_01v8_aM02W1p65L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_aM02W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__nfet_01v8_aM02W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_aM02W3p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
.ENDS sky130_fd_pr__nfet_01v8_aM02W3p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_aM02W3p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
.ENDS sky130_fd_pr__nfet_01v8_aM02W3p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_aM02W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__nfet_01v8_aM02W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_aM02W5p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
.ENDS sky130_fd_pr__nfet_01v8_aM02W5p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_aM02W5p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
.ENDS sky130_fd_pr__nfet_01v8_aM02W5p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_aM04W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
.ENDS sky130_fd_pr__nfet_01v8_aM04W1p65L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_aM04W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
.ENDS sky130_fd_pr__nfet_01v8_aM04W1p65L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_aM04W1p65L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
.ENDS sky130_fd_pr__nfet_01v8_aM04W1p65L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_aM04W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__nfet_01v8_aM04W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_aM04W3p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
.ENDS sky130_fd_pr__nfet_01v8_aM04W3p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_aM04W3p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
.ENDS sky130_fd_pr__nfet_01v8_aM04W3p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_aM04W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__nfet_01v8_aM04W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_aM04W5p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
.ENDS sky130_fd_pr__nfet_01v8_aM04W5p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_aM04W5p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
.ENDS sky130_fd_pr__nfet_01v8_aM04W5p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_hcM04W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__nfet_01v8_hcM04W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_hcM04W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__nfet_01v8_hcM04W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_lvt_aM02W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
.ENDS sky130_fd_pr__nfet_01v8_lvt_aM02W1p65L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_lvt_aM02W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
.ENDS sky130_fd_pr__nfet_01v8_lvt_aM02W1p65L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_lvt_aM02W1p65L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
.ENDS sky130_fd_pr__nfet_01v8_lvt_aM02W1p65L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_lvt_aM02W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__nfet_01v8_lvt_aM02W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_lvt_aM02W3p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
.ENDS sky130_fd_pr__nfet_01v8_lvt_aM02W3p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_lvt_aM02W3p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
.ENDS sky130_fd_pr__nfet_01v8_lvt_aM02W3p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_lvt_aM02W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__nfet_01v8_lvt_aM02W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_lvt_aM02W5p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
.ENDS sky130_fd_pr__nfet_01v8_lvt_aM02W5p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_lvt_aM02W5p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
.ENDS sky130_fd_pr__nfet_01v8_lvt_aM02W5p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_lvt_aM04W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
.ENDS sky130_fd_pr__nfet_01v8_lvt_aM04W1p65L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_lvt_aM04W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
.ENDS sky130_fd_pr__nfet_01v8_lvt_aM04W1p65L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_lvt_aM04W1p65L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
.ENDS sky130_fd_pr__nfet_01v8_lvt_aM04W1p65L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_lvt_aM04W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__nfet_01v8_lvt_aM04W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_lvt_aM04W3p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
.ENDS sky130_fd_pr__nfet_01v8_lvt_aM04W3p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_lvt_aM04W3p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
.ENDS sky130_fd_pr__nfet_01v8_lvt_aM04W3p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_lvt_aM04W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__nfet_01v8_lvt_aM04W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_lvt_aM04W5p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
.ENDS sky130_fd_pr__nfet_01v8_lvt_aM04W5p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_lvt_aM04W5p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
.ENDS sky130_fd_pr__nfet_01v8_lvt_aM04W5p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_lvt_bM02W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM3 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
XM4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
.ENDS sky130_fd_pr__nfet_01v8_lvt_bM02W1p65L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_mcM04W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__nfet_01v8_mcM04W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_01v8_mcM04W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__nfet_01v8_mcM04W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_g5v0d10v5_aM04W3p00L0p50 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
.ENDS sky130_fd_pr__nfet_g5v0d10v5_aM04W3p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_g5v0d10v5_aM04W5p00L0p50 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
.ENDS sky130_fd_pr__nfet_g5v0d10v5_aM04W5p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_g5v0d10v5_aM04W7p00L0p50 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
.ENDS sky130_fd_pr__nfet_g5v0d10v5_aM04W7p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_g5v0d10v5_aM10W3p00L0p50 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM5 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM6 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM7 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM8 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM9 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM10 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
.ENDS sky130_fd_pr__nfet_g5v0d10v5_aM10W3p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_g5v0d10v5_aM10W5p00L0p50 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM5 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM6 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM7 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM8 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM9 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM10 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
.ENDS sky130_fd_pr__nfet_g5v0d10v5_aM10W5p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__nfet_g5v0d10v5_aM10W7p00L0p50 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM5 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM6 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM7 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM8 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM9 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM10 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
.ENDS sky130_fd_pr__nfet_g5v0d10v5_aM10W7p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_aM02W1p65L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.15 m=1
.ENDS sky130_fd_pr__pfet_01v8_aM02W1p65L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_aM02W1p65L0p18 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.18 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.18 m=1
.ENDS sky130_fd_pr__pfet_01v8_aM02W1p65L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_aM02W1p65L0p25 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.25 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.25 m=1
.ENDS sky130_fd_pr__pfet_01v8_aM02W1p65L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_aM02W3p00L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__pfet_01v8_aM02W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_aM02W3p00L0p18 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.18 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.18 m=1
.ENDS sky130_fd_pr__pfet_01v8_aM02W3p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_aM02W3p00L0p25 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.25 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.25 m=1
.ENDS sky130_fd_pr__pfet_01v8_aM02W3p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_aM02W5p00L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__pfet_01v8_aM02W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_aM02W5p00L0p18 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.18 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.18 m=1
.ENDS sky130_fd_pr__pfet_01v8_aM02W5p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_aM02W5p00L0p25 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.25 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.25 m=1
.ENDS sky130_fd_pr__pfet_01v8_aM02W5p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_aM04W1p65L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.15 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.15 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.15 m=1
.ENDS sky130_fd_pr__pfet_01v8_aM04W1p65L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_aM04W1p65L0p18 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.18 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.18 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.18 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.18 m=1
.ENDS sky130_fd_pr__pfet_01v8_aM04W1p65L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_aM04W1p65L0p25 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.25 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.25 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.25 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.25 m=1
.ENDS sky130_fd_pr__pfet_01v8_aM04W1p65L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_aM04W3p00L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__pfet_01v8_aM04W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_aM04W3p00L0p18 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.18 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.18 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.18 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.18 m=1
.ENDS sky130_fd_pr__pfet_01v8_aM04W3p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_aM04W3p00L0p25 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.25 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.25 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.25 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.25 m=1
.ENDS sky130_fd_pr__pfet_01v8_aM04W3p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_aM04W5p00L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__pfet_01v8_aM04W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_aM04W5p00L0p18 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.18 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.18 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.18 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.18 m=1
.ENDS sky130_fd_pr__pfet_01v8_aM04W5p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_aM04W5p00L0p25 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.25 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.25 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.25 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.25 m=1
.ENDS sky130_fd_pr__pfet_01v8_aM04W5p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_hcM04W3p00L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__pfet_01v8_hcM04W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_hcM04W5p00L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__pfet_01v8_hcM04W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_lvt_aM02W3p00L0p35 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.35 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.35 m=1
.ENDS sky130_fd_pr__pfet_01v8_lvt_aM02W3p00L0p35


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_lvt_aM02W3p00L0p50 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.5 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.5 m=1
.ENDS sky130_fd_pr__pfet_01v8_lvt_aM02W3p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_lvt_aM02W5p00L0p35 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.35 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.35 m=1
.ENDS sky130_fd_pr__pfet_01v8_lvt_aM02W5p00L0p35


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_lvt_aM02W5p00L0p50 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.5 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.5 m=1
.ENDS sky130_fd_pr__pfet_01v8_lvt_aM02W5p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_lvt_aM04W3p00L0p35 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.35 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.35 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.35 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.35 m=1
.ENDS sky130_fd_pr__pfet_01v8_lvt_aM04W3p00L0p35


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_lvt_aM04W3p00L0p50 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.5 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.5 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.5 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.5 m=1
.ENDS sky130_fd_pr__pfet_01v8_lvt_aM04W3p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_lvt_aM04W5p00L0p35 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.35 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.35 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.35 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.35 m=1
.ENDS sky130_fd_pr__pfet_01v8_lvt_aM04W5p00L0p35


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_lvt_aM04W5p00L0p50 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.5 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.5 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.5 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.5 m=1
.ENDS sky130_fd_pr__pfet_01v8_lvt_aM04W5p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_mcM04W3p00L0p15 DRAIN GATE SOURCE BULK
*.PININFO DRAIN:? GATE:? SOURCE:? BULK:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__pfet_01v8_mcM04W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_mcM04W5p00L0p15 DRAIN GATE SOURCE BULK
*.PININFO DRAIN:? GATE:? SOURCE:? BULK:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__pfet_01v8_mcM04W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_aM02W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_aM02W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_aM02W3p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_aM02W3p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_aM02W3p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_aM02W3p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_aM04W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_aM04W1p65L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_aM04W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_aM04W1p65L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_aM04W1p65L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_aM04W1p65L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_aM04W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_aM04W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_aM04W3p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_aM04W3p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_aM04W3p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_aM04W3p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM3 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
XM4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM3 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
XM4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM3 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
XM4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM3 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
XM4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM3 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
XM4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM3 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
XM4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM3 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
XM4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM3 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
XM4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM3 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
XM4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM5 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
XM6 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM5 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
XM6 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM5 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
XM6 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM5 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
XM6 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM5 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
XM6 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM5 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
XM6 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM5 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
XM6 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM5 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
XM6 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM5 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
XM6 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_hcM04W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_hcM04W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_hcM04W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_hcM04W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=0.42 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=0.42 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p84L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=0.84 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=0.84 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p84L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aF02W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.0 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.0 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aF02W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aF04W0p84L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=0.84 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=0.84 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=0.84 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=0.84 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aF04W0p84L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aF04W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.0 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.0 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.0 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.0 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aF04W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aF08W0p84L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=0.84 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=0.84 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=0.84 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=0.84 l=0.15 m=1
XM5 DRAIN GATE SOURCE SUBSTRATE model_use_only w=0.84 l=0.15 m=1
XM6 DRAIN GATE SOURCE SUBSTRATE model_use_only w=0.84 l=0.15 m=1
XM7 DRAIN GATE SOURCE SUBSTRATE model_use_only w=0.84 l=0.15 m=1
XM8 DRAIN GATE SOURCE SUBSTRATE model_use_only w=0.84 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aF08W0p84L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.0 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.0 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.0 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.0 l=0.15 m=1
XM5 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.0 l=0.15 m=1
XM6 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.0 l=0.15 m=1
XM7 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.0 l=0.15 m=1
XM8 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.0 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aM02W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aM02W1p65L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aM02W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aM02W1p65L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aM02W1p65L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aM02W1p65L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aM02W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aM02W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aM02W3p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aM02W3p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aM02W3p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aM02W3p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aM02W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aM02W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aM02W5p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aM02W5p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aM02W5p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aM02W5p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aM04W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aM04W1p65L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aM04W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aM04W1p65L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aM04W1p65L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aM04W1p65L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aM04W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aM04W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aM04W3p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aM04W3p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aM04W3p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aM04W3p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aM04W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aM04W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aM04W5p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aM04W5p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_aM04W5p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_aM04W5p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_bM02W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM3 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
XM4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_bM02W1p65L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_bM02W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM3 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
XM4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_bM02W1p65L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_bM02W1p65L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM3 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
XM4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_bM02W1p65L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_bM02W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM3 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
XM4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_bM02W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_bM02W3p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM3 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
XM4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_bM02W3p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_bM02W3p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM3 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
XM4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_bM02W3p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_bM02W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM3 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
XM4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_bM02W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_bM02W5p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM3 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
XM4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_bM02W5p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_bM02W5p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM3 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
XM4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_bM02W5p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_bM04W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15 m=1
XM5 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
XM6 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_bM04W1p65L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_bM04W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.18 m=1
XM5 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
XM6 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_bM04W1p65L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_bM04W1p65L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.25 m=1
XM5 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
XM6 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=1.65 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_bM04W1p65L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_bM04W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM5 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
XM6 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_bM04W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_bM04W3p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.18 m=1
XM5 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
XM6 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_bM04W3p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_bM04W3p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.25 m=1
XM5 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
XM6 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_bM04W3p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_bM04W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM5 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
XM6 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_bM04W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_bM04W5p00L0p18 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.18 m=1
XM5 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
XM6 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_bM04W5p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_lvt_bM04W5p00L0p25 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.25 m=1
XM5 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
XM6 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15
+ m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_lvt_bM04W5p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_mcM04W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_mcM04W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_01v8_mcM04W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__rf_nfet_01v8_mcM04W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_aM04W3p00L0p50 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_aM04W3p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_aM04W5p00L0p50 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_aM04W5p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_aM04W7p00L0p50 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_aM04W7p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W3p00L0p50 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM5 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM6 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM7 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM8 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM9 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM10 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W3p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W5p00L0p50 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM5 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM6 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM7 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM8 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM9 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM10 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W5p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W7p00L0p50 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM5 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM6 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM7 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM8 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM9 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM10 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W7p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_bM02W3p00L0p50 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM3 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5
+ m=1
XM4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5
+ m=1
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_bM02W3p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_bM02W5p00L0p50 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM3 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5
+ m=1
XM4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5
+ m=1
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_bM02W5p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W3p00L0p50 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM5 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5
+ m=1
XM6 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5
+ m=1
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W3p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W5p00L0p50 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM5 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5
+ m=1
XM6 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5
+ m=1
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W5p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W7p00L0p50 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM5 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5
+ m=1
XM6 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5
+ m=1
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W7p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W3p00L0p50 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM5 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM6 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM7 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM8 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM9 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM10 DRAIN GATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5 m=1
XM11 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5
+ m=1
XM12 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=3.01 l=0.5
+ m=1
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W3p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W5p00L0p50 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM5 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM6 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM7 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM8 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM9 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM10 DRAIN GATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5 m=1
XM11 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5
+ m=1
XM12 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=5.05 l=0.5
+ m=1
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W5p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W7p00L0p50 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
XM1 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM2 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM3 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM4 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM5 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM6 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM7 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM8 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM9 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM10 DRAIN GATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
XM11 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5
+ m=1
XM12 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE model_use_only w=7.09 l=0.5
+ m=1
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W7p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=0.84 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=0.84 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aF02W1p68L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=1.68 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=1.68 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aF02W1p68L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aF02W3p00L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.0 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.0 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aF02W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.0 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.0 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=1.68 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=1.68 l=0.15 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=1.68 l=0.15 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=1.68 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aM02W1p65L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aM02W1p65L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aM02W1p65L0p18 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.18 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.18 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aM02W1p65L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aM02W1p65L0p25 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.25 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.25 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aM02W1p65L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aM02W3p00L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aM02W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aM02W3p00L0p18 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.18 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.18 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aM02W3p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aM02W3p00L0p25 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.25 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.25 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aM02W3p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aM02W5p00L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aM02W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aM02W5p00L0p18 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.18 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.18 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aM02W5p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aM02W5p00L0p25 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.25 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.25 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aM02W5p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aM04W1p65L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.15 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.15 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aM04W1p65L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aM04W1p65L0p18 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.18 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.18 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.18 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.18 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aM04W1p65L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aM04W1p65L0p25 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.25 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.25 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.25 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.25 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aM04W1p65L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aM04W3p00L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aM04W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aM04W3p00L0p18 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.18 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.18 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.18 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.18 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aM04W3p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aM04W3p00L0p25 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.25 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.25 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.25 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.25 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aM04W3p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p18 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.18 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.18 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.18 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.18 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p25 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.25 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.25 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.25 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.25 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.15 m=1
XM3 BULK BULK SOURCE BULK model_use_only w=1.65 l=0.15 m=1
XM4 BULK BULK SOURCE BULK model_use_only w=1.65 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p18 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.18 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.18 m=1
XM3 BULK BULK SOURCE BULK model_use_only w=1.65 l=0.15 m=1
XM4 BULK BULK SOURCE BULK model_use_only w=1.65 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p25 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.25 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.25 m=1
XM3 BULK BULK SOURCE BULK model_use_only w=1.65 l=0.15 m=1
XM4 BULK BULK SOURCE BULK model_use_only w=1.65 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM3 BULK BULK SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM4 BULK BULK SOURCE BULK model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p18 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.18 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.18 m=1
XM3 BULK BULK SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM4 BULK BULK SOURCE BULK model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p25 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.25 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.25 m=1
XM3 BULK BULK SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM4 BULK BULK SOURCE BULK model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM3 BULK BULK SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM4 BULK BULK SOURCE BULK model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p18 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.18 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.18 m=1
XM3 BULK BULK SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM4 BULK BULK SOURCE BULK model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p25 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.25 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.25 m=1
XM3 BULK BULK SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM4 BULK BULK SOURCE BULK model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.15 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.15 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.15 m=1
XM5 BULK BULK SOURCE BULK model_use_only w=1.65 l=0.15 m=1
XM6 BULK BULK SOURCE BULK model_use_only w=1.65 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p18 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.18 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.18 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.18 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.18 m=1
XM5 BULK BULK SOURCE BULK model_use_only w=1.65 l=0.15 m=1
XM6 BULK BULK SOURCE BULK model_use_only w=1.65 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p25 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.25 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.25 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.25 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=1.65 l=0.25 m=1
XM5 BULK BULK SOURCE BULK model_use_only w=1.65 l=0.15 m=1
XM6 BULK BULK SOURCE BULK model_use_only w=1.65 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM5 BULK BULK SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM6 BULK BULK SOURCE BULK model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p18 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.18 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.18 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.18 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.18 m=1
XM5 BULK BULK SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM6 BULK BULK SOURCE BULK model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p25 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.25 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.25 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.25 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.25 m=1
XM5 BULK BULK SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM6 BULK BULK SOURCE BULK model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM5 BULK BULK SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM6 BULK BULK SOURCE BULK model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p18 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.18 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.18 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.18 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.18 m=1
XM5 BULK BULK SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM6 BULK BULK SOURCE BULK model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p18


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p25 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.25 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.25 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.25 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.25 m=1
XM5 BULK BULK SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM6 BULK BULK SOURCE BULK model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p25


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_hcM04W3p00L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_hcM04W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_hcM04W5p00L0p15 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_hcM04W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_lvt_aM02W3p00L0p35 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.35 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.35 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_lvt_aM02W3p00L0p35


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_lvt_aM02W3p00L0p50 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.5 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.5 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_lvt_aM02W3p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_lvt_aM02W5p00L0p35 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.35 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.35 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_lvt_aM02W5p00L0p35


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_lvt_aM02W5p00L0p50 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.5 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.5 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_lvt_aM02W5p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_lvt_aM04W3p00L0p35 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.35 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.35 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.35 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.35 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_lvt_aM04W3p00L0p35


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_lvt_aM04W3p00L0p50 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.5 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.5 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.5 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.5 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_lvt_aM04W3p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_lvt_aM04W5p00L0p35 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.35 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.35 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.35 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.35 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_lvt_aM04W5p00L0p35


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_lvt_aM04W5p00L0p50 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.5 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.5 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.5 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.5 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_lvt_aM04W5p00L0p50


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_mcM04W3p00L0p15 DRAIN GATE SOURCE BULK
*.PININFO DRAIN:? GATE:? SOURCE:? BULK:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=3.01 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_mcM04W3p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_mcM04W5p00L0p15 DRAIN GATE SOURCE BULK
*.PININFO DRAIN:? GATE:? SOURCE:? BULK:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM3 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
XM4 DRAIN GATE SOURCE BULK model_use_only w=5.05 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_mcM04W5p00L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_pfet_01v8_mvt_aF02W0p84L0p15 BULK DRAIN GATE SOURCE Name= Formula= techLibCellName=-1 nd= ng= ns= nb= mname= w= l= m=
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
XM1 DRAIN GATE SOURCE BULK model_use_only w=0.84 l=0.15 m=1
XM2 DRAIN GATE SOURCE BULK model_use_only w=0.84 l=0.15 m=1
.ENDS sky130_fd_pr__rf_pfet_01v8_mvt_aF02W0p84L0p15


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__bufbuf_8 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 Abb Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 Abbb Abb VGND VNB sky130_fd_pr__nfet_01v8 m=3 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN4 X Abbb VGND VNB sky130_fd_pr__nfet_01v8 m=8 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP4 X Abbb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 Abb Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 Abbb Abb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=3 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__bufbuf_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__bufbuf_16 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 Abb Ab VGND VNB sky130_fd_pr__nfet_01v8 m=3 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 Abbb Abb VGND VNB sky130_fd_pr__nfet_01v8 m=6 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN4 X Abbb VGND VNB sky130_fd_pr__nfet_01v8 m=16 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP4 X Abbb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=16 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 Abb Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=3 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 Abbb Abb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=6 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__bufbuf_16


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 pndB VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o311ai_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o311ai_0 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 pndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o311ai_0


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 pndB VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o311ai_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 pndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o311ai_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dfsbp_2 CLK D SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
XMXNI36 net128 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI39 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 M1 M0 net111 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net79 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 S0 clkpos net128 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI25 net96 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI26 S0 clkneg net88 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI27 net88 S1 net96 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 M0 clkpos net79 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net111 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 net140 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net140 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI49 Q_N S0 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI40 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI38 S0 clkneg net191 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI37 net191 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M1 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net168 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 M0 clkneg net168 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 net155 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 S0 clkpos net155 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 S0 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 net140 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net140 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI50 Q_N S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dfsbp_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dfsbp_1 CLK D SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
XMXNI36 net129 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI39 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 M1 M0 net112 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net80 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 S0 clkpos net129 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI25 net97 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI26 S0 clkneg net89 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI27 net89 S1 net97 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 M0 clkpos net80 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net112 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 net141 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net141 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI49 Q_N S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI40 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI38 S0 clkneg net192 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI37 net192 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M1 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net169 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 M0 clkneg net169 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 net156 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 S0 clkpos net156 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 S0 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 net141 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net141 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI50 Q_N S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dfsbp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net82 s0 net108 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net108 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 net101 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 M0 clkpos net93 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 net93 M1 net101 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 s0 clkneg net81 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net82 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net81 net82 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI39 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 M1 clkpos s0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net165 net82 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 net82 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 s0 clkpos net165 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net82 s0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI30 net144 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI31 M0 clkneg net144 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI32 net144 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net82 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI40 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 M1 clkneg s0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dfrtp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net82 s0 net108 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net108 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 net101 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 M0 clkpos net93 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 net93 M1 net101 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 s0 clkneg net81 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net82 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net81 net82 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI39 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 M1 clkpos s0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net165 net82 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 net82 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 s0 clkpos net165 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net82 s0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI30 net144 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI31 M0 clkneg net144 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI32 net144 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net82 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI40 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 M1 clkneg s0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dfrtp_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net82 s0 net108 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net108 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 net101 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 M0 clkpos net93 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 net93 M1 net101 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 s0 clkneg net81 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net82 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net81 net82 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI39 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 M1 clkpos s0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net156 net82 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 net82 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 s0 clkpos net156 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net82 s0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI30 net144 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI31 M0 clkneg net144 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI32 net144 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net82 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI40 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 M1 clkneg s0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dfrtp_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sedfxtp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I DE:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI14 net146 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI13 S0 clkneg net146 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 Q S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net114 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI643 net118 q1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI639 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.75 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 S0 clkpos net118 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M0 clkneg net114 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 q1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 net94 deneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 net98 sceneg db VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 VPWR SCD net98 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI31 net95 D net94 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 net95 SCE db VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI40 net87 q1 net95 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI36 deneg DE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI38 VPWR DE net87 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 sceneg SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI641 net222 q1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 S0 clkneg net222 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 Q S0 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net211 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 M0 clkpos net211 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 net95 sceneg db VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 q1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 sceneg SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI32 net95 D net167 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI16 net187 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI15 S0 clkpos net187 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI41 net174 q1 net95 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI39 VGND deneg net174 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI37 deneg DE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 net167 DE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI49 net158 SCE db VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI48 VGND SCD net158 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sedfxtp_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sedfxtp_4 CLK D DE SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I DE:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI14 net146 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI13 S0 clkneg net146 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 Q S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net135 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI643 net118 q1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI639 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.75 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 S0 clkpos net118 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M0 clkneg net135 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 q1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 net107 deneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 net98 sceneg db VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 VPWR SCD net98 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI31 net95 D net107 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 net95 SCE db VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI40 net87 q1 net95 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI36 deneg DE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI38 VPWR DE net87 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 sceneg SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI641 net227 q1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 S0 clkneg net227 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 Q S0 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net206 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 M0 clkpos net206 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 net95 sceneg db VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 q1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 sceneg SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI32 net95 D net190 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI16 net187 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI15 S0 clkpos net187 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI41 net174 q1 net95 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI39 VGND deneg net174 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI37 deneg DE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 net190 DE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI49 net163 SCE db VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI48 VGND SCD net163 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sedfxtp_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sedfxtp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I DE:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI14 net146 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI13 S0 clkneg net146 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 Q S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net114 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI643 net118 q1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI639 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.75 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 S0 clkpos net118 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M0 clkneg net114 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 q1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 net94 deneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 net103 sceneg db VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 VPWR SCD net103 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI31 net95 D net94 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 net95 SCE db VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI40 net87 q1 net95 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI36 deneg DE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI38 VPWR DE net87 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 sceneg SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI641 net222 q1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 S0 clkneg net222 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 Q S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net211 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 M0 clkpos net211 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 net95 sceneg db VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 q1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 sceneg SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI32 net95 D net167 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI16 net187 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI15 S0 clkpos net187 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI41 net179 q1 net95 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI39 VGND deneg net179 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI37 deneg DE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 net167 DE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI49 net158 SCE db VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI48 VGND SCD net158 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sedfxtp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__fahcon_1 A B CI VGND VNB VPB VPWR COUT_N SUM
*.PININFO A:I B:I CI:I VGND:I VNB:I VPB:I VPWR:I COUT_N:O SUM:O
XMXNMIP3 SUM net146 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI32 Bb2 B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI27 Ab Bb1 mid2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI26 Abb B mid2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI22 Abb Bb1 mid1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI23 Ab B mid1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 CIb1 CI VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI13 CIbb2 CIb2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 Abb Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI12 CIb2 CI VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI16 Bb1 B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 CIb2 mid2 net146 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI1 CIbb2 mid1 net146 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI3 Bb2 mid2 COUT_N VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 CIb1 mid1 COUT_N VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 SUM net146 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 CIb1 mid2 COUT_N VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI25 Ab B mid2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 Abb Bb1 mid2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI21 Ab Bb1 mid1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 Abb B mid1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI14 CIb1 CI VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI9 CIbb2 CIb2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI8 CIb2 CI VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 Abb Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 Bb1 B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 CIb2 mid1 net146 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI2 CIbb2 mid2 net146 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI31 Bb2 mid1 COUT_N VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 Bb2 B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__fahcon_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
*.PININFO DIODE:I VGND:I VNB:I VPB:I VPWR:I
XD0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 AREA=0.4347 m=1
.ENDS sky130_fd_sc_hd__diode_2

******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C sndC VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN3 sndC D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand4_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C sndC VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN3 sndC D VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand4_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C sndC VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN3 sndC D VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand4_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMIP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.25 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 net36 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.55 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 Y A net36 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.55 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__clkinvlp_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMIP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.25 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 Y A net31 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.55 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 net35 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.55 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 net31 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.55 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 Y A net35 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.55 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__clkinvlp_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
*.PININFO A:I B:I C_N:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 C C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 y C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN2 C C_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or3b_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
*.PININFO A:I B:I C_N:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 C C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 y C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN2 C C_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or3b_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
*.PININFO A:I B:I C_N:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 C C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 y C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN2 C C_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or3b_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMNnand0 VGND A1_N sndNA1N VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnand1 sndNA1N A2_N inand VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi10 nmid B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi11 nmid B2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi20 Y inand nmid VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand0 inand A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand1 inand A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi10 VPWR B1 sndPB1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi11 sndPB1 B2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi20 Y inand VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o2bb2ai_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMNnand0 VGND A1_N sndNA1N VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnand1 sndNA1N A2_N inand VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi10 nmid B1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi11 nmid B2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi20 Y inand nmid VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand0 inand A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand1 inand A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi10 VPWR B1 sndPB1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi11 sndPB1 B2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi20 Y inand VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o2bb2ai_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMNnand0 VGND A1_N sndNA1N VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnand1 sndNA1N A2_N inand VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi10 nmid B1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi11 nmid B2 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi20 Y inand nmid VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand0 inand A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand1 inand A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi10 VPWR B1 sndPB1 VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi11 sndPB1 B2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi20 Y inand VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o2bb2ai_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 sndA3 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA3 sndA3 A4 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA3 pndA A4 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o41ai_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 sndA3 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA3 sndA3 A4 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA3 pndA A4 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o41ai_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 sndA3 VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA3 sndA3 A4 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA3 pndA A4 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o41ai_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_inputiso1p_1 A SLEEP VGND VNB VPB VPWR X
*.PININFO A:I SLEEP:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR SLEEP sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 sndPA A net36 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI15 VPWR net36 X VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI10 net36 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI16 net36 SLEEP VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI14 X net36 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_inputiso1p_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__clkdlybuf4s25_2 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 A2 Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.25 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 Ab2 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.25 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 X Ab2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 A2 Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.82 l=0.25 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 Ab2 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.82 l=0.25 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 X Ab2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__clkdlybuf4s25_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 A2 Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.25 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 Ab2 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.25 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 X Ab2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 A2 Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.82 l=0.25 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 Ab2 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.82 l=0.25 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 X Ab2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__clkdlybuf4s25_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 Y C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a311oi_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 Y C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a311oi_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 Y C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a311oi_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdfbbn_2 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK_N:I D:I RESET_B:I SCD:I SCE:I SET_B:I VGND:I VNB:I VPB:I
*.PININFO VPWR:I Q:O Q_N:O
XMXNI98 net105 D n0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI103 n1 SCD VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI104 n0 sceb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI120 net105 SCE n1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI46 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 RESET RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI676 M1 M0 net176 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI675 net176 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net213 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI677 M1 RESET net176 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 M0 clkpos net160 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkpos CLK_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 net160 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 S0 clkneg net145 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net145 net117 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 Q_N net117 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 net213 net117 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 net105 clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI668 S0 clkpos net128 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI667 net128 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI630 net117 RESET net116 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI3 net117 S0 net116 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 net116 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI639 sceb SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI94 net105 D p0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI101 net105 sceb p1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI679 M1 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI669 S0 clkneg net265 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net213 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI9 net117 S0 net268 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI670 net265 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI678 net216 RESET VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net257 net117 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 S0 clkpos net257 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI10 net117 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI11 net268 RESET VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 net241 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 net105 clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 M0 clkneg net241 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI643 RESET RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkpos CLK_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI680 M1 M0 net216 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 net213 net117 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI661 Q_N net117 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI640 sceb SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sdfbbn_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdfbbn_1 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK_N:I D:I RESET_B:I SCD:I SCE:I SET_B:I VGND:I VNB:I VPB:I
*.PININFO VPWR:I Q:O Q_N:O
XMXNI98 net105 D n0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI103 n1 SCD VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI104 n0 sceb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI120 net105 SCE n1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI46 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 RESET RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI676 M1 M0 net176 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI675 net176 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net213 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI677 M1 RESET net176 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 M0 clkpos net153 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkpos CLK_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 net153 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 S0 clkneg net145 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net145 net117 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 Q_N net117 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 net213 net117 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 net105 clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI668 S0 clkpos net125 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI667 net125 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI630 net117 RESET net116 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI3 net117 S0 net116 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 net116 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI639 sceb SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI94 net105 D p0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI101 net105 sceb p1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI679 M1 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI669 S0 clkneg net265 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net213 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI9 net117 S0 net268 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI670 net265 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI678 net216 RESET VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net257 net117 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 S0 clkpos net257 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI10 net117 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI11 net268 RESET VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 net241 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 net105 clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 M0 clkneg net241 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI643 RESET RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkpos CLK_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI680 M1 M0 net216 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 net213 net117 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI661 Q_N net117 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI640 sceb SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sdfbbn_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__clkdlybuf4s15_2 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 A2 Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 Ab2 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 X Ab2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 A2 Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.82 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 Ab2 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.82 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 X Ab2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__clkdlybuf4s15_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__clkdlybuf4s15_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 A2 Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 Ab2 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 X Ab2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 A2 Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.82 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 Ab2 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.82 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 X Ab2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__clkdlybuf4s15_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN0 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=16 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 X Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=16 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__clkbuf_16


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN0 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.52 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.52 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.79 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 X Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.79 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__clkbuf_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN0 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=8 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 X Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__clkbuf_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN0 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 X Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__clkbuf_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN0 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 X Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__clkbuf_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_inputiso1n_1 A SLEEP_B VGND VNB VPB VPWR X
*.PININFO A:I SLEEP_B:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNI23 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI8 VPWR net44 X VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 net56 SLEEP_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 sndPA net56 net44 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 net56 SLEEP_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI25 net44 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X net44 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI9 net44 net56 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_inputiso1n_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA3 pndA A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 Y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 sndA3 VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA3 sndA3 A4 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a41oi_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA3 pndA A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 Y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 sndA3 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA3 sndA3 A4 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a41oi_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA3 pndA A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 Y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 sndA3 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA3 sndA3 A4 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a41oi_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMP2 sndPB C sndPC VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMP3 sndPC D Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=0.76
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=0.76
XMXNMN2 Y C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=0.76
XMXNMN3 Y D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=0.76
.ENDS sky130_fd_sc_hd__nor4_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMP2 sndPB C sndPC VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMP3 sndPC D Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=0.76
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=0.76
XMXNMN2 Y C VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=0.76
XMXNMN3 Y D VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=0.76
.ENDS sky130_fd_sc_hd__nor4_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMP2 sndPB C sndPC VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMP3 sndPC D Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=0.76
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=0.76
XMXNMN2 Y C VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=0.76
XMXNMN3 Y D VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=0.76
.ENDS sky130_fd_sc_hd__nor4_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__tapvgnd2_1 VGND VPB VPWR
*.PININFO VGND:I VPB:I VPWR:I
* Notes: substrate is tied to vgnd in the cell and does not appear as
*        a pin.
.ENDS sky130_fd_sc_hd__tapvgnd2_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
*.PININFO A_N:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and3b_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
*.PININFO A_N:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and3b_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
*.PININFO A_N:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and3b_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nor2_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B Y VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=8 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=8 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nor2_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nor2_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nor2_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__macro_sparecell VGND VNB VPB VPWR LO
*.PININFO VGND:I VNB:I VPB:I VPWR:I LO:O
XI1 net59 LO VGND VNB VPB VPWR / sky130_fd_sc_hd__conb_1
XI6 nor2right invright VGND VNB VPB VPWR / sky130_fd_sc_hd__inv_2
XI7 nor2left invleft VGND VNB VPB VPWR / sky130_fd_sc_hd__inv_2
XI4 nd2right nd2right nor2right VGND VNB VPB VPWR /
+ sky130_fd_sc_hd__nor2_2
XI5 nd2left nd2left nor2left VGND VNB VPB VPWR /
+ sky130_fd_sc_hd__nor2_2
XI2 LO LO nd2right VGND VNB VPB VPWR / sky130_fd_sc_hd__nand2_2
XI3 LO LO nd2left VGND VNB VPB VPWR / sky130_fd_sc_hd__nand2_2
.ENDS sky130_fd_sc_hd__macro_sparecell


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
*.PININFO VGND:I VNB:I VPB:I VPWR:I HI:O LO:O
rI12 VGND LO short w=480000u l=45000u
rI11 HI VPWR short w=480000u l=45000u
.ENDS sky130_fd_sc_hd__conb_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__tapvgnd_1 VGND VPB VPWR
*.PININFO VGND:I VPB:I VPWR:I
* Notes: substrate is tied to vgnd in the cell and does not appear as
*        a pin.
.ENDS sky130_fd_sc_hd__tapvgnd_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlymetal6s6s_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab net56 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 net56 net48 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI15 net52 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI9 net48 net44 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI16 net44 net52 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab net56 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 net56 net48 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI8 net48 net44 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 net44 net52 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 net52 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlymetal6s6s_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI657 M0 clkpos net79 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net79 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 Q S1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 S0 clkneg net59 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI641 net59 S1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M1 clkpos S0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M0 clkneg net107 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 S0 clkpos net122 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI639 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.75 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI643 net122 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net107 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 Q S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 M1 clkneg S0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dfxtp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI657 M0 clkpos net79 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net79 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 Q S1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 S0 clkneg net59 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI641 net59 S1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M1 clkpos S0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M0 clkneg net107 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 S0 clkpos net122 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI639 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.75 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI643 net122 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net107 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 Q S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 M1 clkneg S0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dfxtp_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI657 M0 clkpos net79 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net79 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 Q S1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 S0 clkneg net59 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI641 net59 S1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M1 clkpos S0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M0 clkneg net107 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 S0 clkpos net122 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI639 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.75 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI643 net122 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net107 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 Q S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 M1 clkneg S0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dfxtp_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C sndPC VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 sndPC D y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP4 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 y C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN3 y D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN4 X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or4_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C sndPC VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 sndPC D y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP4 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 y C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN3 y D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN4 X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or4_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C sndPC VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 sndPC D y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP4 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 y C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN3 y D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN4 X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or4_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrckapwr_16 A SLEEP KAPWR VGND VNB VPB VPWR X
*.PININFO A:I SLEEP:I KAPWR:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR SLEEP sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA net58 net66 VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 net58 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 Ab net66 KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI9 X Ab KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=16 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 net66 SLEEP VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN1 net66 net58 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 net58 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 Ab net66 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI8 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=16 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_isobufsrckapwr_16


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
*.PININFO VGND:I VNB:I VPB:I VPWR:I
XMXNI1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.55 l=2.89 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI2 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.87 l=2.89 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__decap_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
*.PININFO VGND:I VNB:I VPB:I VPWR:I
XMXNI2 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.87 l=1.05 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.55 l=1.05 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__decap_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
*.PININFO VGND:I VNB:I VPB:I VPWR:I
XMXNI1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.55 l=0.59 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI2 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.87 l=0.59 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__decap_3


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
*.PININFO VGND:I VNB:I VPB:I VPWR:I
XMXNI1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.55 l=4.73 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI2 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.87 l=4.73 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__decap_12


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
*.PININFO VGND:I VNB:I VPB:I VPWR:I
XMXNI1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.55 l=1.97 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI2 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.87 l=1.97 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__decap_6


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 sndB1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 sndB1 B2 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 y B2 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o22a_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 sndB1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 sndB1 B2 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 y B2 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o22a_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 sndB1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 sndB1 B2 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 y B2 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o22a_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdfsbp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I SCD:I SCE:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
*.PININFO Q_N:O
XMXNI101 db sceb p1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI94 db D p0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 sceb SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 net195 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net195 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M1 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net130 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 M0 clkneg net130 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 net122 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI669 S0 clkpos net122 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 S0 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI38 S0 clkneg net107 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI37 net107 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI661 Q_N S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI98 db D n0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=3.1
XMXNI103 n1 SCD VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI120 db SCE n1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI104 n0 sceb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI34 S0 clkpos net219 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI27 net239 S1 net187 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 M0 clkpos net230 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 M1 M0 net199 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net230 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI36 net219 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI26 S0 clkneg net239 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net199 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 net195 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 sceb SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI25 net187 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net195 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 Q_N S0 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sdfsbp_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdfsbp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I SCD:I SCE:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
*.PININFO Q_N:O
XMXNI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI94 db D p0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI101 db sceb p1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net159 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 M0 clkneg net159 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 net138 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI669 S0 clkpos net138 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI661 Q_N S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M1 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 sceb SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 net199 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net199 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 S0 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI38 S0 clkneg net98 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI37 net98 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI120 db SCE n1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI104 n0 sceb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI103 n1 SCD VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI98 db D n0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=3.1
XMXNI27 net243 S1 net215 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 S0 clkpos net230 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net227 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net199 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 sceb SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI25 net215 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 Q_N S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 M0 clkpos net206 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 net199 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 M1 M0 net227 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net206 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI36 net230 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI26 S0 clkneg net243 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sdfsbp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dfxbp_2 CLK D VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
XMXNI657 M0 clkpos net96 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net96 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 Q S1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI669 net88 S1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 S0 clkneg net72 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI641 net72 S1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M1 clkpos S0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI665 Q_N net88 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M0 clkneg net128 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 S0 clkpos net147 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI639 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.75 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI670 net88 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI643 net147 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net128 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 Q S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 M1 clkneg S0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI666 Q_N net88 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dfxbp_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dfxbp_1 CLK D VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
XMXNI657 M0 clkpos net96 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net96 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 Q S1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI669 net88 S1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 S0 clkneg net72 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI641 net72 S1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M1 clkpos S0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI665 Q_N net88 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M0 clkneg net128 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 S0 clkpos net147 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI639 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.75 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI670 net88 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI643 net147 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net128 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 Q S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 M1 clkneg S0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI666 Q_N net88 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dfxbp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMNnor0 inor A1_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnor1 inor A2_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi10 VGND B1 sndNB1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi11 sndNB1 B2 Y VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi20 Y inor VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnor0 VPWR A1_N sndPA1N VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnor1 sndPA1N A2_N inor VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi10 pmid B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi11 pmid B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi20 Y inor pmid VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a2bb2oi_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMNnor0 inor A1_N VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnor1 inor A2_N VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi10 VGND B1 sndNB1 VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi11 sndNB1 B2 Y VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi20 Y inor VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnor0 VPWR A1_N sndPA1N VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnor1 sndPA1N A2_N inor VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi10 pmid B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi11 pmid B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi20 Y inor pmid VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a2bb2oi_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMNnor0 inor A1_N VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnor1 inor A2_N VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi10 VGND B1 sndNB1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi11 sndNB1 B2 Y VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi20 Y inor VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnor0 VPWR A1_N sndPA1N VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnor1 sndPA1N A2_N inor VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi10 pmid B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi11 pmid B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi20 Y inor pmid VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a2bb2oi_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor4bb_2 A B C_N D_N VGND VNB VPB VPWR Y
*.PININFO A:I B:I C_N:I D_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C sndPC VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 sndPC D Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 C C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 D D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 Y C VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN3 Y D VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN2 C C_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 D D_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nor4bb_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor4bb_1 A B C_N D_N VGND VNB VPB VPWR Y
*.PININFO A:I B:I C_N:I D_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C sndPC VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 sndPC D Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 C C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 D D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 Y C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN3 Y D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN2 C C_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 D D_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nor4bb_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor4bb_4 A B C_N D_N VGND VNB VPB VPWR Y
*.PININFO A:I B:I C_N:I D_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C sndPC VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 sndPC D Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 C C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 D D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 Y C VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN3 Y D VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN2 C C_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 D D_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nor4bb_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__ha_4 A B VGND VNB VPB VPWR COUT SUM
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I COUT:O SUM:O
XMXNMIN2 COUT majb VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 SUM sumb VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnand0 VGND A sndNA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnand1 sndNA B majb VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs1 sumb majb nint1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs20 VGND A nint1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs21 VGND B nint1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 COUT majb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 SUM sumb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand0 majb A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand1 majb B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs1 VPWR majb sumb VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs20 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs21 sndPA B sumb VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__ha_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__ha_2 A B VGND VNB VPB VPWR COUT SUM
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I COUT:O SUM:O
XMXNMIN2 COUT majb VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 SUM sumb VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnand0 VGND A sndNA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnand1 sndNA B majb VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs1 sumb majb nint1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs20 VGND A nint1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs21 VGND B nint1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 COUT majb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 SUM sumb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand0 majb A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand1 majb B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs1 VPWR majb sumb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs20 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs21 sndPA B sumb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__ha_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__ha_1 A B VGND VNB VPB VPWR COUT SUM
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I COUT:O SUM:O
XMXNMIN2 COUT majb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 SUM sumb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnand0 VGND A sndNA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnand1 sndNA B majb VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs1 sumb majb nint1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs20 VGND A nint1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs21 VGND B nint1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 COUT majb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 SUM sumb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand0 majb A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand1 majb B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs1 VPWR majb sumb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs20 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs21 sndPA B sumb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__ha_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlclkp_4 CLK GATE VGND VNB VPB VPWR GCLK
*.PININFO CLK:I GATE:I VGND:I VNB:I VPB:I VPWR:I GCLK:O
XMXNI662 net75 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 M0 clkpos net75 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 net63 CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net63 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI38 M0 clkneg net54 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI37 net54 GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkpos CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 GCLK net63 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 m1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 M0 clkneg net110 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net110 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 M0 clkpos net91 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net99 CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net63 m1 net99 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI36 net91 GATE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkpos CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 GCLK net63 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlclkp_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
*.PININFO CLK:I GATE:I VGND:I VNB:I VPB:I VPWR:I GCLK:O
XMXNI662 net75 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 M0 clkpos net75 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 net63 CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net63 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI38 M0 clkneg net54 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI37 net54 GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkpos CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 GCLK net63 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 m1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 M0 clkneg net110 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.39 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net110 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 M0 clkpos net91 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net99 CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net63 m1 net99 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI36 net91 GATE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkpos CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 GCLK net63 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlclkp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlclkp_2 CLK GATE VGND VNB VPB VPWR GCLK
*.PININFO CLK:I GATE:I VGND:I VNB:I VPB:I VPWR:I GCLK:O
XMXNI662 net75 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 M0 clkpos net75 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 net63 CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net63 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI38 M0 clkneg net54 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI37 net54 GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkpos CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 GCLK net63 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 m1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 M0 clkneg net110 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.39 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net110 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 M0 clkpos net91 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net99 CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net63 m1 net99 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI36 net91 GATE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkpos CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 GCLK net63 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlclkp_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN2 X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or2_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN2 X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or2_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or2_0 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN2 X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or2_0


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN2 X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or2_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlymetal6s4s_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab X VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 net59 Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 X net47 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI15 net51 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI9 net47 net43 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI16 net43 net51 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab X VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 net59 Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 X net47 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI8 net47 net43 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 net43 net51 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 net51 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlymetal6s4s_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__xnor3_4 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN3 X net57 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI29 Ab Bb mid2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.6 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI25 Abb Bb mid1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 Bb B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 mid1 Cb net57 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 Cb C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI2 mid2 C net57 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 Abb Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 Ab B mid1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI28 Abb B mid2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 X net57 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 mid1 C net57 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI27 mid2 B Ab VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 Abb Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI23 mid1 B Abb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI26 mid2 Bb Abb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 mid2 Cb net57 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 Cb C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI16 Bb B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 mid1 Bb Ab VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__xnor3_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__xnor3_1 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN3 X net57 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI29 Ab Bb mid2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.6 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI25 Abb Bb mid1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 Bb B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 mid1 Cb net57 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 Cb C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI2 mid2 C net57 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 Abb Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 Ab B mid1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI28 Abb B mid2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 X net57 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 mid1 C net57 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI27 mid2 B Ab VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 Abb Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI23 mid1 B Abb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI26 mid2 Bb Abb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 mid2 Cb net57 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 Cb C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI16 Bb B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 mid1 Bb Ab VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__xnor3_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__xnor3_2 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN3 X net57 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI29 Ab Bb mid2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.6 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI25 Abb Bb mid1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 Bb B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 mid1 Cb net57 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 Cb C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI2 mid2 C net57 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 Abb Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 Ab B mid1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI28 Abb B mid2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 X net57 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 mid1 C net57 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI27 mid2 B Ab VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 Abb Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI23 mid1 B Abb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI26 mid2 Bb Abb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 mid2 Cb net57 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 Cb C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI16 Bb B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 mid1 Bb Ab VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__xnor3_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dfbbn_1 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK_N:I D:I RESET_B:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
*.PININFO Q_N:O
XMXNI46 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 RESET RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI676 M1 M0 net141 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI675 net141 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net162 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI677 M1 RESET net141 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 M0 clkpos net125 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkpos CLK_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 net125 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 S0 clkneg net110 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net110 net82 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 Q_N net82 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 net162 net82 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI668 S0 clkpos net93 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI667 net93 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI630 net82 RESET net81 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI3 net82 S0 net81 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 net81 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI679 M1 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI669 S0 clkneg net218 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net162 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI9 net82 S0 net221 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI670 net218 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI678 net165 RESET VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net210 net82 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 S0 clkpos net210 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI10 net82 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI11 net221 RESET VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 net194 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI665 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 M0 clkneg net194 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI643 RESET RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkpos CLK_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI680 M1 M0 net165 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 net162 net82 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI661 Q_N net82 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dfbbn_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dfbbn_2 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK_N:I D:I RESET_B:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
*.PININFO Q_N:O
XMXNI46 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 RESET RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI676 M1 M0 net141 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI675 net141 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net162 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI677 M1 RESET net141 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 M0 clkpos net125 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkpos CLK_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 net125 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 S0 clkneg net110 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net110 net82 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 Q_N net82 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 net162 net82 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI668 S0 clkpos net93 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI667 net93 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI630 net82 RESET net81 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI3 net82 S0 net81 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 net81 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI679 M1 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI669 S0 clkneg net218 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net162 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI9 net82 S0 net221 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI670 net218 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI678 net165 RESET VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net210 net82 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 S0 clkpos net210 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI10 net82 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI11 net221 RESET VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 net194 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI665 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 M0 clkneg net194 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI643 RESET RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkpos CLK_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI680 M1 M0 net165 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 net162 net82 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI661 Q_N net82 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dfbbn_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab net34 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 net34 net30 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI9 net30 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab net34 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 net34 net30 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI8 net30 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlygate4sd1_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and2_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and2_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and2_0 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and2_0


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and2_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdfstp_4 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SCD:I SCE:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI645 sceb SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 net165 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net165 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M1 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net104 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 M0 clkneg net104 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 net96 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI669 S0 clkpos net96 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 S0 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI38 S0 clkneg net84 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI37 net84 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI101 db sceb p1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI94 db D p0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 S0 clkpos net189 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI27 net209 S1 net157 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 M0 clkpos net200 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 M1 M0 net169 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net200 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI36 net189 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI26 S0 clkneg net209 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net169 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 net165 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 sceb SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI25 net157 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net165 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI98 db D n0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=3.1
XMXNI103 n1 SCD VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI120 db SCE n1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI104 n0 sceb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
.ENDS sky130_fd_sc_hd__sdfstp_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdfstp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SCD:I SCE:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI645 sceb SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 net165 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net165 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M1 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net109 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 M0 clkneg net109 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 net96 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI669 S0 clkpos net96 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 S0 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI38 S0 clkneg net84 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI37 net84 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI101 db sceb p1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI94 db D p0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 S0 clkpos net212 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI27 net209 S1 net157 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 M0 clkpos net200 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 M1 M0 net196 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net200 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI36 net212 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI26 S0 clkneg net209 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net196 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 net165 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 sceb SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI25 net157 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net165 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI98 db D n0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=3.1
XMXNI103 n1 SCD VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI120 db SCE n1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI104 n0 sceb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
.ENDS sky130_fd_sc_hd__sdfstp_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdfstp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SCD:I SCE:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI645 sceb SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 net165 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net165 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M1 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net109 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 M0 clkneg net109 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 net96 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI669 S0 clkpos net96 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 S0 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI38 S0 clkneg net84 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI37 net84 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI101 db sceb p1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI94 db D p0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 S0 clkpos net189 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI27 net209 S1 net157 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 M0 clkpos net200 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 M1 M0 net169 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net200 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI36 net189 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI26 S0 clkneg net209 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net169 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 net165 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 sceb SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI25 net157 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net165 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI98 db D n0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=3.1
XMXNI103 n1 SCD VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI120 db SCE n1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI104 n0 sceb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
.ENDS sky130_fd_sc_hd__sdfstp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI36 net120 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI39 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 M1 M0 net103 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net71 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 S0 clkpos net120 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI25 net88 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI26 S0 clkneg net80 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI27 net80 S1 net88 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 M0 clkpos net71 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net103 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 net128 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net128 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI40 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI38 S0 clkneg net179 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI37 net179 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M1 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net156 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 M0 clkneg net156 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 net143 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 S0 clkpos net143 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 S0 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 net128 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net128 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dfstp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI36 net120 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI39 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 M1 M0 net103 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net71 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 S0 clkpos net120 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI25 net88 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI26 S0 clkneg net80 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI27 net80 S1 net88 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 M0 clkpos net71 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net103 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 net128 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net128 VGND VNB sky130_fd_pr__nfet_01v8 m=5 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI40 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI38 S0 clkneg net179 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI37 net179 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M1 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net156 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 M0 clkneg net156 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 net143 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 S0 clkpos net143 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 S0 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 net128 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net128 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=5 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dfstp_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI36 net120 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI39 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 M1 M0 net103 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net71 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 S0 clkpos net120 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI25 net88 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI26 S0 clkneg net80 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI27 net80 S1 net88 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 M0 clkpos net71 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net103 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 net128 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net128 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI40 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI38 S0 clkneg net179 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI37 net179 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M1 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net156 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 M0 clkneg net156 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 net143 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 S0 clkpos net143 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 S0 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 net128 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net128 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dfstp_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__probec_p_8 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=3 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 net33 Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=3 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 net33 Ab VGND VNB sky130_fd_pr__nfet_01v8 m=8 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
rI112 net33 X sky130_fd_pr__res_generic_po
rI120 VGND met5vgnd sky130_fd_pr__res_generic_po
rI119 VPWR met5vpwr sky130_fd_pr__res_generic_po
.ENDS sky130_fd_sc_hd__probec_p_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdfbbp_1 CLK D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I RESET_B:I SCD:I SCE:I SET_B:I VGND:I VNB:I VPB:I
*.PININFO VPWR:I Q:O Q_N:O
XMXNI98 net105 D n0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI103 n1 SCD VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI104 n0 sceb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI120 net105 SCE n1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 RESET RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI676 M1 M0 net176 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI675 net176 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net213 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI677 M1 RESET net176 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 M0 clkpos net160 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 net160 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 S0 clkneg net145 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net145 net117 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 Q_N net117 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 net213 net117 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 net105 clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI668 S0 clkpos net125 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI667 net125 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI630 net117 RESET net116 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI3 net117 S0 net116 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 net116 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI639 sceb SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI94 net105 D p0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI101 net105 sceb p1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI679 M1 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI669 S0 clkneg net265 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net213 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI9 net117 S0 net268 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI670 net265 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI678 net216 RESET VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net257 net117 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 S0 clkpos net257 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI10 net117 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI11 net268 RESET VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 net241 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 net105 clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 M0 clkneg net241 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI643 RESET RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI680 M1 M0 net216 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 net213 net117 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI661 Q_N net117 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI640 sceb SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sdfbbp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 y B2 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 sndB1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 sndB1 B2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a32o_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 y B2 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 sndB1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 sndB1 B2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a32o_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 y B2 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 sndB1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 sndB1 B2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a32o_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
*.PININFO A_N:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and2b_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
*.PININFO A_N:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and2b_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
*.PININFO A_N:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and2b_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__bufinv_8 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 Abb Ab VGND VNB sky130_fd_pr__nfet_01v8 m=3 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 Y Abb VGND VNB sky130_fd_pr__nfet_01v8 m=8 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 Abb Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=3 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 Y Abb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__bufinv_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=3 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 Abb Ab VGND VNB sky130_fd_pr__nfet_01v8 m=6 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 Y Abb VGND VNB sky130_fd_pr__nfet_01v8 m=16 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=3 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 Abb Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=6 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 Y Abb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=16 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__bufinv_16


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a21o_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a21o_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a21o_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
*.PININFO A_N:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C sndC VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN3 sndC D VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand4b_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
*.PININFO A_N:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C sndC VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN3 sndC D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand4b_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
*.PININFO A_N:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C sndC VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN3 sndC D VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand4b_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMNnor0 inor A VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnor1 inor B VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi10 VGND A sndNA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi11 sndNA B X VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi20 X inor VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnor0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnor1 sndPA B inor VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi10 pmid A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi11 pmid B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi20 X inor pmid VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__xor2_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMNnor0 inor A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnor1 inor B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi10 VGND A sndNA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi11 sndNA B X VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi20 X inor VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnor0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnor1 sndPA B inor VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi10 pmid A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi11 pmid B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi20 X inor pmid VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__xor2_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMNnor0 inor A VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnor1 inor B VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi10 VGND A sndNA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi11 sndNA B X VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi20 X inor VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnor0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnor1 sndPA B inor VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi10 pmid A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi11 pmid B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi20 X inor pmid VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__xor2_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 sndB1 VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 sndB1 B2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 pndB B2 pndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 pndB VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o221ai_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 sndB1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 sndB1 B2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 pndB B2 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 pndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o221ai_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 sndB1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 sndB1 B2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 pndB B2 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 pndB VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o221ai_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 sndA3 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA3 sndA3 A4 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA3 pndA A4 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o41a_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 sndA3 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA3 sndA3 A4 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA3 pndA A4 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o41a_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 sndA3 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA3 sndA3 A4 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA3 pndA A4 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o41a_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
*.PININFO A_N:I B_N:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 B B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C sndC VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN3 sndC D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 B B_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and4bb_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
*.PININFO A_N:I B_N:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 B B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C sndC VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN3 sndC D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 B B_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and4bb_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
*.PININFO A_N:I B_N:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 B B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C sndC VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN3 sndC D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 B B_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and4bb_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
*.PININFO CLK_N:I D:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI46 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net83 net121 net109 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net109 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 net102 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 M0 clkpos net94 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 net94 M1 net102 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 net121 clkneg net82 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net83 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net82 net83 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkpos CLK_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI39 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 M1 clkpos net121 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net166 net83 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 net83 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 net121 clkpos net166 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net83 net121 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI30 net145 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI31 M0 clkneg net145 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI32 net145 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net83 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkpos CLK_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI40 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 M1 clkneg net121 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dfrtn_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I D_N:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C sndPC VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 sndPC D y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 D D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP4 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 y C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN3 y D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN3 D D_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN4 X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or4b_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I D_N:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C sndPC VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 sndPC D y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 D D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP4 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 y C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN3 y D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN3 D D_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN4 X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or4b_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I D_N:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C sndPC VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 sndPC D y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 D D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP4 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 y C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN3 y D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN3 D D_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN4 X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or4b_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 pndB B2 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 y C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 sndB1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 sndB1 B2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a221o_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 pndB B2 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 y C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 sndB1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 sndB1 B2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a221o_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 pndB B2 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 y C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 sndB1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 sndB1 B2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a221o_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMNnand0 VGND A sndNA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnand1 sndNA B inand VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi10 nmid A VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi11 nmid B VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi20 Y inand nmid VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand0 inand A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand1 inand B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi10 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi11 sndPA B Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi20 Y inand VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__xnor2_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMNnand0 VGND A sndNA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnand1 sndNA B inand VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi10 nmid A VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi11 nmid B VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi20 Y inand nmid VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand0 inand A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand1 inand B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi10 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi11 sndPA B Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi20 Y inand VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__xnor2_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMNnand0 VGND A sndNA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnand1 sndNA B inand VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi10 nmid A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi11 nmid B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi20 Y inand nmid VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand0 inand A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand1 inand B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi10 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi11 sndPA B Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi20 Y inand VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__xnor2_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 y C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN3 X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or3_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 y C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN3 X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or3_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 y C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN3 X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or3_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
*.PININFO A_N:I B:I C:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand3b_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
*.PININFO A_N:I B:I C:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand3b_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
*.PININFO A_N:I B:I C:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand3b_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 A2 Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 Ab2 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 X Ab2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 A2 Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.82 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 Ab2 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.82 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 X Ab2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__clkdlybuf4s50_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__clkdlybuf4s50_2 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 A2 Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 Ab2 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 X Ab2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 A2 Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.82 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 Ab2 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.82 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 X Ab2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__clkdlybuf4s50_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__fah_1 A B CI VGND VNB VPB VPWR COUT SUM
*.PININFO A:I B:I CI:I VGND:I VNB:I VPB:I VPWR:I COUT:O SUM:O
XMXNMIN2 COUT net195 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 SUM net123 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 CIb mid2 net195 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 Bb mid1 net195 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI2 CIbb mid2 net123 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 CIb mid1 net123 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 Bb B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 CIbb CIb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 CIb CI VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI8 Ab2 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI9 Abb2 Ab2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI14 Ab1 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 Abb2 B mid1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI21 Ab1 Bb mid1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 Abb2 Bb mid2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI25 Ab1 B mid2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 COUT net195 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 SUM net123 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 CIb mid1 net195 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI3 Bb mid2 net195 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI1 CIbb mid1 net123 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 CIb mid2 net123 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI16 Bb B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 CIbb CIb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 CIb CI VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI12 Ab2 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI13 Abb2 Ab2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 Ab1 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI22 Abb2 Bb mid1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI23 Ab1 B mid1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI26 Abb2 B mid2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI27 Ab1 Bb mid2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__fah_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a222oi_1 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 pndB B2 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 Y C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI8 Y C2 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 sndB1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 sndB1 B2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 net62 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI10 net62 C2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a222oi_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_16 A SLEEP VGND VNB VPB VPWR X
*.PININFO A:I SLEEP:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR Ab sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=16 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt m=16 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 m=16 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN1 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=16 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_isobufsrc_16


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_4 A SLEEP VGND VNB VPB VPWR X
*.PININFO A:I SLEEP:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR SLEEP sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA Ab X VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN1 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_isobufsrc_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_1 A SLEEP VGND VNB VPB VPWR X
*.PININFO A:I SLEEP:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR SLEEP sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA Ab X VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN1 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_isobufsrc_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_2 A SLEEP VGND VNB VPB VPWR X
*.PININFO A:I SLEEP:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR SLEEP sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA Ab X VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN1 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_isobufsrc_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_8 A SLEEP VGND VNB VPB VPWR X
*.PININFO A:I SLEEP:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR Ab sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 m=8 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN1 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=8 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_isobufsrc_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dfbbp_1 CLK D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I RESET_B:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
*.PININFO Q_N:O
XMXNI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 RESET RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI676 M1 M0 net141 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI675 net141 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net162 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI677 M1 RESET net141 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 M0 clkpos net118 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 net118 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 S0 clkneg net110 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net110 net82 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 Q_N net82 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 net162 net82 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI668 S0 clkpos net93 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI667 net93 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI630 net82 RESET net81 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI3 net82 S0 net81 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 net81 SET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI679 M1 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI669 S0 clkneg net218 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net162 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI9 net82 S0 net221 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI670 net218 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI678 net165 RESET VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net210 net82 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 S0 clkpos net210 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI10 net82 SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI11 net221 RESET VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 net194 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI665 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 M0 clkneg net194 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI643 RESET RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI680 M1 M0 net165 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 net162 net82 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI661 Q_N net82 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dfbbp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 y C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a211o_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 y C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a211o_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 y C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a211o_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPD0 VPWR D1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 pndC C1 pndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMND0 y D1 pndC VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o2111a_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPD0 VPWR D1 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 pndC C1 pndB VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMND0 y D1 pndC VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o2111a_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPD0 VPWR D1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 pndC C1 pndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMND0 y D1 pndC VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o2111a_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlrbp_1 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
*.PININFO D:I GATE:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
XMXNI635 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 Q_N net125 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 M0 clkneg net61 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 net125 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 Q m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 clkneg GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 m1 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 net61 db VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 net57 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 M0 clkpos net57 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 clkneg GATE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 Q_N net125 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 Q m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 net125 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net121 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M0 clkneg net116 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net116 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 m1 M0 net121 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 M0 clkpos net96 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 net96 db VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlrbp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlrbp_2 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
*.PININFO D:I GATE:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
XMXNI635 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 Q_N net125 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 M0 clkneg net61 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 net125 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 Q m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 clkneg GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 m1 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 net61 db VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 net57 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 M0 clkpos net57 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 clkneg GATE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 Q_N net125 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 Q m1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 net125 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net108 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M0 clkneg net116 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net116 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 m1 M0 net108 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 M0 clkpos net96 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 net96 db VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlrbp_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 pndB VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o211ai_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 pndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o211ai_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 pndB VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o211ai_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and3_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and3_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and3_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_8 A KAPWR VGND VNB VPB VPWR X
*.PININFO A:I KAPWR:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN0 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=8 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 Ab A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 X Ab KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_clkbufkapwr_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_1 A KAPWR VGND VNB VPB VPWR X
*.PININFO A:I KAPWR:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN0 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.52 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.52 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 Ab A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.79 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 X Ab KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.79 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_clkbufkapwr_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_16 A KAPWR VGND VNB VPB VPWR X
*.PININFO A:I KAPWR:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN0 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=16 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 Ab A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 X Ab KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=16 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_clkbufkapwr_16


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_2 A KAPWR VGND VNB VPB VPWR X
*.PININFO A:I KAPWR:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN0 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 Ab A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 X Ab KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_clkbufkapwr_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_4 A KAPWR VGND VNB VPB VPWR X
*.PININFO A:I KAPWR:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN0 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 Ab A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 X Ab KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_clkbufkapwr_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o31a_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o31a_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o31a_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN2 X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnand0 VGND A1_N sndNA1N VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnand1 sndNA1N A2_N inand VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi10 nmid B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi11 nmid B2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi20 y inand nmid VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand0 inand A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand1 inand A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi10 VPWR B1 sndPB1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi11 sndPB1 B2 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi20 y inand VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o2bb2a_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN2 X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnand0 VGND A1_N sndNA1N VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnand1 sndNA1N A2_N inand VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi10 nmid B1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi11 nmid B2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi20 y inand nmid VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand0 inand A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand1 inand A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi10 VPWR B1 sndPB1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi11 sndPB1 B2 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi20 y inand VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o2bb2a_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN2 X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnand0 VGND A1_N sndNA1N VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnand1 sndNA1N A2_N inand VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi10 nmid B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi11 nmid B2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi20 y inand nmid VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand0 inand A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnand1 inand A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi10 VPWR B1 sndPB1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi11 sndPB1 B2 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi20 y inand VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o2bb2a_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_bleeder_1 sky130_fd_pr__res_generic_po VGND VNB VPB VPWR
*.PININFO sky130_fd_pr__res_generic_po:I VGND:I VNB:I VPB:I VPWR:B
XMXNI2 net29 sky130_fd_pr__res_generic_po net25 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI3 net25 sky130_fd_pr__res_generic_po net24 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI1 VPWR sky130_fd_pr__res_generic_po net29 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 net24 sky130_fd_pr__res_generic_po net16 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 net16 sky130_fd_pr__res_generic_po VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_bleeder_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPB1N B1 B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINB1N B1 B1_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o21bai_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPB1N B1 B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINB1N B1 B1_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o21bai_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPB1N B1 B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINB1N B1 B1_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o21bai_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
*.PININFO A:I B_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 B B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN1 B B_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nor2b_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
*.PININFO A:I B_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 B B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN1 B B_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nor2b_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
*.PININFO A:I B_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 B B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN1 B B_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nor2b_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 sndB1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 sndB1 B2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 Y B2 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o32ai_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 sndB1 VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 sndB1 B2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 Y B2 pndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o32ai_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 sndB1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 sndB1 B2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 Y B2 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o32ai_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 pndC C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPD0 Y D1 pndC VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMND0 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a2111oi_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a2111oi_0 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 pndC C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPD0 Y D1 pndC VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMND0 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a2111oi_0


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 pndC C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPD0 Y D1 pndC VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMND0 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a2111oi_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 pndC C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPD0 Y D1 pndC VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMND0 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a2111oi_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_16 A KAPWR VGND VNB VPB VPWR Y
*.PININFO A:I KAPWR:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMIN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=16 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=24 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_clkinvkapwr_16


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_2 A KAPWR VGND VNB VPB VPWR Y
*.PININFO A:I KAPWR:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMIN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=3 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_clkinvkapwr_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_8 A KAPWR VGND VNB VPB VPWR Y
*.PININFO A:I KAPWR:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMIN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=8 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=12 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_clkinvkapwr_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_4 A KAPWR VGND VNB VPB VPWR Y
*.PININFO A:I KAPWR:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMIN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=6 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_clkinvkapwr_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_1 A KAPWR VGND VNB VPB VPWR Y
*.PININFO A:I KAPWR:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMIN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_clkinvkapwr_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
*.PININFO D:I GATE:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
XMXNI635 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 Q_N net114 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 M0 clkneg net58 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 net114 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 Q m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 clkneg GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 net58 db VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 net54 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 M0 clkpos net54 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 clkneg GATE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 Q_N net114 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 Q m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 net114 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M0 clkneg net109 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net109 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 m1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 M0 clkpos net89 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 net89 db VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlxbp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
*.PININFO D:I GATE_N:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI635 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 M0 clkneg net53 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 Q m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 clkpos GATE_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 net53 db VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 net44 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 M0 clkpos net44 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 clkpos GATE_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 Q m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M0 clkneg net96 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net96 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 m1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 M0 clkpos net76 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 net76 db VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlxtn_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlxtn_4 D GATE_N VGND VNB VPB VPWR Q
*.PININFO D:I GATE_N:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI635 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 M0 clkneg net51 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 Q m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 clkpos GATE_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 net51 db VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 net47 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 M0 clkpos net47 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 clkpos GATE_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 Q m1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M0 clkneg net94 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net94 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 m1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 M0 clkpos net74 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 net74 db VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlxtn_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
*.PININFO D:I GATE_N:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI635 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 M0 clkneg net51 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 Q m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 clkpos GATE_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 net51 db VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 net47 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 M0 clkpos net47 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 clkpos GATE_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 Q m1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M0 clkneg net94 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net94 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 m1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 M0 clkpos net74 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 net74 db VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlxtn_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 y C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a311o_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 y C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a311o_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 y C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a311o_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand3_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand3_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand3_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
*.PININFO A:I B_N:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 B B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN1 B B_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or2b_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
*.PININFO A:I B_N:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 B B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN1 B B_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or2b_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
*.PININFO A:I B_N:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 B B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN1 B B_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or2b_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
*.PININFO A_N:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand2b_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
*.PININFO A_N:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand2b_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
*.PININFO A_N:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand2b_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 pndB B2 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 Y C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 sndB1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 sndB1 B2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a221oi_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 pndB B2 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 Y C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 sndB1 VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 sndB1 B2 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a221oi_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 pndB B2 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 Y C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 sndB1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 sndB1 B2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a221oi_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
XMXNI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net99 s0 net125 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net125 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 net118 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 M0 clkpos net110 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 net110 M1 net118 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 s0 clkneg net98 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net99 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net98 net99 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI39 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 M1 clkpos s0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI53 net142 net99 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI50 Q_N net142 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net190 net99 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 net99 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 s0 clkpos net190 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net99 s0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI30 net169 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI31 M0 clkneg net169 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI32 net169 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net99 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI40 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 M1 clkneg s0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI52 net142 net99 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI51 Q_N net142 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dfrbp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
XMXNI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net99 s0 net125 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net125 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 net118 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 M0 clkpos net110 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 net110 M1 net118 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 s0 clkneg net98 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net99 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net98 net99 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI39 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 M1 clkpos s0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI53 net142 net99 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI50 Q_N net142 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net181 net99 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 net99 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 s0 clkpos net181 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net99 s0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI30 net169 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI31 M0 clkneg net169 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI32 net169 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net99 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI40 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 M1 clkneg s0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI52 net142 net99 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI51 Q_N net142 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dfrbp_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
*.PININFO VGND:I VNB:I VPB:I VPWR:I
* Notes: Cell contains no devices
.ENDS sky130_fd_sc_hd__fill_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__fill_4 VGND VNB VPB VPWR
*.PININFO VGND:I VNB:I VPB:I VPWR:I
* Notes: Cell contains no devices
.ENDS sky130_fd_sc_hd__fill_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
*.PININFO VGND:I VNB:I VPB:I VPWR:I
* Notes: Cell contains no devices
.ENDS sky130_fd_sc_hd__fill_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__fill_8 VGND VNB VPB VPWR
*.PININFO VGND:I VNB:I VPB:I VPWR:I
* Notes: Cell contains no devices
.ENDS sky130_fd_sc_hd__fill_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab net34 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 net34 net30 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI9 net30 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab net34 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 net34 net30 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI8 net30 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlygate4sd3_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 y C1 pndB VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o211a_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 y C1 pndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o211a_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 y C1 pndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o211a_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlygate4sd2_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab net34 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.18 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 net34 net30 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.18 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI9 net30 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab net34 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.18
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 net34 net30 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.18
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI8 net30 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlygate4sd2_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdfxtp_1 CLK D SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI652 M1 clkpos S0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI639 sceb SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 M0 clkpos net78 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net78 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI641 net54 S1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 Q S1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 S0 clkneg net54 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI98 db D n0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=3.1
XMXNI103 n1 SCD VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI120 db SCE n1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI104 n0 sceb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI643 net122 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI640 sceb SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net155 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 Q S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 M1 clkneg S0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M0 clkneg net155 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 S0 clkpos net122 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.75 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI94 db D p0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI101 db sceb p1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sdfxtp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdfxtp_4 CLK D SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI652 M1 clkpos S0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI639 sceb SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 M0 clkpos net78 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net78 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI641 net54 S1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 Q S1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 S0 clkneg net54 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI98 db D n0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=3.1
XMXNI103 n1 SCD VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI120 db SCE n1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI104 n0 sceb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI643 net163 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI640 sceb SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net155 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 Q S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 M1 clkneg S0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M0 clkneg net155 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 S0 clkpos net163 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.75 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI94 db D p0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI101 db sceb p1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sdfxtp_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdfxtp_2 CLK D SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI652 M1 clkpos S0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI639 sceb SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 M0 clkpos net78 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net78 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI641 net54 S1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 Q S1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 S0 clkneg net54 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI98 db D n0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=3.1
XMXNI103 n1 SCD VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI120 db SCE n1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI104 n0 sceb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI643 net163 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI640 sceb SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net138 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 Q S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 M1 clkneg S0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M0 clkneg net138 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 S0 clkpos net163 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.75 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI94 db D p0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI101 db sceb p1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sdfxtp_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__maj3_1 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN2 X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN10 y B sndNBa VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN11 sndNBa A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN20 y B sndNBc VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN21 sndNBc C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN30 y C sndNCa VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN31 sndNCa A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP10 VPWR A sndPAb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP11 sndPAb B y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP20 VPWR C sndPCb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP21 sndPCb B y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP30 VPWR A sndPAc VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP31 sndPAc C y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__maj3_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__maj3_2 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN2 X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN10 y B sndNBa VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN11 sndNBa A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN20 y B sndNBc VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN21 sndNBc C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN30 y C sndNCa VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN31 sndNCa A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP10 VPWR A sndPAb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP11 sndPAb B y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP20 VPWR C sndPCb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP21 sndPCb B y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP30 VPWR A sndPAc VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP31 sndPAc C y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__maj3_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__maj3_4 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN2 X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN10 y B sndNBa VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN11 sndNBa A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN20 y B sndNBc VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN21 sndNBc C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN30 y C sndNCa VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN31 sndNCa A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP10 VPWR A sndPAb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP11 sndPAb B y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP20 VPWR C sndPCb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP21 sndPCb B y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP30 VPWR A sndPAc VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP31 sndPAc C y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__maj3_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
*.PININFO A_N:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C sndC VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN3 sndC D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and4b_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
*.PININFO A_N:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C sndC VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN3 sndC D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and4b_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
*.PININFO A_N:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C sndC VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN3 sndC D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and4b_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a31o_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a31o_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a31o_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
*.PININFO A_N:I B_N:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 B B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C sndC VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN3 sndC D VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 B B_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand4bb_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
*.PININFO A_N:I B_N:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 B B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C sndC VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN3 sndC D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 B B_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand4bb_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
*.PININFO A_N:I B_N:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 A A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 B B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C sndC VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN3 sndC D VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 A A_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 B B_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand4bb_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 y B2 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 sndB1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 sndB1 B2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a22o_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 y B2 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 sndB1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 sndB1 B2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a22o_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 y B2 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 sndB1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 sndB1 B2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a22o_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlrtn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q
*.PININFO D:I GATE_N:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI635 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 M0 clkneg net54 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 Q m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 clkpos GATE_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 m1 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 net54 db VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 net50 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 M0 clkpos net50 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 clkpos GATE_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 Q m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net93 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M0 clkneg net101 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net101 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 m1 M0 net93 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 M0 clkpos net81 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 net81 db VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlrtn_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlrtn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q
*.PININFO D:I GATE_N:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI635 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 M0 clkneg net54 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 Q m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 clkpos GATE_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 m1 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 net54 db VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 net50 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 M0 clkpos net50 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 clkpos GATE_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 Q m1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net93 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M0 clkneg net101 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net101 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 m1 M0 net93 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 M0 clkpos net81 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 net81 db VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlrtn_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlrtn_4 D GATE_N RESET_B VGND VNB VPB VPWR Q
*.PININFO D:I GATE_N:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI635 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 M0 clkneg net55 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 Q m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 clkpos GATE_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 m1 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 net55 db VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 net51 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 M0 clkpos net51 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 clkpos GATE_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 Q m1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net94 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M0 clkneg net102 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net102 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 m1 M0 net94 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 M0 clkpos net82 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 net82 db VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlrtn_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__edfxbp_1 CLK D DE VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I DE:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
XMXNI14 net124 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI13 S0 clkneg net124 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 net68 deneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 Q S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net109 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI643 net92 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI639 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.75 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 S0 clkpos net92 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M0 clkneg net109 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI10 net85 DE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI9 db S1 net85 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 deneg DE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI8 db D net68 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI21 Q_N S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI641 net193 S1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 S0 clkneg net193 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net148 DE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 Q S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net168 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 M0 clkpos net168 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI16 net161 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI15 S0 clkpos net161 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 deneg DE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 db D net148 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI11 db S1 net141 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI12 net141 deneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI22 Q_N S1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__edfxbp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN2 X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnor0 inor A1_N VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnor1 inor A2_N VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi10 VGND B1 sndNB1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi11 sndNB1 B2 y VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi20 y inor VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi20 y inor pmid VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnor0 VPWR A1_N sndPA1N VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnor1 sndPA1N A2_N inor VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi10 pmid B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi11 pmid B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a2bb2o_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN2 X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnor0 inor A1_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnor1 inor A2_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi10 VGND B1 sndNB1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi11 sndNB1 B2 y VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi20 y inor VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi20 y inor pmid VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnor0 VPWR A1_N sndPA1N VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnor1 sndPA1N A2_N inor VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi10 pmid B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi11 pmid B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a2bb2o_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN2 X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnor0 inor A1_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNnor1 inor A2_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi10 VGND B1 sndNB1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi11 sndNB1 B2 y VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNaoi20 y inor VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi20 y inor pmid VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnor0 VPWR A1_N sndPA1N VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPnor1 sndPA1N A2_N inor VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi10 pmid B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPaoi11 pmid B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a2bb2o_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdfxbp_1 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
XMXNI98 db D n0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=3.1
XMXNI103 n1 SCD VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI120 db SCE n1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI104 n0 sceb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI657 M0 clkpos net129 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net129 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI641 net120 S1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 S0 clkneg net120 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 Q S1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI639 sceb SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M1 clkpos S0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI661 Q_N net153 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net153 S1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI94 db D p0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI101 db sceb p1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 S0 clkpos net177 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.75 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net160 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 Q S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q_N net153 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI643 net177 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 M1 clkneg S0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI640 sceb SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M0 clkneg net160 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 net153 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sdfxbp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdfxbp_2 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
XMXNI98 db D n0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=3.1
XMXNI103 n1 SCD VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI120 db SCE n1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI104 n0 sceb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI657 M0 clkpos net129 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net129 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI641 net120 S1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 S0 clkneg net120 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 Q S1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI639 sceb SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M1 clkpos S0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI661 Q_N net153 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net153 S1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI94 db D p0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI101 db sceb p1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 S0 clkpos net196 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.75 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net189 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 Q S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q_N net153 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI643 net196 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 M1 clkneg S0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI640 sceb SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M0 clkneg net189 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 net153 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sdfxbp_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPB1N B1 B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINB1N B1 B1_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a21bo_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPB1N B1 B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINB1N B1 B1_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a21bo_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPB1N B1 B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINB1N B1 B1_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a21bo_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 Y C VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nor3_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 Y C VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nor3_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 Y C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nor3_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__einvp_4 A TE VGND VNB VPB VPWR Z
*.PININFO A:I TE:I VGND:I VNB:I VPB:I VPWR:I Z:O
XMXNMN0 Z A sndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA TE VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 TEB TE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP0 VPWR TEB sndTEB VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=0.94 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndTEB A Z VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 TEB TE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__einvp_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
*.PININFO A:I TE:I VGND:I VNB:I VPB:I VPWR:I Z:O
XMXNMN0 Z A sndA VNB sky130_fd_pr__nfet_01v8 m=8 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA TE VGND VNB sky130_fd_pr__nfet_01v8 m=8 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 TEB TE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP0 VPWR TEB sndTEB VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=0.94 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndTEB A Z VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 TEB TE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__einvp_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__einvp_1 A TE VGND VNB VPB VPWR Z
*.PININFO A:I TE:I VGND:I VNB:I VPB:I VPWR:I Z:O
XMXNMN0 Z A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA TE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 TEB TE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP0 VPWR TEB sndTEB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndTEB A Z VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 TEB TE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__einvp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__einvp_2 A TE VGND VNB VPB VPWR Z
*.PININFO A:I TE:I VGND:I VNB:I VPB:I VPWR:I Z:O
XMXNMN0 Z A sndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA TE VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 TEB TE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP0 VPWR TEB sndTEB VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=0.94 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndTEB A Z VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 TEB TE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__einvp_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 Y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a21oi_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 Y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a21oi_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 Y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a21oi_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdlclkp_1 CLK GATE SCE VGND VNB VPB VPWR GCLK
*.PININFO CLK:I GATE:I SCE:I VGND:I VNB:I VPB:I VPWR:I GCLK:O
XMXNI662 net88 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 M0 clkpos net88 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 net76 CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net76 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI22 net63 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI21 net116 GATE net63 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkpos CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 GCLK net76 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 net116 clkneg M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 net116 clkpos M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 m1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 M0 clkneg net123 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net123 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 net116 SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net112 CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net76 m1 net112 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI23 net116 GATE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkpos CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 GCLK net76 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sdlclkp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdlclkp_2 CLK GATE SCE VGND VNB VPB VPWR GCLK
*.PININFO CLK:I GATE:I SCE:I VGND:I VNB:I VPB:I VPWR:I GCLK:O
XMXNI662 net88 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 M0 clkpos net88 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 net76 CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net76 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI22 net63 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI21 net116 GATE net63 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkpos CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 GCLK net76 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 net116 clkneg M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 net116 clkpos M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 m1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 M0 clkneg net123 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net123 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 net116 SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net112 CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net76 m1 net112 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI23 net116 GATE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkpos CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 GCLK net76 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sdlclkp_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdlclkp_4 CLK GATE SCE VGND VNB VPB VPWR GCLK
*.PININFO CLK:I GATE:I SCE:I VGND:I VNB:I VPB:I VPWR:I GCLK:O
XMXNI662 net88 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 M0 clkpos net88 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 net76 CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net76 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI22 net63 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI21 net116 GATE net63 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 clkpos CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 GCLK net76 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 net116 clkneg M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 net116 clkpos M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 m1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 M0 clkneg net123 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net123 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 net116 SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net112 CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net76 m1 net112 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI23 net116 GATE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 clkpos CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 GCLK net76 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sdlclkp_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlrtp_1 D GATE RESET_B VGND VNB VPB VPWR Q
*.PININFO D:I GATE:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI635 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 M0 clkneg net54 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.36 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 Q m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 clkneg GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 m1 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 net54 db VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 net50 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 M0 clkpos net50 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.36 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 clkneg GATE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 Q m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net93 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M0 clkneg net101 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net101 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 m1 M0 net93 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 M0 clkpos net81 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 net81 db VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlrtp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlrtp_4 D GATE RESET_B VGND VNB VPB VPWR Q
*.PININFO D:I GATE:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI635 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 M0 clkneg net55 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 Q m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 clkneg GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 m1 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 net55 db VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 net51 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 M0 clkpos net51 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 clkneg GATE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 Q m1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net94 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M0 clkneg net102 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net102 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 m1 M0 net94 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 M0 clkpos net82 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 net82 db VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlrtp_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlrtp_2 D GATE RESET_B VGND VNB VPB VPWR Q
*.PININFO D:I GATE:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI635 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 M0 clkneg net54 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 Q m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 clkneg GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 m1 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 net54 db VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 net50 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 M0 clkpos net50 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 clkneg GATE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 Q m1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net93 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M0 clkneg net101 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net101 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 m1 M0 net93 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 M0 clkpos net81 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 net81 db VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlrtp_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 pndC C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPD0 y D1 pndC VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMND0 y D1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a2111o_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 pndC C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPD0 y D1 pndC VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMND0 y D1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a2111o_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 pndC C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPD0 y D1 pndC VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMND0 y D1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a2111o_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__fahcin_1 A B CIN VGND VNB VPB VPWR COUT SUM
*.PININFO A:I B:I CIN:I VGND:I VNB:I VPB:I VPWR:I COUT:O SUM:O
XMXNMIP3 SUM net144 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI32 Bbb Bb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI27 Ab Bb mid2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI26 Abb B mid2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI22 Abb Bb mid1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI23 Ab B mid1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 CINb1 CIN VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI13 CINbb2 CINb2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 Abb Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI12 CINb2 CIN VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI16 Bb B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 CINbb2 mid2 net144 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI1 CINb2 mid1 net144 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI3 Bbb mid2 COUT VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 CINb1 mid1 COUT VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 SUM net144 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 CINb1 mid2 COUT VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI25 Ab B mid2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 Abb Bb mid2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI21 Ab Bb mid1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 Abb B mid1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI14 CINb1 CIN VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI9 CINbb2 CINb2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI8 CINb2 CIN VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 Abb Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 Bb B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 CINbb2 mid1 net144 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI2 CINb2 mid2 net144 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI31 Bbb mid1 COUT VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 Bbb Bb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__fahcin_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_6 KAPWR VGND VNB VPB VPWR
*.PININFO KAPWR:I VGND:I VNB:I VPB:I VPWR:I
XMXNI1 VGND KAPWR VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.55 l=1.97 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI2 KAPWR VGND KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.87 l=1.97
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_decapkapwr_6


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_3 KAPWR VGND VNB VPB VPWR
*.PININFO KAPWR:I VGND:I VNB:I VPB:I VPWR:I
XMXNI1 VGND KAPWR VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.55 l=0.59 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI2 KAPWR VGND KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.87 l=0.59
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_decapkapwr_3


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_12 KAPWR VGND VNB VPB VPWR
*.PININFO KAPWR:I VGND:I VNB:I VPB:I VPWR:I
XMXNI1 VGND KAPWR VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.55 l=4.73 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI2 KAPWR VGND KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.87 l=4.73
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_decapkapwr_12


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_8 KAPWR VGND VNB VPB VPWR
*.PININFO KAPWR:I VGND:I VNB:I VPB:I VPWR:I
XMXNI1 VGND KAPWR VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.55 l=2.89 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI2 KAPWR VGND KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.87 l=2.89
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_decapkapwr_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_4 KAPWR VGND VNB VPB VPWR
*.PININFO KAPWR:I VGND:I VNB:I VPB:I VPWR:I
XMXNI1 VGND KAPWR VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.55 l=1.05 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI2 KAPWR VGND KAPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.87 l=1.05
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_decapkapwr_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 y C1 pndB VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o311a_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 y C1 pndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o311a_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 y C1 pndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o311a_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdfrtn_1 CLK_N D RESET_B SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK_N:I D:I RESET_B:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I
*.PININFO Q:O
XMXNI642 clkpos CLK_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net87 net153 net117 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net117 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 net110 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 sceb SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 M0 clkpos net98 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 net98 M1 net110 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 net153 clkneg net93 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 Q net87 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net93 net87 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 M1 clkpos net153 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI98 db D n0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=3.1
XMXNI103 n1 SCD VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.18 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI120 db SCE n1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI104 n0 sceb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI643 clkpos CLK_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net190 net87 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 net87 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 net153 clkpos net190 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net87 net153 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI30 net169 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI31 M0 clkneg net169 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI32 net169 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI660 Q net87 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 M1 clkneg net153 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 sceb SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI101 db sceb p1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI94 db D p0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sdfrtn_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sedfxbp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I DE:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O
*.PININFO Q_N:O
XMXNI14 net155 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI13 S0 clkneg net155 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 Q S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net144 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI643 net127 q1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI639 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.75 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 S0 clkpos net127 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M0 clkneg net144 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 q1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 net116 deneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 net107 sceneg db VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 VPWR SCD net107 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI31 net104 D net116 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 net104 SCE db VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI40 net87 q1 net104 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI36 deneg DE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI38 VPWR DE net87 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 sceneg SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI52 Q_N q1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI641 net240 q1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 S0 clkneg net240 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 Q S0 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net224 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 M0 clkpos net224 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 net104 sceneg db VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 q1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 sceneg SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI32 net104 D net180 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI16 net200 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI15 S0 clkpos net200 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI41 net192 q1 net104 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI39 VGND deneg net192 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI37 deneg DE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 net180 DE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI49 net176 SCE db VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI48 VGND SCD net176 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI53 Q_N q1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sedfxbp_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sedfxbp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I DE:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O
*.PININFO Q_N:O
XMXNI14 net155 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI13 S0 clkneg net155 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 Q S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net123 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI643 net127 q1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI639 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.75 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 S0 clkpos net127 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M0 clkneg net123 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 q1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 net116 deneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 net107 sceneg db VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 VPWR SCD net107 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI31 net104 D net116 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 net104 SCE db VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI40 net87 q1 net104 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI36 deneg DE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI38 VPWR DE net87 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 sceneg SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI52 Q_N q1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI641 net235 q1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 S0 clkneg net235 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 Q S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net224 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 M0 clkpos net224 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 net104 sceneg db VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 q1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 sceneg SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI32 net104 D net203 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI16 net200 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI15 S0 clkpos net200 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI41 net192 q1 net104 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI39 VGND deneg net192 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI37 deneg DE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 net203 DE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI49 net176 SCE db VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI48 VGND SCD net176 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI53 Q_N q1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sedfxbp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 Y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a31oi_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 Y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a31oi_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 Y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a31oi_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
*.PININFO D:I GATE:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI635 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 M0 clkneg net51 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 Q m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 clkneg GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 net51 db VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 net47 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 M0 clkpos net47 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 clkneg GATE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 Q m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M0 clkneg net94 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net94 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 m1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 M0 clkpos net74 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 net74 db VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlxtp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__clkdlybuf4s18_2 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 A2 Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.18 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 Ab2 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.18 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 X Ab2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 A2 Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.82 l=0.18 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 Ab2 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.82 l=0.18 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 X Ab2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__clkdlybuf4s18_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__clkdlybuf4s18_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 A2 Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.18 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 Ab2 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.18 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 X Ab2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 A2 Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.82 l=0.18 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 Ab2 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.82 l=0.18 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 X Ab2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__clkdlybuf4s18_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C sndC VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN3 sndC D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and4_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C sndC VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN3 sndC D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and4_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B sndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN2 sndB C sndC VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN3 sndC D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN0 X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__and4_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o21a_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o21a_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o21a_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__probe_p_8 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=3 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 net29 Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=3 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 net29 Ab VGND VNB sky130_fd_pr__nfet_01v8 m=8 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
rI112 net29 X sky130_fd_pr__res_generic_po
.ENDS sky130_fd_sc_hd__probe_p_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMIN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=6 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__clkinv_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMIN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=3 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__clkinv_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMIN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__clkinv_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMIN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=8 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=12 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__clkinv_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMIN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=16 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=24 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__clkinv_16


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdfrtp_4 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I RESET_B:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I
*.PININFO Q:O
XMXNI642 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net84 S0 net114 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net114 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 net107 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 sceb SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 M0 clkpos net95 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 net95 M1 net107 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 S0 clkneg net90 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 Q net84 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net90 net84 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 M1 clkpos S0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI98 db D n0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=3.1
XMXNI103 n1 SCD VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.18 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI120 db SCE n1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI104 n0 sceb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI643 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net187 net84 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 net84 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 S0 clkpos net187 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net84 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI30 net166 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI31 M0 clkneg net166 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI32 net166 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 Q net84 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 M1 clkneg S0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 sceb SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI101 db sceb p1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI94 db D p0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sdfrtp_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I RESET_B:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I
*.PININFO Q:O
XMXNI642 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net84 S0 net114 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net114 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 net107 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 sceb SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 M0 clkpos net95 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 net95 M1 net107 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 S0 clkneg net90 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 Q net84 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net90 net84 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 M1 clkpos S0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI98 db D n0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=3.1
XMXNI103 n1 SCD VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.18 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI120 db SCE n1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI104 n0 sceb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI643 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net187 net84 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 net84 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 S0 clkpos net187 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net84 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI30 net166 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI31 M0 clkneg net166 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI32 net166 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 Q net84 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 M1 clkneg S0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 sceb SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI101 db sceb p1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI94 db D p0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sdfrtp_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I RESET_B:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I
*.PININFO Q:O
XMXNI642 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net84 S0 net114 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net114 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 net107 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 sceb SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 M0 clkpos net95 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 net95 M1 net107 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 S0 clkneg net83 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 Q net84 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net83 net84 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 M1 clkpos S0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI98 db D n0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=3.1
XMXNI103 n1 SCD VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.18 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI120 db SCE n1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI104 n0 sceb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI643 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net187 net84 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 net84 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 S0 clkpos net187 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net84 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI30 net166 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI31 M0 clkneg net166 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI32 net166 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 Q net84 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 M1 clkneg S0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 sceb SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI101 db sceb p1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI94 db D p0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sdfrtp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__xor3_4 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIP3 X net117 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 mid1 Cb net117 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI1 mid2 C net117 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 Cb C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 Abb Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 mid1 Bb Ab VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI16 Bb B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI23 mid1 B Abb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI26 mid2 Bb Abb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI27 mid2 B Ab VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 X net117 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 Cb C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 mid1 C net117 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI2 mid2 Cb net117 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 Abb Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 Bb B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 Ab B mid1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI25 Abb Bb mid1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI28 Abb B mid2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI29 Ab Bb mid2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.6 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__xor3_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__xor3_2 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIP3 X net117 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 mid1 Cb net117 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI1 mid2 C net117 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 Cb C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 Abb Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 mid1 Bb Ab VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI16 Bb B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI23 mid1 B Abb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI26 mid2 Bb Abb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI27 mid2 B Ab VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 X net117 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 Cb C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 mid1 C net117 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI2 mid2 Cb net117 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 Abb Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 Bb B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 Ab B mid1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI25 Abb Bb mid1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI28 Abb B mid2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI29 Ab Bb mid2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.6 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__xor3_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__xor3_1 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIP3 X net117 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 mid1 Cb net117 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI1 mid2 C net117 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 Cb C VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI45 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI47 Abb Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 mid1 Bb Ab VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI16 Bb B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI23 mid1 B Abb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI26 mid2 Bb Abb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI27 mid2 B Ab VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 X net117 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 Cb C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 mid1 C net117 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI2 mid2 Cb net117 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI44 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI46 Abb Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 Bb B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 Ab B mid1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI25 Abb Bb mid1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI28 Abb B mid2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI29 Ab Bb mid2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.6 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__xor3_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 sndB1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 sndB1 B2 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 pndB B2 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 y C1 pndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o221a_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 sndB1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 sndB1 B2 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 pndB B2 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 y C1 pndB VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o221a_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 sndB1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 sndB1 B2 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 pndB B2 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 y C1 pndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o221a_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
*.PININFO A0:I A1:I A2:I A3:I S0:I S1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMNA00 sndNS0ba0 S0b xlowb VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNA01 VGND A0 sndNS0ba0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNA10 sndNS0a1 S0 xlowb VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNA11 VGND A1 sndNS0a1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNA20 sndNS0ba2 S0b xhib VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNA21 VGND A2 sndNS0ba2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNA30 sndNS0a3 S0 xhib VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNA31 VGND A3 sndNS0a3 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNs1o xb S1b xlowb VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNs2o xb S1 xhib VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMIN1 VGND S1 S1b VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMIN2 VGND S0 S0b VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMIN4 VGND xb X VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA00 sndPA0a0 A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA01 xlowb S0 sndPA0a0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA10 sndPA1a1 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA11 xlowb S0b sndPA1a1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA20 sndPA2a2 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA21 xhib S0 sndPA2a2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA30 sndPA3a3 A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA31 xhib S0b sndPA3a3 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPs1o xb S1 xlowb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPs2o xb S1b xhib VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMIP1 VPWR S1 S1b VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMIP2 VPWR S0 S0b VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMIP4 VPWR xb X VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
.ENDS sky130_fd_sc_hd__mux4_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__mux4_4 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
*.PININFO A0:I A1:I A2:I A3:I S0:I S1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMNA00 sndNS0ba0 S0b xlowb VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNA01 VGND A0 sndNS0ba0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNA10 sndNS0a1 S0 xlowb VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNA11 VGND A1 sndNS0a1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNA20 sndNS0ba2 S0b xhib VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNA21 VGND A2 sndNS0ba2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNA30 sndNS0a3 S0 xhib VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNA31 VGND A3 sndNS0a3 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNs1o xb S1b xlowb VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNs2o xb S1 xhib VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMIN1 VGND S1 S1b VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMIN2 VGND S0 S0b VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMIN4 VGND xb X VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA00 sndPA0a0 A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA01 xlowb S0 sndPA0a0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA10 sndPA1a1 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA11 xlowb S0b sndPA1a1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA20 sndPA2a2 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA21 xhib S0 sndPA2a2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA30 sndPA3a3 A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA31 xhib S0b sndPA3a3 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPs1o xb S1 xlowb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPs2o xb S1b xhib VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMIP1 VPWR S1 S1b VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMIP2 VPWR S0 S0b VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMIP4 VPWR xb X VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
.ENDS sky130_fd_sc_hd__mux4_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
*.PININFO A0:I A1:I A2:I A3:I S0:I S1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMNA00 sndNS0ba0 S0b xlowb VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNA01 VGND A0 sndNS0ba0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNA10 sndNS0a1 S0 xlowb VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNA11 VGND A1 sndNS0a1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNA20 sndNS0ba2 S0b xhib VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNA21 VGND A2 sndNS0ba2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNA30 sndNS0a3 S0 xhib VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNA31 VGND A3 sndNS0a3 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNs1o xb S1b xlowb VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMNs2o xb S1 xhib VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMIN1 VGND S1 S1b VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMIN2 VGND S0 S0b VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMIN4 VGND xb X VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA00 sndPA0a0 A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA01 xlowb S0 sndPA0a0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA10 sndPA1a1 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA11 xlowb S0b sndPA1a1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA20 sndPA2a2 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA21 xhib S0 sndPA2a2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA30 sndPA3a3 A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPA31 xhib S0b sndPA3a3 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPs1o xb S1 xlowb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMPs2o xb S1b xhib VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMIP1 VPWR S1 S1b VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMIP2 VPWR S0 S0b VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXNMIP4 VPWR xb X VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
.ENDS sky130_fd_sc_hd__mux4_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__fa_2 A B CIN VGND VNB VPB VPWR COUT SUM
*.PININFO A:I B:I CIN:I VGND:I VNB:I VPB:I VPWR:I COUT:O SUM:O
XMXNMNs1s nint1 majb sumb VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 COUT majb VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 SUM sumb VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNmaj10 majb B sndNAp1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNmaj11 sndNAp1 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNmaj30 majb CIN nmajmid VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNmaj21 nmajmid A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNmaj20 VGND B nmajmid VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs2s0 VGND A sndNAn4 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs2s1 sndNAn4 B sndNBn4 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs2s2 sndNBn4 CIN sumb VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs3s0 nint1 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs3s1 nint1 B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs3s2 nint1 CIN VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 COUT majb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 SUM sumb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPmaj10 VPWR A sndPAp1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.63 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPmaj11 sndPAp1 B majb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.63 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPmaj20 VPWR B pmajmid VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.63 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPmaj30 pmajmid CIN majb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.63 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPmaj21 pmajmid A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.63 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs2s0 VPWR A sndPAp4 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.63 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs2s1 sndPAp4 B sndPBp4 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.63 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs2s2 sndPBp4 CIN sumb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs3s0 pint1 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs3s1 pint1 B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs3s2 pint1 CIN VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs1s pint1 majb sumb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__fa_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM
*.PININFO A:I B:I CIN:I VGND:I VNB:I VPB:I VPWR:I COUT:O SUM:O
XMXNMNs1s nint1 majb sumb VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 COUT majb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 SUM sumb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNmaj10 majb B sndNAp1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNmaj11 sndNAp1 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNmaj30 majb CIN sndNCINn3 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNmaj31 sndNCINn3 B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNmaj20 VGND A sndNCINn3 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs2s0 VGND A sndNAn4 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs2s1 sndNAn4 B sndNBn4 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs2s2 sndNBn4 CIN sumb VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs3s0 nint1 B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs3s1 nint1 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs3s2 nint1 CIN VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 COUT majb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 SUM sumb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPmaj10 VPWR A sndPAp1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPmaj11 sndPAp1 B majb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPmaj20 VPWR A sndPCINp3 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPmaj21 sndPCINp3 CIN majb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPmaj31 sndPCINp3 B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs2s0 VPWR A sndPAp4 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs2s1 sndPAp4 B sndPBp4 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs2s2 sndPBp4 CIN sumb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs3s0 pint1 B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs3s1 pint1 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs3s2 pint1 CIN VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs1s pint1 majb sumb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__fa_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__fa_4 A B CIN VGND VNB VPB VPWR COUT SUM
*.PININFO A:I B:I CIN:I VGND:I VNB:I VPB:I VPWR:I COUT:O SUM:O
XMXNMNs1s nint1 majb sumb VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 COUT majb VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 SUM sumb VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNmaj10 majb B sndNAp1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNmaj11 sndNAp1 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNmaj30 majb CIN nmajmid VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNmaj21 nmajmid A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNmaj20 VGND B nmajmid VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs2s0 VGND A sndNAn4 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs2s1 sndNAn4 B sndNBn4 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs2s2 sndNBn4 CIN sumb VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs3s0 nint1 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs3s1 nint1 B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNs3s2 nint1 CIN VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 COUT majb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 SUM sumb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPmaj10 VPWR A sndPAp1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.63 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPmaj11 sndPAp1 B majb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.63 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPmaj20 VPWR B pmajmid VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPmaj30 pmajmid CIN majb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPmaj21 pmajmid A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs2s0 VPWR A sndPAp4 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.63 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs2s1 sndPAp4 B sndPBp4 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.63 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs2s2 sndPBp4 CIN sumb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs3s0 pint1 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs3s1 pint1 B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs3s2 pint1 CIN VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPs1s pint1 majb sumb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__fa_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__mux2i_1 A0 A1 S VGND VNB VPB VPWR Y
*.PININFO A0:I A1:I S:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMNA00 Y A0 smdNA0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA01 smdNA0 Sb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA10 Y A1 sndNA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA11 sndNA1 S VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 Sb S VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA00 VPWR S sndPS VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA01 sndPS A0 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA10 VPWR Sb sndPSb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA11 sndPSb A1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Sb S VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__mux2i_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__mux2i_4 A0 A1 S VGND VNB VPB VPWR Y
*.PININFO A0:I A1:I S:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMNA00 Y A0 smdNA0 VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA01 smdNA0 Sb VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA10 Y A1 sndNA1 VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA11 sndNA1 S VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 Sb S VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA00 VPWR S sndPS VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA01 sndPS A0 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA10 VPWR Sb sndPSb VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA11 sndPSb A1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Sb S VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__mux2i_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__mux2i_2 A0 A1 S VGND VNB VPB VPWR Y
*.PININFO A0:I A1:I S:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMNA00 Y A0 smdNA0 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA01 smdNA0 Sb VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA10 Y A1 sndNA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA11 sndNA1 S VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 Sb S VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA00 VPWR S sndPS VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA01 sndPS A0 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA10 VPWR Sb sndPSb VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA11 sndPSb A1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Sb S VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__mux2i_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand2_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand2_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=8 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B VGND VNB sky130_fd_pr__nfet_01v8 m=8 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand2_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA B VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nand2_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 Y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 Y B2 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 sndB1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 sndB1 B2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a32oi_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 Y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 Y B2 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 sndB1 VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 sndB1 B2 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a32oi_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 Y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 Y B2 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 sndB1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 sndB1 B2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a32oi_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_inputisolatch_1 D SLEEP_B VGND VNB VPB VPWR Q
*.PININFO D:I SLEEP_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI677 Q s0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 sleepneg sleeppos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI674 net39 s0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 s0 sleepneg net49 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 net49 D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 s0 sleeppos net38 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net38 net39 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI670 sleeppos SLEEP_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI643 sleeppos SLEEP_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.55 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 sleepneg sleeppos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.55 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal
+ perim=1.14
XMXNI662 net86 net39 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 s0 sleepneg net86 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net39 s0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 Q s0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 s0 sleeppos net69 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 net69 D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_inputisolatch_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o21ai_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o21ai_0 A1 A2 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o21ai_0


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o21ai_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.7 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o21ai_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlrbn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
*.PININFO D:I GATE_N:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
XMXNI635 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 Q_N net125 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 M0 clkneg net61 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 net125 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 Q m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 clkpos GATE_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 m1 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 net61 db VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 net57 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 M0 clkpos net57 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 clkpos GATE_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 Q_N net125 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 Q m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 net125 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net108 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M0 clkneg net116 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net116 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 m1 M0 net108 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 M0 clkpos net96 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 net96 db VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlrbn_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlrbn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
*.PININFO D:I GATE_N:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
XMXNI635 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 Q_N net125 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 M0 clkneg net61 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 net125 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 Q m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 clkpos GATE_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 m1 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 net61 db VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 net57 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 M0 clkpos net57 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 clkpos GATE_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 Q_N net125 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 Q m1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 net125 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net108 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M0 clkneg net116 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net116 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 m1 M0 net108 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 M0 clkpos net96 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 net96 db VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlrbn_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_inputiso0p_1 A SLEEP VGND VNB VPB VPWR X
*.PININFO A:I SLEEP:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNI8 net36 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 net36 sleepb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 X net36 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 sleepb SLEEP VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI10 net36 sleepb sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI21 X net36 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 sleepb SLEEP VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI11 sndA A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_inputiso0p_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMIP1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=8 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__inv_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMIN1 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=16 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=16 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__inv_16


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMIP1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__inv_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMIN1 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__inv_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMIN1 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=6 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=6 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__inv_6


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMIN1 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__inv_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMIN1 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=12 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=12 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__inv_12


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 sndB1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 sndB1 B2 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 y B2 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o32a_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 sndB1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 sndB1 B2 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 y B2 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o32a_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 sndB1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 sndB1 B2 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 y B2 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o32a_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__tap_1 VGND VNB VPB VPWR
*.PININFO VGND:I VNB:I VPB:I VPWR:I
* Notes: Tap pins in this cell are not connected to power buses.
.ENDS sky130_fd_sc_hd__tap_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__tap_2 VGND VNB VPB VPWR
*.PININFO VGND:I VNB:I VPB:I VPWR:I
* Notes: Tap pins in this cell are not connected to power buses.
.ENDS sky130_fd_sc_hd__tap_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlxbn_1 D GATE_N VGND VNB VPB VPWR Q Q_N
*.PININFO D:I GATE_N:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
XMXNI635 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 Q_N net112 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 M0 clkneg net56 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 net112 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 Q m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 clkpos GATE_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 net56 db VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 net52 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 M0 clkpos net52 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 clkpos GATE_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 Q_N net112 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 Q m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 net112 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M0 clkneg net107 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net107 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 m1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 M0 clkpos net87 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 net87 db VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlxbn_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlxbn_2 D GATE_N VGND VNB VPB VPWR Q Q_N
*.PININFO D:I GATE_N:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
XMXNI635 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 Q_N net114 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 M0 clkneg net58 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 net114 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 Q m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 clkpos GATE_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 net58 db VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI653 net54 m1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 M0 clkpos net54 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 m1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 db D VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 clkpos GATE_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 Q_N net114 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 Q m1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 net114 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 M0 clkneg net109 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net109 m1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 m1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkneg clkpos VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 db D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 M0 clkpos net89 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 net89 db VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlxbn_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__buf_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=3 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=8 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=3 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__buf_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=6 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=6 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__buf_6


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.52 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.52 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.79 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.79 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__buf_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__buf_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__buf_16 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=6 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=16 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=6 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=16 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__buf_16


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X Ab VGND VNB sky130_fd_pr__nfet_01v8 m=12 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=12 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__buf_12


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPB1N B1 B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINB1N B1 B1_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o21ba_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPB1N B1 B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINB1N B1 B1_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o21ba_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPB1N B1 B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINB1N B1 B1_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o21ba_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4 A LOWLVPWR VGND VNB VPB VPWR X
*.PININFO A:I LOWLVPWR:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNI2 net72 cross1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.79 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI3 cross1 net72 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.79 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI20 Ab A LOWLVPWR LOWLVPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI24 X net60 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI28 net60 cross1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.79 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 cross1 Ab VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 net72 A VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI23 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI25 X net60 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI29 net60 cross1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMIN1 Ab net55 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 net59 Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 net55 net47 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI15 net51 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI9 net47 X VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI16 X net51 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Ab net55 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 net59 Ab VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 net55 net47 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI8 net47 X VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 X net51 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 net51 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__dlymetal6s2s_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPD0 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 pndC C1 pndB VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMND0 Y D1 pndC VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o2111ai_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPD0 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 pndC C1 pndB VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMND0 Y D1 pndC VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o2111ai_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPD0 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 pndB B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 pndC C1 pndB VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMND0 Y D1 pndC VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o2111ai_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I D_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C sndPC VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 sndPC D Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 D D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 Y C VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN3 Y D VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN3 D D_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nor4b_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I D_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C sndPC VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 sndPC D Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 D D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 Y C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN3 Y D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN3 D D_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nor4b_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I D_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C sndPC VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 sndPC D Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 D D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 Y C VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN3 Y D VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN3 D D_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nor4b_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2 A VGND VPB VPWRIN VPWR X
*.PININFO A:I VGND:I VPB:I VPWRIN:I VPWR:I X:O
XMXN1000 VPWR a_620_911# a_714_47# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
+ ad=8.352e+11p pd=7.41e+06u as=2.1725e+11p ps=2.13e+06u
XMXN1001 a_1032_911# a_620_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
XMXN1002 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.62905e+12p ps=1.514e+07u
XMXN1003 a_714_47# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
XMXN1004 a_714_47# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
XMXN1005 X a_1032_911# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=2.405e+11p pd=2.04e+06u as=0p ps=0u
XMXN1006 VPWR a_1032_911# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=3.7e+11p ps=2.74e+06u
XMXN1007 VGND A a_714_47# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
XMXN1008 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
XMXN1009 a_1032_911# a_620_911# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
XMXN1010 VGND A a_714_47# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
XMXN1011 a_505_297# A VPWRIN VPWRIN sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
XMXN1012 a_505_297# A VGND VGND sky130_fd_pr__nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
XMXN1013 X a_1032_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
XMXN1014 VGND a_1032_911# X VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
XMXN1015 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
XMXN1016 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
XMXN1017 VPWR a_714_47# a_620_911# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1 A VGND VPB VPWRIN VPWR X
*.PININFO A:I VGND:I VPB:I VPWRIN:I VPWR:I X:O
XMXN1000 X a_1028_32# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
+ ad=2.1725e+11p pd=2.13e+06u as=4.7795e+11p ps=4.37e+06u
XMXN1001 VPWR a_620_911# a_714_58# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
XMXN1002 a_1028_32# a_620_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
+ ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
XMXN1003 X a_1028_32# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=1.8525e+11p pd=1.87e+06u as=1.4178e+12p ps=1.319e+07u
XMXN1004 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=0p ps=0u
XMXN1005 a_714_58# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
XMXN1006 a_714_58# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
XMXN1007 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
XMXN1008 a_1028_32# a_620_911# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
XMXN1009 a_505_297# A VPWRIN VPWRIN sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
XMXN1010 a_505_297# A VGND VGND sky130_fd_pr__nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
XMXN1011 VGND A a_714_58# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
XMXN1012 VGND A a_714_58# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
XMXN1013 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
XMXN1014 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
XMXN1015 VPWR a_714_58# a_620_911# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4 A VGND VPB VPWRIN VPWR X
*.PININFO A:I VGND:I VPB:I VPWRIN:I VPWR:I X:O
XMXN1000 VPWR a_620_911# a_714_47# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
+ ad=1.1152e+12p pd=9.97e+06u as=2.1725e+11p ps=2.13e+06u
XMXN1001 a_1032_911# a_620_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
XMXN1002 X a_1032_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
+ ad=6.5e+11p pd=5.3e+06u as=0p ps=0u
XMXN1003 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.81105e+12p ps=1.7e+07u
XMXN1004 a_714_47# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
XMXN1005 a_714_47# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
XMXN1006 X a_1032_911# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=4.225e+11p pd=3.9e+06u as=0p ps=0u
XMXN1007 X a_1032_911# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
XMXN1008 VPWR a_1032_911# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
XMXN1009 VGND A a_714_47# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
XMXN1010 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
XMXN1011 a_1032_911# a_620_911# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
XMXN1012 VGND A a_714_47# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
XMXN1013 a_505_297# A VPWRIN VPWRIN sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
XMXN1014 a_505_297# A VGND VGND sky130_fd_pr__nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
XMXN1015 X a_1032_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
XMXN1016 VPWR a_1032_911# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
XMXN1017 VGND a_1032_911# X VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
XMXN1018 VGND a_1032_911# X VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
XMXN1019 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
XMXN1020 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
XMXN1021 VPWR a_714_47# a_620_911# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 sndB1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 sndB1 B2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 Y B2 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o22ai_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 sndB1 VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 sndB1 B2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 Y B2 pndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o22ai_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 sndB1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 sndB1 B2 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 Y B2 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o22ai_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__edfxtp_1 CLK D DE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I DE:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXNI14 net115 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI13 S0 clkneg net115 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 net59 deneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI651 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI645 Q S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net79 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI643 net83 S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI639 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.75 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI644 S0 clkpos net83 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 M0 clkneg net79 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI10 net76 DE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 S1 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI9 db S1 net76 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 deneg DE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI8 db D net59 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI641 net175 S1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI642 S0 clkneg net175 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net172 DE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI646 Q S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net160 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 M0 clkpos net160 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI18 S1 S0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI16 net148 M1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI15 S0 clkpos net148 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 deneg DE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI7 db D net172 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI11 db S1 net128 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI12 net128 deneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__edfxtp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
*.PININFO A:I TE_B:I VGND:I VNB:I VPB:I VPWR:I Z:O
XMXNMN0 Z net35 sndA VNB sky130_fd_pr__nfet_01v8 m=8 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA net39 VGND VNB sky130_fd_pr__nfet_01v8 m=8 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 net39 TE_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 net35 A VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP0 VPWR TE_B sndTEB VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=0.94 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndTEB net35 Z VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 net39 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 net35 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__ebufn_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
*.PININFO A:I TE_B:I VGND:I VNB:I VPB:I VPWR:I Z:O
XMXNMN0 Z net35 sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA net39 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 net39 TE_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 net35 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP0 VPWR TE_B sndTEB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndTEB net35 Z VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 net39 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 net35 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__ebufn_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
*.PININFO A:I TE_B:I VGND:I VNB:I VPB:I VPWR:I Z:O
XMXNMN0 Z net35 sndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA net39 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 net39 TE_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 net35 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP0 VPWR TE_B sndTEB VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=0.94 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndTEB net35 Z VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 net39 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 net35 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__ebufn_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__ebufn_4 A TE_B VGND VNB VPB VPWR Z
*.PININFO A:I TE_B:I VGND:I VNB:I VPB:I VPWR:I Z:O
XMXNMN0 Z net35 sndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA net39 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 net39 TE_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI6 net35 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP0 VPWR TE_B sndTEB VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=0.94 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndTEB net35 Z VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 net39 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI5 net35 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__ebufn_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
*.PININFO A:I B:I C_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 C C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 Y C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN2 C C_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nor3b_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
*.PININFO A:I B:I C_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 C C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 Y C VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN2 C C_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nor3b_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
*.PININFO A:I B:I C_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 C C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 Y C VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN2 C C_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__nor3b_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__einvn_0 A TE_B VGND VNB VPB VPWR Z
*.PININFO A:I TE_B:I VGND:I VNB:I VPB:I VPWR:I Z:O
XMXNMN0 Z A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA net25 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 net25 TE_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP0 VPWR TE_B sndTEB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndTEB A Z VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 net25 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__einvn_0


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__einvn_8 A TE_B VGND VNB VPB VPWR Z
*.PININFO A:I TE_B:I VGND:I VNB:I VPB:I VPWR:I Z:O
XMXNMN0 Z A sndA VNB sky130_fd_pr__nfet_01v8 m=8 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA TE VGND VNB sky130_fd_pr__nfet_01v8 m=8 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 TE TE_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP0 VPWR TE_B sndTEB VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=0.94 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndTEB A Z VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 TE TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__einvn_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__einvn_4 A TE_B VGND VNB VPB VPWR Z
*.PININFO A:I TE_B:I VGND:I VNB:I VPB:I VPWR:I Z:O
XMXNMN0 Z A sndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA TE VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 TE TE_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP0 VPWR TE_B sndTEB VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=0.94 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndTEB A Z VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 TE TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__einvn_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__einvn_2 A TE_B VGND VNB VPB VPWR Z
*.PININFO A:I TE_B:I VGND:I VNB:I VPB:I VPWR:I Z:O
XMXNMN0 Z A sndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA TE VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 TE TE_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP0 VPWR TE_B sndTEB VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=0.94 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndTEB A Z VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 TE TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__einvn_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__einvn_1 A TE_B VGND VNB VPB VPWR Z
*.PININFO A:I TE_B:I VGND:I VNB:I VPB:I VPWR:I Z:O
XMXNMN0 Z A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 sndA net25 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 net25 TE_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP0 VPWR TE_B sndTEB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndTEB A Z VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 net25 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__einvn_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2 A LOWLVPWR VGND VPB VPWR X
*.PININFO A:I LOWLVPWR:I VGND:I VPB:I VPWR:I X:O
XMXN1000 VPWR a_620_911# a_714_47# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
+ ad=8.352e+11p pd=7.41e+06u as=2.1725e+11p ps=2.13e+06u
XMXN1001 a_1032_911# a_620_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
XMXN1002 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.62905e+12p ps=1.514e+07u
XMXN1003 a_714_47# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
XMXN1004 a_714_47# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
XMXN1005 X a_1032_911# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=2.405e+11p pd=2.04e+06u as=0p ps=0u
XMXN1006 VPWR a_1032_911# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=3.7e+11p ps=2.74e+06u
XMXN1007 VGND A a_714_47# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
XMXN1008 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
XMXN1009 a_1032_911# a_620_911# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
XMXN1010 VGND A a_714_47# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
XMXN1011 a_505_297# A LOWLVPWR LOWLVPWR sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
XMXN1012 a_505_297# A VGND VGND sky130_fd_pr__nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
XMXN1013 X a_1032_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
XMXN1014 VGND a_1032_911# X VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
XMXN1015 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
XMXN1016 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
XMXN1017 VPWR a_714_47# a_620_911# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4 A LOWLVPWR VGND VPB VPWR X
*.PININFO A:I LOWLVPWR:I VGND:I VPB:I VPWR:I X:O
XMXN1000 VPWR a_620_911# a_714_47# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
+ ad=1.1152e+12p pd=9.97e+06u as=2.1725e+11p ps=2.13e+06u
XMXN1001 a_1032_911# a_620_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
XMXN1002 X a_1032_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
+ ad=6.5e+11p pd=5.3e+06u as=0p ps=0u
XMXN1003 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.81105e+12p ps=1.7e+07u
XMXN1004 a_714_47# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
XMXN1005 a_714_47# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
XMXN1006 X a_1032_911# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=4.225e+11p pd=3.9e+06u as=0p ps=0u
XMXN1007 X a_1032_911# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
XMXN1008 VPWR a_1032_911# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
XMXN1009 VGND A a_714_47# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
XMXN1010 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
XMXN1011 a_1032_911# a_620_911# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
XMXN1012 VGND A a_714_47# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
XMXN1013 a_505_297# A LOWLVPWR LOWLVPWR sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
XMXN1014 a_505_297# A VGND VGND sky130_fd_pr__nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
XMXN1015 X a_1032_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
XMXN1016 VPWR a_1032_911# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
XMXN1017 VGND a_1032_911# X VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
XMXN1018 VGND a_1032_911# X VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
XMXN1019 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
XMXN1020 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
XMXN1021 VPWR a_714_47# a_620_911# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1 A LOWLVPWR VGND VPB VPWR X
*.PININFO A:I LOWLVPWR:I VGND:I VPB:I VPWR:I X:O
XMXN1000 X a_1028_32# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
+ ad=2.1725e+11p pd=2.13e+06u as=4.7795e+11p ps=4.37e+06u
XMXN1001 VPWR a_620_911# a_714_58# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
XMXN1002 a_1028_32# a_620_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
+ ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
XMXN1003 X a_1028_32# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=1.8525e+11p pd=1.87e+06u as=1.4178e+12p ps=1.319e+07u
XMXN1004 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=0p ps=0u
XMXN1005 a_714_58# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
XMXN1006 a_714_58# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
XMXN1007 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
XMXN1008 a_1028_32# a_620_911# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
XMXN1009 a_505_297# A LOWLVPWR LOWLVPWR sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
XMXN1010 a_505_297# A VGND VGND sky130_fd_pr__nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
XMXN1011 VGND A a_714_58# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
XMXN1012 VGND A a_714_58# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
XMXN1013 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
XMXN1014 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
XMXN1015 VPWR a_714_58# a_620_911# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA3 pndA A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 sndA3 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA3 sndA3 A4 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a41o_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA3 pndA A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 sndA3 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA3 sndA3 A4 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a41o_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 pndA A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA3 pndA A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPX X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 sndA2 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 sndA2 A3 sndA3 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA3 sndA3 A4 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINX X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a41o_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 net40 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 net40 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 Y B1 net40 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPB1N B1 B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINB1N B1 B1_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a21boi_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 net40 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 net40 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 Y B1 net40 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPB1N B1 B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINB1N B1 B1_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a21boi_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a21boi_0 A1 A2 B1_N VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 net40 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 net40 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 Y B1 net40 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPB1N B1 B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINB1N B1 B1_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a21boi_0


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 net40 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 net40 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 Y B1 net40 VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIPB1N B1 B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMINB1N B1 B1_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a21boi_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 Y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 Y B2 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 sndB1 VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 sndB1 B2 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a22oi_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 Y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 Y B2 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 sndB1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 sndB1 B2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a22oi_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 Y B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB1 Y B2 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 sndB1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB1 sndB1 B2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a22oi_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
*.PININFO VGND:I VPWR:I
* Notes: substrate is tied to vgnd and well is tied to vpwr in the
*        cell and do not appear as pins.
.ENDS sky130_fd_sc_hd__tapvpwrvgnd_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__lpflow_inputiso0n_1 A SLEEP_B VGND VNB VPB VPWR X
*.PININFO A:I SLEEP_B:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNI14 X net36 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 net36 A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI13 sndA SLEEP_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 net36 SLEEP_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI19 X net36 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI17 net36 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__lpflow_inputiso0n_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
*.PININFO A:I B:I C_N:I D_N:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C sndPC VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 sndPC D y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 C C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 D D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP4 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 y C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN3 y D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN2 C C_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 D D_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN4 X y VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or4bb_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
*.PININFO A:I B:I C_N:I D_N:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C sndPC VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 sndPC D y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 C C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 D D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP4 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 y C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN3 y D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN2 C C_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 D D_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN4 X y VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or4bb_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
*.PININFO A:I B:I C_N:I D_N:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP2 sndPB C sndPC VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMP3 sndPC D y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 C C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP3 D D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP4 X y VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMN0 y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN1 y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN2 y C VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMN3 y D VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=1.14
XMXNMIN2 C C_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN3 D D_N VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN4 X y VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__or4bb_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
*.PININFO A0:I A1:I S:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMNA00 xb A0 smdNA0 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA01 smdNA0 Sb VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA10 xb A1 sndNA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA11 sndNA1 S VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 Sb S VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X xb VGND VNB sky130_fd_pr__nfet_01v8 m=8 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA00 VPWR S sndPS VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA01 sndPS A0 xb VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA10 VPWR Sb sndPSb VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA11 sndPSb A1 xb VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Sb S VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X xb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=8 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__mux2_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
*.PININFO A0:I A1:I S:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMNA00 xb A0 smdNA0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA01 smdNA0 Sb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA10 xb A1 sndNA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA11 sndNA1 S VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 Sb S VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X xb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA00 VPWR S sndPS VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA01 sndPS A0 xb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA10 VPWR Sb sndPSb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA11 sndPSb A1 xb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Sb S VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X xb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__mux2_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
*.PININFO A0:I A1:I S:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMNA00 xb A0 smdNA0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA01 smdNA0 Sb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA10 xb A1 sndNA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA11 sndNA1 S VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 Sb S VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X xb VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA00 VPWR S sndPS VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA01 sndPS A0 xb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA10 VPWR Sb sndPSb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA11 sndPSb A1 xb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Sb S VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X xb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__mux2_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
*.PININFO A0:I A1:I S:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXNMNA00 xb A0 smdNA0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA01 smdNA0 Sb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA10 xb A1 sndNA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA11 sndNA1 S VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN1 Sb S VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIN2 X xb VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA00 VPWR S sndPS VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA01 sndPS A0 xb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA10 VPWR Sb sndPSb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA11 sndPSb A1 xb VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP1 Sb S VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMIP2 X xb VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__mux2_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdfrbp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I RESET_B:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I
*.PININFO Q:O Q_N:O
XMXNI642 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net92 S0 net134 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net134 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 net127 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 sceb SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 M0 clkpos net115 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 net115 M1 net127 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 S0 clkneg net110 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 Q net92 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net110 net92 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 M1 clkpos S0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI672 net171 net92 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI670 Q_N net171 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI98 db D n0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=3.1
XMXNI103 n1 SCD VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.18 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI120 db SCE n1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI104 n0 sceb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI643 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net215 net92 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 net92 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 S0 clkpos net215 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net92 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI30 net194 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI31 M0 clkneg net194 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI32 net194 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 Q net92 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 M1 clkneg S0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 sceb SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI673 net171 net92 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.64 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI671 Q_N net171 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI101 db sceb p1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI94 db D p0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sdfrbp_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__sdfrbp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I RESET_B:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I
*.PININFO Q:O Q_N:O
XMXNI642 clkneg CLK VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI42 db clkneg M0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI656 net92 S0 net134 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI657 net134 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI33 net127 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI634 sceb SCE VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI4 M0 clkpos net115 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI34 net115 M1 net127 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI655 S0 clkneg net103 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI652 Q net92 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI654 net103 net92 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI647 M1 M0 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.64 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI649 M1 clkpos S0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI672 net171 net92 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.52 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI670 Q_N net171 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.52 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI98 db D n0 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265 sb=0.265
+ sd=0.28 topography=normal perim=3.1
XMXNI103 n1 SCD VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.18 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI120 db SCE n1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI104 n0 sceb VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXNI643 clkneg CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI635 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI43 db clkpos M0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI662 net215 net92 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI659 net92 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI664 S0 clkpos net215 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI658 net92 S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI30 net194 M1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI31 M0 clkneg net194 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI32 net194 RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI663 Q net92 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI648 M1 M0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI650 M1 clkneg S0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.42 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI633 sceb SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI673 net171 net92 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.79 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI671 Q_N net171 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.79 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI101 db sceb p1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI94 db D p0 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=0.54 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__sdfrbp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 Y C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a211oi_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 Y C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a211oi_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 pndB B1 pndA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPC0 Y C1 pndB VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNC0 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__a211oi_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=4 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=4 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o31ai_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o31ai_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__o31ai_2  A1 A2 A3 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXNMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA1 sndA1 A2 sndA2 VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPA2 sndA2 A3 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt m=2 w=1.0 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNA2 pndA A3 VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXNMNB0 Y B1 pndA VNB sky130_fd_pr__nfet_01v8 m=2 w=0.65 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hd__o31ai_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__dfsbp_1 CLK D SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
XMXMI36 net060 M0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI42 db clkneg M0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI39 db D VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI656 M1 M0 net0107 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI654 net0104 M1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI34 S0 clkpos net060 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI25 net52 SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI26 S0 clkneg net44 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI27 net44 S1 net52 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI647 S1 S0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI655 M0 clkpos net0104 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI657 net0107 SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI651 Q_N S0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI652 net072 S0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI653 Q net072 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI40 db D VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI38 S0 clkneg net0127 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI37 net0127 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI43 db clkpos M0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI659 M1 SET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI662 net0172 M1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI664 M0 clkneg net0172 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI6 net55 S1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI5 S0 clkpos net55 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI24 S0 SET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI648 S1 S0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI658 M1 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI663 net072 S0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI660 Q net072 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI661 Q_N S0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__dfsbp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXMI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI42 db clkneg M0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI656 net062 s0 net052 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI657 net052 RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI33 net51 RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI4 M0 clkpos net43 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI34 net43 M1 net51 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI655 s0 clkneg net061 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI652 net069 s0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI653 Q net069 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI654 net061 net062 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI647 M1 M0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI39 db D net098 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI38 net098 RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI649 M1 clkpos s0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI43 db clkpos M0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI662 net089 net062 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI659 net062 RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI664 s0 clkpos net089 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI658 net062 s0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI30 net54 M1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI31 M0 clkneg net54 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI32 M0 RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI663 net069 s0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI660 Q net069 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI648 M1 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI41 db RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI40 db D VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI650 M1 clkneg s0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__dfrtp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__diode_2 DIODE VGND VNB VPB VPWR
*.PININFO DIODE:I VGND:I VNB:I VPB:I VPWR:I
XD0 VNB DIODE sky130_fd_pr__diode_pw2nd_11v0
* Notes: Tap diode is not represented here.
.ENDS sky130_fd_sc_hvl__diode_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__lsbufhv2lv_simple_1 A LVPWR VGND VNB VPB VPWR X
*.PININFO A:I LVPWR:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMMIN1 Ab A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN2 X Ab VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP1 Ab A LVPWR LVPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP2 X Ab LVPWR LVPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__lsbufhv2lv_simple_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__nor2_1 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXMMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMP1 sndPA B Y VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN0 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN1 Y B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__nor2_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__conb_1 VGND VNB VPB VPWR HI LO
*.PININFO VGND:I VNB:I VPB:I VPWR:I HI:O LO:O
rI12 VGND LO short
rI11 HI VPWR short
.ENDS sky130_fd_sc_hvl__conb_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__dfxtp_1 CLK D VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXMI657 M0 clkpos net72 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI656 net72 M1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI646 Q S1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI648 db clkneg M0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI654 db D VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI642 S0 clkneg net48 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI641 net48 S1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI652 M1 clkpos S0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI649 S1 S0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI634 M1 M0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI659 M0 clkneg net100 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI650 S1 S0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI644 S0 clkpos net119 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI639 M1 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI643 net119 S1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI658 net100 M1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI645 Q S1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI651 db clkpos M0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI655 db D VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI653 M1 clkneg S0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__dfxtp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

********.SUBCKT sky130_fd_sc_hvl__decap_8 VGND VNB VPB VPWR

.SUBCKT sky130_fd_sc_hvl__decap_8 VNB VPB VGND VPWR

*.PININFO VGND:I VNB:I VPB:I VPWR:I
XMXMI1 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=0.75 l=1.0 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI2 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=1.0 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__decap_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__decap_4 VGND VNB VPB VPWR
*.PININFO VGND:I VNB:I VPB:I VPWR:I
XMXMI1 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.0 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI2 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=1.0 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__decap_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPA1 sndA1 A2 y VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPB0 VPWR B1 sndB1 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPB1 sndB1 B2 y VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIPX X y VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNB0 y B1 pndA VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNB1 y B2 pndA VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMINX X y VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__o22a_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__sdfsbp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I SCD:I SCE:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
*.PININFO Q_N:O
XMXMI104 db sceb n0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI98 n0 D VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI120 db SCE n1 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI103 n1 SCD VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI36 net125 M0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI42 db clkneg M0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI656 M1 M0 net136 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI654 net141 M1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI34 S0 clkpos net125 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI25 net153 SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI26 S0 clkneg net161 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI27 net161 S1 net153 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI647 S1 S0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI655 M0 clkpos net141 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI657 net136 SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI651 Q_N S0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI652 net265 S0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI653 Q net265 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI49 sceb SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI101 db sceb p1 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI94 db D p0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI38 S0 clkneg net212 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI37 net212 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI43 db clkpos M0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI659 M1 SET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI662 net237 M1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI664 M0 clkneg net237 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI6 net248 S1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI5 S0 clkpos net248 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI24 S0 SET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI648 S1 S0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI658 M1 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI663 net265 S0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI660 Q net265 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI661 Q_N S0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI50 sceb SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__sdfsbp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__dfxbp_1 CLK D VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
XMXMI657 M0 clkpos net72 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI656 net72 M1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI646 Q S1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI662 net116 S1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI648 db clkneg M0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI654 db D VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI642 S0 clkneg net48 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI641 net48 S1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI661 Q_N net116 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI652 M1 clkpos S0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI649 S1 S0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI634 M1 M0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI659 M0 clkneg net100 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI660 Q_N net116 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI650 S1 S0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI644 S0 clkpos net119 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI647 net116 S1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI639 M1 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI643 net119 S1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI658 net100 M1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI645 Q S1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI651 db clkpos M0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI655 db D VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI653 M1 clkneg S0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__dfxbp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
*.PININFO CLK:I GATE:I VGND:I VNB:I VPB:I VPWR:I GCLK:O
XMXMI635 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI22 M1 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI29 net048 M1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI28 net048 CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI650 GCLK net048 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI633 clkpos CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI653 net59 M1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI651 M0 clkpos net59 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI638 net043 GATE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI27 M0 clkneg net043 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI634 clkpos CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI649 GCLK net048 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI31 net084 CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI652 M0 clkneg net102 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI654 net102 M1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI26 net076 GATE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI636 clkneg clkpos VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI637 M0 clkpos net076 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI30 net048 M1 net084 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI23 M1 M0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__dlclkp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__lsbufhv2hv_lh_1 A LOWHVPWR VGND VNB VPB VPWR X
*.PININFO A:I LOWHVPWR:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMI18 cross2 cross1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI7 Abb Ab LOWHVPWR LOWHVPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI15 X cross2 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI19 cross1 cross2 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI27 Ab A LOWHVPWR LOWHVPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI8 Abb Ab VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI16 X cross2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI21 cross2 Abb VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=4 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI22 cross1 Ab VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=4 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI28 Ab A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__lsbufhv2hv_lh_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__or2_1 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMP1 sndPA B y VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP2 X y VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN0 y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN1 y B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN2 X y VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__or2_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__and2_1 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMMP0 y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMP1 y B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP0 X y VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN0 y A sndA VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN1 sndA B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN0 X y VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__and2_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__sdfstp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SCD:I SCE:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXMI104 db sceb n0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI98 n0 D VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI120 db SCE n1 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI103 n1 SCD VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI36 net125 M0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI42 db clkneg M0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI656 M1 M0 net136 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI654 net141 M1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI34 S0 clkpos net125 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI25 net153 SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI26 S0 clkneg net161 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI27 net161 S1 net153 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI647 S1 S0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI655 M0 clkpos net141 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI657 net136 SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI652 net265 S0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI653 Q net265 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI49 sceb SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI101 db sceb p1 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI94 db D p0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI38 S0 clkneg net212 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI37 net212 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI43 db clkpos M0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI659 M1 SET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI662 net237 M1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI664 M0 clkneg net237 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI6 net248 S1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI5 S0 clkpos net248 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI24 S0 SET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI648 S1 S0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI658 M1 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI663 net265 S0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI660 Q net265 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI50 sceb SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__sdfstp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXMI36 net060 M0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI42 db clkneg M0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI39 db D VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI656 M1 M0 net0107 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI654 net0104 M1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI34 S0 clkpos net060 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI25 net52 SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI26 S0 clkneg net44 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI27 net44 S1 net52 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI647 S1 S0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI655 M0 clkpos net0104 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI657 net0107 SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI652 net072 S0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI653 Q net072 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI40 db D VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI38 S0 clkneg net0127 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI37 net0127 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI43 db clkpos M0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI659 M1 SET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI662 net0172 M1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI664 M0 clkneg net0172 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI6 net55 S1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI5 S0 clkpos net55 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI24 S0 SET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI648 S1 S0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI658 M1 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI663 net072 S0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI660 Q net072 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__dfstp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__probec_p_8 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
rI112 net34 X sky130_fd_pr__res_generic_po
XMXMMIN1 Ab A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=3 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN2 net34 Ab VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=8 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP2 net34 Ab VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=8 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__probec_p_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPB0 y B1 pndA VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIPX X y VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNB0 y B1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMINX X y VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__a21o_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__xor2_1 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMMNnor0 inor A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNnor1 inor B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNaoi10 VGND A sndNA VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNaoi11 sndNA B X VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNaoi20 X inor VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPnor0 VPWR A sndPA VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPnor1 sndPA B inor VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPaoi10 pmid A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPaoi11 pmid B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPaoi20 X inor pmid VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__xor2_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__xnor2_1 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXMMNnand0 VGND A sndNA VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNnand1 sndNA B inand VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNaoi10 nmid A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNaoi11 nmid B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNaoi20 Y inand nmid VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPnand0 inand A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPnand1 inand B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPaoi10 VPWR A sndPA VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPaoi11 sndPA B Y VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPaoi20 Y inand VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__xnor2_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__or3_1 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMP2 sndPB C y VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP3 X y VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN0 y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN1 y B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN2 y C VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN3 X y VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__or3_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1 A SLEEP_B LVPWR VGND VNB VPB VPWR X
*.PININFO A:I SLEEP_B:I LVPWR:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMM8 X t1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMM3 t1 t2 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=2.0 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI7 isolate_ahv SLEEP_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI33 t4 t3 LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP1 t3 A LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMM4 t2 t1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=2.0 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMM9 t2 isolate_ahv VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.8
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI34 t4 t3 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMM7 X t1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI16 t2 t3 net54 VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI15 t1 t4 net54 VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN1 t3 A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI6 isolate_ahv SLEEP_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal
+ perim=1.14
XMXMI23 net54 SLEEP_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.6
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1 A LVPWR VGND VNB VPB VPWR X
*.PININFO A:I LVPWR:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMI33 cross2 X_n VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI31 cross1 X_n VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI18 cross2 cross1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI7 Abb Ab LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI30 X_n cross1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI15 X X_n VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI19 cross1 cross2 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI27 Ab A LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI8 Abb Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI16 X X_n VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI21 net81 Abb VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI22 cross1 Ab VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI32 cross2 X_n net81 VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI28 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI29 X_n cross1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__and3_1 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMMP0 y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMP1 y B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMP2 y C VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP0 X y VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN0 y A sndA VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN1 sndA B sndB VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN2 sndB C VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN0 X y VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__and3_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

********.SUBCKT sky130_fd_sc_hvl__lsbufhv2lv_1 A LVPWR VGND VNB VPB VPWR X

.SUBCKT sky130_fd_sc_hvl__lsbufhv2lv_1 VNB VPB LVPWR A VPWR X VGND


*.PININFO A:I LVPWR:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMI7 Abb Ab VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI35 cross1 cross2 LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI36 cross2 cross1 LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI34 X cross2 LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI27 Ab A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI8 Abb Ab VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI21 cross2 Abb VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=4 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI22 cross1 Ab VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=4 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI28 Ab A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI29 X cross2 VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__lsbufhv2lv_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__nand3_1 A B C VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXMMP0 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMP1 Y B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMP2 Y C VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN0 Y A sndA VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN1 sndA B sndB VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN2 sndB C VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__nand3_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__sdlxtp_1 D GATE SCD SCE VGND VNB VPB VPWR Q
*.PININFO D:I GATE:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXMI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI101 db sceb p1 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI94 db D p0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI635 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI22 net069 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI25 db clkneg M0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI650 Q M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI633 clkneg GATE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI653 net59 net069 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI651 M0 clkpos net59 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI50 sceb SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI103 n1 SCD VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI120 db SCE n1 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI104 db sceb n0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI98 n0 D VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI634 clkneg GATE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI649 Q M0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI652 M0 clkneg net102 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI654 net102 net069 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI24 db clkpos M0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI23 net069 M0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI49 sceb SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__sdlxtp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
XMXMI651 Q_N s0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI42 db clkneg M0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI656 net062 s0 net052 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI657 net052 RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI33 net51 RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI4 M0 clkpos net43 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI34 net43 M1 net51 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI655 s0 clkneg net061 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI652 net069 s0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI653 Q net069 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI654 net061 net062 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI647 M1 M0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI39 db D net098 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI38 net098 RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI649 M1 clkpos s0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI43 db clkpos M0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI662 net089 net062 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI659 net062 RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI664 s0 clkpos net089 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI658 net062 s0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI30 net54 M1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI31 M0 clkneg net54 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI32 M0 RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI663 net069 s0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI660 Q net069 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI661 Q_N s0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI648 M1 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI41 db RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI40 db D VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI650 M1 clkneg s0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__dfrbp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__fill_4 VGND VNB VPB VPWR
*.PININFO VGND:I VNB:I VPB:I VPWR:I
* Notes: Cell contains no devices
.ENDS sky130_fd_sc_hvl__fill_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__fill_1 VGND VNB VPB VPWR
*.PININFO VGND:I VNB:I VPB:I VPWR:I
* Notes: Cell contains no devices
.ENDS sky130_fd_sc_hvl__fill_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__fill_8 VGND VNB VPB VPWR
*.PININFO VGND:I VNB:I VPB:I VPWR:I
* Notes: Cell contains no devices
.ENDS sky130_fd_sc_hvl__fill_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__fill_2 VGND VNB VPB VPWR
*.PININFO VGND:I VNB:I VPB:I VPWR:I
* Notes: Cell contains no devices
.ENDS sky130_fd_sc_hvl__fill_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__schmittbuf_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
rI39 net069 VGND sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=1.355 isHV=TRUE
rI38 VPWR net32 sky130_fd_pr__res_generic_pd__hv m=1 w=0.29 l=3.11 isHV=TRUE
XMXMI5 net32 net36 net40 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN0 net36 A net40 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN1 net40 A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN1 X net36 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI6 net069 net36 net56 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMP0 VPWR A net56 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMP1 net56 A net36 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP1 X net36 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__schmittbuf_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__sdfxtp_1 CLK D SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXMI120 db SCE n1 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI103 n1 SCD VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI104 db sceb n0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI98 n0 D VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI657 M0 clkpos net72 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI656 net72 M1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI49 sceb SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI646 Q S1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI648 db clkneg M0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI642 S0 clkneg net48 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI641 net48 S1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI652 M1 clkpos S0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI649 S1 S0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI634 M1 M0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI101 db sceb p1 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI94 db D p0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI659 M0 clkneg net100 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI50 sceb SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI650 S1 S0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI644 S0 clkpos net119 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI639 M1 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI643 net119 S1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI658 net100 M1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI645 Q S1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI651 db clkpos M0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI653 M1 clkneg S0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__sdfxtp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__lsbufhv2hv_hl_1 A LOWHVPWR VGND VNB VPB VPWR X
*.PININFO A:I LOWHVPWR:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMMIN1 Ab A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN2 X Ab VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP1 Ab A LOWHVPWR LOWHVPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP2 X Ab LOWHVPWR LOWHVPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__lsbufhv2hv_hl_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPB0 y B1 pndA VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPB1 y B2 pndA VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIPX X y VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNA0 y A1 sndA1 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNB0 y B1 sndB1 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNB1 sndB1 B2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMINX X y VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__a22o_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__sdfxbp_1 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
XMXMI120 db SCE n1 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI103 n1 SCD VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI104 db sceb n0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI98 n0 D VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI657 M0 clkpos net72 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI656 net72 M1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI49 sceb SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI646 Q S1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI662 net116 S1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI648 db clkneg M0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI642 S0 clkneg net48 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI641 net48 S1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI661 Q_N net116 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI652 M1 clkpos S0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI649 S1 S0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI635 clkneg CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI634 M1 M0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI101 db sceb p1 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI94 db D p0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI659 M0 clkneg net100 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI50 sceb SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI660 Q_N net116 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI650 S1 S0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI644 S0 clkpos net119 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI647 net116 S1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI639 M1 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI643 net119 S1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI638 clkneg CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI658 net100 M1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI645 Q S1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI651 db clkpos M0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI653 M1 clkneg S0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI637 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__sdfxbp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__nor3_1 A B C VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXMMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMP1 sndPA B sndPB VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMP2 sndPB C Y VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN0 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN1 Y B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN2 Y C VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__nor3_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__einvp_1 A TE VGND VNB VPB VPWR Z
*.PININFO A:I TE:I VGND:I VNB:I VPB:I VPWR:I Z:O
XMXMMN0 Z A sndA VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN1 sndA TE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN1 TEB TE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMP0 VPWR TEB sndTEB VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMP1 sndTEB A Z VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP1 TEB TE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__einvp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXMMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPB0 Y B1 pndA VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNB0 Y B1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__a21oi_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__sdlclkp_1 CLK GATE SCE VGND VNB VPB VPWR GCLK
*.PININFO CLK:I GATE:I SCE:I VGND:I VNB:I VPB:I VPWR:I GCLK:O
XMXMI635 clkneg clkpos VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI22 M1 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI29 net048 M1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI28 net048 CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI650 GCLK net048 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI633 clkpos CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI653 net59 M1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI651 M0 clkpos net59 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI638 net043 GATE net037 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI27 M0 clkneg net043 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI33 net037 SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI634 clkpos CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI649 GCLK net048 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI31 net084 CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI652 M0 clkneg net102 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI654 net102 M1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI32 net043 GATE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI26 net043 SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI636 clkneg clkpos VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI637 net043 clkpos M0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI30 net048 M1 net084 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI23 M1 M0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__sdlclkp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__dlrtp_1 D GATE RESET_B VGND VNB VPB VPWR Q
*.PININFO D:I GATE:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXMI635 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI22 M0 clkpos net79 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI25 net76 clkneg M0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI650 Q net96 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI633 clkneg GATE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI638 db D VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI30 VPWR db net76 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI32 net96 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI29 net79 net96 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI26 net96 RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI634 clkneg GATE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI649 Q net96 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI652 net116 net96 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI24 net99 clkpos M0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI637 db D VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI31 VGND db net99 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI33 net96 M0 net95 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI27 net95 RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI23 M0 clkneg net116 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__dlrtp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__dlxtp_1 D GATE VGND VNB VPB VPWR Q
*.PININFO D:I GATE:I VGND:I VNB:I VPB:I VPWR:I Q:O
XMXMI635 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI22 net069 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI25 db clkneg M0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI650 Q M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI633 clkneg GATE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI653 net59 net069 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI651 M0 clkpos net59 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI638 db D VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI634 clkneg GATE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI649 Q M0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI652 M0 clkneg net102 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI654 net102 net069 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI24 db clkpos M0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI636 clkpos clkneg VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI637 db D VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI23 net069 M0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__dlxtp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPA1 sndA1 A2 y VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPB0 VPWR B1 y VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIPX X y VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNB0 y B1 pndA VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMINX X y VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__o21a_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__probe_p_8 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
rI112 net23 X sky130_fd_pr__res_generic_po
XMXMMIN1 Ab A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=3 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN2 net23 Ab VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=8 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP2 net23 Ab VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=8 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__probe_p_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I RESET_B:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I
*.PININFO Q:O
XMXMI98 n0 D net076 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI14 net076 RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI104 db sceb n0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI120 db SCE n1 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI103 n1 SCD net076 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI42 db clkneg M0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI656 net062 s0 net052 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI657 net052 RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI33 net51 RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI4 M0 clkpos net43 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI34 net43 M1 net51 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI655 s0 clkneg net061 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI652 net069 s0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI49 sceb SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI653 Q net069 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI654 net061 net062 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI647 M1 M0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI649 M1 clkpos s0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI94 db D p0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI15 db RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI101 db sceb p1 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI43 db clkpos M0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI662 net089 net062 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI659 net062 RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI664 s0 clkpos net089 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI658 net062 s0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI30 net54 M1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI31 M0 clkneg net54 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI32 M0 RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI663 net069 s0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI660 Q net069 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI50 sceb SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI648 M1 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI650 M1 clkneg s0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__sdfrtp_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
*.PININFO A0:I A1:I A2:I A3:I S0:I S1:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMMNA00 sndNS0ba0 S0b xlowb VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMNA01 VGND A0 sndNS0ba0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMNA10 sndNS0a1 S0 xlowb VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMNA11 VGND A1 sndNS0a1 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMNA20 sndNS0ba2 S0b xhib VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMNA21 VGND A2 sndNS0ba2 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMNA30 sndNS0a3 S0 xhib VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMNA31 VGND A3 sndNS0a3 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMNs1o xb S1b xlowb VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMNs2o xb S1 xhib VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMIN1 VGND S1 S1b VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMIN2 VGND S0 S0b VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMIN4 VGND xb X VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMPA00 sndPA0a0 A0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMPA01 xlowb S0 sndPA0a0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMPA10 sndPA1a1 A1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMPA11 xlowb S0b sndPA1a1 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMPA20 sndPA2a2 A2 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMPA21 xhib S0 sndPA2a2 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMPA30 sndPA3a3 A3 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMPA31 xhib S0b sndPA3a3 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMPs1o xb S1 xlowb VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMPs2o xb S1b xhib VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMIP1 VPWR S1 S1b VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMIP2 VPWR S0 S0b VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
XMXMMIP4 VPWR xb X VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=0.76
.ENDS sky130_fd_sc_hvl__mux4_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__nand2_1 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXMMP0 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMP1 Y B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN0 Y A sndA VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN1 sndA B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__nand2_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXMMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPA1 sndA1 A2 Y VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPB0 VPWR B1 Y VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNB0 Y B1 pndA VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__o21ai_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__inv_16 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXMMIP1 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=16 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=16 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__inv_16


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__inv_8 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXMMIP1 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=8 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=8 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__inv_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__inv_1 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXMMIP1 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__inv_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__inv_2 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXMMIP1 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__inv_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__inv_4 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXMMIP1 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=4 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__inv_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__buf_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMMIN1 Ab A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN2 X Ab VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP2 X Ab VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__buf_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__buf_8 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMMIN1 Ab A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=3 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN2 X Ab VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=8 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP2 X Ab VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=8 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__buf_8


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__buf_32 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMMIN1 Ab A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=10 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN2 X Ab VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=32 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=10 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP2 X Ab VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=32 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__buf_32


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__buf_4 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMMIN1 Ab A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN2 X Ab VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=4 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP2 X Ab VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__buf_4


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__buf_2 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMMIN1 Ab A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN2 X Ab VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP2 X Ab VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__buf_2


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__buf_16 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMMIN1 Ab A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=6 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN2 X Ab VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=16 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP1 Ab A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=6 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP2 X Ab VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=16 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__buf_16


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXMMPA0 VPWR A1 sndA1 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPA1 sndA1 A2 Y VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPB0 VPWR B1 sndB1 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPB1 sndB1 B2 Y VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNA0 pndA A1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNA1 pndA A2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNB0 Y B1 pndA VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNB1 Y B2 pndA VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__o22ai_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__einvn_1 A TE_B VGND VNB VPB VPWR Z
*.PININFO A:I TE_B:I VGND:I VNB:I VPB:I VPWR:I Z:O
XMXMMN0 Z A sndA VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMN1 sndA TE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN1 TE TE_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMP0 VPWR TE_B sndTEB VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMP1 sndTEB A Z VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP1 TE TE_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__einvn_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
XMXMMPA0 pndA A1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPA1 pndA A2 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPB0 Y B1 pndA VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPB1 Y B2 pndA VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNA0 Y A1 sndA1 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNA1 sndA1 A2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNB0 Y B1 sndB1 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNB1 sndB1 B2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__a22oi_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__lsbuflv2hv_1 A LVPWR VGND VNB VPB VPWR X
*.PININFO A:I LVPWR:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMI18 net81 cross1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI7 Abb Ab LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI30 net65 cross1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI15 X net65 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI19 cross1 net81 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI27 Ab A LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI8 Abb Ab VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI16 X net65 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI21 net81 Abb VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=5 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI22 cross1 Ab VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=5 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI28 Ab A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.84 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI29 net65 cross1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__lsbuflv2hv_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3 A SLEEP_B LVPWR VGND VNB VPB VPWR X
*.PININFO A:I SLEEP_B:I LVPWR:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMM9 t1 isolate_ahv VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI44 t2 VGND VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI16 t2 t3 VGND VNB sky130_fd_pr__nfet_05v0_nvt m=4 w=1.0 l=0.9 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN1 net065 A VGND VNB sky130_fd_pr__nfet_01v8 m=2 w=0.74 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI47 X t8 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI63 t4 t3 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.74 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI15 t1 t4 VGND VNB sky130_fd_pr__nfet_05v0_nvt m=4 w=1.0 l=0.9 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI35 isolate_ahv SLEEP_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal
+ perim=1.14
XMXMI45 t8 t1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI58 t3 net065 VGND VNB sky130_fd_pr__nfet_01v8 m=4 w=0.74 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMM3 t1 t2 net128 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMM4 t2 t1 net128 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI53 net128 isolate_ahv VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.0 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI46 t8 t1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP1 net065 A LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt m=2 w=1.12 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI36 isolate_ahv SLEEP_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal
+ perim=1.14
XMXMI64 t4 t3 LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt m=4 w=1.12 l=0.15 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI57 t3 net065 LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt m=4 w=1.12 l=0.15
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI48 X t8 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=3 w=3.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__mux2_1 A0 A1 S VGND VNB VPB VPWR X
*.PININFO A0:I A1:I S:I VGND:I VNB:I VPB:I VPWR:I X:O
XMXMMNA00 xb A0 smdNA0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNA01 smdNA0 Sb VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNA10 xb A1 sndNA1 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMNA11 sndNA1 S VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN1 Sb S VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIN2 X xb VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPA00 VPWR S sndPS VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPA01 sndPS A0 xb VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPA10 VPWR Sb sndPSb VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMPA11 sndPSb A1 xb VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP1 Sb S VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMMIP2 X xb VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__mux2_1


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__sdfrbp_1  CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I RESET_B:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I
*.PININFO Q:O Q_N:O
XMXMI98 n0 D net076 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI14 net076 RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI104 db sceb n0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI120 db SCE n1 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI103 n1 SCD net076 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=3.1
XMXMI651 Q_N s0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI46 clkpos clkneg VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI42 db clkneg M0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI656 net062 s0 net052 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI657 net052 RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI33 net51 RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI4 M0 clkpos net43 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI34 net43 M1 net51 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI655 s0 clkneg net061 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI652 net069 s0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI49 sceb SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI653 Q net069 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI654 net061 net062 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI44 clkneg CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI647 M1 M0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI649 M1 clkpos s0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI94 db D p0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI15 db RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI101 db sceb p1 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI107 p0 SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI108 p1 SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI47 clkpos clkneg VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI43 db clkpos M0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI662 net089 net062 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI659 net062 RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI664 s0 clkpos net089 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI658 net062 s0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI30 net54 M1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI31 M0 clkneg net54 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI32 M0 RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI663 net069 s0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI660 Q net069 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI661 Q_N s0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI50 sceb SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI45 clkneg CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ sa=0.265 sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI648 M1 M0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
XMXMI650 M1 clkneg s0 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 sa=0.265
+ sb=0.265 sd=0.28 topography=normal perim=1.14
.ENDS sky130_fd_sc_hvl__sdfrbp_1


******* EOF

**************************************************
* OpenRAM generated memory.
* Words: 256
* Data bits: 32
* Banks: 1
* Column mux: 2:1
**************************************************
* SPICE3 file created from dff.ext - technology: EFS8A

.subckt dff D Q clk vdd gnd
XM1000 a_511_725# a_n8_115# VDD VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15 m=1
XM1001 a_353_115# CLK a_11_624# GND sky130_fd_pr__nfet_01v8 W=1 L=0.15 m=1
XM1002 a_353_725# a_203_89# a_11_624# VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15 m=1
XM1003 a_11_624# a_203_89# a_161_115# GND sky130_fd_pr__nfet_01v8 W=1 L=0.15 m=1
XM1004 a_11_624# CLK a_161_725# VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15 m=1
XM1005 GND Q a_703_115# GND sky130_fd_pr__nfet_01v8 W=1 L=0.15 m=1
XM1006 VDD Q a_703_725# VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15 m=1
XM1007 a_203_89# CLK GND GND sky130_fd_pr__nfet_01v8 W=1 L=0.15 m=1
XM1008 a_203_89# CLK VDD VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15 m=1
XM1009 a_161_115# D GND GND sky130_fd_pr__nfet_01v8 W=1 L=0.15 m=1
XM1010 a_161_725# D VDD VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15 m=1
XM1011 GND a_11_624# a_n8_115# GND sky130_fd_pr__nfet_01v8 W=1 L=0.15 m=1
XM1012 a_703_115# a_203_89# ON GND sky130_fd_pr__nfet_01v8 W=1 L=0.15 m=1
XM1013 VDD a_11_624# a_n8_115# VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15 m=1
XM1014 a_703_725# CLK ON VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15 m=1
XM1015 Q ON VDD VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15 m=1
XM1016 Q ON GND GND sky130_fd_pr__nfet_01v8 W=1 L=0.15 m=1
XM1017 ON a_203_89# a_511_725# VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15 m=1
XM1018 ON CLK a_511_115# GND sky130_fd_pr__nfet_01v8 W=1 L=0.15 m=1
XM1019 GND a_n8_115# a_353_115# GND sky130_fd_pr__nfet_01v8 W=1 L=0.15 m=1
XM1020 VDD a_n8_115# a_353_725# VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15 m=1
XM1021 a_511_115# a_n8_115# GND GND sky130_fd_pr__nfet_01v8 W=1 L=0.15 m=1
.ends

.SUBCKT row_addr_dff din_0 din_1 din_2 din_3 din_4 din_5 din_6 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5 dout_6 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 7 cols: 1
Xdff_r0_c0 din_0 dout_0 clk vdd gnd dff
Xdff_r1_c0 din_1 dout_1 clk vdd gnd dff
Xdff_r2_c0 din_2 dout_2 clk vdd gnd dff
Xdff_r3_c0 din_3 dout_3 clk vdd gnd dff
Xdff_r4_c0 din_4 dout_4 clk vdd gnd dff
Xdff_r5_c0 din_5 dout_5 clk vdd gnd dff
Xdff_r6_c0 din_6 dout_6 clk vdd gnd dff
.ENDS row_addr_dff

.SUBCKT col_addr_dff din_0 dout_0 clk vdd gnd
* INPUT : din_0 
* OUTPUT: dout_0 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 1
Xdff_r0_c0 din_0 dout_0 clk vdd gnd dff
.ENDS col_addr_dff

.SUBCKT data_dff din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10 din_11 din_12 din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20 din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30 din_31 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5 dout_6 dout_7 dout_8 dout_9 dout_10 dout_11 dout_12 dout_13 dout_14 dout_15 dout_16 dout_17 dout_18 dout_19 dout_20 dout_21 dout_22 dout_23 dout_24 dout_25 dout_26 dout_27 dout_28 dout_29 dout_30 dout_31 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* INPUT : din_7 
* INPUT : din_8 
* INPUT : din_9 
* INPUT : din_10 
* INPUT : din_11 
* INPUT : din_12 
* INPUT : din_13 
* INPUT : din_14 
* INPUT : din_15 
* INPUT : din_16 
* INPUT : din_17 
* INPUT : din_18 
* INPUT : din_19 
* INPUT : din_20 
* INPUT : din_21 
* INPUT : din_22 
* INPUT : din_23 
* INPUT : din_24 
* INPUT : din_25 
* INPUT : din_26 
* INPUT : din_27 
* INPUT : din_28 
* INPUT : din_29 
* INPUT : din_30 
* INPUT : din_31 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* OUTPUT: dout_7 
* OUTPUT: dout_8 
* OUTPUT: dout_9 
* OUTPUT: dout_10 
* OUTPUT: dout_11 
* OUTPUT: dout_12 
* OUTPUT: dout_13 
* OUTPUT: dout_14 
* OUTPUT: dout_15 
* OUTPUT: dout_16 
* OUTPUT: dout_17 
* OUTPUT: dout_18 
* OUTPUT: dout_19 
* OUTPUT: dout_20 
* OUTPUT: dout_21 
* OUTPUT: dout_22 
* OUTPUT: dout_23 
* OUTPUT: dout_24 
* OUTPUT: dout_25 
* OUTPUT: dout_26 
* OUTPUT: dout_27 
* OUTPUT: dout_28 
* OUTPUT: dout_29 
* OUTPUT: dout_30 
* OUTPUT: dout_31 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 32
Xdff_r0_c0 din_0 dout_0 clk vdd gnd dff
Xdff_r0_c1 din_1 dout_1 clk vdd gnd dff
Xdff_r0_c2 din_2 dout_2 clk vdd gnd dff
Xdff_r0_c3 din_3 dout_3 clk vdd gnd dff
Xdff_r0_c4 din_4 dout_4 clk vdd gnd dff
Xdff_r0_c5 din_5 dout_5 clk vdd gnd dff
Xdff_r0_c6 din_6 dout_6 clk vdd gnd dff
Xdff_r0_c7 din_7 dout_7 clk vdd gnd dff
Xdff_r0_c8 din_8 dout_8 clk vdd gnd dff
Xdff_r0_c9 din_9 dout_9 clk vdd gnd dff
Xdff_r0_c10 din_10 dout_10 clk vdd gnd dff
Xdff_r0_c11 din_11 dout_11 clk vdd gnd dff
Xdff_r0_c12 din_12 dout_12 clk vdd gnd dff
Xdff_r0_c13 din_13 dout_13 clk vdd gnd dff
Xdff_r0_c14 din_14 dout_14 clk vdd gnd dff
Xdff_r0_c15 din_15 dout_15 clk vdd gnd dff
Xdff_r0_c16 din_16 dout_16 clk vdd gnd dff
Xdff_r0_c17 din_17 dout_17 clk vdd gnd dff
Xdff_r0_c18 din_18 dout_18 clk vdd gnd dff
Xdff_r0_c19 din_19 dout_19 clk vdd gnd dff
Xdff_r0_c20 din_20 dout_20 clk vdd gnd dff
Xdff_r0_c21 din_21 dout_21 clk vdd gnd dff
Xdff_r0_c22 din_22 dout_22 clk vdd gnd dff
Xdff_r0_c23 din_23 dout_23 clk vdd gnd dff
Xdff_r0_c24 din_24 dout_24 clk vdd gnd dff
Xdff_r0_c25 din_25 dout_25 clk vdd gnd dff
Xdff_r0_c26 din_26 dout_26 clk vdd gnd dff
Xdff_r0_c27 din_27 dout_27 clk vdd gnd dff
Xdff_r0_c28 din_28 dout_28 clk vdd gnd dff
Xdff_r0_c29 din_29 dout_29 clk vdd gnd dff
Xdff_r0_c30 din_30 dout_30 clk vdd gnd dff
Xdff_r0_c31 din_31 dout_31 clk vdd gnd dff
.ENDS data_dff

.SUBCKT wmask_dff din_0 din_1 din_2 din_3 dout_0 dout_1 dout_2 dout_3 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 4
Xdff_r0_c0 din_0 dout_0 clk vdd gnd dff
Xdff_r0_c1 din_1 dout_1 clk vdd gnd dff
Xdff_r0_c2 din_2 dout_2 clk vdd gnd dff
Xdff_r0_c3 din_3 dout_3 clk vdd gnd dff
.ENDS wmask_dff

* ptx M{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=0.15 pd=1.40 ps=1.40 as=0.21u ad=0.21u

.SUBCKT precharge_0 bl br en_bar vdd
* OUTPUT: bl 
* OUTPUT: br 
* INPUT : en_bar 
* POWER : vdd 
XMlower_pmos bl en_bar br vdd sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=0.15 pd=1.40 ps=1.40 as=0.21u ad=0.21u
XMupper_pmos1 bl en_bar vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=0.15 pd=1.40 ps=1.40 as=0.21u ad=0.21u
XMupper_pmos2 br en_bar vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=0.15 pd=1.40 ps=1.40 as=0.21u ad=0.21u
.ENDS precharge_0

.SUBCKT precharge_array bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 en_bar vdd
* OUTPUT: bl_0 
* OUTPUT: br_0 
* OUTPUT: bl_1 
* OUTPUT: br_1 
* OUTPUT: bl_2 
* OUTPUT: br_2 
* OUTPUT: bl_3 
* OUTPUT: br_3 
* OUTPUT: bl_4 
* OUTPUT: br_4 
* OUTPUT: bl_5 
* OUTPUT: br_5 
* OUTPUT: bl_6 
* OUTPUT: br_6 
* OUTPUT: bl_7 
* OUTPUT: br_7 
* OUTPUT: bl_8 
* OUTPUT: br_8 
* OUTPUT: bl_9 
* OUTPUT: br_9 
* OUTPUT: bl_10 
* OUTPUT: br_10 
* OUTPUT: bl_11 
* OUTPUT: br_11 
* OUTPUT: bl_12 
* OUTPUT: br_12 
* OUTPUT: bl_13 
* OUTPUT: br_13 
* OUTPUT: bl_14 
* OUTPUT: br_14 
* OUTPUT: bl_15 
* OUTPUT: br_15 
* OUTPUT: bl_16 
* OUTPUT: br_16 
* OUTPUT: bl_17 
* OUTPUT: br_17 
* OUTPUT: bl_18 
* OUTPUT: br_18 
* OUTPUT: bl_19 
* OUTPUT: br_19 
* OUTPUT: bl_20 
* OUTPUT: br_20 
* OUTPUT: bl_21 
* OUTPUT: br_21 
* OUTPUT: bl_22 
* OUTPUT: br_22 
* OUTPUT: bl_23 
* OUTPUT: br_23 
* OUTPUT: bl_24 
* OUTPUT: br_24 
* OUTPUT: bl_25 
* OUTPUT: br_25 
* OUTPUT: bl_26 
* OUTPUT: br_26 
* OUTPUT: bl_27 
* OUTPUT: br_27 
* OUTPUT: bl_28 
* OUTPUT: br_28 
* OUTPUT: bl_29 
* OUTPUT: br_29 
* OUTPUT: bl_30 
* OUTPUT: br_30 
* OUTPUT: bl_31 
* OUTPUT: br_31 
* OUTPUT: bl_32 
* OUTPUT: br_32 
* OUTPUT: bl_33 
* OUTPUT: br_33 
* OUTPUT: bl_34 
* OUTPUT: br_34 
* OUTPUT: bl_35 
* OUTPUT: br_35 
* OUTPUT: bl_36 
* OUTPUT: br_36 
* OUTPUT: bl_37 
* OUTPUT: br_37 
* OUTPUT: bl_38 
* OUTPUT: br_38 
* OUTPUT: bl_39 
* OUTPUT: br_39 
* OUTPUT: bl_40 
* OUTPUT: br_40 
* OUTPUT: bl_41 
* OUTPUT: br_41 
* OUTPUT: bl_42 
* OUTPUT: br_42 
* OUTPUT: bl_43 
* OUTPUT: br_43 
* OUTPUT: bl_44 
* OUTPUT: br_44 
* OUTPUT: bl_45 
* OUTPUT: br_45 
* OUTPUT: bl_46 
* OUTPUT: br_46 
* OUTPUT: bl_47 
* OUTPUT: br_47 
* OUTPUT: bl_48 
* OUTPUT: br_48 
* OUTPUT: bl_49 
* OUTPUT: br_49 
* OUTPUT: bl_50 
* OUTPUT: br_50 
* OUTPUT: bl_51 
* OUTPUT: br_51 
* OUTPUT: bl_52 
* OUTPUT: br_52 
* OUTPUT: bl_53 
* OUTPUT: br_53 
* OUTPUT: bl_54 
* OUTPUT: br_54 
* OUTPUT: bl_55 
* OUTPUT: br_55 
* OUTPUT: bl_56 
* OUTPUT: br_56 
* OUTPUT: bl_57 
* OUTPUT: br_57 
* OUTPUT: bl_58 
* OUTPUT: br_58 
* OUTPUT: bl_59 
* OUTPUT: br_59 
* OUTPUT: bl_60 
* OUTPUT: br_60 
* OUTPUT: bl_61 
* OUTPUT: br_61 
* OUTPUT: bl_62 
* OUTPUT: br_62 
* OUTPUT: bl_63 
* OUTPUT: br_63 
* OUTPUT: bl_64 
* OUTPUT: br_64 
* INPUT : en_bar 
* POWER : vdd 
* cols: 65 size: 1 bl: bl0 br: br0
Xpre_column_0 bl_0 br_0 en_bar vdd precharge_0
Xpre_column_1 bl_1 br_1 en_bar vdd precharge_0
Xpre_column_2 bl_2 br_2 en_bar vdd precharge_0
Xpre_column_3 bl_3 br_3 en_bar vdd precharge_0
Xpre_column_4 bl_4 br_4 en_bar vdd precharge_0
Xpre_column_5 bl_5 br_5 en_bar vdd precharge_0
Xpre_column_6 bl_6 br_6 en_bar vdd precharge_0
Xpre_column_7 bl_7 br_7 en_bar vdd precharge_0
Xpre_column_8 bl_8 br_8 en_bar vdd precharge_0
Xpre_column_9 bl_9 br_9 en_bar vdd precharge_0
Xpre_column_10 bl_10 br_10 en_bar vdd precharge_0
Xpre_column_11 bl_11 br_11 en_bar vdd precharge_0
Xpre_column_12 bl_12 br_12 en_bar vdd precharge_0
Xpre_column_13 bl_13 br_13 en_bar vdd precharge_0
Xpre_column_14 bl_14 br_14 en_bar vdd precharge_0
Xpre_column_15 bl_15 br_15 en_bar vdd precharge_0
Xpre_column_16 bl_16 br_16 en_bar vdd precharge_0
Xpre_column_17 bl_17 br_17 en_bar vdd precharge_0
Xpre_column_18 bl_18 br_18 en_bar vdd precharge_0
Xpre_column_19 bl_19 br_19 en_bar vdd precharge_0
Xpre_column_20 bl_20 br_20 en_bar vdd precharge_0
Xpre_column_21 bl_21 br_21 en_bar vdd precharge_0
Xpre_column_22 bl_22 br_22 en_bar vdd precharge_0
Xpre_column_23 bl_23 br_23 en_bar vdd precharge_0
Xpre_column_24 bl_24 br_24 en_bar vdd precharge_0
Xpre_column_25 bl_25 br_25 en_bar vdd precharge_0
Xpre_column_26 bl_26 br_26 en_bar vdd precharge_0
Xpre_column_27 bl_27 br_27 en_bar vdd precharge_0
Xpre_column_28 bl_28 br_28 en_bar vdd precharge_0
Xpre_column_29 bl_29 br_29 en_bar vdd precharge_0
Xpre_column_30 bl_30 br_30 en_bar vdd precharge_0
Xpre_column_31 bl_31 br_31 en_bar vdd precharge_0
Xpre_column_32 bl_32 br_32 en_bar vdd precharge_0
Xpre_column_33 bl_33 br_33 en_bar vdd precharge_0
Xpre_column_34 bl_34 br_34 en_bar vdd precharge_0
Xpre_column_35 bl_35 br_35 en_bar vdd precharge_0
Xpre_column_36 bl_36 br_36 en_bar vdd precharge_0
Xpre_column_37 bl_37 br_37 en_bar vdd precharge_0
Xpre_column_38 bl_38 br_38 en_bar vdd precharge_0
Xpre_column_39 bl_39 br_39 en_bar vdd precharge_0
Xpre_column_40 bl_40 br_40 en_bar vdd precharge_0
Xpre_column_41 bl_41 br_41 en_bar vdd precharge_0
Xpre_column_42 bl_42 br_42 en_bar vdd precharge_0
Xpre_column_43 bl_43 br_43 en_bar vdd precharge_0
Xpre_column_44 bl_44 br_44 en_bar vdd precharge_0
Xpre_column_45 bl_45 br_45 en_bar vdd precharge_0
Xpre_column_46 bl_46 br_46 en_bar vdd precharge_0
Xpre_column_47 bl_47 br_47 en_bar vdd precharge_0
Xpre_column_48 bl_48 br_48 en_bar vdd precharge_0
Xpre_column_49 bl_49 br_49 en_bar vdd precharge_0
Xpre_column_50 bl_50 br_50 en_bar vdd precharge_0
Xpre_column_51 bl_51 br_51 en_bar vdd precharge_0
Xpre_column_52 bl_52 br_52 en_bar vdd precharge_0
Xpre_column_53 bl_53 br_53 en_bar vdd precharge_0
Xpre_column_54 bl_54 br_54 en_bar vdd precharge_0
Xpre_column_55 bl_55 br_55 en_bar vdd precharge_0
Xpre_column_56 bl_56 br_56 en_bar vdd precharge_0
Xpre_column_57 bl_57 br_57 en_bar vdd precharge_0
Xpre_column_58 bl_58 br_58 en_bar vdd precharge_0
Xpre_column_59 bl_59 br_59 en_bar vdd precharge_0
Xpre_column_60 bl_60 br_60 en_bar vdd precharge_0
Xpre_column_61 bl_61 br_61 en_bar vdd precharge_0
Xpre_column_62 bl_62 br_62 en_bar vdd precharge_0
Xpre_column_63 bl_63 br_63 en_bar vdd precharge_0
Xpre_column_64 bl_64 br_64 en_bar vdd precharge_0
.ENDS precharge_array
*********************** "sense_amp" ******************************

.SUBCKT sense_amp bl br dout en vdd gnd
XM1000 gnd en a_56_432# gnd sky130_fd_pr__nfet_01v8 W=0.65 L=0.15 m=1
XM1001 a_56_432# dint_bar dint gnd sky130_fd_pr__nfet_01v8 W=0.65 L=0.15 m=1
XM1002 dint_bar dint a_56_432# gnd sky130_fd_pr__nfet_01v8 W=0.65 L=0.15 m=1

XM1003 vdd dint_bar dint vdd sky130_fd_pr__pfet_01v8 W=1.26 L=0.15 m=1
XM1004 dint_bar dint vdd vdd sky130_fd_pr__pfet_01v8 W=1.26 L=0.15 m=1

XM1005 bl en dint vdd sky130_fd_pr__pfet_01v8 W=2 L=0.15 m=1
XM1006 dint_bar en br vdd sky130_fd_pr__pfet_01v8 W=2 L=0.15 m=1

XM1007 vdd dint_bar dout vdd sky130_fd_pr__pfet_01v8 W=1.26 L=0.15 m=1
XM1008 dout dint_bar gnd gnd sky130_fd_pr__nfet_01v8 W=0.65 L=0.15 m=1

.ENDS sense_amp

.SUBCKT sense_amp_array data_0 bl_0 br_0 data_1 bl_1 br_1 data_2 bl_2 br_2 data_3 bl_3 br_3 data_4 bl_4 br_4 data_5 bl_5 br_5 data_6 bl_6 br_6 data_7 bl_7 br_7 data_8 bl_8 br_8 data_9 bl_9 br_9 data_10 bl_10 br_10 data_11 bl_11 br_11 data_12 bl_12 br_12 data_13 bl_13 br_13 data_14 bl_14 br_14 data_15 bl_15 br_15 data_16 bl_16 br_16 data_17 bl_17 br_17 data_18 bl_18 br_18 data_19 bl_19 br_19 data_20 bl_20 br_20 data_21 bl_21 br_21 data_22 bl_22 br_22 data_23 bl_23 br_23 data_24 bl_24 br_24 data_25 bl_25 br_25 data_26 bl_26 br_26 data_27 bl_27 br_27 data_28 bl_28 br_28 data_29 bl_29 br_29 data_30 bl_30 br_30 data_31 bl_31 br_31 en vdd gnd
* OUTPUT: data_0 
* INPUT : bl_0 
* INPUT : br_0 
* OUTPUT: data_1 
* INPUT : bl_1 
* INPUT : br_1 
* OUTPUT: data_2 
* INPUT : bl_2 
* INPUT : br_2 
* OUTPUT: data_3 
* INPUT : bl_3 
* INPUT : br_3 
* OUTPUT: data_4 
* INPUT : bl_4 
* INPUT : br_4 
* OUTPUT: data_5 
* INPUT : bl_5 
* INPUT : br_5 
* OUTPUT: data_6 
* INPUT : bl_6 
* INPUT : br_6 
* OUTPUT: data_7 
* INPUT : bl_7 
* INPUT : br_7 
* OUTPUT: data_8 
* INPUT : bl_8 
* INPUT : br_8 
* OUTPUT: data_9 
* INPUT : bl_9 
* INPUT : br_9 
* OUTPUT: data_10 
* INPUT : bl_10 
* INPUT : br_10 
* OUTPUT: data_11 
* INPUT : bl_11 
* INPUT : br_11 
* OUTPUT: data_12 
* INPUT : bl_12 
* INPUT : br_12 
* OUTPUT: data_13 
* INPUT : bl_13 
* INPUT : br_13 
* OUTPUT: data_14 
* INPUT : bl_14 
* INPUT : br_14 
* OUTPUT: data_15 
* INPUT : bl_15 
* INPUT : br_15 
* OUTPUT: data_16 
* INPUT : bl_16 
* INPUT : br_16 
* OUTPUT: data_17 
* INPUT : bl_17 
* INPUT : br_17 
* OUTPUT: data_18 
* INPUT : bl_18 
* INPUT : br_18 
* OUTPUT: data_19 
* INPUT : bl_19 
* INPUT : br_19 
* OUTPUT: data_20 
* INPUT : bl_20 
* INPUT : br_20 
* OUTPUT: data_21 
* INPUT : bl_21 
* INPUT : br_21 
* OUTPUT: data_22 
* INPUT : bl_22 
* INPUT : br_22 
* OUTPUT: data_23 
* INPUT : bl_23 
* INPUT : br_23 
* OUTPUT: data_24 
* INPUT : bl_24 
* INPUT : br_24 
* OUTPUT: data_25 
* INPUT : bl_25 
* INPUT : br_25 
* OUTPUT: data_26 
* INPUT : bl_26 
* INPUT : br_26 
* OUTPUT: data_27 
* INPUT : bl_27 
* INPUT : br_27 
* OUTPUT: data_28 
* INPUT : bl_28 
* INPUT : br_28 
* OUTPUT: data_29 
* INPUT : bl_29 
* INPUT : br_29 
* OUTPUT: data_30 
* INPUT : bl_30 
* INPUT : br_30 
* OUTPUT: data_31 
* INPUT : bl_31 
* INPUT : br_31 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* words_per_row: 2
Xsa_d0 bl_0 br_0 data_0 en vdd gnd sense_amp
Xsa_d1 bl_1 br_1 data_1 en vdd gnd sense_amp
Xsa_d2 bl_2 br_2 data_2 en vdd gnd sense_amp
Xsa_d3 bl_3 br_3 data_3 en vdd gnd sense_amp
Xsa_d4 bl_4 br_4 data_4 en vdd gnd sense_amp
Xsa_d5 bl_5 br_5 data_5 en vdd gnd sense_amp
Xsa_d6 bl_6 br_6 data_6 en vdd gnd sense_amp
Xsa_d7 bl_7 br_7 data_7 en vdd gnd sense_amp
Xsa_d8 bl_8 br_8 data_8 en vdd gnd sense_amp
Xsa_d9 bl_9 br_9 data_9 en vdd gnd sense_amp
Xsa_d10 bl_10 br_10 data_10 en vdd gnd sense_amp
Xsa_d11 bl_11 br_11 data_11 en vdd gnd sense_amp
Xsa_d12 bl_12 br_12 data_12 en vdd gnd sense_amp
Xsa_d13 bl_13 br_13 data_13 en vdd gnd sense_amp
Xsa_d14 bl_14 br_14 data_14 en vdd gnd sense_amp
Xsa_d15 bl_15 br_15 data_15 en vdd gnd sense_amp
Xsa_d16 bl_16 br_16 data_16 en vdd gnd sense_amp
Xsa_d17 bl_17 br_17 data_17 en vdd gnd sense_amp
Xsa_d18 bl_18 br_18 data_18 en vdd gnd sense_amp
Xsa_d19 bl_19 br_19 data_19 en vdd gnd sense_amp
Xsa_d20 bl_20 br_20 data_20 en vdd gnd sense_amp
Xsa_d21 bl_21 br_21 data_21 en vdd gnd sense_amp
Xsa_d22 bl_22 br_22 data_22 en vdd gnd sense_amp
Xsa_d23 bl_23 br_23 data_23 en vdd gnd sense_amp
Xsa_d24 bl_24 br_24 data_24 en vdd gnd sense_amp
Xsa_d25 bl_25 br_25 data_25 en vdd gnd sense_amp
Xsa_d26 bl_26 br_26 data_26 en vdd gnd sense_amp
Xsa_d27 bl_27 br_27 data_27 en vdd gnd sense_amp
Xsa_d28 bl_28 br_28 data_28 en vdd gnd sense_amp
Xsa_d29 bl_29 br_29 data_29 en vdd gnd sense_amp
Xsa_d30 bl_30 br_30 data_30 en vdd gnd sense_amp
Xsa_d31 bl_31 br_31 data_31 en vdd gnd sense_amp
.ENDS sense_amp_array

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=3.0 l=0.15 pd=6.06 ps=6.06 as=1.08u ad=1.08u

.SUBCKT single_level_column_mux bl br bl_out br_out sel gnd
* INOUT : bl 
* INOUT : br 
* INOUT : bl_out 
* INOUT : br_out 
* INOUT : sel 
* INOUT : gnd 
XMmux_tx1 bl sel bl_out gnd sky130_fd_pr__nfet_01v8 m=1 w=3.0 l=0.15 pd=6.06 ps=6.06 as=1.08u ad=1.08u
XMmux_tx2 br sel br_out gnd sky130_fd_pr__nfet_01v8 m=1 w=3.0 l=0.15 pd=6.06 ps=6.06 as=1.08u ad=1.08u
.ENDS single_level_column_mux

.SUBCKT single_level_column_mux_array bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 sel_0 sel_1 bl_out_0 br_out_0 bl_out_1 br_out_1 bl_out_2 br_out_2 bl_out_3 br_out_3 bl_out_4 br_out_4 bl_out_5 br_out_5 bl_out_6 br_out_6 bl_out_7 br_out_7 bl_out_8 br_out_8 bl_out_9 br_out_9 bl_out_10 br_out_10 bl_out_11 br_out_11 bl_out_12 br_out_12 bl_out_13 br_out_13 bl_out_14 br_out_14 bl_out_15 br_out_15 bl_out_16 br_out_16 bl_out_17 br_out_17 bl_out_18 br_out_18 bl_out_19 br_out_19 bl_out_20 br_out_20 bl_out_21 br_out_21 bl_out_22 br_out_22 bl_out_23 br_out_23 bl_out_24 br_out_24 bl_out_25 br_out_25 bl_out_26 br_out_26 bl_out_27 br_out_27 bl_out_28 br_out_28 bl_out_29 br_out_29 bl_out_30 br_out_30 bl_out_31 br_out_31 gnd
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : sel_0 
* INOUT : sel_1 
* INOUT : bl_out_0 
* INOUT : br_out_0 
* INOUT : bl_out_1 
* INOUT : br_out_1 
* INOUT : bl_out_2 
* INOUT : br_out_2 
* INOUT : bl_out_3 
* INOUT : br_out_3 
* INOUT : bl_out_4 
* INOUT : br_out_4 
* INOUT : bl_out_5 
* INOUT : br_out_5 
* INOUT : bl_out_6 
* INOUT : br_out_6 
* INOUT : bl_out_7 
* INOUT : br_out_7 
* INOUT : bl_out_8 
* INOUT : br_out_8 
* INOUT : bl_out_9 
* INOUT : br_out_9 
* INOUT : bl_out_10 
* INOUT : br_out_10 
* INOUT : bl_out_11 
* INOUT : br_out_11 
* INOUT : bl_out_12 
* INOUT : br_out_12 
* INOUT : bl_out_13 
* INOUT : br_out_13 
* INOUT : bl_out_14 
* INOUT : br_out_14 
* INOUT : bl_out_15 
* INOUT : br_out_15 
* INOUT : bl_out_16 
* INOUT : br_out_16 
* INOUT : bl_out_17 
* INOUT : br_out_17 
* INOUT : bl_out_18 
* INOUT : br_out_18 
* INOUT : bl_out_19 
* INOUT : br_out_19 
* INOUT : bl_out_20 
* INOUT : br_out_20 
* INOUT : bl_out_21 
* INOUT : br_out_21 
* INOUT : bl_out_22 
* INOUT : br_out_22 
* INOUT : bl_out_23 
* INOUT : br_out_23 
* INOUT : bl_out_24 
* INOUT : br_out_24 
* INOUT : bl_out_25 
* INOUT : br_out_25 
* INOUT : bl_out_26 
* INOUT : br_out_26 
* INOUT : bl_out_27 
* INOUT : br_out_27 
* INOUT : bl_out_28 
* INOUT : br_out_28 
* INOUT : bl_out_29 
* INOUT : br_out_29 
* INOUT : bl_out_30 
* INOUT : br_out_30 
* INOUT : bl_out_31 
* INOUT : br_out_31 
* INOUT : gnd 
* cols: 64 word_size: 32 bl: bl0 br: br0
XXMUX0 bl_0 br_0 bl_out_0 br_out_0 sel_0 gnd single_level_column_mux
XXMUX1 bl_1 br_1 bl_out_0 br_out_0 sel_1 gnd single_level_column_mux
XXMUX2 bl_2 br_2 bl_out_1 br_out_1 sel_0 gnd single_level_column_mux
XXMUX3 bl_3 br_3 bl_out_1 br_out_1 sel_1 gnd single_level_column_mux
XXMUX4 bl_4 br_4 bl_out_2 br_out_2 sel_0 gnd single_level_column_mux
XXMUX5 bl_5 br_5 bl_out_2 br_out_2 sel_1 gnd single_level_column_mux
XXMUX6 bl_6 br_6 bl_out_3 br_out_3 sel_0 gnd single_level_column_mux
XXMUX7 bl_7 br_7 bl_out_3 br_out_3 sel_1 gnd single_level_column_mux
XXMUX8 bl_8 br_8 bl_out_4 br_out_4 sel_0 gnd single_level_column_mux
XXMUX9 bl_9 br_9 bl_out_4 br_out_4 sel_1 gnd single_level_column_mux
XXMUX10 bl_10 br_10 bl_out_5 br_out_5 sel_0 gnd single_level_column_mux
XXMUX11 bl_11 br_11 bl_out_5 br_out_5 sel_1 gnd single_level_column_mux
XXMUX12 bl_12 br_12 bl_out_6 br_out_6 sel_0 gnd single_level_column_mux
XXMUX13 bl_13 br_13 bl_out_6 br_out_6 sel_1 gnd single_level_column_mux
XXMUX14 bl_14 br_14 bl_out_7 br_out_7 sel_0 gnd single_level_column_mux
XXMUX15 bl_15 br_15 bl_out_7 br_out_7 sel_1 gnd single_level_column_mux
XXMUX16 bl_16 br_16 bl_out_8 br_out_8 sel_0 gnd single_level_column_mux
XXMUX17 bl_17 br_17 bl_out_8 br_out_8 sel_1 gnd single_level_column_mux
XXMUX18 bl_18 br_18 bl_out_9 br_out_9 sel_0 gnd single_level_column_mux
XXMUX19 bl_19 br_19 bl_out_9 br_out_9 sel_1 gnd single_level_column_mux
XXMUX20 bl_20 br_20 bl_out_10 br_out_10 sel_0 gnd single_level_column_mux
XXMUX21 bl_21 br_21 bl_out_10 br_out_10 sel_1 gnd single_level_column_mux
XXMUX22 bl_22 br_22 bl_out_11 br_out_11 sel_0 gnd single_level_column_mux
XXMUX23 bl_23 br_23 bl_out_11 br_out_11 sel_1 gnd single_level_column_mux
XXMUX24 bl_24 br_24 bl_out_12 br_out_12 sel_0 gnd single_level_column_mux
XXMUX25 bl_25 br_25 bl_out_12 br_out_12 sel_1 gnd single_level_column_mux
XXMUX26 bl_26 br_26 bl_out_13 br_out_13 sel_0 gnd single_level_column_mux
XXMUX27 bl_27 br_27 bl_out_13 br_out_13 sel_1 gnd single_level_column_mux
XXMUX28 bl_28 br_28 bl_out_14 br_out_14 sel_0 gnd single_level_column_mux
XXMUX29 bl_29 br_29 bl_out_14 br_out_14 sel_1 gnd single_level_column_mux
XXMUX30 bl_30 br_30 bl_out_15 br_out_15 sel_0 gnd single_level_column_mux
XXMUX31 bl_31 br_31 bl_out_15 br_out_15 sel_1 gnd single_level_column_mux
XXMUX32 bl_32 br_32 bl_out_16 br_out_16 sel_0 gnd single_level_column_mux
XXMUX33 bl_33 br_33 bl_out_16 br_out_16 sel_1 gnd single_level_column_mux
XXMUX34 bl_34 br_34 bl_out_17 br_out_17 sel_0 gnd single_level_column_mux
XXMUX35 bl_35 br_35 bl_out_17 br_out_17 sel_1 gnd single_level_column_mux
XXMUX36 bl_36 br_36 bl_out_18 br_out_18 sel_0 gnd single_level_column_mux
XXMUX37 bl_37 br_37 bl_out_18 br_out_18 sel_1 gnd single_level_column_mux
XXMUX38 bl_38 br_38 bl_out_19 br_out_19 sel_0 gnd single_level_column_mux
XXMUX39 bl_39 br_39 bl_out_19 br_out_19 sel_1 gnd single_level_column_mux
XXMUX40 bl_40 br_40 bl_out_20 br_out_20 sel_0 gnd single_level_column_mux
XXMUX41 bl_41 br_41 bl_out_20 br_out_20 sel_1 gnd single_level_column_mux
XXMUX42 bl_42 br_42 bl_out_21 br_out_21 sel_0 gnd single_level_column_mux
XXMUX43 bl_43 br_43 bl_out_21 br_out_21 sel_1 gnd single_level_column_mux
XXMUX44 bl_44 br_44 bl_out_22 br_out_22 sel_0 gnd single_level_column_mux
XXMUX45 bl_45 br_45 bl_out_22 br_out_22 sel_1 gnd single_level_column_mux
XXMUX46 bl_46 br_46 bl_out_23 br_out_23 sel_0 gnd single_level_column_mux
XXMUX47 bl_47 br_47 bl_out_23 br_out_23 sel_1 gnd single_level_column_mux
XXMUX48 bl_48 br_48 bl_out_24 br_out_24 sel_0 gnd single_level_column_mux
XXMUX49 bl_49 br_49 bl_out_24 br_out_24 sel_1 gnd single_level_column_mux
XXMUX50 bl_50 br_50 bl_out_25 br_out_25 sel_0 gnd single_level_column_mux
XXMUX51 bl_51 br_51 bl_out_25 br_out_25 sel_1 gnd single_level_column_mux
XXMUX52 bl_52 br_52 bl_out_26 br_out_26 sel_0 gnd single_level_column_mux
XXMUX53 bl_53 br_53 bl_out_26 br_out_26 sel_1 gnd single_level_column_mux
XXMUX54 bl_54 br_54 bl_out_27 br_out_27 sel_0 gnd single_level_column_mux
XXMUX55 bl_55 br_55 bl_out_27 br_out_27 sel_1 gnd single_level_column_mux
XXMUX56 bl_56 br_56 bl_out_28 br_out_28 sel_0 gnd single_level_column_mux
XXMUX57 bl_57 br_57 bl_out_28 br_out_28 sel_1 gnd single_level_column_mux
XXMUX58 bl_58 br_58 bl_out_29 br_out_29 sel_0 gnd single_level_column_mux
XXMUX59 bl_59 br_59 bl_out_29 br_out_29 sel_1 gnd single_level_column_mux
XXMUX60 bl_60 br_60 bl_out_30 br_out_30 sel_0 gnd single_level_column_mux
XXMUX61 bl_61 br_61 bl_out_30 br_out_30 sel_1 gnd single_level_column_mux
XXMUX62 bl_62 br_62 bl_out_31 br_out_31 sel_0 gnd single_level_column_mux
XXMUX63 bl_63 br_63 bl_out_31 br_out_31 sel_1 gnd single_level_column_mux
.ENDS single_level_column_mux_array
*********************** "write_driver" ******************************

.SUBCKT write_driver din bl br en vdd gnd

**** Inverter to conver Data_in to data_in_bar ******
* din_bar = sky130_fd_pr__model__typical__inv(din)
XM_1 din_bar din gnd gnd sky130_fd_pr__nfet_01v8 W=0.36 L=0.15 m=1
XM_2 din_bar din vdd vdd sky130_fd_pr__pfet_01v8 W=0.55 L=0.15 m=1

**** 2input nand gate follwed by inverter to drive BL ******
* din_bar_gated = nand(en, din)
XM_3 din_bar_gated en net_7 gnd sky130_fd_pr__nfet_01v8 W=0.55 L=0.15 m=1
XM_4 net_7 din gnd gnd sky130_fd_pr__nfet_01v8 W=0.55 L=0.15 m=1
XM_5 din_bar_gated en vdd vdd sky130_fd_pr__pfet_01v8 W=0.55 L=0.15 m=1
XM_6 din_bar_gated din vdd vdd sky130_fd_pr__pfet_01v8 W=0.55 L=0.15 m=1
* din_bar_gated_bar = sky130_fd_pr__model__typical__inv(din_bar_gated)
XM_7 din_bar_gated_bar din_bar_gated vdd vdd sky130_fd_pr__pfet_01v8 W=0.55 L=0.15 m=1
XM_8 din_bar_gated_bar din_bar_gated gnd gnd sky130_fd_pr__nfet_01v8 W=0.36 L=0.15 m=1

**** 2input nand gate follwed by inverter to drive BR******
* din_gated = nand(en, din_bar)
XM_9 din_gated en vdd vdd sky130_fd_pr__pfet_01v8 W=0.55 L=0.15 m=1
XM_10 din_gated en net_8 gnd sky130_fd_pr__nfet_01v8 W=0.55 L=0.15 m=1
XM_11 net_8 din_bar gnd gnd sky130_fd_pr__nfet_01v8 W=0.55 L=0.15 m=1
XM_12 din_gated din_bar vdd vdd sky130_fd_pr__pfet_01v8 W=0.55 L=0.15 m=1
* din_gated_bar = sky130_fd_pr__model__typical__inv(din_gated)
XM_13 din_gated_bar din_gated vdd vdd sky130_fd_pr__pfet_01v8 W=0.55 L=0.15 m=1
XM_14 din_gated_bar din_gated gnd gnd sky130_fd_pr__nfet_01v8 W=0.36 L=0.15 m=1

************************************************
* pull down with en enable
XM_15 bl din_gated_bar gnd gnd sky130_fd_pr__nfet_01v8 W=1 L=0.15 m=1
XM_16 br din_bar_gated_bar gnd gnd sky130_fd_pr__nfet_01v8 W=1 L=0.15 m=1

.ENDS write_driver

.SUBCKT write_driver_array data_0 data_1 data_2 data_3 data_4 data_5 data_6 data_7 data_8 data_9 data_10 data_11 data_12 data_13 data_14 data_15 data_16 data_17 data_18 data_19 data_20 data_21 data_22 data_23 data_24 data_25 data_26 data_27 data_28 data_29 data_30 data_31 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 en_0 en_1 en_2 en_3 vdd gnd
* INPUT : data_0 
* INPUT : data_1 
* INPUT : data_2 
* INPUT : data_3 
* INPUT : data_4 
* INPUT : data_5 
* INPUT : data_6 
* INPUT : data_7 
* INPUT : data_8 
* INPUT : data_9 
* INPUT : data_10 
* INPUT : data_11 
* INPUT : data_12 
* INPUT : data_13 
* INPUT : data_14 
* INPUT : data_15 
* INPUT : data_16 
* INPUT : data_17 
* INPUT : data_18 
* INPUT : data_19 
* INPUT : data_20 
* INPUT : data_21 
* INPUT : data_22 
* INPUT : data_23 
* INPUT : data_24 
* INPUT : data_25 
* INPUT : data_26 
* INPUT : data_27 
* INPUT : data_28 
* INPUT : data_29 
* INPUT : data_30 
* INPUT : data_31 
* OUTPUT: bl_0 
* OUTPUT: br_0 
* OUTPUT: bl_1 
* OUTPUT: br_1 
* OUTPUT: bl_2 
* OUTPUT: br_2 
* OUTPUT: bl_3 
* OUTPUT: br_3 
* OUTPUT: bl_4 
* OUTPUT: br_4 
* OUTPUT: bl_5 
* OUTPUT: br_5 
* OUTPUT: bl_6 
* OUTPUT: br_6 
* OUTPUT: bl_7 
* OUTPUT: br_7 
* OUTPUT: bl_8 
* OUTPUT: br_8 
* OUTPUT: bl_9 
* OUTPUT: br_9 
* OUTPUT: bl_10 
* OUTPUT: br_10 
* OUTPUT: bl_11 
* OUTPUT: br_11 
* OUTPUT: bl_12 
* OUTPUT: br_12 
* OUTPUT: bl_13 
* OUTPUT: br_13 
* OUTPUT: bl_14 
* OUTPUT: br_14 
* OUTPUT: bl_15 
* OUTPUT: br_15 
* OUTPUT: bl_16 
* OUTPUT: br_16 
* OUTPUT: bl_17 
* OUTPUT: br_17 
* OUTPUT: bl_18 
* OUTPUT: br_18 
* OUTPUT: bl_19 
* OUTPUT: br_19 
* OUTPUT: bl_20 
* OUTPUT: br_20 
* OUTPUT: bl_21 
* OUTPUT: br_21 
* OUTPUT: bl_22 
* OUTPUT: br_22 
* OUTPUT: bl_23 
* OUTPUT: br_23 
* OUTPUT: bl_24 
* OUTPUT: br_24 
* OUTPUT: bl_25 
* OUTPUT: br_25 
* OUTPUT: bl_26 
* OUTPUT: br_26 
* OUTPUT: bl_27 
* OUTPUT: br_27 
* OUTPUT: bl_28 
* OUTPUT: br_28 
* OUTPUT: bl_29 
* OUTPUT: br_29 
* OUTPUT: bl_30 
* OUTPUT: br_30 
* OUTPUT: bl_31 
* OUTPUT: br_31 
* INPUT : en_0 
* INPUT : en_1 
* INPUT : en_2 
* INPUT : en_3 
* POWER : vdd 
* GROUND: gnd 
* word_size 32
Xwrite_driver0 data_0 bl_0 br_0 en_0 vdd gnd write_driver
Xwrite_driver2 data_1 bl_1 br_1 en_0 vdd gnd write_driver
Xwrite_driver4 data_2 bl_2 br_2 en_0 vdd gnd write_driver
Xwrite_driver6 data_3 bl_3 br_3 en_0 vdd gnd write_driver
Xwrite_driver8 data_4 bl_4 br_4 en_0 vdd gnd write_driver
Xwrite_driver10 data_5 bl_5 br_5 en_0 vdd gnd write_driver
Xwrite_driver12 data_6 bl_6 br_6 en_0 vdd gnd write_driver
Xwrite_driver14 data_7 bl_7 br_7 en_0 vdd gnd write_driver
Xwrite_driver16 data_8 bl_8 br_8 en_1 vdd gnd write_driver
Xwrite_driver18 data_9 bl_9 br_9 en_1 vdd gnd write_driver
Xwrite_driver20 data_10 bl_10 br_10 en_1 vdd gnd write_driver
Xwrite_driver22 data_11 bl_11 br_11 en_1 vdd gnd write_driver
Xwrite_driver24 data_12 bl_12 br_12 en_1 vdd gnd write_driver
Xwrite_driver26 data_13 bl_13 br_13 en_1 vdd gnd write_driver
Xwrite_driver28 data_14 bl_14 br_14 en_1 vdd gnd write_driver
Xwrite_driver30 data_15 bl_15 br_15 en_1 vdd gnd write_driver
Xwrite_driver32 data_16 bl_16 br_16 en_2 vdd gnd write_driver
Xwrite_driver34 data_17 bl_17 br_17 en_2 vdd gnd write_driver
Xwrite_driver36 data_18 bl_18 br_18 en_2 vdd gnd write_driver
Xwrite_driver38 data_19 bl_19 br_19 en_2 vdd gnd write_driver
Xwrite_driver40 data_20 bl_20 br_20 en_2 vdd gnd write_driver
Xwrite_driver42 data_21 bl_21 br_21 en_2 vdd gnd write_driver
Xwrite_driver44 data_22 bl_22 br_22 en_2 vdd gnd write_driver
Xwrite_driver46 data_23 bl_23 br_23 en_2 vdd gnd write_driver
Xwrite_driver48 data_24 bl_24 br_24 en_3 vdd gnd write_driver
Xwrite_driver50 data_25 bl_25 br_25 en_3 vdd gnd write_driver
Xwrite_driver52 data_26 bl_26 br_26 en_3 vdd gnd write_driver
Xwrite_driver54 data_27 bl_27 br_27 en_3 vdd gnd write_driver
Xwrite_driver56 data_28 bl_28 br_28 en_3 vdd gnd write_driver
Xwrite_driver58 data_29 bl_29 br_29 en_3 vdd gnd write_driver
Xwrite_driver60 data_30 bl_30 br_30 en_3 vdd gnd write_driver
Xwrite_driver62 data_31 bl_31 br_31 en_3 vdd gnd write_driver
.ENDS write_driver_array

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u

* ptx M{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u

.SUBCKT pnand2 A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpnand2_pmos1 vdd A Z vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
XMpnand2_pmos2 Z B vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
XMpnand2_nmos1 Z B net1 gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
XMpnand2_nmos2 net1 A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS pnand2

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u

* ptx M{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u

.SUBCKT pinv A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS pinv

.SUBCKT pdriver A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [2.0]
Xbuf_inv1 A Z vdd gnd pinv
.ENDS pdriver

.SUBCKT pand2 A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpand2_nand A B zb_int vdd gnd pnand2
Xpand2_inv zb_int Z vdd gnd pdriver
.ENDS pand2

.SUBCKT write_mask_and_array wmask_in_0 wmask_in_1 wmask_in_2 wmask_in_3 en wmask_out_0 wmask_out_1 wmask_out_2 wmask_out_3 vdd gnd
* INPUT : wmask_in_0 
* INPUT : wmask_in_1 
* INPUT : wmask_in_2 
* INPUT : wmask_in_3 
* INPUT : en 
* OUTPUT: wmask_out_0 
* OUTPUT: wmask_out_1 
* OUTPUT: wmask_out_2 
* OUTPUT: wmask_out_3 
* POWER : vdd 
* GROUND: gnd 
* write_size 8
Xand2_0 wmask_in_0 en wmask_out_0 vdd gnd pand2
Xand2_1 wmask_in_1 en wmask_out_1 vdd gnd pand2
Xand2_2 wmask_in_2 en wmask_out_2 vdd gnd pand2
Xand2_3 wmask_in_3 en wmask_out_3 vdd gnd pand2
.ENDS write_mask_and_array

.SUBCKT port_data rbl_bl rbl_br bl0_0 br0_0 bl0_1 br0_1 bl0_2 br0_2 bl0_3 br0_3 bl0_4 br0_4 bl0_5 br0_5 bl0_6 br0_6 bl0_7 br0_7 bl0_8 br0_8 bl0_9 br0_9 bl0_10 br0_10 bl0_11 br0_11 bl0_12 br0_12 bl0_13 br0_13 bl0_14 br0_14 bl0_15 br0_15 bl0_16 br0_16 bl0_17 br0_17 bl0_18 br0_18 bl0_19 br0_19 bl0_20 br0_20 bl0_21 br0_21 bl0_22 br0_22 bl0_23 br0_23 bl0_24 br0_24 bl0_25 br0_25 bl0_26 br0_26 bl0_27 br0_27 bl0_28 br0_28 bl0_29 br0_29 bl0_30 br0_30 bl0_31 br0_31 bl0_32 br0_32 bl0_33 br0_33 bl0_34 br0_34 bl0_35 br0_35 bl0_36 br0_36 bl0_37 br0_37 bl0_38 br0_38 bl0_39 br0_39 bl0_40 br0_40 bl0_41 br0_41 bl0_42 br0_42 bl0_43 br0_43 bl0_44 br0_44 bl0_45 br0_45 bl0_46 br0_46 bl0_47 br0_47 bl0_48 br0_48 bl0_49 br0_49 bl0_50 br0_50 bl0_51 br0_51 bl0_52 br0_52 bl0_53 br0_53 bl0_54 br0_54 bl0_55 br0_55 bl0_56 br0_56 bl0_57 br0_57 bl0_58 br0_58 bl0_59 br0_59 bl0_60 br0_60 bl0_61 br0_61 bl0_62 br0_62 bl0_63 br0_63 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5 dout_6 dout_7 dout_8 dout_9 dout_10 dout_11 dout_12 dout_13 dout_14 dout_15 dout_16 dout_17 dout_18 dout_19 dout_20 dout_21 dout_22 dout_23 dout_24 dout_25 dout_26 dout_27 dout_28 dout_29 dout_30 dout_31 din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10 din_11 din_12 din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20 din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30 din_31 sel_0 sel_1 s_en p_en_bar w_en bank_wmask_0 bank_wmask_1 bank_wmask_2 bank_wmask_3 vdd gnd
* INOUT : rbl_bl 
* INOUT : rbl_br 
* INOUT : bl0_0 
* INOUT : br0_0 
* INOUT : bl0_1 
* INOUT : br0_1 
* INOUT : bl0_2 
* INOUT : br0_2 
* INOUT : bl0_3 
* INOUT : br0_3 
* INOUT : bl0_4 
* INOUT : br0_4 
* INOUT : bl0_5 
* INOUT : br0_5 
* INOUT : bl0_6 
* INOUT : br0_6 
* INOUT : bl0_7 
* INOUT : br0_7 
* INOUT : bl0_8 
* INOUT : br0_8 
* INOUT : bl0_9 
* INOUT : br0_9 
* INOUT : bl0_10 
* INOUT : br0_10 
* INOUT : bl0_11 
* INOUT : br0_11 
* INOUT : bl0_12 
* INOUT : br0_12 
* INOUT : bl0_13 
* INOUT : br0_13 
* INOUT : bl0_14 
* INOUT : br0_14 
* INOUT : bl0_15 
* INOUT : br0_15 
* INOUT : bl0_16 
* INOUT : br0_16 
* INOUT : bl0_17 
* INOUT : br0_17 
* INOUT : bl0_18 
* INOUT : br0_18 
* INOUT : bl0_19 
* INOUT : br0_19 
* INOUT : bl0_20 
* INOUT : br0_20 
* INOUT : bl0_21 
* INOUT : br0_21 
* INOUT : bl0_22 
* INOUT : br0_22 
* INOUT : bl0_23 
* INOUT : br0_23 
* INOUT : bl0_24 
* INOUT : br0_24 
* INOUT : bl0_25 
* INOUT : br0_25 
* INOUT : bl0_26 
* INOUT : br0_26 
* INOUT : bl0_27 
* INOUT : br0_27 
* INOUT : bl0_28 
* INOUT : br0_28 
* INOUT : bl0_29 
* INOUT : br0_29 
* INOUT : bl0_30 
* INOUT : br0_30 
* INOUT : bl0_31 
* INOUT : br0_31 
* INOUT : bl0_32 
* INOUT : br0_32 
* INOUT : bl0_33 
* INOUT : br0_33 
* INOUT : bl0_34 
* INOUT : br0_34 
* INOUT : bl0_35 
* INOUT : br0_35 
* INOUT : bl0_36 
* INOUT : br0_36 
* INOUT : bl0_37 
* INOUT : br0_37 
* INOUT : bl0_38 
* INOUT : br0_38 
* INOUT : bl0_39 
* INOUT : br0_39 
* INOUT : bl0_40 
* INOUT : br0_40 
* INOUT : bl0_41 
* INOUT : br0_41 
* INOUT : bl0_42 
* INOUT : br0_42 
* INOUT : bl0_43 
* INOUT : br0_43 
* INOUT : bl0_44 
* INOUT : br0_44 
* INOUT : bl0_45 
* INOUT : br0_45 
* INOUT : bl0_46 
* INOUT : br0_46 
* INOUT : bl0_47 
* INOUT : br0_47 
* INOUT : bl0_48 
* INOUT : br0_48 
* INOUT : bl0_49 
* INOUT : br0_49 
* INOUT : bl0_50 
* INOUT : br0_50 
* INOUT : bl0_51 
* INOUT : br0_51 
* INOUT : bl0_52 
* INOUT : br0_52 
* INOUT : bl0_53 
* INOUT : br0_53 
* INOUT : bl0_54 
* INOUT : br0_54 
* INOUT : bl0_55 
* INOUT : br0_55 
* INOUT : bl0_56 
* INOUT : br0_56 
* INOUT : bl0_57 
* INOUT : br0_57 
* INOUT : bl0_58 
* INOUT : br0_58 
* INOUT : bl0_59 
* INOUT : br0_59 
* INOUT : bl0_60 
* INOUT : br0_60 
* INOUT : bl0_61 
* INOUT : br0_61 
* INOUT : bl0_62 
* INOUT : br0_62 
* INOUT : bl0_63 
* INOUT : br0_63 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* OUTPUT: dout_7 
* OUTPUT: dout_8 
* OUTPUT: dout_9 
* OUTPUT: dout_10 
* OUTPUT: dout_11 
* OUTPUT: dout_12 
* OUTPUT: dout_13 
* OUTPUT: dout_14 
* OUTPUT: dout_15 
* OUTPUT: dout_16 
* OUTPUT: dout_17 
* OUTPUT: dout_18 
* OUTPUT: dout_19 
* OUTPUT: dout_20 
* OUTPUT: dout_21 
* OUTPUT: dout_22 
* OUTPUT: dout_23 
* OUTPUT: dout_24 
* OUTPUT: dout_25 
* OUTPUT: dout_26 
* OUTPUT: dout_27 
* OUTPUT: dout_28 
* OUTPUT: dout_29 
* OUTPUT: dout_30 
* OUTPUT: dout_31 
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* INPUT : din_7 
* INPUT : din_8 
* INPUT : din_9 
* INPUT : din_10 
* INPUT : din_11 
* INPUT : din_12 
* INPUT : din_13 
* INPUT : din_14 
* INPUT : din_15 
* INPUT : din_16 
* INPUT : din_17 
* INPUT : din_18 
* INPUT : din_19 
* INPUT : din_20 
* INPUT : din_21 
* INPUT : din_22 
* INPUT : din_23 
* INPUT : din_24 
* INPUT : din_25 
* INPUT : din_26 
* INPUT : din_27 
* INPUT : din_28 
* INPUT : din_29 
* INPUT : din_30 
* INPUT : din_31 
* INPUT : sel_0 
* INPUT : sel_1 
* INPUT : s_en 
* INPUT : p_en_bar 
* INPUT : w_en 
* INPUT : bank_wmask_0 
* INPUT : bank_wmask_1 
* INPUT : bank_wmask_2 
* INPUT : bank_wmask_3 
* POWER : vdd 
* GROUND: gnd 
Xprecharge_array0 rbl_bl rbl_br bl0_0 br0_0 bl0_1 br0_1 bl0_2 br0_2 bl0_3 br0_3 bl0_4 br0_4 bl0_5 br0_5 bl0_6 br0_6 bl0_7 br0_7 bl0_8 br0_8 bl0_9 br0_9 bl0_10 br0_10 bl0_11 br0_11 bl0_12 br0_12 bl0_13 br0_13 bl0_14 br0_14 bl0_15 br0_15 bl0_16 br0_16 bl0_17 br0_17 bl0_18 br0_18 bl0_19 br0_19 bl0_20 br0_20 bl0_21 br0_21 bl0_22 br0_22 bl0_23 br0_23 bl0_24 br0_24 bl0_25 br0_25 bl0_26 br0_26 bl0_27 br0_27 bl0_28 br0_28 bl0_29 br0_29 bl0_30 br0_30 bl0_31 br0_31 bl0_32 br0_32 bl0_33 br0_33 bl0_34 br0_34 bl0_35 br0_35 bl0_36 br0_36 bl0_37 br0_37 bl0_38 br0_38 bl0_39 br0_39 bl0_40 br0_40 bl0_41 br0_41 bl0_42 br0_42 bl0_43 br0_43 bl0_44 br0_44 bl0_45 br0_45 bl0_46 br0_46 bl0_47 br0_47 bl0_48 br0_48 bl0_49 br0_49 bl0_50 br0_50 bl0_51 br0_51 bl0_52 br0_52 bl0_53 br0_53 bl0_54 br0_54 bl0_55 br0_55 bl0_56 br0_56 bl0_57 br0_57 bl0_58 br0_58 bl0_59 br0_59 bl0_60 br0_60 bl0_61 br0_61 bl0_62 br0_62 bl0_63 br0_63 p_en_bar vdd precharge_array
Xsense_amp_array0 dout_0 bl0_out_0 br0_out_0 dout_1 bl0_out_1 br0_out_1 dout_2 bl0_out_2 br0_out_2 dout_3 bl0_out_3 br0_out_3 dout_4 bl0_out_4 br0_out_4 dout_5 bl0_out_5 br0_out_5 dout_6 bl0_out_6 br0_out_6 dout_7 bl0_out_7 br0_out_7 dout_8 bl0_out_8 br0_out_8 dout_9 bl0_out_9 br0_out_9 dout_10 bl0_out_10 br0_out_10 dout_11 bl0_out_11 br0_out_11 dout_12 bl0_out_12 br0_out_12 dout_13 bl0_out_13 br0_out_13 dout_14 bl0_out_14 br0_out_14 dout_15 bl0_out_15 br0_out_15 dout_16 bl0_out_16 br0_out_16 dout_17 bl0_out_17 br0_out_17 dout_18 bl0_out_18 br0_out_18 dout_19 bl0_out_19 br0_out_19 dout_20 bl0_out_20 br0_out_20 dout_21 bl0_out_21 br0_out_21 dout_22 bl0_out_22 br0_out_22 dout_23 bl0_out_23 br0_out_23 dout_24 bl0_out_24 br0_out_24 dout_25 bl0_out_25 br0_out_25 dout_26 bl0_out_26 br0_out_26 dout_27 bl0_out_27 br0_out_27 dout_28 bl0_out_28 br0_out_28 dout_29 bl0_out_29 br0_out_29 dout_30 bl0_out_30 br0_out_30 dout_31 bl0_out_31 br0_out_31 s_en vdd gnd sense_amp_array
Xwrite_driver_array0 din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10 din_11 din_12 din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20 din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30 din_31 bl0_out_0 br0_out_0 bl0_out_1 br0_out_1 bl0_out_2 br0_out_2 bl0_out_3 br0_out_3 bl0_out_4 br0_out_4 bl0_out_5 br0_out_5 bl0_out_6 br0_out_6 bl0_out_7 br0_out_7 bl0_out_8 br0_out_8 bl0_out_9 br0_out_9 bl0_out_10 br0_out_10 bl0_out_11 br0_out_11 bl0_out_12 br0_out_12 bl0_out_13 br0_out_13 bl0_out_14 br0_out_14 bl0_out_15 br0_out_15 bl0_out_16 br0_out_16 bl0_out_17 br0_out_17 bl0_out_18 br0_out_18 bl0_out_19 br0_out_19 bl0_out_20 br0_out_20 bl0_out_21 br0_out_21 bl0_out_22 br0_out_22 bl0_out_23 br0_out_23 bl0_out_24 br0_out_24 bl0_out_25 br0_out_25 bl0_out_26 br0_out_26 bl0_out_27 br0_out_27 bl0_out_28 br0_out_28 bl0_out_29 br0_out_29 bl0_out_30 br0_out_30 bl0_out_31 br0_out_31 wdriver_sel_0 wdriver_sel_1 wdriver_sel_2 wdriver_sel_3 vdd gnd write_driver_array
Xwrite_mask_and_array0 bank_wmask_0 bank_wmask_1 bank_wmask_2 bank_wmask_3 w_en wdriver_sel_0 wdriver_sel_1 wdriver_sel_2 wdriver_sel_3 vdd gnd write_mask_and_array
Xcolumn_mux_array0 bl0_0 br0_0 bl0_1 br0_1 bl0_2 br0_2 bl0_3 br0_3 bl0_4 br0_4 bl0_5 br0_5 bl0_6 br0_6 bl0_7 br0_7 bl0_8 br0_8 bl0_9 br0_9 bl0_10 br0_10 bl0_11 br0_11 bl0_12 br0_12 bl0_13 br0_13 bl0_14 br0_14 bl0_15 br0_15 bl0_16 br0_16 bl0_17 br0_17 bl0_18 br0_18 bl0_19 br0_19 bl0_20 br0_20 bl0_21 br0_21 bl0_22 br0_22 bl0_23 br0_23 bl0_24 br0_24 bl0_25 br0_25 bl0_26 br0_26 bl0_27 br0_27 bl0_28 br0_28 bl0_29 br0_29 bl0_30 br0_30 bl0_31 br0_31 bl0_32 br0_32 bl0_33 br0_33 bl0_34 br0_34 bl0_35 br0_35 bl0_36 br0_36 bl0_37 br0_37 bl0_38 br0_38 bl0_39 br0_39 bl0_40 br0_40 bl0_41 br0_41 bl0_42 br0_42 bl0_43 br0_43 bl0_44 br0_44 bl0_45 br0_45 bl0_46 br0_46 bl0_47 br0_47 bl0_48 br0_48 bl0_49 br0_49 bl0_50 br0_50 bl0_51 br0_51 bl0_52 br0_52 bl0_53 br0_53 bl0_54 br0_54 bl0_55 br0_55 bl0_56 br0_56 bl0_57 br0_57 bl0_58 br0_58 bl0_59 br0_59 bl0_60 br0_60 bl0_61 br0_61 bl0_62 br0_62 bl0_63 br0_63 sel_0 sel_1 bl0_out_0 br0_out_0 bl0_out_1 br0_out_1 bl0_out_2 br0_out_2 bl0_out_3 br0_out_3 bl0_out_4 br0_out_4 bl0_out_5 br0_out_5 bl0_out_6 br0_out_6 bl0_out_7 br0_out_7 bl0_out_8 br0_out_8 bl0_out_9 br0_out_9 bl0_out_10 br0_out_10 bl0_out_11 br0_out_11 bl0_out_12 br0_out_12 bl0_out_13 br0_out_13 bl0_out_14 br0_out_14 bl0_out_15 br0_out_15 bl0_out_16 br0_out_16 bl0_out_17 br0_out_17 bl0_out_18 br0_out_18 bl0_out_19 br0_out_19 bl0_out_20 br0_out_20 bl0_out_21 br0_out_21 bl0_out_22 br0_out_22 bl0_out_23 br0_out_23 bl0_out_24 br0_out_24 bl0_out_25 br0_out_25 bl0_out_26 br0_out_26 bl0_out_27 br0_out_27 bl0_out_28 br0_out_28 bl0_out_29 br0_out_29 bl0_out_30 br0_out_30 bl0_out_31 br0_out_31 gnd single_level_column_mux_array
.ENDS port_data

.SUBCKT precharge_1 bl br en_bar vdd
* OUTPUT: bl 
* OUTPUT: br 
* INPUT : en_bar 
* POWER : vdd 
XMlower_pmos bl en_bar br vdd sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=0.15 pd=1.40 ps=1.40 as=0.21u ad=0.21u
XMupper_pmos1 bl en_bar vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=0.15 pd=1.40 ps=1.40 as=0.21u ad=0.21u
XMupper_pmos2 br en_bar vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=0.15 pd=1.40 ps=1.40 as=0.21u ad=0.21u
.ENDS precharge_1

.SUBCKT precharge_array_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 en_bar vdd
* OUTPUT: bl_0 
* OUTPUT: br_0 
* OUTPUT: bl_1 
* OUTPUT: br_1 
* OUTPUT: bl_2 
* OUTPUT: br_2 
* OUTPUT: bl_3 
* OUTPUT: br_3 
* OUTPUT: bl_4 
* OUTPUT: br_4 
* OUTPUT: bl_5 
* OUTPUT: br_5 
* OUTPUT: bl_6 
* OUTPUT: br_6 
* OUTPUT: bl_7 
* OUTPUT: br_7 
* OUTPUT: bl_8 
* OUTPUT: br_8 
* OUTPUT: bl_9 
* OUTPUT: br_9 
* OUTPUT: bl_10 
* OUTPUT: br_10 
* OUTPUT: bl_11 
* OUTPUT: br_11 
* OUTPUT: bl_12 
* OUTPUT: br_12 
* OUTPUT: bl_13 
* OUTPUT: br_13 
* OUTPUT: bl_14 
* OUTPUT: br_14 
* OUTPUT: bl_15 
* OUTPUT: br_15 
* OUTPUT: bl_16 
* OUTPUT: br_16 
* OUTPUT: bl_17 
* OUTPUT: br_17 
* OUTPUT: bl_18 
* OUTPUT: br_18 
* OUTPUT: bl_19 
* OUTPUT: br_19 
* OUTPUT: bl_20 
* OUTPUT: br_20 
* OUTPUT: bl_21 
* OUTPUT: br_21 
* OUTPUT: bl_22 
* OUTPUT: br_22 
* OUTPUT: bl_23 
* OUTPUT: br_23 
* OUTPUT: bl_24 
* OUTPUT: br_24 
* OUTPUT: bl_25 
* OUTPUT: br_25 
* OUTPUT: bl_26 
* OUTPUT: br_26 
* OUTPUT: bl_27 
* OUTPUT: br_27 
* OUTPUT: bl_28 
* OUTPUT: br_28 
* OUTPUT: bl_29 
* OUTPUT: br_29 
* OUTPUT: bl_30 
* OUTPUT: br_30 
* OUTPUT: bl_31 
* OUTPUT: br_31 
* OUTPUT: bl_32 
* OUTPUT: br_32 
* OUTPUT: bl_33 
* OUTPUT: br_33 
* OUTPUT: bl_34 
* OUTPUT: br_34 
* OUTPUT: bl_35 
* OUTPUT: br_35 
* OUTPUT: bl_36 
* OUTPUT: br_36 
* OUTPUT: bl_37 
* OUTPUT: br_37 
* OUTPUT: bl_38 
* OUTPUT: br_38 
* OUTPUT: bl_39 
* OUTPUT: br_39 
* OUTPUT: bl_40 
* OUTPUT: br_40 
* OUTPUT: bl_41 
* OUTPUT: br_41 
* OUTPUT: bl_42 
* OUTPUT: br_42 
* OUTPUT: bl_43 
* OUTPUT: br_43 
* OUTPUT: bl_44 
* OUTPUT: br_44 
* OUTPUT: bl_45 
* OUTPUT: br_45 
* OUTPUT: bl_46 
* OUTPUT: br_46 
* OUTPUT: bl_47 
* OUTPUT: br_47 
* OUTPUT: bl_48 
* OUTPUT: br_48 
* OUTPUT: bl_49 
* OUTPUT: br_49 
* OUTPUT: bl_50 
* OUTPUT: br_50 
* OUTPUT: bl_51 
* OUTPUT: br_51 
* OUTPUT: bl_52 
* OUTPUT: br_52 
* OUTPUT: bl_53 
* OUTPUT: br_53 
* OUTPUT: bl_54 
* OUTPUT: br_54 
* OUTPUT: bl_55 
* OUTPUT: br_55 
* OUTPUT: bl_56 
* OUTPUT: br_56 
* OUTPUT: bl_57 
* OUTPUT: br_57 
* OUTPUT: bl_58 
* OUTPUT: br_58 
* OUTPUT: bl_59 
* OUTPUT: br_59 
* OUTPUT: bl_60 
* OUTPUT: br_60 
* OUTPUT: bl_61 
* OUTPUT: br_61 
* OUTPUT: bl_62 
* OUTPUT: br_62 
* OUTPUT: bl_63 
* OUTPUT: br_63 
* OUTPUT: bl_64 
* OUTPUT: br_64 
* INPUT : en_bar 
* POWER : vdd 
* cols: 65 size: 1 bl: bl1 br: br1
Xpre_column_0 bl_0 br_0 en_bar vdd precharge_1
Xpre_column_1 bl_1 br_1 en_bar vdd precharge_1
Xpre_column_2 bl_2 br_2 en_bar vdd precharge_1
Xpre_column_3 bl_3 br_3 en_bar vdd precharge_1
Xpre_column_4 bl_4 br_4 en_bar vdd precharge_1
Xpre_column_5 bl_5 br_5 en_bar vdd precharge_1
Xpre_column_6 bl_6 br_6 en_bar vdd precharge_1
Xpre_column_7 bl_7 br_7 en_bar vdd precharge_1
Xpre_column_8 bl_8 br_8 en_bar vdd precharge_1
Xpre_column_9 bl_9 br_9 en_bar vdd precharge_1
Xpre_column_10 bl_10 br_10 en_bar vdd precharge_1
Xpre_column_11 bl_11 br_11 en_bar vdd precharge_1
Xpre_column_12 bl_12 br_12 en_bar vdd precharge_1
Xpre_column_13 bl_13 br_13 en_bar vdd precharge_1
Xpre_column_14 bl_14 br_14 en_bar vdd precharge_1
Xpre_column_15 bl_15 br_15 en_bar vdd precharge_1
Xpre_column_16 bl_16 br_16 en_bar vdd precharge_1
Xpre_column_17 bl_17 br_17 en_bar vdd precharge_1
Xpre_column_18 bl_18 br_18 en_bar vdd precharge_1
Xpre_column_19 bl_19 br_19 en_bar vdd precharge_1
Xpre_column_20 bl_20 br_20 en_bar vdd precharge_1
Xpre_column_21 bl_21 br_21 en_bar vdd precharge_1
Xpre_column_22 bl_22 br_22 en_bar vdd precharge_1
Xpre_column_23 bl_23 br_23 en_bar vdd precharge_1
Xpre_column_24 bl_24 br_24 en_bar vdd precharge_1
Xpre_column_25 bl_25 br_25 en_bar vdd precharge_1
Xpre_column_26 bl_26 br_26 en_bar vdd precharge_1
Xpre_column_27 bl_27 br_27 en_bar vdd precharge_1
Xpre_column_28 bl_28 br_28 en_bar vdd precharge_1
Xpre_column_29 bl_29 br_29 en_bar vdd precharge_1
Xpre_column_30 bl_30 br_30 en_bar vdd precharge_1
Xpre_column_31 bl_31 br_31 en_bar vdd precharge_1
Xpre_column_32 bl_32 br_32 en_bar vdd precharge_1
Xpre_column_33 bl_33 br_33 en_bar vdd precharge_1
Xpre_column_34 bl_34 br_34 en_bar vdd precharge_1
Xpre_column_35 bl_35 br_35 en_bar vdd precharge_1
Xpre_column_36 bl_36 br_36 en_bar vdd precharge_1
Xpre_column_37 bl_37 br_37 en_bar vdd precharge_1
Xpre_column_38 bl_38 br_38 en_bar vdd precharge_1
Xpre_column_39 bl_39 br_39 en_bar vdd precharge_1
Xpre_column_40 bl_40 br_40 en_bar vdd precharge_1
Xpre_column_41 bl_41 br_41 en_bar vdd precharge_1
Xpre_column_42 bl_42 br_42 en_bar vdd precharge_1
Xpre_column_43 bl_43 br_43 en_bar vdd precharge_1
Xpre_column_44 bl_44 br_44 en_bar vdd precharge_1
Xpre_column_45 bl_45 br_45 en_bar vdd precharge_1
Xpre_column_46 bl_46 br_46 en_bar vdd precharge_1
Xpre_column_47 bl_47 br_47 en_bar vdd precharge_1
Xpre_column_48 bl_48 br_48 en_bar vdd precharge_1
Xpre_column_49 bl_49 br_49 en_bar vdd precharge_1
Xpre_column_50 bl_50 br_50 en_bar vdd precharge_1
Xpre_column_51 bl_51 br_51 en_bar vdd precharge_1
Xpre_column_52 bl_52 br_52 en_bar vdd precharge_1
Xpre_column_53 bl_53 br_53 en_bar vdd precharge_1
Xpre_column_54 bl_54 br_54 en_bar vdd precharge_1
Xpre_column_55 bl_55 br_55 en_bar vdd precharge_1
Xpre_column_56 bl_56 br_56 en_bar vdd precharge_1
Xpre_column_57 bl_57 br_57 en_bar vdd precharge_1
Xpre_column_58 bl_58 br_58 en_bar vdd precharge_1
Xpre_column_59 bl_59 br_59 en_bar vdd precharge_1
Xpre_column_60 bl_60 br_60 en_bar vdd precharge_1
Xpre_column_61 bl_61 br_61 en_bar vdd precharge_1
Xpre_column_62 bl_62 br_62 en_bar vdd precharge_1
Xpre_column_63 bl_63 br_63 en_bar vdd precharge_1
Xpre_column_64 bl_64 br_64 en_bar vdd precharge_1
.ENDS precharge_array_0

.SUBCKT single_level_column_mux_0 bl br bl_out br_out sel gnd
* INOUT : bl 
* INOUT : br 
* INOUT : bl_out 
* INOUT : br_out 
* INOUT : sel 
* INOUT : gnd 
XMmux_tx1 bl sel bl_out gnd sky130_fd_pr__nfet_01v8 m=1 w=3.0 l=0.15 pd=6.06 ps=6.06 as=1.08u ad=1.08u
XMmux_tx2 br sel br_out gnd sky130_fd_pr__nfet_01v8 m=1 w=3.0 l=0.15 pd=6.06 ps=6.06 as=1.08u ad=1.08u
.ENDS single_level_column_mux_0

.SUBCKT single_level_column_mux_array_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 sel_0 sel_1 bl_out_0 br_out_0 bl_out_1 br_out_1 bl_out_2 br_out_2 bl_out_3 br_out_3 bl_out_4 br_out_4 bl_out_5 br_out_5 bl_out_6 br_out_6 bl_out_7 br_out_7 bl_out_8 br_out_8 bl_out_9 br_out_9 bl_out_10 br_out_10 bl_out_11 br_out_11 bl_out_12 br_out_12 bl_out_13 br_out_13 bl_out_14 br_out_14 bl_out_15 br_out_15 bl_out_16 br_out_16 bl_out_17 br_out_17 bl_out_18 br_out_18 bl_out_19 br_out_19 bl_out_20 br_out_20 bl_out_21 br_out_21 bl_out_22 br_out_22 bl_out_23 br_out_23 bl_out_24 br_out_24 bl_out_25 br_out_25 bl_out_26 br_out_26 bl_out_27 br_out_27 bl_out_28 br_out_28 bl_out_29 br_out_29 bl_out_30 br_out_30 bl_out_31 br_out_31 gnd
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : sel_0 
* INOUT : sel_1 
* INOUT : bl_out_0 
* INOUT : br_out_0 
* INOUT : bl_out_1 
* INOUT : br_out_1 
* INOUT : bl_out_2 
* INOUT : br_out_2 
* INOUT : bl_out_3 
* INOUT : br_out_3 
* INOUT : bl_out_4 
* INOUT : br_out_4 
* INOUT : bl_out_5 
* INOUT : br_out_5 
* INOUT : bl_out_6 
* INOUT : br_out_6 
* INOUT : bl_out_7 
* INOUT : br_out_7 
* INOUT : bl_out_8 
* INOUT : br_out_8 
* INOUT : bl_out_9 
* INOUT : br_out_9 
* INOUT : bl_out_10 
* INOUT : br_out_10 
* INOUT : bl_out_11 
* INOUT : br_out_11 
* INOUT : bl_out_12 
* INOUT : br_out_12 
* INOUT : bl_out_13 
* INOUT : br_out_13 
* INOUT : bl_out_14 
* INOUT : br_out_14 
* INOUT : bl_out_15 
* INOUT : br_out_15 
* INOUT : bl_out_16 
* INOUT : br_out_16 
* INOUT : bl_out_17 
* INOUT : br_out_17 
* INOUT : bl_out_18 
* INOUT : br_out_18 
* INOUT : bl_out_19 
* INOUT : br_out_19 
* INOUT : bl_out_20 
* INOUT : br_out_20 
* INOUT : bl_out_21 
* INOUT : br_out_21 
* INOUT : bl_out_22 
* INOUT : br_out_22 
* INOUT : bl_out_23 
* INOUT : br_out_23 
* INOUT : bl_out_24 
* INOUT : br_out_24 
* INOUT : bl_out_25 
* INOUT : br_out_25 
* INOUT : bl_out_26 
* INOUT : br_out_26 
* INOUT : bl_out_27 
* INOUT : br_out_27 
* INOUT : bl_out_28 
* INOUT : br_out_28 
* INOUT : bl_out_29 
* INOUT : br_out_29 
* INOUT : bl_out_30 
* INOUT : br_out_30 
* INOUT : bl_out_31 
* INOUT : br_out_31 
* INOUT : gnd 
* cols: 64 word_size: 32 bl: bl1 br: br1
XXMUX0 bl_0 br_0 bl_out_0 br_out_0 sel_0 gnd single_level_column_mux_0
XXMUX1 bl_1 br_1 bl_out_0 br_out_0 sel_1 gnd single_level_column_mux_0
XXMUX2 bl_2 br_2 bl_out_1 br_out_1 sel_0 gnd single_level_column_mux_0
XXMUX3 bl_3 br_3 bl_out_1 br_out_1 sel_1 gnd single_level_column_mux_0
XXMUX4 bl_4 br_4 bl_out_2 br_out_2 sel_0 gnd single_level_column_mux_0
XXMUX5 bl_5 br_5 bl_out_2 br_out_2 sel_1 gnd single_level_column_mux_0
XXMUX6 bl_6 br_6 bl_out_3 br_out_3 sel_0 gnd single_level_column_mux_0
XXMUX7 bl_7 br_7 bl_out_3 br_out_3 sel_1 gnd single_level_column_mux_0
XXMUX8 bl_8 br_8 bl_out_4 br_out_4 sel_0 gnd single_level_column_mux_0
XXMUX9 bl_9 br_9 bl_out_4 br_out_4 sel_1 gnd single_level_column_mux_0
XXMUX10 bl_10 br_10 bl_out_5 br_out_5 sel_0 gnd single_level_column_mux_0
XXMUX11 bl_11 br_11 bl_out_5 br_out_5 sel_1 gnd single_level_column_mux_0
XXMUX12 bl_12 br_12 bl_out_6 br_out_6 sel_0 gnd single_level_column_mux_0
XXMUX13 bl_13 br_13 bl_out_6 br_out_6 sel_1 gnd single_level_column_mux_0
XXMUX14 bl_14 br_14 bl_out_7 br_out_7 sel_0 gnd single_level_column_mux_0
XXMUX15 bl_15 br_15 bl_out_7 br_out_7 sel_1 gnd single_level_column_mux_0
XXMUX16 bl_16 br_16 bl_out_8 br_out_8 sel_0 gnd single_level_column_mux_0
XXMUX17 bl_17 br_17 bl_out_8 br_out_8 sel_1 gnd single_level_column_mux_0
XXMUX18 bl_18 br_18 bl_out_9 br_out_9 sel_0 gnd single_level_column_mux_0
XXMUX19 bl_19 br_19 bl_out_9 br_out_9 sel_1 gnd single_level_column_mux_0
XXMUX20 bl_20 br_20 bl_out_10 br_out_10 sel_0 gnd single_level_column_mux_0
XXMUX21 bl_21 br_21 bl_out_10 br_out_10 sel_1 gnd single_level_column_mux_0
XXMUX22 bl_22 br_22 bl_out_11 br_out_11 sel_0 gnd single_level_column_mux_0
XXMUX23 bl_23 br_23 bl_out_11 br_out_11 sel_1 gnd single_level_column_mux_0
XXMUX24 bl_24 br_24 bl_out_12 br_out_12 sel_0 gnd single_level_column_mux_0
XXMUX25 bl_25 br_25 bl_out_12 br_out_12 sel_1 gnd single_level_column_mux_0
XXMUX26 bl_26 br_26 bl_out_13 br_out_13 sel_0 gnd single_level_column_mux_0
XXMUX27 bl_27 br_27 bl_out_13 br_out_13 sel_1 gnd single_level_column_mux_0
XXMUX28 bl_28 br_28 bl_out_14 br_out_14 sel_0 gnd single_level_column_mux_0
XXMUX29 bl_29 br_29 bl_out_14 br_out_14 sel_1 gnd single_level_column_mux_0
XXMUX30 bl_30 br_30 bl_out_15 br_out_15 sel_0 gnd single_level_column_mux_0
XXMUX31 bl_31 br_31 bl_out_15 br_out_15 sel_1 gnd single_level_column_mux_0
XXMUX32 bl_32 br_32 bl_out_16 br_out_16 sel_0 gnd single_level_column_mux_0
XXMUX33 bl_33 br_33 bl_out_16 br_out_16 sel_1 gnd single_level_column_mux_0
XXMUX34 bl_34 br_34 bl_out_17 br_out_17 sel_0 gnd single_level_column_mux_0
XXMUX35 bl_35 br_35 bl_out_17 br_out_17 sel_1 gnd single_level_column_mux_0
XXMUX36 bl_36 br_36 bl_out_18 br_out_18 sel_0 gnd single_level_column_mux_0
XXMUX37 bl_37 br_37 bl_out_18 br_out_18 sel_1 gnd single_level_column_mux_0
XXMUX38 bl_38 br_38 bl_out_19 br_out_19 sel_0 gnd single_level_column_mux_0
XXMUX39 bl_39 br_39 bl_out_19 br_out_19 sel_1 gnd single_level_column_mux_0
XXMUX40 bl_40 br_40 bl_out_20 br_out_20 sel_0 gnd single_level_column_mux_0
XXMUX41 bl_41 br_41 bl_out_20 br_out_20 sel_1 gnd single_level_column_mux_0
XXMUX42 bl_42 br_42 bl_out_21 br_out_21 sel_0 gnd single_level_column_mux_0
XXMUX43 bl_43 br_43 bl_out_21 br_out_21 sel_1 gnd single_level_column_mux_0
XXMUX44 bl_44 br_44 bl_out_22 br_out_22 sel_0 gnd single_level_column_mux_0
XXMUX45 bl_45 br_45 bl_out_22 br_out_22 sel_1 gnd single_level_column_mux_0
XXMUX46 bl_46 br_46 bl_out_23 br_out_23 sel_0 gnd single_level_column_mux_0
XXMUX47 bl_47 br_47 bl_out_23 br_out_23 sel_1 gnd single_level_column_mux_0
XXMUX48 bl_48 br_48 bl_out_24 br_out_24 sel_0 gnd single_level_column_mux_0
XXMUX49 bl_49 br_49 bl_out_24 br_out_24 sel_1 gnd single_level_column_mux_0
XXMUX50 bl_50 br_50 bl_out_25 br_out_25 sel_0 gnd single_level_column_mux_0
XXMUX51 bl_51 br_51 bl_out_25 br_out_25 sel_1 gnd single_level_column_mux_0
XXMUX52 bl_52 br_52 bl_out_26 br_out_26 sel_0 gnd single_level_column_mux_0
XXMUX53 bl_53 br_53 bl_out_26 br_out_26 sel_1 gnd single_level_column_mux_0
XXMUX54 bl_54 br_54 bl_out_27 br_out_27 sel_0 gnd single_level_column_mux_0
XXMUX55 bl_55 br_55 bl_out_27 br_out_27 sel_1 gnd single_level_column_mux_0
XXMUX56 bl_56 br_56 bl_out_28 br_out_28 sel_0 gnd single_level_column_mux_0
XXMUX57 bl_57 br_57 bl_out_28 br_out_28 sel_1 gnd single_level_column_mux_0
XXMUX58 bl_58 br_58 bl_out_29 br_out_29 sel_0 gnd single_level_column_mux_0
XXMUX59 bl_59 br_59 bl_out_29 br_out_29 sel_1 gnd single_level_column_mux_0
XXMUX60 bl_60 br_60 bl_out_30 br_out_30 sel_0 gnd single_level_column_mux_0
XXMUX61 bl_61 br_61 bl_out_30 br_out_30 sel_1 gnd single_level_column_mux_0
XXMUX62 bl_62 br_62 bl_out_31 br_out_31 sel_0 gnd single_level_column_mux_0
XXMUX63 bl_63 br_63 bl_out_31 br_out_31 sel_1 gnd single_level_column_mux_0
.ENDS single_level_column_mux_array_0

.SUBCKT port_data_0 rbl_bl rbl_br bl1_0 br1_0 bl1_1 br1_1 bl1_2 br1_2 bl1_3 br1_3 bl1_4 br1_4 bl1_5 br1_5 bl1_6 br1_6 bl1_7 br1_7 bl1_8 br1_8 bl1_9 br1_9 bl1_10 br1_10 bl1_11 br1_11 bl1_12 br1_12 bl1_13 br1_13 bl1_14 br1_14 bl1_15 br1_15 bl1_16 br1_16 bl1_17 br1_17 bl1_18 br1_18 bl1_19 br1_19 bl1_20 br1_20 bl1_21 br1_21 bl1_22 br1_22 bl1_23 br1_23 bl1_24 br1_24 bl1_25 br1_25 bl1_26 br1_26 bl1_27 br1_27 bl1_28 br1_28 bl1_29 br1_29 bl1_30 br1_30 bl1_31 br1_31 bl1_32 br1_32 bl1_33 br1_33 bl1_34 br1_34 bl1_35 br1_35 bl1_36 br1_36 bl1_37 br1_37 bl1_38 br1_38 bl1_39 br1_39 bl1_40 br1_40 bl1_41 br1_41 bl1_42 br1_42 bl1_43 br1_43 bl1_44 br1_44 bl1_45 br1_45 bl1_46 br1_46 bl1_47 br1_47 bl1_48 br1_48 bl1_49 br1_49 bl1_50 br1_50 bl1_51 br1_51 bl1_52 br1_52 bl1_53 br1_53 bl1_54 br1_54 bl1_55 br1_55 bl1_56 br1_56 bl1_57 br1_57 bl1_58 br1_58 bl1_59 br1_59 bl1_60 br1_60 bl1_61 br1_61 bl1_62 br1_62 bl1_63 br1_63 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5 dout_6 dout_7 dout_8 dout_9 dout_10 dout_11 dout_12 dout_13 dout_14 dout_15 dout_16 dout_17 dout_18 dout_19 dout_20 dout_21 dout_22 dout_23 dout_24 dout_25 dout_26 dout_27 dout_28 dout_29 dout_30 dout_31 sel_0 sel_1 s_en p_en_bar vdd gnd
* INOUT : rbl_bl 
* INOUT : rbl_br 
* INOUT : bl1_0 
* INOUT : br1_0 
* INOUT : bl1_1 
* INOUT : br1_1 
* INOUT : bl1_2 
* INOUT : br1_2 
* INOUT : bl1_3 
* INOUT : br1_3 
* INOUT : bl1_4 
* INOUT : br1_4 
* INOUT : bl1_5 
* INOUT : br1_5 
* INOUT : bl1_6 
* INOUT : br1_6 
* INOUT : bl1_7 
* INOUT : br1_7 
* INOUT : bl1_8 
* INOUT : br1_8 
* INOUT : bl1_9 
* INOUT : br1_9 
* INOUT : bl1_10 
* INOUT : br1_10 
* INOUT : bl1_11 
* INOUT : br1_11 
* INOUT : bl1_12 
* INOUT : br1_12 
* INOUT : bl1_13 
* INOUT : br1_13 
* INOUT : bl1_14 
* INOUT : br1_14 
* INOUT : bl1_15 
* INOUT : br1_15 
* INOUT : bl1_16 
* INOUT : br1_16 
* INOUT : bl1_17 
* INOUT : br1_17 
* INOUT : bl1_18 
* INOUT : br1_18 
* INOUT : bl1_19 
* INOUT : br1_19 
* INOUT : bl1_20 
* INOUT : br1_20 
* INOUT : bl1_21 
* INOUT : br1_21 
* INOUT : bl1_22 
* INOUT : br1_22 
* INOUT : bl1_23 
* INOUT : br1_23 
* INOUT : bl1_24 
* INOUT : br1_24 
* INOUT : bl1_25 
* INOUT : br1_25 
* INOUT : bl1_26 
* INOUT : br1_26 
* INOUT : bl1_27 
* INOUT : br1_27 
* INOUT : bl1_28 
* INOUT : br1_28 
* INOUT : bl1_29 
* INOUT : br1_29 
* INOUT : bl1_30 
* INOUT : br1_30 
* INOUT : bl1_31 
* INOUT : br1_31 
* INOUT : bl1_32 
* INOUT : br1_32 
* INOUT : bl1_33 
* INOUT : br1_33 
* INOUT : bl1_34 
* INOUT : br1_34 
* INOUT : bl1_35 
* INOUT : br1_35 
* INOUT : bl1_36 
* INOUT : br1_36 
* INOUT : bl1_37 
* INOUT : br1_37 
* INOUT : bl1_38 
* INOUT : br1_38 
* INOUT : bl1_39 
* INOUT : br1_39 
* INOUT : bl1_40 
* INOUT : br1_40 
* INOUT : bl1_41 
* INOUT : br1_41 
* INOUT : bl1_42 
* INOUT : br1_42 
* INOUT : bl1_43 
* INOUT : br1_43 
* INOUT : bl1_44 
* INOUT : br1_44 
* INOUT : bl1_45 
* INOUT : br1_45 
* INOUT : bl1_46 
* INOUT : br1_46 
* INOUT : bl1_47 
* INOUT : br1_47 
* INOUT : bl1_48 
* INOUT : br1_48 
* INOUT : bl1_49 
* INOUT : br1_49 
* INOUT : bl1_50 
* INOUT : br1_50 
* INOUT : bl1_51 
* INOUT : br1_51 
* INOUT : bl1_52 
* INOUT : br1_52 
* INOUT : bl1_53 
* INOUT : br1_53 
* INOUT : bl1_54 
* INOUT : br1_54 
* INOUT : bl1_55 
* INOUT : br1_55 
* INOUT : bl1_56 
* INOUT : br1_56 
* INOUT : bl1_57 
* INOUT : br1_57 
* INOUT : bl1_58 
* INOUT : br1_58 
* INOUT : bl1_59 
* INOUT : br1_59 
* INOUT : bl1_60 
* INOUT : br1_60 
* INOUT : bl1_61 
* INOUT : br1_61 
* INOUT : bl1_62 
* INOUT : br1_62 
* INOUT : bl1_63 
* INOUT : br1_63 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* OUTPUT: dout_7 
* OUTPUT: dout_8 
* OUTPUT: dout_9 
* OUTPUT: dout_10 
* OUTPUT: dout_11 
* OUTPUT: dout_12 
* OUTPUT: dout_13 
* OUTPUT: dout_14 
* OUTPUT: dout_15 
* OUTPUT: dout_16 
* OUTPUT: dout_17 
* OUTPUT: dout_18 
* OUTPUT: dout_19 
* OUTPUT: dout_20 
* OUTPUT: dout_21 
* OUTPUT: dout_22 
* OUTPUT: dout_23 
* OUTPUT: dout_24 
* OUTPUT: dout_25 
* OUTPUT: dout_26 
* OUTPUT: dout_27 
* OUTPUT: dout_28 
* OUTPUT: dout_29 
* OUTPUT: dout_30 
* OUTPUT: dout_31 
* INPUT : sel_0 
* INPUT : sel_1 
* INPUT : s_en 
* INPUT : p_en_bar 
* POWER : vdd 
* GROUND: gnd 
Xprecharge_array1 bl1_0 br1_0 bl1_1 br1_1 bl1_2 br1_2 bl1_3 br1_3 bl1_4 br1_4 bl1_5 br1_5 bl1_6 br1_6 bl1_7 br1_7 bl1_8 br1_8 bl1_9 br1_9 bl1_10 br1_10 bl1_11 br1_11 bl1_12 br1_12 bl1_13 br1_13 bl1_14 br1_14 bl1_15 br1_15 bl1_16 br1_16 bl1_17 br1_17 bl1_18 br1_18 bl1_19 br1_19 bl1_20 br1_20 bl1_21 br1_21 bl1_22 br1_22 bl1_23 br1_23 bl1_24 br1_24 bl1_25 br1_25 bl1_26 br1_26 bl1_27 br1_27 bl1_28 br1_28 bl1_29 br1_29 bl1_30 br1_30 bl1_31 br1_31 bl1_32 br1_32 bl1_33 br1_33 bl1_34 br1_34 bl1_35 br1_35 bl1_36 br1_36 bl1_37 br1_37 bl1_38 br1_38 bl1_39 br1_39 bl1_40 br1_40 bl1_41 br1_41 bl1_42 br1_42 bl1_43 br1_43 bl1_44 br1_44 bl1_45 br1_45 bl1_46 br1_46 bl1_47 br1_47 bl1_48 br1_48 bl1_49 br1_49 bl1_50 br1_50 bl1_51 br1_51 bl1_52 br1_52 bl1_53 br1_53 bl1_54 br1_54 bl1_55 br1_55 bl1_56 br1_56 bl1_57 br1_57 bl1_58 br1_58 bl1_59 br1_59 bl1_60 br1_60 bl1_61 br1_61 bl1_62 br1_62 bl1_63 br1_63 rbl_bl rbl_br p_en_bar vdd precharge_array_0
Xsense_amp_array1 dout_0 bl1_out_0 br1_out_0 dout_1 bl1_out_1 br1_out_1 dout_2 bl1_out_2 br1_out_2 dout_3 bl1_out_3 br1_out_3 dout_4 bl1_out_4 br1_out_4 dout_5 bl1_out_5 br1_out_5 dout_6 bl1_out_6 br1_out_6 dout_7 bl1_out_7 br1_out_7 dout_8 bl1_out_8 br1_out_8 dout_9 bl1_out_9 br1_out_9 dout_10 bl1_out_10 br1_out_10 dout_11 bl1_out_11 br1_out_11 dout_12 bl1_out_12 br1_out_12 dout_13 bl1_out_13 br1_out_13 dout_14 bl1_out_14 br1_out_14 dout_15 bl1_out_15 br1_out_15 dout_16 bl1_out_16 br1_out_16 dout_17 bl1_out_17 br1_out_17 dout_18 bl1_out_18 br1_out_18 dout_19 bl1_out_19 br1_out_19 dout_20 bl1_out_20 br1_out_20 dout_21 bl1_out_21 br1_out_21 dout_22 bl1_out_22 br1_out_22 dout_23 bl1_out_23 br1_out_23 dout_24 bl1_out_24 br1_out_24 dout_25 bl1_out_25 br1_out_25 dout_26 bl1_out_26 br1_out_26 dout_27 bl1_out_27 br1_out_27 dout_28 bl1_out_28 br1_out_28 dout_29 bl1_out_29 br1_out_29 dout_30 bl1_out_30 br1_out_30 dout_31 bl1_out_31 br1_out_31 s_en vdd gnd sense_amp_array
Xcolumn_mux_array1 bl1_0 br1_0 bl1_1 br1_1 bl1_2 br1_2 bl1_3 br1_3 bl1_4 br1_4 bl1_5 br1_5 bl1_6 br1_6 bl1_7 br1_7 bl1_8 br1_8 bl1_9 br1_9 bl1_10 br1_10 bl1_11 br1_11 bl1_12 br1_12 bl1_13 br1_13 bl1_14 br1_14 bl1_15 br1_15 bl1_16 br1_16 bl1_17 br1_17 bl1_18 br1_18 bl1_19 br1_19 bl1_20 br1_20 bl1_21 br1_21 bl1_22 br1_22 bl1_23 br1_23 bl1_24 br1_24 bl1_25 br1_25 bl1_26 br1_26 bl1_27 br1_27 bl1_28 br1_28 bl1_29 br1_29 bl1_30 br1_30 bl1_31 br1_31 bl1_32 br1_32 bl1_33 br1_33 bl1_34 br1_34 bl1_35 br1_35 bl1_36 br1_36 bl1_37 br1_37 bl1_38 br1_38 bl1_39 br1_39 bl1_40 br1_40 bl1_41 br1_41 bl1_42 br1_42 bl1_43 br1_43 bl1_44 br1_44 bl1_45 br1_45 bl1_46 br1_46 bl1_47 br1_47 bl1_48 br1_48 bl1_49 br1_49 bl1_50 br1_50 bl1_51 br1_51 bl1_52 br1_52 bl1_53 br1_53 bl1_54 br1_54 bl1_55 br1_55 bl1_56 br1_56 bl1_57 br1_57 bl1_58 br1_58 bl1_59 br1_59 bl1_60 br1_60 bl1_61 br1_61 bl1_62 br1_62 bl1_63 br1_63 sel_0 sel_1 bl1_out_0 br1_out_0 bl1_out_1 br1_out_1 bl1_out_2 br1_out_2 bl1_out_3 br1_out_3 bl1_out_4 br1_out_4 bl1_out_5 br1_out_5 bl1_out_6 br1_out_6 bl1_out_7 br1_out_7 bl1_out_8 br1_out_8 bl1_out_9 br1_out_9 bl1_out_10 br1_out_10 bl1_out_11 br1_out_11 bl1_out_12 br1_out_12 bl1_out_13 br1_out_13 bl1_out_14 br1_out_14 bl1_out_15 br1_out_15 bl1_out_16 br1_out_16 bl1_out_17 br1_out_17 bl1_out_18 br1_out_18 bl1_out_19 br1_out_19 bl1_out_20 br1_out_20 bl1_out_21 br1_out_21 bl1_out_22 br1_out_22 bl1_out_23 br1_out_23 bl1_out_24 br1_out_24 bl1_out_25 br1_out_25 bl1_out_26 br1_out_26 bl1_out_27 br1_out_27 bl1_out_28 br1_out_28 bl1_out_29 br1_out_29 bl1_out_30 br1_out_30 bl1_out_31 br1_out_31 gnd single_level_column_mux_array_0
.ENDS port_data_0
* NGSPICE file created from nand2_dec.ext - technology: EFS8A


* Top level circuit nand2_dec
.subckt nand2_dec A B Z vdd gnd

XM1001 Z B vdd vdd sky130_fd_pr__pfet_01v8 W=1.12 L=0.15 m=1
XM1002 vdd A Z vdd sky130_fd_pr__pfet_01v8 W=1.12 L=0.15 m=1
XM1000 Z A a_n722_276# gnd sky130_fd_pr__nfet_01v8 W=0.74 L=0.15 m=1
XM1003 a_n722_276# B gnd gnd sky130_fd_pr__nfet_01v8 W=0.74 L=0.15 m=1
.ends


* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u

* ptx M{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u

.SUBCKT pinv_dec A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u
.ENDS pinv_dec

.SUBCKT and2_dec A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpand2_dec_nand A B zb_int vdd gnd nand2_dec
Xpand2_dec_inv zb_int Z vdd gnd pinv_dec
.ENDS and2_dec
* NGSPICE file created from nand3_dec.ext - technology: EFS8A


* Top level circuit nand3_dec
.subckt nand3_dec A B C Z vdd gnd

XM1001 Z A a_n346_328# gnd sky130_fd_pr__nfet_01v8 W=0.74 L=0.15 m=1
XM1002 a_n346_256# C gnd gnd sky130_fd_pr__nfet_01v8 W=0.74 L=0.15 m=1
XM1003 a_n346_328# B a_n346_256# gnd sky130_fd_pr__nfet_01v8 W=0.74 L=0.15 m=1
XM1000 Z B vdd vdd sky130_fd_pr__pfet_01v8 W=1.12 L=0.15 m=1
XM1004 Z A vdd vdd sky130_fd_pr__pfet_01v8 W=1.12 L=0.15 m=1
XM1005 Z C vdd vdd sky130_fd_pr__pfet_01v8 W=1.12 L=0.15 m=1
.ends


.SUBCKT and3_dec A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpand3_dec_nand A B C zb_int vdd gnd nand3_dec
Xpand3_dec_inv zb_int Z vdd gnd pinv_dec
.ENDS and3_dec

.SUBCKT hierarchical_predecode2x4 in_0 in_1 out_0 out_1 out_2 out_3 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0 in_0 inbar_0 vdd gnd pinv_dec
Xpre_inv_1 in_1 inbar_1 vdd gnd pinv_dec
XXpre2x4_and_0 inbar_0 inbar_1 out_0 vdd gnd and2_dec
XXpre2x4_and_1 in_0 inbar_1 out_1 vdd gnd and2_dec
XXpre2x4_and_2 inbar_0 in_1 out_2 vdd gnd and2_dec
XXpre2x4_and_3 in_0 in_1 out_3 vdd gnd and2_dec
.ENDS hierarchical_predecode2x4

.SUBCKT hierarchical_predecode3x8 in_0 in_1 in_2 out_0 out_1 out_2 out_3 out_4 out_5 out_6 out_7 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* OUTPUT: out_4 
* OUTPUT: out_5 
* OUTPUT: out_6 
* OUTPUT: out_7 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0 in_0 inbar_0 vdd gnd pinv_dec
Xpre_inv_1 in_1 inbar_1 vdd gnd pinv_dec
Xpre_inv_2 in_2 inbar_2 vdd gnd pinv_dec
XXpre3x8_and_0 inbar_0 inbar_1 inbar_2 out_0 vdd gnd and3_dec
XXpre3x8_and_1 in_0 inbar_1 inbar_2 out_1 vdd gnd and3_dec
XXpre3x8_and_2 inbar_0 in_1 inbar_2 out_2 vdd gnd and3_dec
XXpre3x8_and_3 in_0 in_1 inbar_2 out_3 vdd gnd and3_dec
XXpre3x8_and_4 inbar_0 inbar_1 in_2 out_4 vdd gnd and3_dec
XXpre3x8_and_5 in_0 inbar_1 in_2 out_5 vdd gnd and3_dec
XXpre3x8_and_6 inbar_0 in_1 in_2 out_6 vdd gnd and3_dec
XXpre3x8_and_7 in_0 in_1 in_2 out_7 vdd gnd and3_dec
.ENDS hierarchical_predecode3x8

.SUBCKT hierarchical_decoder addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 addr_6 decode_0 decode_1 decode_2 decode_3 decode_4 decode_5 decode_6 decode_7 decode_8 decode_9 decode_10 decode_11 decode_12 decode_13 decode_14 decode_15 decode_16 decode_17 decode_18 decode_19 decode_20 decode_21 decode_22 decode_23 decode_24 decode_25 decode_26 decode_27 decode_28 decode_29 decode_30 decode_31 decode_32 decode_33 decode_34 decode_35 decode_36 decode_37 decode_38 decode_39 decode_40 decode_41 decode_42 decode_43 decode_44 decode_45 decode_46 decode_47 decode_48 decode_49 decode_50 decode_51 decode_52 decode_53 decode_54 decode_55 decode_56 decode_57 decode_58 decode_59 decode_60 decode_61 decode_62 decode_63 decode_64 decode_65 decode_66 decode_67 decode_68 decode_69 decode_70 decode_71 decode_72 decode_73 decode_74 decode_75 decode_76 decode_77 decode_78 decode_79 decode_80 decode_81 decode_82 decode_83 decode_84 decode_85 decode_86 decode_87 decode_88 decode_89 decode_90 decode_91 decode_92 decode_93 decode_94 decode_95 decode_96 decode_97 decode_98 decode_99 decode_100 decode_101 decode_102 decode_103 decode_104 decode_105 decode_106 decode_107 decode_108 decode_109 decode_110 decode_111 decode_112 decode_113 decode_114 decode_115 decode_116 decode_117 decode_118 decode_119 decode_120 decode_121 decode_122 decode_123 decode_124 decode_125 decode_126 decode_127 vdd gnd
* INPUT : addr_0 
* INPUT : addr_1 
* INPUT : addr_2 
* INPUT : addr_3 
* INPUT : addr_4 
* INPUT : addr_5 
* INPUT : addr_6 
* OUTPUT: decode_0 
* OUTPUT: decode_1 
* OUTPUT: decode_2 
* OUTPUT: decode_3 
* OUTPUT: decode_4 
* OUTPUT: decode_5 
* OUTPUT: decode_6 
* OUTPUT: decode_7 
* OUTPUT: decode_8 
* OUTPUT: decode_9 
* OUTPUT: decode_10 
* OUTPUT: decode_11 
* OUTPUT: decode_12 
* OUTPUT: decode_13 
* OUTPUT: decode_14 
* OUTPUT: decode_15 
* OUTPUT: decode_16 
* OUTPUT: decode_17 
* OUTPUT: decode_18 
* OUTPUT: decode_19 
* OUTPUT: decode_20 
* OUTPUT: decode_21 
* OUTPUT: decode_22 
* OUTPUT: decode_23 
* OUTPUT: decode_24 
* OUTPUT: decode_25 
* OUTPUT: decode_26 
* OUTPUT: decode_27 
* OUTPUT: decode_28 
* OUTPUT: decode_29 
* OUTPUT: decode_30 
* OUTPUT: decode_31 
* OUTPUT: decode_32 
* OUTPUT: decode_33 
* OUTPUT: decode_34 
* OUTPUT: decode_35 
* OUTPUT: decode_36 
* OUTPUT: decode_37 
* OUTPUT: decode_38 
* OUTPUT: decode_39 
* OUTPUT: decode_40 
* OUTPUT: decode_41 
* OUTPUT: decode_42 
* OUTPUT: decode_43 
* OUTPUT: decode_44 
* OUTPUT: decode_45 
* OUTPUT: decode_46 
* OUTPUT: decode_47 
* OUTPUT: decode_48 
* OUTPUT: decode_49 
* OUTPUT: decode_50 
* OUTPUT: decode_51 
* OUTPUT: decode_52 
* OUTPUT: decode_53 
* OUTPUT: decode_54 
* OUTPUT: decode_55 
* OUTPUT: decode_56 
* OUTPUT: decode_57 
* OUTPUT: decode_58 
* OUTPUT: decode_59 
* OUTPUT: decode_60 
* OUTPUT: decode_61 
* OUTPUT: decode_62 
* OUTPUT: decode_63 
* OUTPUT: decode_64 
* OUTPUT: decode_65 
* OUTPUT: decode_66 
* OUTPUT: decode_67 
* OUTPUT: decode_68 
* OUTPUT: decode_69 
* OUTPUT: decode_70 
* OUTPUT: decode_71 
* OUTPUT: decode_72 
* OUTPUT: decode_73 
* OUTPUT: decode_74 
* OUTPUT: decode_75 
* OUTPUT: decode_76 
* OUTPUT: decode_77 
* OUTPUT: decode_78 
* OUTPUT: decode_79 
* OUTPUT: decode_80 
* OUTPUT: decode_81 
* OUTPUT: decode_82 
* OUTPUT: decode_83 
* OUTPUT: decode_84 
* OUTPUT: decode_85 
* OUTPUT: decode_86 
* OUTPUT: decode_87 
* OUTPUT: decode_88 
* OUTPUT: decode_89 
* OUTPUT: decode_90 
* OUTPUT: decode_91 
* OUTPUT: decode_92 
* OUTPUT: decode_93 
* OUTPUT: decode_94 
* OUTPUT: decode_95 
* OUTPUT: decode_96 
* OUTPUT: decode_97 
* OUTPUT: decode_98 
* OUTPUT: decode_99 
* OUTPUT: decode_100 
* OUTPUT: decode_101 
* OUTPUT: decode_102 
* OUTPUT: decode_103 
* OUTPUT: decode_104 
* OUTPUT: decode_105 
* OUTPUT: decode_106 
* OUTPUT: decode_107 
* OUTPUT: decode_108 
* OUTPUT: decode_109 
* OUTPUT: decode_110 
* OUTPUT: decode_111 
* OUTPUT: decode_112 
* OUTPUT: decode_113 
* OUTPUT: decode_114 
* OUTPUT: decode_115 
* OUTPUT: decode_116 
* OUTPUT: decode_117 
* OUTPUT: decode_118 
* OUTPUT: decode_119 
* OUTPUT: decode_120 
* OUTPUT: decode_121 
* OUTPUT: decode_122 
* OUTPUT: decode_123 
* OUTPUT: decode_124 
* OUTPUT: decode_125 
* OUTPUT: decode_126 
* OUTPUT: decode_127 
* POWER : vdd 
* GROUND: gnd 
Xpre_0 addr_0 addr_1 out_0 out_1 out_2 out_3 vdd gnd hierarchical_predecode2x4
Xpre_1 addr_2 addr_3 out_4 out_5 out_6 out_7 vdd gnd hierarchical_predecode2x4
Xpre3x8_0 addr_4 addr_5 addr_6 out_8 out_9 out_10 out_11 out_12 out_13 out_14 out_15 vdd gnd hierarchical_predecode3x8
XDEC_AND_0 out_0 out_4 out_8 decode_0 vdd gnd and3_dec
XDEC_AND_16 out_0 out_4 out_9 decode_16 vdd gnd and3_dec
XDEC_AND_32 out_0 out_4 out_10 decode_32 vdd gnd and3_dec
XDEC_AND_48 out_0 out_4 out_11 decode_48 vdd gnd and3_dec
XDEC_AND_64 out_0 out_4 out_12 decode_64 vdd gnd and3_dec
XDEC_AND_80 out_0 out_4 out_13 decode_80 vdd gnd and3_dec
XDEC_AND_96 out_0 out_4 out_14 decode_96 vdd gnd and3_dec
XDEC_AND_112 out_0 out_4 out_15 decode_112 vdd gnd and3_dec
XDEC_AND_4 out_0 out_5 out_8 decode_4 vdd gnd and3_dec
XDEC_AND_20 out_0 out_5 out_9 decode_20 vdd gnd and3_dec
XDEC_AND_36 out_0 out_5 out_10 decode_36 vdd gnd and3_dec
XDEC_AND_52 out_0 out_5 out_11 decode_52 vdd gnd and3_dec
XDEC_AND_68 out_0 out_5 out_12 decode_68 vdd gnd and3_dec
XDEC_AND_84 out_0 out_5 out_13 decode_84 vdd gnd and3_dec
XDEC_AND_100 out_0 out_5 out_14 decode_100 vdd gnd and3_dec
XDEC_AND_116 out_0 out_5 out_15 decode_116 vdd gnd and3_dec
XDEC_AND_8 out_0 out_6 out_8 decode_8 vdd gnd and3_dec
XDEC_AND_24 out_0 out_6 out_9 decode_24 vdd gnd and3_dec
XDEC_AND_40 out_0 out_6 out_10 decode_40 vdd gnd and3_dec
XDEC_AND_56 out_0 out_6 out_11 decode_56 vdd gnd and3_dec
XDEC_AND_72 out_0 out_6 out_12 decode_72 vdd gnd and3_dec
XDEC_AND_88 out_0 out_6 out_13 decode_88 vdd gnd and3_dec
XDEC_AND_104 out_0 out_6 out_14 decode_104 vdd gnd and3_dec
XDEC_AND_120 out_0 out_6 out_15 decode_120 vdd gnd and3_dec
XDEC_AND_12 out_0 out_7 out_8 decode_12 vdd gnd and3_dec
XDEC_AND_28 out_0 out_7 out_9 decode_28 vdd gnd and3_dec
XDEC_AND_44 out_0 out_7 out_10 decode_44 vdd gnd and3_dec
XDEC_AND_60 out_0 out_7 out_11 decode_60 vdd gnd and3_dec
XDEC_AND_76 out_0 out_7 out_12 decode_76 vdd gnd and3_dec
XDEC_AND_92 out_0 out_7 out_13 decode_92 vdd gnd and3_dec
XDEC_AND_108 out_0 out_7 out_14 decode_108 vdd gnd and3_dec
XDEC_AND_124 out_0 out_7 out_15 decode_124 vdd gnd and3_dec
XDEC_AND_1 out_1 out_4 out_8 decode_1 vdd gnd and3_dec
XDEC_AND_17 out_1 out_4 out_9 decode_17 vdd gnd and3_dec
XDEC_AND_33 out_1 out_4 out_10 decode_33 vdd gnd and3_dec
XDEC_AND_49 out_1 out_4 out_11 decode_49 vdd gnd and3_dec
XDEC_AND_65 out_1 out_4 out_12 decode_65 vdd gnd and3_dec
XDEC_AND_81 out_1 out_4 out_13 decode_81 vdd gnd and3_dec
XDEC_AND_97 out_1 out_4 out_14 decode_97 vdd gnd and3_dec
XDEC_AND_113 out_1 out_4 out_15 decode_113 vdd gnd and3_dec
XDEC_AND_5 out_1 out_5 out_8 decode_5 vdd gnd and3_dec
XDEC_AND_21 out_1 out_5 out_9 decode_21 vdd gnd and3_dec
XDEC_AND_37 out_1 out_5 out_10 decode_37 vdd gnd and3_dec
XDEC_AND_53 out_1 out_5 out_11 decode_53 vdd gnd and3_dec
XDEC_AND_69 out_1 out_5 out_12 decode_69 vdd gnd and3_dec
XDEC_AND_85 out_1 out_5 out_13 decode_85 vdd gnd and3_dec
XDEC_AND_101 out_1 out_5 out_14 decode_101 vdd gnd and3_dec
XDEC_AND_117 out_1 out_5 out_15 decode_117 vdd gnd and3_dec
XDEC_AND_9 out_1 out_6 out_8 decode_9 vdd gnd and3_dec
XDEC_AND_25 out_1 out_6 out_9 decode_25 vdd gnd and3_dec
XDEC_AND_41 out_1 out_6 out_10 decode_41 vdd gnd and3_dec
XDEC_AND_57 out_1 out_6 out_11 decode_57 vdd gnd and3_dec
XDEC_AND_73 out_1 out_6 out_12 decode_73 vdd gnd and3_dec
XDEC_AND_89 out_1 out_6 out_13 decode_89 vdd gnd and3_dec
XDEC_AND_105 out_1 out_6 out_14 decode_105 vdd gnd and3_dec
XDEC_AND_121 out_1 out_6 out_15 decode_121 vdd gnd and3_dec
XDEC_AND_13 out_1 out_7 out_8 decode_13 vdd gnd and3_dec
XDEC_AND_29 out_1 out_7 out_9 decode_29 vdd gnd and3_dec
XDEC_AND_45 out_1 out_7 out_10 decode_45 vdd gnd and3_dec
XDEC_AND_61 out_1 out_7 out_11 decode_61 vdd gnd and3_dec
XDEC_AND_77 out_1 out_7 out_12 decode_77 vdd gnd and3_dec
XDEC_AND_93 out_1 out_7 out_13 decode_93 vdd gnd and3_dec
XDEC_AND_109 out_1 out_7 out_14 decode_109 vdd gnd and3_dec
XDEC_AND_125 out_1 out_7 out_15 decode_125 vdd gnd and3_dec
XDEC_AND_2 out_2 out_4 out_8 decode_2 vdd gnd and3_dec
XDEC_AND_18 out_2 out_4 out_9 decode_18 vdd gnd and3_dec
XDEC_AND_34 out_2 out_4 out_10 decode_34 vdd gnd and3_dec
XDEC_AND_50 out_2 out_4 out_11 decode_50 vdd gnd and3_dec
XDEC_AND_66 out_2 out_4 out_12 decode_66 vdd gnd and3_dec
XDEC_AND_82 out_2 out_4 out_13 decode_82 vdd gnd and3_dec
XDEC_AND_98 out_2 out_4 out_14 decode_98 vdd gnd and3_dec
XDEC_AND_114 out_2 out_4 out_15 decode_114 vdd gnd and3_dec
XDEC_AND_6 out_2 out_5 out_8 decode_6 vdd gnd and3_dec
XDEC_AND_22 out_2 out_5 out_9 decode_22 vdd gnd and3_dec
XDEC_AND_38 out_2 out_5 out_10 decode_38 vdd gnd and3_dec
XDEC_AND_54 out_2 out_5 out_11 decode_54 vdd gnd and3_dec
XDEC_AND_70 out_2 out_5 out_12 decode_70 vdd gnd and3_dec
XDEC_AND_86 out_2 out_5 out_13 decode_86 vdd gnd and3_dec
XDEC_AND_102 out_2 out_5 out_14 decode_102 vdd gnd and3_dec
XDEC_AND_118 out_2 out_5 out_15 decode_118 vdd gnd and3_dec
XDEC_AND_10 out_2 out_6 out_8 decode_10 vdd gnd and3_dec
XDEC_AND_26 out_2 out_6 out_9 decode_26 vdd gnd and3_dec
XDEC_AND_42 out_2 out_6 out_10 decode_42 vdd gnd and3_dec
XDEC_AND_58 out_2 out_6 out_11 decode_58 vdd gnd and3_dec
XDEC_AND_74 out_2 out_6 out_12 decode_74 vdd gnd and3_dec
XDEC_AND_90 out_2 out_6 out_13 decode_90 vdd gnd and3_dec
XDEC_AND_106 out_2 out_6 out_14 decode_106 vdd gnd and3_dec
XDEC_AND_122 out_2 out_6 out_15 decode_122 vdd gnd and3_dec
XDEC_AND_14 out_2 out_7 out_8 decode_14 vdd gnd and3_dec
XDEC_AND_30 out_2 out_7 out_9 decode_30 vdd gnd and3_dec
XDEC_AND_46 out_2 out_7 out_10 decode_46 vdd gnd and3_dec
XDEC_AND_62 out_2 out_7 out_11 decode_62 vdd gnd and3_dec
XDEC_AND_78 out_2 out_7 out_12 decode_78 vdd gnd and3_dec
XDEC_AND_94 out_2 out_7 out_13 decode_94 vdd gnd and3_dec
XDEC_AND_110 out_2 out_7 out_14 decode_110 vdd gnd and3_dec
XDEC_AND_126 out_2 out_7 out_15 decode_126 vdd gnd and3_dec
XDEC_AND_3 out_3 out_4 out_8 decode_3 vdd gnd and3_dec
XDEC_AND_19 out_3 out_4 out_9 decode_19 vdd gnd and3_dec
XDEC_AND_35 out_3 out_4 out_10 decode_35 vdd gnd and3_dec
XDEC_AND_51 out_3 out_4 out_11 decode_51 vdd gnd and3_dec
XDEC_AND_67 out_3 out_4 out_12 decode_67 vdd gnd and3_dec
XDEC_AND_83 out_3 out_4 out_13 decode_83 vdd gnd and3_dec
XDEC_AND_99 out_3 out_4 out_14 decode_99 vdd gnd and3_dec
XDEC_AND_115 out_3 out_4 out_15 decode_115 vdd gnd and3_dec
XDEC_AND_7 out_3 out_5 out_8 decode_7 vdd gnd and3_dec
XDEC_AND_23 out_3 out_5 out_9 decode_23 vdd gnd and3_dec
XDEC_AND_39 out_3 out_5 out_10 decode_39 vdd gnd and3_dec
XDEC_AND_55 out_3 out_5 out_11 decode_55 vdd gnd and3_dec
XDEC_AND_71 out_3 out_5 out_12 decode_71 vdd gnd and3_dec
XDEC_AND_87 out_3 out_5 out_13 decode_87 vdd gnd and3_dec
XDEC_AND_103 out_3 out_5 out_14 decode_103 vdd gnd and3_dec
XDEC_AND_119 out_3 out_5 out_15 decode_119 vdd gnd and3_dec
XDEC_AND_11 out_3 out_6 out_8 decode_11 vdd gnd and3_dec
XDEC_AND_27 out_3 out_6 out_9 decode_27 vdd gnd and3_dec
XDEC_AND_43 out_3 out_6 out_10 decode_43 vdd gnd and3_dec
XDEC_AND_59 out_3 out_6 out_11 decode_59 vdd gnd and3_dec
XDEC_AND_75 out_3 out_6 out_12 decode_75 vdd gnd and3_dec
XDEC_AND_91 out_3 out_6 out_13 decode_91 vdd gnd and3_dec
XDEC_AND_107 out_3 out_6 out_14 decode_107 vdd gnd and3_dec
XDEC_AND_123 out_3 out_6 out_15 decode_123 vdd gnd and3_dec
XDEC_AND_15 out_3 out_7 out_8 decode_15 vdd gnd and3_dec
XDEC_AND_31 out_3 out_7 out_9 decode_31 vdd gnd and3_dec
XDEC_AND_47 out_3 out_7 out_10 decode_47 vdd gnd and3_dec
XDEC_AND_63 out_3 out_7 out_11 decode_63 vdd gnd and3_dec
XDEC_AND_79 out_3 out_7 out_12 decode_79 vdd gnd and3_dec
XDEC_AND_95 out_3 out_7 out_13 decode_95 vdd gnd and3_dec
XDEC_AND_111 out_3 out_7 out_14 decode_111 vdd gnd and3_dec
XDEC_AND_127 out_3 out_7 out_15 decode_127 vdd gnd and3_dec
.ENDS hierarchical_decoder

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u

* ptx M{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u

.SUBCKT pinv_dec_0 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u
.ENDS pinv_dec_0

.SUBCKT wordline_driver A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xwld_nand A B zb_int vdd gnd nand2_dec
Xwl_driver zb_int Z vdd gnd pinv_dec_0
.ENDS wordline_driver

.SUBCKT wordline_driver_array in_0 in_1 in_2 in_3 in_4 in_5 in_6 in_7 in_8 in_9 in_10 in_11 in_12 in_13 in_14 in_15 in_16 in_17 in_18 in_19 in_20 in_21 in_22 in_23 in_24 in_25 in_26 in_27 in_28 in_29 in_30 in_31 in_32 in_33 in_34 in_35 in_36 in_37 in_38 in_39 in_40 in_41 in_42 in_43 in_44 in_45 in_46 in_47 in_48 in_49 in_50 in_51 in_52 in_53 in_54 in_55 in_56 in_57 in_58 in_59 in_60 in_61 in_62 in_63 in_64 in_65 in_66 in_67 in_68 in_69 in_70 in_71 in_72 in_73 in_74 in_75 in_76 in_77 in_78 in_79 in_80 in_81 in_82 in_83 in_84 in_85 in_86 in_87 in_88 in_89 in_90 in_91 in_92 in_93 in_94 in_95 in_96 in_97 in_98 in_99 in_100 in_101 in_102 in_103 in_104 in_105 in_106 in_107 in_108 in_109 in_110 in_111 in_112 in_113 in_114 in_115 in_116 in_117 in_118 in_119 in_120 in_121 in_122 in_123 in_124 in_125 in_126 in_127 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 en vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* INPUT : in_3 
* INPUT : in_4 
* INPUT : in_5 
* INPUT : in_6 
* INPUT : in_7 
* INPUT : in_8 
* INPUT : in_9 
* INPUT : in_10 
* INPUT : in_11 
* INPUT : in_12 
* INPUT : in_13 
* INPUT : in_14 
* INPUT : in_15 
* INPUT : in_16 
* INPUT : in_17 
* INPUT : in_18 
* INPUT : in_19 
* INPUT : in_20 
* INPUT : in_21 
* INPUT : in_22 
* INPUT : in_23 
* INPUT : in_24 
* INPUT : in_25 
* INPUT : in_26 
* INPUT : in_27 
* INPUT : in_28 
* INPUT : in_29 
* INPUT : in_30 
* INPUT : in_31 
* INPUT : in_32 
* INPUT : in_33 
* INPUT : in_34 
* INPUT : in_35 
* INPUT : in_36 
* INPUT : in_37 
* INPUT : in_38 
* INPUT : in_39 
* INPUT : in_40 
* INPUT : in_41 
* INPUT : in_42 
* INPUT : in_43 
* INPUT : in_44 
* INPUT : in_45 
* INPUT : in_46 
* INPUT : in_47 
* INPUT : in_48 
* INPUT : in_49 
* INPUT : in_50 
* INPUT : in_51 
* INPUT : in_52 
* INPUT : in_53 
* INPUT : in_54 
* INPUT : in_55 
* INPUT : in_56 
* INPUT : in_57 
* INPUT : in_58 
* INPUT : in_59 
* INPUT : in_60 
* INPUT : in_61 
* INPUT : in_62 
* INPUT : in_63 
* INPUT : in_64 
* INPUT : in_65 
* INPUT : in_66 
* INPUT : in_67 
* INPUT : in_68 
* INPUT : in_69 
* INPUT : in_70 
* INPUT : in_71 
* INPUT : in_72 
* INPUT : in_73 
* INPUT : in_74 
* INPUT : in_75 
* INPUT : in_76 
* INPUT : in_77 
* INPUT : in_78 
* INPUT : in_79 
* INPUT : in_80 
* INPUT : in_81 
* INPUT : in_82 
* INPUT : in_83 
* INPUT : in_84 
* INPUT : in_85 
* INPUT : in_86 
* INPUT : in_87 
* INPUT : in_88 
* INPUT : in_89 
* INPUT : in_90 
* INPUT : in_91 
* INPUT : in_92 
* INPUT : in_93 
* INPUT : in_94 
* INPUT : in_95 
* INPUT : in_96 
* INPUT : in_97 
* INPUT : in_98 
* INPUT : in_99 
* INPUT : in_100 
* INPUT : in_101 
* INPUT : in_102 
* INPUT : in_103 
* INPUT : in_104 
* INPUT : in_105 
* INPUT : in_106 
* INPUT : in_107 
* INPUT : in_108 
* INPUT : in_109 
* INPUT : in_110 
* INPUT : in_111 
* INPUT : in_112 
* INPUT : in_113 
* INPUT : in_114 
* INPUT : in_115 
* INPUT : in_116 
* INPUT : in_117 
* INPUT : in_118 
* INPUT : in_119 
* INPUT : in_120 
* INPUT : in_121 
* INPUT : in_122 
* INPUT : in_123 
* INPUT : in_124 
* INPUT : in_125 
* INPUT : in_126 
* INPUT : in_127 
* OUTPUT: wl_0 
* OUTPUT: wl_1 
* OUTPUT: wl_2 
* OUTPUT: wl_3 
* OUTPUT: wl_4 
* OUTPUT: wl_5 
* OUTPUT: wl_6 
* OUTPUT: wl_7 
* OUTPUT: wl_8 
* OUTPUT: wl_9 
* OUTPUT: wl_10 
* OUTPUT: wl_11 
* OUTPUT: wl_12 
* OUTPUT: wl_13 
* OUTPUT: wl_14 
* OUTPUT: wl_15 
* OUTPUT: wl_16 
* OUTPUT: wl_17 
* OUTPUT: wl_18 
* OUTPUT: wl_19 
* OUTPUT: wl_20 
* OUTPUT: wl_21 
* OUTPUT: wl_22 
* OUTPUT: wl_23 
* OUTPUT: wl_24 
* OUTPUT: wl_25 
* OUTPUT: wl_26 
* OUTPUT: wl_27 
* OUTPUT: wl_28 
* OUTPUT: wl_29 
* OUTPUT: wl_30 
* OUTPUT: wl_31 
* OUTPUT: wl_32 
* OUTPUT: wl_33 
* OUTPUT: wl_34 
* OUTPUT: wl_35 
* OUTPUT: wl_36 
* OUTPUT: wl_37 
* OUTPUT: wl_38 
* OUTPUT: wl_39 
* OUTPUT: wl_40 
* OUTPUT: wl_41 
* OUTPUT: wl_42 
* OUTPUT: wl_43 
* OUTPUT: wl_44 
* OUTPUT: wl_45 
* OUTPUT: wl_46 
* OUTPUT: wl_47 
* OUTPUT: wl_48 
* OUTPUT: wl_49 
* OUTPUT: wl_50 
* OUTPUT: wl_51 
* OUTPUT: wl_52 
* OUTPUT: wl_53 
* OUTPUT: wl_54 
* OUTPUT: wl_55 
* OUTPUT: wl_56 
* OUTPUT: wl_57 
* OUTPUT: wl_58 
* OUTPUT: wl_59 
* OUTPUT: wl_60 
* OUTPUT: wl_61 
* OUTPUT: wl_62 
* OUTPUT: wl_63 
* OUTPUT: wl_64 
* OUTPUT: wl_65 
* OUTPUT: wl_66 
* OUTPUT: wl_67 
* OUTPUT: wl_68 
* OUTPUT: wl_69 
* OUTPUT: wl_70 
* OUTPUT: wl_71 
* OUTPUT: wl_72 
* OUTPUT: wl_73 
* OUTPUT: wl_74 
* OUTPUT: wl_75 
* OUTPUT: wl_76 
* OUTPUT: wl_77 
* OUTPUT: wl_78 
* OUTPUT: wl_79 
* OUTPUT: wl_80 
* OUTPUT: wl_81 
* OUTPUT: wl_82 
* OUTPUT: wl_83 
* OUTPUT: wl_84 
* OUTPUT: wl_85 
* OUTPUT: wl_86 
* OUTPUT: wl_87 
* OUTPUT: wl_88 
* OUTPUT: wl_89 
* OUTPUT: wl_90 
* OUTPUT: wl_91 
* OUTPUT: wl_92 
* OUTPUT: wl_93 
* OUTPUT: wl_94 
* OUTPUT: wl_95 
* OUTPUT: wl_96 
* OUTPUT: wl_97 
* OUTPUT: wl_98 
* OUTPUT: wl_99 
* OUTPUT: wl_100 
* OUTPUT: wl_101 
* OUTPUT: wl_102 
* OUTPUT: wl_103 
* OUTPUT: wl_104 
* OUTPUT: wl_105 
* OUTPUT: wl_106 
* OUTPUT: wl_107 
* OUTPUT: wl_108 
* OUTPUT: wl_109 
* OUTPUT: wl_110 
* OUTPUT: wl_111 
* OUTPUT: wl_112 
* OUTPUT: wl_113 
* OUTPUT: wl_114 
* OUTPUT: wl_115 
* OUTPUT: wl_116 
* OUTPUT: wl_117 
* OUTPUT: wl_118 
* OUTPUT: wl_119 
* OUTPUT: wl_120 
* OUTPUT: wl_121 
* OUTPUT: wl_122 
* OUTPUT: wl_123 
* OUTPUT: wl_124 
* OUTPUT: wl_125 
* OUTPUT: wl_126 
* OUTPUT: wl_127 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* rows: 128 cols: 64
Xwl_driver_and0 in_0 en wl_0 vdd gnd wordline_driver
Xwl_driver_and1 in_1 en wl_1 vdd gnd wordline_driver
Xwl_driver_and2 in_2 en wl_2 vdd gnd wordline_driver
Xwl_driver_and3 in_3 en wl_3 vdd gnd wordline_driver
Xwl_driver_and4 in_4 en wl_4 vdd gnd wordline_driver
Xwl_driver_and5 in_5 en wl_5 vdd gnd wordline_driver
Xwl_driver_and6 in_6 en wl_6 vdd gnd wordline_driver
Xwl_driver_and7 in_7 en wl_7 vdd gnd wordline_driver
Xwl_driver_and8 in_8 en wl_8 vdd gnd wordline_driver
Xwl_driver_and9 in_9 en wl_9 vdd gnd wordline_driver
Xwl_driver_and10 in_10 en wl_10 vdd gnd wordline_driver
Xwl_driver_and11 in_11 en wl_11 vdd gnd wordline_driver
Xwl_driver_and12 in_12 en wl_12 vdd gnd wordline_driver
Xwl_driver_and13 in_13 en wl_13 vdd gnd wordline_driver
Xwl_driver_and14 in_14 en wl_14 vdd gnd wordline_driver
Xwl_driver_and15 in_15 en wl_15 vdd gnd wordline_driver
Xwl_driver_and16 in_16 en wl_16 vdd gnd wordline_driver
Xwl_driver_and17 in_17 en wl_17 vdd gnd wordline_driver
Xwl_driver_and18 in_18 en wl_18 vdd gnd wordline_driver
Xwl_driver_and19 in_19 en wl_19 vdd gnd wordline_driver
Xwl_driver_and20 in_20 en wl_20 vdd gnd wordline_driver
Xwl_driver_and21 in_21 en wl_21 vdd gnd wordline_driver
Xwl_driver_and22 in_22 en wl_22 vdd gnd wordline_driver
Xwl_driver_and23 in_23 en wl_23 vdd gnd wordline_driver
Xwl_driver_and24 in_24 en wl_24 vdd gnd wordline_driver
Xwl_driver_and25 in_25 en wl_25 vdd gnd wordline_driver
Xwl_driver_and26 in_26 en wl_26 vdd gnd wordline_driver
Xwl_driver_and27 in_27 en wl_27 vdd gnd wordline_driver
Xwl_driver_and28 in_28 en wl_28 vdd gnd wordline_driver
Xwl_driver_and29 in_29 en wl_29 vdd gnd wordline_driver
Xwl_driver_and30 in_30 en wl_30 vdd gnd wordline_driver
Xwl_driver_and31 in_31 en wl_31 vdd gnd wordline_driver
Xwl_driver_and32 in_32 en wl_32 vdd gnd wordline_driver
Xwl_driver_and33 in_33 en wl_33 vdd gnd wordline_driver
Xwl_driver_and34 in_34 en wl_34 vdd gnd wordline_driver
Xwl_driver_and35 in_35 en wl_35 vdd gnd wordline_driver
Xwl_driver_and36 in_36 en wl_36 vdd gnd wordline_driver
Xwl_driver_and37 in_37 en wl_37 vdd gnd wordline_driver
Xwl_driver_and38 in_38 en wl_38 vdd gnd wordline_driver
Xwl_driver_and39 in_39 en wl_39 vdd gnd wordline_driver
Xwl_driver_and40 in_40 en wl_40 vdd gnd wordline_driver
Xwl_driver_and41 in_41 en wl_41 vdd gnd wordline_driver
Xwl_driver_and42 in_42 en wl_42 vdd gnd wordline_driver
Xwl_driver_and43 in_43 en wl_43 vdd gnd wordline_driver
Xwl_driver_and44 in_44 en wl_44 vdd gnd wordline_driver
Xwl_driver_and45 in_45 en wl_45 vdd gnd wordline_driver
Xwl_driver_and46 in_46 en wl_46 vdd gnd wordline_driver
Xwl_driver_and47 in_47 en wl_47 vdd gnd wordline_driver
Xwl_driver_and48 in_48 en wl_48 vdd gnd wordline_driver
Xwl_driver_and49 in_49 en wl_49 vdd gnd wordline_driver
Xwl_driver_and50 in_50 en wl_50 vdd gnd wordline_driver
Xwl_driver_and51 in_51 en wl_51 vdd gnd wordline_driver
Xwl_driver_and52 in_52 en wl_52 vdd gnd wordline_driver
Xwl_driver_and53 in_53 en wl_53 vdd gnd wordline_driver
Xwl_driver_and54 in_54 en wl_54 vdd gnd wordline_driver
Xwl_driver_and55 in_55 en wl_55 vdd gnd wordline_driver
Xwl_driver_and56 in_56 en wl_56 vdd gnd wordline_driver
Xwl_driver_and57 in_57 en wl_57 vdd gnd wordline_driver
Xwl_driver_and58 in_58 en wl_58 vdd gnd wordline_driver
Xwl_driver_and59 in_59 en wl_59 vdd gnd wordline_driver
Xwl_driver_and60 in_60 en wl_60 vdd gnd wordline_driver
Xwl_driver_and61 in_61 en wl_61 vdd gnd wordline_driver
Xwl_driver_and62 in_62 en wl_62 vdd gnd wordline_driver
Xwl_driver_and63 in_63 en wl_63 vdd gnd wordline_driver
Xwl_driver_and64 in_64 en wl_64 vdd gnd wordline_driver
Xwl_driver_and65 in_65 en wl_65 vdd gnd wordline_driver
Xwl_driver_and66 in_66 en wl_66 vdd gnd wordline_driver
Xwl_driver_and67 in_67 en wl_67 vdd gnd wordline_driver
Xwl_driver_and68 in_68 en wl_68 vdd gnd wordline_driver
Xwl_driver_and69 in_69 en wl_69 vdd gnd wordline_driver
Xwl_driver_and70 in_70 en wl_70 vdd gnd wordline_driver
Xwl_driver_and71 in_71 en wl_71 vdd gnd wordline_driver
Xwl_driver_and72 in_72 en wl_72 vdd gnd wordline_driver
Xwl_driver_and73 in_73 en wl_73 vdd gnd wordline_driver
Xwl_driver_and74 in_74 en wl_74 vdd gnd wordline_driver
Xwl_driver_and75 in_75 en wl_75 vdd gnd wordline_driver
Xwl_driver_and76 in_76 en wl_76 vdd gnd wordline_driver
Xwl_driver_and77 in_77 en wl_77 vdd gnd wordline_driver
Xwl_driver_and78 in_78 en wl_78 vdd gnd wordline_driver
Xwl_driver_and79 in_79 en wl_79 vdd gnd wordline_driver
Xwl_driver_and80 in_80 en wl_80 vdd gnd wordline_driver
Xwl_driver_and81 in_81 en wl_81 vdd gnd wordline_driver
Xwl_driver_and82 in_82 en wl_82 vdd gnd wordline_driver
Xwl_driver_and83 in_83 en wl_83 vdd gnd wordline_driver
Xwl_driver_and84 in_84 en wl_84 vdd gnd wordline_driver
Xwl_driver_and85 in_85 en wl_85 vdd gnd wordline_driver
Xwl_driver_and86 in_86 en wl_86 vdd gnd wordline_driver
Xwl_driver_and87 in_87 en wl_87 vdd gnd wordline_driver
Xwl_driver_and88 in_88 en wl_88 vdd gnd wordline_driver
Xwl_driver_and89 in_89 en wl_89 vdd gnd wordline_driver
Xwl_driver_and90 in_90 en wl_90 vdd gnd wordline_driver
Xwl_driver_and91 in_91 en wl_91 vdd gnd wordline_driver
Xwl_driver_and92 in_92 en wl_92 vdd gnd wordline_driver
Xwl_driver_and93 in_93 en wl_93 vdd gnd wordline_driver
Xwl_driver_and94 in_94 en wl_94 vdd gnd wordline_driver
Xwl_driver_and95 in_95 en wl_95 vdd gnd wordline_driver
Xwl_driver_and96 in_96 en wl_96 vdd gnd wordline_driver
Xwl_driver_and97 in_97 en wl_97 vdd gnd wordline_driver
Xwl_driver_and98 in_98 en wl_98 vdd gnd wordline_driver
Xwl_driver_and99 in_99 en wl_99 vdd gnd wordline_driver
Xwl_driver_and100 in_100 en wl_100 vdd gnd wordline_driver
Xwl_driver_and101 in_101 en wl_101 vdd gnd wordline_driver
Xwl_driver_and102 in_102 en wl_102 vdd gnd wordline_driver
Xwl_driver_and103 in_103 en wl_103 vdd gnd wordline_driver
Xwl_driver_and104 in_104 en wl_104 vdd gnd wordline_driver
Xwl_driver_and105 in_105 en wl_105 vdd gnd wordline_driver
Xwl_driver_and106 in_106 en wl_106 vdd gnd wordline_driver
Xwl_driver_and107 in_107 en wl_107 vdd gnd wordline_driver
Xwl_driver_and108 in_108 en wl_108 vdd gnd wordline_driver
Xwl_driver_and109 in_109 en wl_109 vdd gnd wordline_driver
Xwl_driver_and110 in_110 en wl_110 vdd gnd wordline_driver
Xwl_driver_and111 in_111 en wl_111 vdd gnd wordline_driver
Xwl_driver_and112 in_112 en wl_112 vdd gnd wordline_driver
Xwl_driver_and113 in_113 en wl_113 vdd gnd wordline_driver
Xwl_driver_and114 in_114 en wl_114 vdd gnd wordline_driver
Xwl_driver_and115 in_115 en wl_115 vdd gnd wordline_driver
Xwl_driver_and116 in_116 en wl_116 vdd gnd wordline_driver
Xwl_driver_and117 in_117 en wl_117 vdd gnd wordline_driver
Xwl_driver_and118 in_118 en wl_118 vdd gnd wordline_driver
Xwl_driver_and119 in_119 en wl_119 vdd gnd wordline_driver
Xwl_driver_and120 in_120 en wl_120 vdd gnd wordline_driver
Xwl_driver_and121 in_121 en wl_121 vdd gnd wordline_driver
Xwl_driver_and122 in_122 en wl_122 vdd gnd wordline_driver
Xwl_driver_and123 in_123 en wl_123 vdd gnd wordline_driver
Xwl_driver_and124 in_124 en wl_124 vdd gnd wordline_driver
Xwl_driver_and125 in_125 en wl_125 vdd gnd wordline_driver
Xwl_driver_and126 in_126 en wl_126 vdd gnd wordline_driver
Xwl_driver_and127 in_127 en wl_127 vdd gnd wordline_driver
.ENDS wordline_driver_array

.SUBCKT port_address addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 addr_6 wl_en wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 vdd gnd
* INPUT : addr_0 
* INPUT : addr_1 
* INPUT : addr_2 
* INPUT : addr_3 
* INPUT : addr_4 
* INPUT : addr_5 
* INPUT : addr_6 
* INPUT : wl_en 
* OUTPUT: wl_0 
* OUTPUT: wl_1 
* OUTPUT: wl_2 
* OUTPUT: wl_3 
* OUTPUT: wl_4 
* OUTPUT: wl_5 
* OUTPUT: wl_6 
* OUTPUT: wl_7 
* OUTPUT: wl_8 
* OUTPUT: wl_9 
* OUTPUT: wl_10 
* OUTPUT: wl_11 
* OUTPUT: wl_12 
* OUTPUT: wl_13 
* OUTPUT: wl_14 
* OUTPUT: wl_15 
* OUTPUT: wl_16 
* OUTPUT: wl_17 
* OUTPUT: wl_18 
* OUTPUT: wl_19 
* OUTPUT: wl_20 
* OUTPUT: wl_21 
* OUTPUT: wl_22 
* OUTPUT: wl_23 
* OUTPUT: wl_24 
* OUTPUT: wl_25 
* OUTPUT: wl_26 
* OUTPUT: wl_27 
* OUTPUT: wl_28 
* OUTPUT: wl_29 
* OUTPUT: wl_30 
* OUTPUT: wl_31 
* OUTPUT: wl_32 
* OUTPUT: wl_33 
* OUTPUT: wl_34 
* OUTPUT: wl_35 
* OUTPUT: wl_36 
* OUTPUT: wl_37 
* OUTPUT: wl_38 
* OUTPUT: wl_39 
* OUTPUT: wl_40 
* OUTPUT: wl_41 
* OUTPUT: wl_42 
* OUTPUT: wl_43 
* OUTPUT: wl_44 
* OUTPUT: wl_45 
* OUTPUT: wl_46 
* OUTPUT: wl_47 
* OUTPUT: wl_48 
* OUTPUT: wl_49 
* OUTPUT: wl_50 
* OUTPUT: wl_51 
* OUTPUT: wl_52 
* OUTPUT: wl_53 
* OUTPUT: wl_54 
* OUTPUT: wl_55 
* OUTPUT: wl_56 
* OUTPUT: wl_57 
* OUTPUT: wl_58 
* OUTPUT: wl_59 
* OUTPUT: wl_60 
* OUTPUT: wl_61 
* OUTPUT: wl_62 
* OUTPUT: wl_63 
* OUTPUT: wl_64 
* OUTPUT: wl_65 
* OUTPUT: wl_66 
* OUTPUT: wl_67 
* OUTPUT: wl_68 
* OUTPUT: wl_69 
* OUTPUT: wl_70 
* OUTPUT: wl_71 
* OUTPUT: wl_72 
* OUTPUT: wl_73 
* OUTPUT: wl_74 
* OUTPUT: wl_75 
* OUTPUT: wl_76 
* OUTPUT: wl_77 
* OUTPUT: wl_78 
* OUTPUT: wl_79 
* OUTPUT: wl_80 
* OUTPUT: wl_81 
* OUTPUT: wl_82 
* OUTPUT: wl_83 
* OUTPUT: wl_84 
* OUTPUT: wl_85 
* OUTPUT: wl_86 
* OUTPUT: wl_87 
* OUTPUT: wl_88 
* OUTPUT: wl_89 
* OUTPUT: wl_90 
* OUTPUT: wl_91 
* OUTPUT: wl_92 
* OUTPUT: wl_93 
* OUTPUT: wl_94 
* OUTPUT: wl_95 
* OUTPUT: wl_96 
* OUTPUT: wl_97 
* OUTPUT: wl_98 
* OUTPUT: wl_99 
* OUTPUT: wl_100 
* OUTPUT: wl_101 
* OUTPUT: wl_102 
* OUTPUT: wl_103 
* OUTPUT: wl_104 
* OUTPUT: wl_105 
* OUTPUT: wl_106 
* OUTPUT: wl_107 
* OUTPUT: wl_108 
* OUTPUT: wl_109 
* OUTPUT: wl_110 
* OUTPUT: wl_111 
* OUTPUT: wl_112 
* OUTPUT: wl_113 
* OUTPUT: wl_114 
* OUTPUT: wl_115 
* OUTPUT: wl_116 
* OUTPUT: wl_117 
* OUTPUT: wl_118 
* OUTPUT: wl_119 
* OUTPUT: wl_120 
* OUTPUT: wl_121 
* OUTPUT: wl_122 
* OUTPUT: wl_123 
* OUTPUT: wl_124 
* OUTPUT: wl_125 
* OUTPUT: wl_126 
* OUTPUT: wl_127 
* POWER : vdd 
* GROUND: gnd 
Xrow_decoder addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 addr_6 dec_out_0 dec_out_1 dec_out_2 dec_out_3 dec_out_4 dec_out_5 dec_out_6 dec_out_7 dec_out_8 dec_out_9 dec_out_10 dec_out_11 dec_out_12 dec_out_13 dec_out_14 dec_out_15 dec_out_16 dec_out_17 dec_out_18 dec_out_19 dec_out_20 dec_out_21 dec_out_22 dec_out_23 dec_out_24 dec_out_25 dec_out_26 dec_out_27 dec_out_28 dec_out_29 dec_out_30 dec_out_31 dec_out_32 dec_out_33 dec_out_34 dec_out_35 dec_out_36 dec_out_37 dec_out_38 dec_out_39 dec_out_40 dec_out_41 dec_out_42 dec_out_43 dec_out_44 dec_out_45 dec_out_46 dec_out_47 dec_out_48 dec_out_49 dec_out_50 dec_out_51 dec_out_52 dec_out_53 dec_out_54 dec_out_55 dec_out_56 dec_out_57 dec_out_58 dec_out_59 dec_out_60 dec_out_61 dec_out_62 dec_out_63 dec_out_64 dec_out_65 dec_out_66 dec_out_67 dec_out_68 dec_out_69 dec_out_70 dec_out_71 dec_out_72 dec_out_73 dec_out_74 dec_out_75 dec_out_76 dec_out_77 dec_out_78 dec_out_79 dec_out_80 dec_out_81 dec_out_82 dec_out_83 dec_out_84 dec_out_85 dec_out_86 dec_out_87 dec_out_88 dec_out_89 dec_out_90 dec_out_91 dec_out_92 dec_out_93 dec_out_94 dec_out_95 dec_out_96 dec_out_97 dec_out_98 dec_out_99 dec_out_100 dec_out_101 dec_out_102 dec_out_103 dec_out_104 dec_out_105 dec_out_106 dec_out_107 dec_out_108 dec_out_109 dec_out_110 dec_out_111 dec_out_112 dec_out_113 dec_out_114 dec_out_115 dec_out_116 dec_out_117 dec_out_118 dec_out_119 dec_out_120 dec_out_121 dec_out_122 dec_out_123 dec_out_124 dec_out_125 dec_out_126 dec_out_127 vdd gnd hierarchical_decoder
Xwordline_driver dec_out_0 dec_out_1 dec_out_2 dec_out_3 dec_out_4 dec_out_5 dec_out_6 dec_out_7 dec_out_8 dec_out_9 dec_out_10 dec_out_11 dec_out_12 dec_out_13 dec_out_14 dec_out_15 dec_out_16 dec_out_17 dec_out_18 dec_out_19 dec_out_20 dec_out_21 dec_out_22 dec_out_23 dec_out_24 dec_out_25 dec_out_26 dec_out_27 dec_out_28 dec_out_29 dec_out_30 dec_out_31 dec_out_32 dec_out_33 dec_out_34 dec_out_35 dec_out_36 dec_out_37 dec_out_38 dec_out_39 dec_out_40 dec_out_41 dec_out_42 dec_out_43 dec_out_44 dec_out_45 dec_out_46 dec_out_47 dec_out_48 dec_out_49 dec_out_50 dec_out_51 dec_out_52 dec_out_53 dec_out_54 dec_out_55 dec_out_56 dec_out_57 dec_out_58 dec_out_59 dec_out_60 dec_out_61 dec_out_62 dec_out_63 dec_out_64 dec_out_65 dec_out_66 dec_out_67 dec_out_68 dec_out_69 dec_out_70 dec_out_71 dec_out_72 dec_out_73 dec_out_74 dec_out_75 dec_out_76 dec_out_77 dec_out_78 dec_out_79 dec_out_80 dec_out_81 dec_out_82 dec_out_83 dec_out_84 dec_out_85 dec_out_86 dec_out_87 dec_out_88 dec_out_89 dec_out_90 dec_out_91 dec_out_92 dec_out_93 dec_out_94 dec_out_95 dec_out_96 dec_out_97 dec_out_98 dec_out_99 dec_out_100 dec_out_101 dec_out_102 dec_out_103 dec_out_104 dec_out_105 dec_out_106 dec_out_107 dec_out_108 dec_out_109 dec_out_110 dec_out_111 dec_out_112 dec_out_113 dec_out_114 dec_out_115 dec_out_116 dec_out_117 dec_out_118 dec_out_119 dec_out_120 dec_out_121 dec_out_122 dec_out_123 dec_out_124 dec_out_125 dec_out_126 dec_out_127 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_en vdd gnd wordline_driver_array
.ENDS port_address

.SUBCKT sky130_fd_bd_sram__openram_dp_cell bl0 br0 bl1 br1 wl0 wl1 vdd gnd
**
*.SEEDPROM

* Bitcell Core
XM0 Q wl1 bl1 gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM1 gnd Q_bar Q gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM2 gnd Q_bar Q gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM3 bl0 wl0 Q gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM4 Q_bar wl1 br1 gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM5 gnd Q Q_bar gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM6 gnd Q Q_bar gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM7 br0 wl0 Q_bar gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM8 vdd Q Q_bar vdd sky130_fd_pr__special_pfet_pass W=0.14 L=0.15 m=1
XM9 Q Q_bar vdd vdd sky130_fd_pr__special_pfet_pass W=0.14 L=0.15 m=1

* drainOnly PMOS
XM10 Q_bar wl1 Q_bar vdd sky130_fd_pr__special_pfet_pass L=0.08 W=0.14 m=1
XM11 Q wl0 Q vdd sky130_fd_pr__special_pfet_pass L=0.08 W=0.14 m=1

* drainOnly NMOS
XM12 bl1 gnd bl1 gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.08 m=1
XM14 br1 gnd br1 gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.08 m=1

.ENDS

.SUBCKT bitcell_array bl0_0 br0_0 bl1_0 br1_0 bl0_1 br0_1 bl1_1 br1_1 bl0_2 br0_2 bl1_2 br1_2 bl0_3 br0_3 bl1_3 br1_3 bl0_4 br0_4 bl1_4 br1_4 bl0_5 br0_5 bl1_5 br1_5 bl0_6 br0_6 bl1_6 br1_6 bl0_7 br0_7 bl1_7 br1_7 bl0_8 br0_8 bl1_8 br1_8 bl0_9 br0_9 bl1_9 br1_9 bl0_10 br0_10 bl1_10 br1_10 bl0_11 br0_11 bl1_11 br1_11 bl0_12 br0_12 bl1_12 br1_12 bl0_13 br0_13 bl1_13 br1_13 bl0_14 br0_14 bl1_14 br1_14 bl0_15 br0_15 bl1_15 br1_15 bl0_16 br0_16 bl1_16 br1_16 bl0_17 br0_17 bl1_17 br1_17 bl0_18 br0_18 bl1_18 br1_18 bl0_19 br0_19 bl1_19 br1_19 bl0_20 br0_20 bl1_20 br1_20 bl0_21 br0_21 bl1_21 br1_21 bl0_22 br0_22 bl1_22 br1_22 bl0_23 br0_23 bl1_23 br1_23 bl0_24 br0_24 bl1_24 br1_24 bl0_25 br0_25 bl1_25 br1_25 bl0_26 br0_26 bl1_26 br1_26 bl0_27 br0_27 bl1_27 br1_27 bl0_28 br0_28 bl1_28 br1_28 bl0_29 br0_29 bl1_29 br1_29 bl0_30 br0_30 bl1_30 br1_30 bl0_31 br0_31 bl1_31 br1_31 bl0_32 br0_32 bl1_32 br1_32 bl0_33 br0_33 bl1_33 br1_33 bl0_34 br0_34 bl1_34 br1_34 bl0_35 br0_35 bl1_35 br1_35 bl0_36 br0_36 bl1_36 br1_36 bl0_37 br0_37 bl1_37 br1_37 bl0_38 br0_38 bl1_38 br1_38 bl0_39 br0_39 bl1_39 br1_39 bl0_40 br0_40 bl1_40 br1_40 bl0_41 br0_41 bl1_41 br1_41 bl0_42 br0_42 bl1_42 br1_42 bl0_43 br0_43 bl1_43 br1_43 bl0_44 br0_44 bl1_44 br1_44 bl0_45 br0_45 bl1_45 br1_45 bl0_46 br0_46 bl1_46 br1_46 bl0_47 br0_47 bl1_47 br1_47 bl0_48 br0_48 bl1_48 br1_48 bl0_49 br0_49 bl1_49 br1_49 bl0_50 br0_50 bl1_50 br1_50 bl0_51 br0_51 bl1_51 br1_51 bl0_52 br0_52 bl1_52 br1_52 bl0_53 br0_53 bl1_53 br1_53 bl0_54 br0_54 bl1_54 br1_54 bl0_55 br0_55 bl1_55 br1_55 bl0_56 br0_56 bl1_56 br1_56 bl0_57 br0_57 bl1_57 br1_57 bl0_58 br0_58 bl1_58 br1_58 bl0_59 br0_59 bl1_59 br1_59 bl0_60 br0_60 bl1_60 br1_60 bl0_61 br0_61 bl1_61 br1_61 bl0_62 br0_62 bl1_62 br1_62 bl0_63 br0_63 bl1_63 br1_63 wl0_0 wl1_0 wl0_1 wl1_1 wl0_2 wl1_2 wl0_3 wl1_3 wl0_4 wl1_4 wl0_5 wl1_5 wl0_6 wl1_6 wl0_7 wl1_7 wl0_8 wl1_8 wl0_9 wl1_9 wl0_10 wl1_10 wl0_11 wl1_11 wl0_12 wl1_12 wl0_13 wl1_13 wl0_14 wl1_14 wl0_15 wl1_15 wl0_16 wl1_16 wl0_17 wl1_17 wl0_18 wl1_18 wl0_19 wl1_19 wl0_20 wl1_20 wl0_21 wl1_21 wl0_22 wl1_22 wl0_23 wl1_23 wl0_24 wl1_24 wl0_25 wl1_25 wl0_26 wl1_26 wl0_27 wl1_27 wl0_28 wl1_28 wl0_29 wl1_29 wl0_30 wl1_30 wl0_31 wl1_31 wl0_32 wl1_32 wl0_33 wl1_33 wl0_34 wl1_34 wl0_35 wl1_35 wl0_36 wl1_36 wl0_37 wl1_37 wl0_38 wl1_38 wl0_39 wl1_39 wl0_40 wl1_40 wl0_41 wl1_41 wl0_42 wl1_42 wl0_43 wl1_43 wl0_44 wl1_44 wl0_45 wl1_45 wl0_46 wl1_46 wl0_47 wl1_47 wl0_48 wl1_48 wl0_49 wl1_49 wl0_50 wl1_50 wl0_51 wl1_51 wl0_52 wl1_52 wl0_53 wl1_53 wl0_54 wl1_54 wl0_55 wl1_55 wl0_56 wl1_56 wl0_57 wl1_57 wl0_58 wl1_58 wl0_59 wl1_59 wl0_60 wl1_60 wl0_61 wl1_61 wl0_62 wl1_62 wl0_63 wl1_63 wl0_64 wl1_64 wl0_65 wl1_65 wl0_66 wl1_66 wl0_67 wl1_67 wl0_68 wl1_68 wl0_69 wl1_69 wl0_70 wl1_70 wl0_71 wl1_71 wl0_72 wl1_72 wl0_73 wl1_73 wl0_74 wl1_74 wl0_75 wl1_75 wl0_76 wl1_76 wl0_77 wl1_77 wl0_78 wl1_78 wl0_79 wl1_79 wl0_80 wl1_80 wl0_81 wl1_81 wl0_82 wl1_82 wl0_83 wl1_83 wl0_84 wl1_84 wl0_85 wl1_85 wl0_86 wl1_86 wl0_87 wl1_87 wl0_88 wl1_88 wl0_89 wl1_89 wl0_90 wl1_90 wl0_91 wl1_91 wl0_92 wl1_92 wl0_93 wl1_93 wl0_94 wl1_94 wl0_95 wl1_95 wl0_96 wl1_96 wl0_97 wl1_97 wl0_98 wl1_98 wl0_99 wl1_99 wl0_100 wl1_100 wl0_101 wl1_101 wl0_102 wl1_102 wl0_103 wl1_103 wl0_104 wl1_104 wl0_105 wl1_105 wl0_106 wl1_106 wl0_107 wl1_107 wl0_108 wl1_108 wl0_109 wl1_109 wl0_110 wl1_110 wl0_111 wl1_111 wl0_112 wl1_112 wl0_113 wl1_113 wl0_114 wl1_114 wl0_115 wl1_115 wl0_116 wl1_116 wl0_117 wl1_117 wl0_118 wl1_118 wl0_119 wl1_119 wl0_120 wl1_120 wl0_121 wl1_121 wl0_122 wl1_122 wl0_123 wl1_123 wl0_124 wl1_124 wl0_125 wl1_125 wl0_126 wl1_126 wl0_127 wl1_127 vdd gnd
* INOUT : bl0_0 
* INOUT : br0_0 
* INOUT : bl1_0 
* INOUT : br1_0 
* INOUT : bl0_1 
* INOUT : br0_1 
* INOUT : bl1_1 
* INOUT : br1_1 
* INOUT : bl0_2 
* INOUT : br0_2 
* INOUT : bl1_2 
* INOUT : br1_2 
* INOUT : bl0_3 
* INOUT : br0_3 
* INOUT : bl1_3 
* INOUT : br1_3 
* INOUT : bl0_4 
* INOUT : br0_4 
* INOUT : bl1_4 
* INOUT : br1_4 
* INOUT : bl0_5 
* INOUT : br0_5 
* INOUT : bl1_5 
* INOUT : br1_5 
* INOUT : bl0_6 
* INOUT : br0_6 
* INOUT : bl1_6 
* INOUT : br1_6 
* INOUT : bl0_7 
* INOUT : br0_7 
* INOUT : bl1_7 
* INOUT : br1_7 
* INOUT : bl0_8 
* INOUT : br0_8 
* INOUT : bl1_8 
* INOUT : br1_8 
* INOUT : bl0_9 
* INOUT : br0_9 
* INOUT : bl1_9 
* INOUT : br1_9 
* INOUT : bl0_10 
* INOUT : br0_10 
* INOUT : bl1_10 
* INOUT : br1_10 
* INOUT : bl0_11 
* INOUT : br0_11 
* INOUT : bl1_11 
* INOUT : br1_11 
* INOUT : bl0_12 
* INOUT : br0_12 
* INOUT : bl1_12 
* INOUT : br1_12 
* INOUT : bl0_13 
* INOUT : br0_13 
* INOUT : bl1_13 
* INOUT : br1_13 
* INOUT : bl0_14 
* INOUT : br0_14 
* INOUT : bl1_14 
* INOUT : br1_14 
* INOUT : bl0_15 
* INOUT : br0_15 
* INOUT : bl1_15 
* INOUT : br1_15 
* INOUT : bl0_16 
* INOUT : br0_16 
* INOUT : bl1_16 
* INOUT : br1_16 
* INOUT : bl0_17 
* INOUT : br0_17 
* INOUT : bl1_17 
* INOUT : br1_17 
* INOUT : bl0_18 
* INOUT : br0_18 
* INOUT : bl1_18 
* INOUT : br1_18 
* INOUT : bl0_19 
* INOUT : br0_19 
* INOUT : bl1_19 
* INOUT : br1_19 
* INOUT : bl0_20 
* INOUT : br0_20 
* INOUT : bl1_20 
* INOUT : br1_20 
* INOUT : bl0_21 
* INOUT : br0_21 
* INOUT : bl1_21 
* INOUT : br1_21 
* INOUT : bl0_22 
* INOUT : br0_22 
* INOUT : bl1_22 
* INOUT : br1_22 
* INOUT : bl0_23 
* INOUT : br0_23 
* INOUT : bl1_23 
* INOUT : br1_23 
* INOUT : bl0_24 
* INOUT : br0_24 
* INOUT : bl1_24 
* INOUT : br1_24 
* INOUT : bl0_25 
* INOUT : br0_25 
* INOUT : bl1_25 
* INOUT : br1_25 
* INOUT : bl0_26 
* INOUT : br0_26 
* INOUT : bl1_26 
* INOUT : br1_26 
* INOUT : bl0_27 
* INOUT : br0_27 
* INOUT : bl1_27 
* INOUT : br1_27 
* INOUT : bl0_28 
* INOUT : br0_28 
* INOUT : bl1_28 
* INOUT : br1_28 
* INOUT : bl0_29 
* INOUT : br0_29 
* INOUT : bl1_29 
* INOUT : br1_29 
* INOUT : bl0_30 
* INOUT : br0_30 
* INOUT : bl1_30 
* INOUT : br1_30 
* INOUT : bl0_31 
* INOUT : br0_31 
* INOUT : bl1_31 
* INOUT : br1_31 
* INOUT : bl0_32 
* INOUT : br0_32 
* INOUT : bl1_32 
* INOUT : br1_32 
* INOUT : bl0_33 
* INOUT : br0_33 
* INOUT : bl1_33 
* INOUT : br1_33 
* INOUT : bl0_34 
* INOUT : br0_34 
* INOUT : bl1_34 
* INOUT : br1_34 
* INOUT : bl0_35 
* INOUT : br0_35 
* INOUT : bl1_35 
* INOUT : br1_35 
* INOUT : bl0_36 
* INOUT : br0_36 
* INOUT : bl1_36 
* INOUT : br1_36 
* INOUT : bl0_37 
* INOUT : br0_37 
* INOUT : bl1_37 
* INOUT : br1_37 
* INOUT : bl0_38 
* INOUT : br0_38 
* INOUT : bl1_38 
* INOUT : br1_38 
* INOUT : bl0_39 
* INOUT : br0_39 
* INOUT : bl1_39 
* INOUT : br1_39 
* INOUT : bl0_40 
* INOUT : br0_40 
* INOUT : bl1_40 
* INOUT : br1_40 
* INOUT : bl0_41 
* INOUT : br0_41 
* INOUT : bl1_41 
* INOUT : br1_41 
* INOUT : bl0_42 
* INOUT : br0_42 
* INOUT : bl1_42 
* INOUT : br1_42 
* INOUT : bl0_43 
* INOUT : br0_43 
* INOUT : bl1_43 
* INOUT : br1_43 
* INOUT : bl0_44 
* INOUT : br0_44 
* INOUT : bl1_44 
* INOUT : br1_44 
* INOUT : bl0_45 
* INOUT : br0_45 
* INOUT : bl1_45 
* INOUT : br1_45 
* INOUT : bl0_46 
* INOUT : br0_46 
* INOUT : bl1_46 
* INOUT : br1_46 
* INOUT : bl0_47 
* INOUT : br0_47 
* INOUT : bl1_47 
* INOUT : br1_47 
* INOUT : bl0_48 
* INOUT : br0_48 
* INOUT : bl1_48 
* INOUT : br1_48 
* INOUT : bl0_49 
* INOUT : br0_49 
* INOUT : bl1_49 
* INOUT : br1_49 
* INOUT : bl0_50 
* INOUT : br0_50 
* INOUT : bl1_50 
* INOUT : br1_50 
* INOUT : bl0_51 
* INOUT : br0_51 
* INOUT : bl1_51 
* INOUT : br1_51 
* INOUT : bl0_52 
* INOUT : br0_52 
* INOUT : bl1_52 
* INOUT : br1_52 
* INOUT : bl0_53 
* INOUT : br0_53 
* INOUT : bl1_53 
* INOUT : br1_53 
* INOUT : bl0_54 
* INOUT : br0_54 
* INOUT : bl1_54 
* INOUT : br1_54 
* INOUT : bl0_55 
* INOUT : br0_55 
* INOUT : bl1_55 
* INOUT : br1_55 
* INOUT : bl0_56 
* INOUT : br0_56 
* INOUT : bl1_56 
* INOUT : br1_56 
* INOUT : bl0_57 
* INOUT : br0_57 
* INOUT : bl1_57 
* INOUT : br1_57 
* INOUT : bl0_58 
* INOUT : br0_58 
* INOUT : bl1_58 
* INOUT : br1_58 
* INOUT : bl0_59 
* INOUT : br0_59 
* INOUT : bl1_59 
* INOUT : br1_59 
* INOUT : bl0_60 
* INOUT : br0_60 
* INOUT : bl1_60 
* INOUT : br1_60 
* INOUT : bl0_61 
* INOUT : br0_61 
* INOUT : bl1_61 
* INOUT : br1_61 
* INOUT : bl0_62 
* INOUT : br0_62 
* INOUT : bl1_62 
* INOUT : br1_62 
* INOUT : bl0_63 
* INOUT : br0_63 
* INOUT : bl1_63 
* INOUT : br1_63 
* INPUT : wl0_0 
* INPUT : wl1_0 
* INPUT : wl0_1 
* INPUT : wl1_1 
* INPUT : wl0_2 
* INPUT : wl1_2 
* INPUT : wl0_3 
* INPUT : wl1_3 
* INPUT : wl0_4 
* INPUT : wl1_4 
* INPUT : wl0_5 
* INPUT : wl1_5 
* INPUT : wl0_6 
* INPUT : wl1_6 
* INPUT : wl0_7 
* INPUT : wl1_7 
* INPUT : wl0_8 
* INPUT : wl1_8 
* INPUT : wl0_9 
* INPUT : wl1_9 
* INPUT : wl0_10 
* INPUT : wl1_10 
* INPUT : wl0_11 
* INPUT : wl1_11 
* INPUT : wl0_12 
* INPUT : wl1_12 
* INPUT : wl0_13 
* INPUT : wl1_13 
* INPUT : wl0_14 
* INPUT : wl1_14 
* INPUT : wl0_15 
* INPUT : wl1_15 
* INPUT : wl0_16 
* INPUT : wl1_16 
* INPUT : wl0_17 
* INPUT : wl1_17 
* INPUT : wl0_18 
* INPUT : wl1_18 
* INPUT : wl0_19 
* INPUT : wl1_19 
* INPUT : wl0_20 
* INPUT : wl1_20 
* INPUT : wl0_21 
* INPUT : wl1_21 
* INPUT : wl0_22 
* INPUT : wl1_22 
* INPUT : wl0_23 
* INPUT : wl1_23 
* INPUT : wl0_24 
* INPUT : wl1_24 
* INPUT : wl0_25 
* INPUT : wl1_25 
* INPUT : wl0_26 
* INPUT : wl1_26 
* INPUT : wl0_27 
* INPUT : wl1_27 
* INPUT : wl0_28 
* INPUT : wl1_28 
* INPUT : wl0_29 
* INPUT : wl1_29 
* INPUT : wl0_30 
* INPUT : wl1_30 
* INPUT : wl0_31 
* INPUT : wl1_31 
* INPUT : wl0_32 
* INPUT : wl1_32 
* INPUT : wl0_33 
* INPUT : wl1_33 
* INPUT : wl0_34 
* INPUT : wl1_34 
* INPUT : wl0_35 
* INPUT : wl1_35 
* INPUT : wl0_36 
* INPUT : wl1_36 
* INPUT : wl0_37 
* INPUT : wl1_37 
* INPUT : wl0_38 
* INPUT : wl1_38 
* INPUT : wl0_39 
* INPUT : wl1_39 
* INPUT : wl0_40 
* INPUT : wl1_40 
* INPUT : wl0_41 
* INPUT : wl1_41 
* INPUT : wl0_42 
* INPUT : wl1_42 
* INPUT : wl0_43 
* INPUT : wl1_43 
* INPUT : wl0_44 
* INPUT : wl1_44 
* INPUT : wl0_45 
* INPUT : wl1_45 
* INPUT : wl0_46 
* INPUT : wl1_46 
* INPUT : wl0_47 
* INPUT : wl1_47 
* INPUT : wl0_48 
* INPUT : wl1_48 
* INPUT : wl0_49 
* INPUT : wl1_49 
* INPUT : wl0_50 
* INPUT : wl1_50 
* INPUT : wl0_51 
* INPUT : wl1_51 
* INPUT : wl0_52 
* INPUT : wl1_52 
* INPUT : wl0_53 
* INPUT : wl1_53 
* INPUT : wl0_54 
* INPUT : wl1_54 
* INPUT : wl0_55 
* INPUT : wl1_55 
* INPUT : wl0_56 
* INPUT : wl1_56 
* INPUT : wl0_57 
* INPUT : wl1_57 
* INPUT : wl0_58 
* INPUT : wl1_58 
* INPUT : wl0_59 
* INPUT : wl1_59 
* INPUT : wl0_60 
* INPUT : wl1_60 
* INPUT : wl0_61 
* INPUT : wl1_61 
* INPUT : wl0_62 
* INPUT : wl1_62 
* INPUT : wl0_63 
* INPUT : wl1_63 
* INPUT : wl0_64 
* INPUT : wl1_64 
* INPUT : wl0_65 
* INPUT : wl1_65 
* INPUT : wl0_66 
* INPUT : wl1_66 
* INPUT : wl0_67 
* INPUT : wl1_67 
* INPUT : wl0_68 
* INPUT : wl1_68 
* INPUT : wl0_69 
* INPUT : wl1_69 
* INPUT : wl0_70 
* INPUT : wl1_70 
* INPUT : wl0_71 
* INPUT : wl1_71 
* INPUT : wl0_72 
* INPUT : wl1_72 
* INPUT : wl0_73 
* INPUT : wl1_73 
* INPUT : wl0_74 
* INPUT : wl1_74 
* INPUT : wl0_75 
* INPUT : wl1_75 
* INPUT : wl0_76 
* INPUT : wl1_76 
* INPUT : wl0_77 
* INPUT : wl1_77 
* INPUT : wl0_78 
* INPUT : wl1_78 
* INPUT : wl0_79 
* INPUT : wl1_79 
* INPUT : wl0_80 
* INPUT : wl1_80 
* INPUT : wl0_81 
* INPUT : wl1_81 
* INPUT : wl0_82 
* INPUT : wl1_82 
* INPUT : wl0_83 
* INPUT : wl1_83 
* INPUT : wl0_84 
* INPUT : wl1_84 
* INPUT : wl0_85 
* INPUT : wl1_85 
* INPUT : wl0_86 
* INPUT : wl1_86 
* INPUT : wl0_87 
* INPUT : wl1_87 
* INPUT : wl0_88 
* INPUT : wl1_88 
* INPUT : wl0_89 
* INPUT : wl1_89 
* INPUT : wl0_90 
* INPUT : wl1_90 
* INPUT : wl0_91 
* INPUT : wl1_91 
* INPUT : wl0_92 
* INPUT : wl1_92 
* INPUT : wl0_93 
* INPUT : wl1_93 
* INPUT : wl0_94 
* INPUT : wl1_94 
* INPUT : wl0_95 
* INPUT : wl1_95 
* INPUT : wl0_96 
* INPUT : wl1_96 
* INPUT : wl0_97 
* INPUT : wl1_97 
* INPUT : wl0_98 
* INPUT : wl1_98 
* INPUT : wl0_99 
* INPUT : wl1_99 
* INPUT : wl0_100 
* INPUT : wl1_100 
* INPUT : wl0_101 
* INPUT : wl1_101 
* INPUT : wl0_102 
* INPUT : wl1_102 
* INPUT : wl0_103 
* INPUT : wl1_103 
* INPUT : wl0_104 
* INPUT : wl1_104 
* INPUT : wl0_105 
* INPUT : wl1_105 
* INPUT : wl0_106 
* INPUT : wl1_106 
* INPUT : wl0_107 
* INPUT : wl1_107 
* INPUT : wl0_108 
* INPUT : wl1_108 
* INPUT : wl0_109 
* INPUT : wl1_109 
* INPUT : wl0_110 
* INPUT : wl1_110 
* INPUT : wl0_111 
* INPUT : wl1_111 
* INPUT : wl0_112 
* INPUT : wl1_112 
* INPUT : wl0_113 
* INPUT : wl1_113 
* INPUT : wl0_114 
* INPUT : wl1_114 
* INPUT : wl0_115 
* INPUT : wl1_115 
* INPUT : wl0_116 
* INPUT : wl1_116 
* INPUT : wl0_117 
* INPUT : wl1_117 
* INPUT : wl0_118 
* INPUT : wl1_118 
* INPUT : wl0_119 
* INPUT : wl1_119 
* INPUT : wl0_120 
* INPUT : wl1_120 
* INPUT : wl0_121 
* INPUT : wl1_121 
* INPUT : wl0_122 
* INPUT : wl1_122 
* INPUT : wl0_123 
* INPUT : wl1_123 
* INPUT : wl0_124 
* INPUT : wl1_124 
* INPUT : wl0_125 
* INPUT : wl1_125 
* INPUT : wl0_126 
* INPUT : wl1_126 
* INPUT : wl0_127 
* INPUT : wl1_127 
* POWER : vdd 
* GROUND: gnd 
* rows: 128 cols: 64
Xbit_r0_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r0_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r1_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r2_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r3_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r4_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r5_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r6_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r7_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r8_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r9_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r10_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r11_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r12_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r13_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r14_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r15_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r16_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r17_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r18_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r19_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r20_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r21_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r22_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r23_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r24_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r25_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r26_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r27_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r28_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r29_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r30_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r31_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r32_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r33_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r34_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r35_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r36_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r37_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r38_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r39_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r40_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r41_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r42_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r43_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r44_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r45_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r46_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r47_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r48_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r49_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r50_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r51_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r52_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r53_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r54_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r55_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r56_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r57_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r58_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r59_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r60_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r61_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r62_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r63_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r64_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r65_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r66_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r67_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r68_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r69_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r70_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r71_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r72_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r73_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r74_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r75_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r76_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r77_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r78_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r79_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r80_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r81_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r82_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r83_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r84_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r85_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r86_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r87_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r88_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r89_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r90_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r91_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r92_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r93_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r94_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r95_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r96_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r97_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r98_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r99_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r100_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r101_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r102_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r103_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r104_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r105_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r106_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r107_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r108_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r109_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r110_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r111_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r112_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r113_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r114_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r115_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r116_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r117_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r118_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r119_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r120_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r121_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r122_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r123_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r124_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r125_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r126_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell
Xbit_r127_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell
.ENDS bitcell_array

.SUBCKT sky130_fd_bd_sram__openram_dp_cell_replica bl0 br0 bl1 br1 wl0 wl1 vdd gnd
**
*.SEEDPROM

* Bitcell Core
XM0 Q wl1 bl1 gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM1 gnd vdd Q gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM2 gnd vdd Q gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM3 bl0 wl0 Q gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM4 vdd wl1 br1 gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM5 gnd Q vdd gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM6 gnd Q vdd gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM7 br0 wl0 vdd gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM8 vdd Q vdd vdd sky130_fd_pr__special_pfet_pass W=0.14 L=0.15 m=1
XM9 Q vdd vdd vdd sky130_fd_pr__special_pfet_pass W=0.14 L=0.15 m=1

* drainOnly PMOS
XM10 vdd wl1 vdd vdd sky130_fd_pr__special_pfet_pass L=0.08 W=0.14 m=1
XM11 Q wl0 Q vdd sky130_fd_pr__special_pfet_pass L=0.08 W=0.14 m=1

* drainOnly NMOS
XM12 bl1 gnd bl1 gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.08 m=1
XM14 br1 gnd br1 gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.08 m=1

.ENDS

.SUBCKT sky130_fd_bd_sram__openram_dp_cell_dummy bl0 br0 bl1 br1 wl0 wl1 vdd gnd
**
*.SEEDPROM

* Bitcell Core
XM1 1 gnd gnd gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM2 1 wl1 bl1 gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM3 2 gnd gnd gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM4 2 wl1 br1 gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM5 3 gnd gnd gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM6 3 wl0 bl0 gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM7 4 gnd gnd gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1
XM8 4 wl0 br0 gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.15 m=1

* drainOnly NMOS
XM9 bl1 gnd bl1 gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.08 m=1
XM10 br1 gnd br1 gnd sky130_fd_pr__special_nfet_latch W=0.21 L=0.08 m=1

.ENDS

.SUBCKT replica_column bl0_0 br0_0 bl1_0 br1_0 wl0_0 wl1_0 wl0_1 wl1_1 wl0_2 wl1_2 wl0_3 wl1_3 wl0_4 wl1_4 wl0_5 wl1_5 wl0_6 wl1_6 wl0_7 wl1_7 wl0_8 wl1_8 wl0_9 wl1_9 wl0_10 wl1_10 wl0_11 wl1_11 wl0_12 wl1_12 wl0_13 wl1_13 wl0_14 wl1_14 wl0_15 wl1_15 wl0_16 wl1_16 wl0_17 wl1_17 wl0_18 wl1_18 wl0_19 wl1_19 wl0_20 wl1_20 wl0_21 wl1_21 wl0_22 wl1_22 wl0_23 wl1_23 wl0_24 wl1_24 wl0_25 wl1_25 wl0_26 wl1_26 wl0_27 wl1_27 wl0_28 wl1_28 wl0_29 wl1_29 wl0_30 wl1_30 wl0_31 wl1_31 wl0_32 wl1_32 wl0_33 wl1_33 wl0_34 wl1_34 wl0_35 wl1_35 wl0_36 wl1_36 wl0_37 wl1_37 wl0_38 wl1_38 wl0_39 wl1_39 wl0_40 wl1_40 wl0_41 wl1_41 wl0_42 wl1_42 wl0_43 wl1_43 wl0_44 wl1_44 wl0_45 wl1_45 wl0_46 wl1_46 wl0_47 wl1_47 wl0_48 wl1_48 wl0_49 wl1_49 wl0_50 wl1_50 wl0_51 wl1_51 wl0_52 wl1_52 wl0_53 wl1_53 wl0_54 wl1_54 wl0_55 wl1_55 wl0_56 wl1_56 wl0_57 wl1_57 wl0_58 wl1_58 wl0_59 wl1_59 wl0_60 wl1_60 wl0_61 wl1_61 wl0_62 wl1_62 wl0_63 wl1_63 wl0_64 wl1_64 wl0_65 wl1_65 wl0_66 wl1_66 wl0_67 wl1_67 wl0_68 wl1_68 wl0_69 wl1_69 wl0_70 wl1_70 wl0_71 wl1_71 wl0_72 wl1_72 wl0_73 wl1_73 wl0_74 wl1_74 wl0_75 wl1_75 wl0_76 wl1_76 wl0_77 wl1_77 wl0_78 wl1_78 wl0_79 wl1_79 wl0_80 wl1_80 wl0_81 wl1_81 wl0_82 wl1_82 wl0_83 wl1_83 wl0_84 wl1_84 wl0_85 wl1_85 wl0_86 wl1_86 wl0_87 wl1_87 wl0_88 wl1_88 wl0_89 wl1_89 wl0_90 wl1_90 wl0_91 wl1_91 wl0_92 wl1_92 wl0_93 wl1_93 wl0_94 wl1_94 wl0_95 wl1_95 wl0_96 wl1_96 wl0_97 wl1_97 wl0_98 wl1_98 wl0_99 wl1_99 wl0_100 wl1_100 wl0_101 wl1_101 wl0_102 wl1_102 wl0_103 wl1_103 wl0_104 wl1_104 wl0_105 wl1_105 wl0_106 wl1_106 wl0_107 wl1_107 wl0_108 wl1_108 wl0_109 wl1_109 wl0_110 wl1_110 wl0_111 wl1_111 wl0_112 wl1_112 wl0_113 wl1_113 wl0_114 wl1_114 wl0_115 wl1_115 wl0_116 wl1_116 wl0_117 wl1_117 wl0_118 wl1_118 wl0_119 wl1_119 wl0_120 wl1_120 wl0_121 wl1_121 wl0_122 wl1_122 wl0_123 wl1_123 wl0_124 wl1_124 wl0_125 wl1_125 wl0_126 wl1_126 wl0_127 wl1_127 wl0_128 wl1_128 wl0_129 wl1_129 wl0_130 wl1_130 wl0_131 wl1_131 vdd gnd
* OUTPUT: bl0_0 
* OUTPUT: br0_0 
* OUTPUT: bl1_0 
* OUTPUT: br1_0 
* INPUT : wl0_0 
* INPUT : wl1_0 
* INPUT : wl0_1 
* INPUT : wl1_1 
* INPUT : wl0_2 
* INPUT : wl1_2 
* INPUT : wl0_3 
* INPUT : wl1_3 
* INPUT : wl0_4 
* INPUT : wl1_4 
* INPUT : wl0_5 
* INPUT : wl1_5 
* INPUT : wl0_6 
* INPUT : wl1_6 
* INPUT : wl0_7 
* INPUT : wl1_7 
* INPUT : wl0_8 
* INPUT : wl1_8 
* INPUT : wl0_9 
* INPUT : wl1_9 
* INPUT : wl0_10 
* INPUT : wl1_10 
* INPUT : wl0_11 
* INPUT : wl1_11 
* INPUT : wl0_12 
* INPUT : wl1_12 
* INPUT : wl0_13 
* INPUT : wl1_13 
* INPUT : wl0_14 
* INPUT : wl1_14 
* INPUT : wl0_15 
* INPUT : wl1_15 
* INPUT : wl0_16 
* INPUT : wl1_16 
* INPUT : wl0_17 
* INPUT : wl1_17 
* INPUT : wl0_18 
* INPUT : wl1_18 
* INPUT : wl0_19 
* INPUT : wl1_19 
* INPUT : wl0_20 
* INPUT : wl1_20 
* INPUT : wl0_21 
* INPUT : wl1_21 
* INPUT : wl0_22 
* INPUT : wl1_22 
* INPUT : wl0_23 
* INPUT : wl1_23 
* INPUT : wl0_24 
* INPUT : wl1_24 
* INPUT : wl0_25 
* INPUT : wl1_25 
* INPUT : wl0_26 
* INPUT : wl1_26 
* INPUT : wl0_27 
* INPUT : wl1_27 
* INPUT : wl0_28 
* INPUT : wl1_28 
* INPUT : wl0_29 
* INPUT : wl1_29 
* INPUT : wl0_30 
* INPUT : wl1_30 
* INPUT : wl0_31 
* INPUT : wl1_31 
* INPUT : wl0_32 
* INPUT : wl1_32 
* INPUT : wl0_33 
* INPUT : wl1_33 
* INPUT : wl0_34 
* INPUT : wl1_34 
* INPUT : wl0_35 
* INPUT : wl1_35 
* INPUT : wl0_36 
* INPUT : wl1_36 
* INPUT : wl0_37 
* INPUT : wl1_37 
* INPUT : wl0_38 
* INPUT : wl1_38 
* INPUT : wl0_39 
* INPUT : wl1_39 
* INPUT : wl0_40 
* INPUT : wl1_40 
* INPUT : wl0_41 
* INPUT : wl1_41 
* INPUT : wl0_42 
* INPUT : wl1_42 
* INPUT : wl0_43 
* INPUT : wl1_43 
* INPUT : wl0_44 
* INPUT : wl1_44 
* INPUT : wl0_45 
* INPUT : wl1_45 
* INPUT : wl0_46 
* INPUT : wl1_46 
* INPUT : wl0_47 
* INPUT : wl1_47 
* INPUT : wl0_48 
* INPUT : wl1_48 
* INPUT : wl0_49 
* INPUT : wl1_49 
* INPUT : wl0_50 
* INPUT : wl1_50 
* INPUT : wl0_51 
* INPUT : wl1_51 
* INPUT : wl0_52 
* INPUT : wl1_52 
* INPUT : wl0_53 
* INPUT : wl1_53 
* INPUT : wl0_54 
* INPUT : wl1_54 
* INPUT : wl0_55 
* INPUT : wl1_55 
* INPUT : wl0_56 
* INPUT : wl1_56 
* INPUT : wl0_57 
* INPUT : wl1_57 
* INPUT : wl0_58 
* INPUT : wl1_58 
* INPUT : wl0_59 
* INPUT : wl1_59 
* INPUT : wl0_60 
* INPUT : wl1_60 
* INPUT : wl0_61 
* INPUT : wl1_61 
* INPUT : wl0_62 
* INPUT : wl1_62 
* INPUT : wl0_63 
* INPUT : wl1_63 
* INPUT : wl0_64 
* INPUT : wl1_64 
* INPUT : wl0_65 
* INPUT : wl1_65 
* INPUT : wl0_66 
* INPUT : wl1_66 
* INPUT : wl0_67 
* INPUT : wl1_67 
* INPUT : wl0_68 
* INPUT : wl1_68 
* INPUT : wl0_69 
* INPUT : wl1_69 
* INPUT : wl0_70 
* INPUT : wl1_70 
* INPUT : wl0_71 
* INPUT : wl1_71 
* INPUT : wl0_72 
* INPUT : wl1_72 
* INPUT : wl0_73 
* INPUT : wl1_73 
* INPUT : wl0_74 
* INPUT : wl1_74 
* INPUT : wl0_75 
* INPUT : wl1_75 
* INPUT : wl0_76 
* INPUT : wl1_76 
* INPUT : wl0_77 
* INPUT : wl1_77 
* INPUT : wl0_78 
* INPUT : wl1_78 
* INPUT : wl0_79 
* INPUT : wl1_79 
* INPUT : wl0_80 
* INPUT : wl1_80 
* INPUT : wl0_81 
* INPUT : wl1_81 
* INPUT : wl0_82 
* INPUT : wl1_82 
* INPUT : wl0_83 
* INPUT : wl1_83 
* INPUT : wl0_84 
* INPUT : wl1_84 
* INPUT : wl0_85 
* INPUT : wl1_85 
* INPUT : wl0_86 
* INPUT : wl1_86 
* INPUT : wl0_87 
* INPUT : wl1_87 
* INPUT : wl0_88 
* INPUT : wl1_88 
* INPUT : wl0_89 
* INPUT : wl1_89 
* INPUT : wl0_90 
* INPUT : wl1_90 
* INPUT : wl0_91 
* INPUT : wl1_91 
* INPUT : wl0_92 
* INPUT : wl1_92 
* INPUT : wl0_93 
* INPUT : wl1_93 
* INPUT : wl0_94 
* INPUT : wl1_94 
* INPUT : wl0_95 
* INPUT : wl1_95 
* INPUT : wl0_96 
* INPUT : wl1_96 
* INPUT : wl0_97 
* INPUT : wl1_97 
* INPUT : wl0_98 
* INPUT : wl1_98 
* INPUT : wl0_99 
* INPUT : wl1_99 
* INPUT : wl0_100 
* INPUT : wl1_100 
* INPUT : wl0_101 
* INPUT : wl1_101 
* INPUT : wl0_102 
* INPUT : wl1_102 
* INPUT : wl0_103 
* INPUT : wl1_103 
* INPUT : wl0_104 
* INPUT : wl1_104 
* INPUT : wl0_105 
* INPUT : wl1_105 
* INPUT : wl0_106 
* INPUT : wl1_106 
* INPUT : wl0_107 
* INPUT : wl1_107 
* INPUT : wl0_108 
* INPUT : wl1_108 
* INPUT : wl0_109 
* INPUT : wl1_109 
* INPUT : wl0_110 
* INPUT : wl1_110 
* INPUT : wl0_111 
* INPUT : wl1_111 
* INPUT : wl0_112 
* INPUT : wl1_112 
* INPUT : wl0_113 
* INPUT : wl1_113 
* INPUT : wl0_114 
* INPUT : wl1_114 
* INPUT : wl0_115 
* INPUT : wl1_115 
* INPUT : wl0_116 
* INPUT : wl1_116 
* INPUT : wl0_117 
* INPUT : wl1_117 
* INPUT : wl0_118 
* INPUT : wl1_118 
* INPUT : wl0_119 
* INPUT : wl1_119 
* INPUT : wl0_120 
* INPUT : wl1_120 
* INPUT : wl0_121 
* INPUT : wl1_121 
* INPUT : wl0_122 
* INPUT : wl1_122 
* INPUT : wl0_123 
* INPUT : wl1_123 
* INPUT : wl0_124 
* INPUT : wl1_124 
* INPUT : wl0_125 
* INPUT : wl1_125 
* INPUT : wl0_126 
* INPUT : wl1_126 
* INPUT : wl0_127 
* INPUT : wl1_127 
* INPUT : wl0_128 
* INPUT : wl1_128 
* INPUT : wl0_129 
* INPUT : wl1_129 
* INPUT : wl0_130 
* INPUT : wl1_130 
* INPUT : wl0_131 
* INPUT : wl1_131 
* POWER : vdd 
* GROUND: gnd 
Xrbc_1 bl0_0 br0_0 bl1_0 br1_0 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_2 bl0_0 br0_0 bl1_0 br1_0 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_3 bl0_0 br0_0 bl1_0 br1_0 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_4 bl0_0 br0_0 bl1_0 br1_0 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_5 bl0_0 br0_0 bl1_0 br1_0 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_6 bl0_0 br0_0 bl1_0 br1_0 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_7 bl0_0 br0_0 bl1_0 br1_0 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_8 bl0_0 br0_0 bl1_0 br1_0 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_9 bl0_0 br0_0 bl1_0 br1_0 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_10 bl0_0 br0_0 bl1_0 br1_0 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_11 bl0_0 br0_0 bl1_0 br1_0 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_12 bl0_0 br0_0 bl1_0 br1_0 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_13 bl0_0 br0_0 bl1_0 br1_0 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_14 bl0_0 br0_0 bl1_0 br1_0 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_15 bl0_0 br0_0 bl1_0 br1_0 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_16 bl0_0 br0_0 bl1_0 br1_0 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_17 bl0_0 br0_0 bl1_0 br1_0 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_18 bl0_0 br0_0 bl1_0 br1_0 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_19 bl0_0 br0_0 bl1_0 br1_0 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_20 bl0_0 br0_0 bl1_0 br1_0 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_21 bl0_0 br0_0 bl1_0 br1_0 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_22 bl0_0 br0_0 bl1_0 br1_0 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_23 bl0_0 br0_0 bl1_0 br1_0 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_24 bl0_0 br0_0 bl1_0 br1_0 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_25 bl0_0 br0_0 bl1_0 br1_0 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_26 bl0_0 br0_0 bl1_0 br1_0 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_27 bl0_0 br0_0 bl1_0 br1_0 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_28 bl0_0 br0_0 bl1_0 br1_0 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_29 bl0_0 br0_0 bl1_0 br1_0 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_30 bl0_0 br0_0 bl1_0 br1_0 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_31 bl0_0 br0_0 bl1_0 br1_0 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_32 bl0_0 br0_0 bl1_0 br1_0 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_33 bl0_0 br0_0 bl1_0 br1_0 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_34 bl0_0 br0_0 bl1_0 br1_0 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_35 bl0_0 br0_0 bl1_0 br1_0 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_36 bl0_0 br0_0 bl1_0 br1_0 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_37 bl0_0 br0_0 bl1_0 br1_0 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_38 bl0_0 br0_0 bl1_0 br1_0 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_39 bl0_0 br0_0 bl1_0 br1_0 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_40 bl0_0 br0_0 bl1_0 br1_0 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_41 bl0_0 br0_0 bl1_0 br1_0 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_42 bl0_0 br0_0 bl1_0 br1_0 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_43 bl0_0 br0_0 bl1_0 br1_0 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_44 bl0_0 br0_0 bl1_0 br1_0 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_45 bl0_0 br0_0 bl1_0 br1_0 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_46 bl0_0 br0_0 bl1_0 br1_0 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_47 bl0_0 br0_0 bl1_0 br1_0 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_48 bl0_0 br0_0 bl1_0 br1_0 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_49 bl0_0 br0_0 bl1_0 br1_0 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_50 bl0_0 br0_0 bl1_0 br1_0 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_51 bl0_0 br0_0 bl1_0 br1_0 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_52 bl0_0 br0_0 bl1_0 br1_0 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_53 bl0_0 br0_0 bl1_0 br1_0 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_54 bl0_0 br0_0 bl1_0 br1_0 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_55 bl0_0 br0_0 bl1_0 br1_0 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_56 bl0_0 br0_0 bl1_0 br1_0 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_57 bl0_0 br0_0 bl1_0 br1_0 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_58 bl0_0 br0_0 bl1_0 br1_0 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_59 bl0_0 br0_0 bl1_0 br1_0 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_60 bl0_0 br0_0 bl1_0 br1_0 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_61 bl0_0 br0_0 bl1_0 br1_0 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_62 bl0_0 br0_0 bl1_0 br1_0 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_63 bl0_0 br0_0 bl1_0 br1_0 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_64 bl0_0 br0_0 bl1_0 br1_0 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_65 bl0_0 br0_0 bl1_0 br1_0 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_66 bl0_0 br0_0 bl1_0 br1_0 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_67 bl0_0 br0_0 bl1_0 br1_0 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_68 bl0_0 br0_0 bl1_0 br1_0 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_69 bl0_0 br0_0 bl1_0 br1_0 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_70 bl0_0 br0_0 bl1_0 br1_0 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_71 bl0_0 br0_0 bl1_0 br1_0 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_72 bl0_0 br0_0 bl1_0 br1_0 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_73 bl0_0 br0_0 bl1_0 br1_0 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_74 bl0_0 br0_0 bl1_0 br1_0 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_75 bl0_0 br0_0 bl1_0 br1_0 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_76 bl0_0 br0_0 bl1_0 br1_0 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_77 bl0_0 br0_0 bl1_0 br1_0 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_78 bl0_0 br0_0 bl1_0 br1_0 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_79 bl0_0 br0_0 bl1_0 br1_0 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_80 bl0_0 br0_0 bl1_0 br1_0 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_81 bl0_0 br0_0 bl1_0 br1_0 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_82 bl0_0 br0_0 bl1_0 br1_0 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_83 bl0_0 br0_0 bl1_0 br1_0 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_84 bl0_0 br0_0 bl1_0 br1_0 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_85 bl0_0 br0_0 bl1_0 br1_0 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_86 bl0_0 br0_0 bl1_0 br1_0 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_87 bl0_0 br0_0 bl1_0 br1_0 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_88 bl0_0 br0_0 bl1_0 br1_0 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_89 bl0_0 br0_0 bl1_0 br1_0 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_90 bl0_0 br0_0 bl1_0 br1_0 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_91 bl0_0 br0_0 bl1_0 br1_0 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_92 bl0_0 br0_0 bl1_0 br1_0 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_93 bl0_0 br0_0 bl1_0 br1_0 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_94 bl0_0 br0_0 bl1_0 br1_0 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_95 bl0_0 br0_0 bl1_0 br1_0 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_96 bl0_0 br0_0 bl1_0 br1_0 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_97 bl0_0 br0_0 bl1_0 br1_0 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_98 bl0_0 br0_0 bl1_0 br1_0 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_99 bl0_0 br0_0 bl1_0 br1_0 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_100 bl0_0 br0_0 bl1_0 br1_0 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_101 bl0_0 br0_0 bl1_0 br1_0 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_102 bl0_0 br0_0 bl1_0 br1_0 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_103 bl0_0 br0_0 bl1_0 br1_0 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_104 bl0_0 br0_0 bl1_0 br1_0 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_105 bl0_0 br0_0 bl1_0 br1_0 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_106 bl0_0 br0_0 bl1_0 br1_0 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_107 bl0_0 br0_0 bl1_0 br1_0 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_108 bl0_0 br0_0 bl1_0 br1_0 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_109 bl0_0 br0_0 bl1_0 br1_0 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_110 bl0_0 br0_0 bl1_0 br1_0 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_111 bl0_0 br0_0 bl1_0 br1_0 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_112 bl0_0 br0_0 bl1_0 br1_0 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_113 bl0_0 br0_0 bl1_0 br1_0 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_114 bl0_0 br0_0 bl1_0 br1_0 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_115 bl0_0 br0_0 bl1_0 br1_0 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_116 bl0_0 br0_0 bl1_0 br1_0 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_117 bl0_0 br0_0 bl1_0 br1_0 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_118 bl0_0 br0_0 bl1_0 br1_0 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_119 bl0_0 br0_0 bl1_0 br1_0 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_120 bl0_0 br0_0 bl1_0 br1_0 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_121 bl0_0 br0_0 bl1_0 br1_0 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_122 bl0_0 br0_0 bl1_0 br1_0 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_123 bl0_0 br0_0 bl1_0 br1_0 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_124 bl0_0 br0_0 bl1_0 br1_0 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_125 bl0_0 br0_0 bl1_0 br1_0 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_126 bl0_0 br0_0 bl1_0 br1_0 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_127 bl0_0 br0_0 bl1_0 br1_0 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_128 bl0_0 br0_0 bl1_0 br1_0 wl0_128 wl1_128 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_129 bl0_0 br0_0 bl1_0 br1_0 wl0_129 wl1_129 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_130 bl0_0 br0_0 bl1_0 br1_0 wl0_130 wl1_130 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
.ENDS replica_column

.SUBCKT replica_column_0 bl0_0 br0_0 bl1_0 br1_0 wl0_0 wl1_0 wl0_1 wl1_1 wl0_2 wl1_2 wl0_3 wl1_3 wl0_4 wl1_4 wl0_5 wl1_5 wl0_6 wl1_6 wl0_7 wl1_7 wl0_8 wl1_8 wl0_9 wl1_9 wl0_10 wl1_10 wl0_11 wl1_11 wl0_12 wl1_12 wl0_13 wl1_13 wl0_14 wl1_14 wl0_15 wl1_15 wl0_16 wl1_16 wl0_17 wl1_17 wl0_18 wl1_18 wl0_19 wl1_19 wl0_20 wl1_20 wl0_21 wl1_21 wl0_22 wl1_22 wl0_23 wl1_23 wl0_24 wl1_24 wl0_25 wl1_25 wl0_26 wl1_26 wl0_27 wl1_27 wl0_28 wl1_28 wl0_29 wl1_29 wl0_30 wl1_30 wl0_31 wl1_31 wl0_32 wl1_32 wl0_33 wl1_33 wl0_34 wl1_34 wl0_35 wl1_35 wl0_36 wl1_36 wl0_37 wl1_37 wl0_38 wl1_38 wl0_39 wl1_39 wl0_40 wl1_40 wl0_41 wl1_41 wl0_42 wl1_42 wl0_43 wl1_43 wl0_44 wl1_44 wl0_45 wl1_45 wl0_46 wl1_46 wl0_47 wl1_47 wl0_48 wl1_48 wl0_49 wl1_49 wl0_50 wl1_50 wl0_51 wl1_51 wl0_52 wl1_52 wl0_53 wl1_53 wl0_54 wl1_54 wl0_55 wl1_55 wl0_56 wl1_56 wl0_57 wl1_57 wl0_58 wl1_58 wl0_59 wl1_59 wl0_60 wl1_60 wl0_61 wl1_61 wl0_62 wl1_62 wl0_63 wl1_63 wl0_64 wl1_64 wl0_65 wl1_65 wl0_66 wl1_66 wl0_67 wl1_67 wl0_68 wl1_68 wl0_69 wl1_69 wl0_70 wl1_70 wl0_71 wl1_71 wl0_72 wl1_72 wl0_73 wl1_73 wl0_74 wl1_74 wl0_75 wl1_75 wl0_76 wl1_76 wl0_77 wl1_77 wl0_78 wl1_78 wl0_79 wl1_79 wl0_80 wl1_80 wl0_81 wl1_81 wl0_82 wl1_82 wl0_83 wl1_83 wl0_84 wl1_84 wl0_85 wl1_85 wl0_86 wl1_86 wl0_87 wl1_87 wl0_88 wl1_88 wl0_89 wl1_89 wl0_90 wl1_90 wl0_91 wl1_91 wl0_92 wl1_92 wl0_93 wl1_93 wl0_94 wl1_94 wl0_95 wl1_95 wl0_96 wl1_96 wl0_97 wl1_97 wl0_98 wl1_98 wl0_99 wl1_99 wl0_100 wl1_100 wl0_101 wl1_101 wl0_102 wl1_102 wl0_103 wl1_103 wl0_104 wl1_104 wl0_105 wl1_105 wl0_106 wl1_106 wl0_107 wl1_107 wl0_108 wl1_108 wl0_109 wl1_109 wl0_110 wl1_110 wl0_111 wl1_111 wl0_112 wl1_112 wl0_113 wl1_113 wl0_114 wl1_114 wl0_115 wl1_115 wl0_116 wl1_116 wl0_117 wl1_117 wl0_118 wl1_118 wl0_119 wl1_119 wl0_120 wl1_120 wl0_121 wl1_121 wl0_122 wl1_122 wl0_123 wl1_123 wl0_124 wl1_124 wl0_125 wl1_125 wl0_126 wl1_126 wl0_127 wl1_127 wl0_128 wl1_128 wl0_129 wl1_129 wl0_130 wl1_130 wl0_131 wl1_131 vdd gnd
* OUTPUT: bl0_0 
* OUTPUT: br0_0 
* OUTPUT: bl1_0 
* OUTPUT: br1_0 
* INPUT : wl0_0 
* INPUT : wl1_0 
* INPUT : wl0_1 
* INPUT : wl1_1 
* INPUT : wl0_2 
* INPUT : wl1_2 
* INPUT : wl0_3 
* INPUT : wl1_3 
* INPUT : wl0_4 
* INPUT : wl1_4 
* INPUT : wl0_5 
* INPUT : wl1_5 
* INPUT : wl0_6 
* INPUT : wl1_6 
* INPUT : wl0_7 
* INPUT : wl1_7 
* INPUT : wl0_8 
* INPUT : wl1_8 
* INPUT : wl0_9 
* INPUT : wl1_9 
* INPUT : wl0_10 
* INPUT : wl1_10 
* INPUT : wl0_11 
* INPUT : wl1_11 
* INPUT : wl0_12 
* INPUT : wl1_12 
* INPUT : wl0_13 
* INPUT : wl1_13 
* INPUT : wl0_14 
* INPUT : wl1_14 
* INPUT : wl0_15 
* INPUT : wl1_15 
* INPUT : wl0_16 
* INPUT : wl1_16 
* INPUT : wl0_17 
* INPUT : wl1_17 
* INPUT : wl0_18 
* INPUT : wl1_18 
* INPUT : wl0_19 
* INPUT : wl1_19 
* INPUT : wl0_20 
* INPUT : wl1_20 
* INPUT : wl0_21 
* INPUT : wl1_21 
* INPUT : wl0_22 
* INPUT : wl1_22 
* INPUT : wl0_23 
* INPUT : wl1_23 
* INPUT : wl0_24 
* INPUT : wl1_24 
* INPUT : wl0_25 
* INPUT : wl1_25 
* INPUT : wl0_26 
* INPUT : wl1_26 
* INPUT : wl0_27 
* INPUT : wl1_27 
* INPUT : wl0_28 
* INPUT : wl1_28 
* INPUT : wl0_29 
* INPUT : wl1_29 
* INPUT : wl0_30 
* INPUT : wl1_30 
* INPUT : wl0_31 
* INPUT : wl1_31 
* INPUT : wl0_32 
* INPUT : wl1_32 
* INPUT : wl0_33 
* INPUT : wl1_33 
* INPUT : wl0_34 
* INPUT : wl1_34 
* INPUT : wl0_35 
* INPUT : wl1_35 
* INPUT : wl0_36 
* INPUT : wl1_36 
* INPUT : wl0_37 
* INPUT : wl1_37 
* INPUT : wl0_38 
* INPUT : wl1_38 
* INPUT : wl0_39 
* INPUT : wl1_39 
* INPUT : wl0_40 
* INPUT : wl1_40 
* INPUT : wl0_41 
* INPUT : wl1_41 
* INPUT : wl0_42 
* INPUT : wl1_42 
* INPUT : wl0_43 
* INPUT : wl1_43 
* INPUT : wl0_44 
* INPUT : wl1_44 
* INPUT : wl0_45 
* INPUT : wl1_45 
* INPUT : wl0_46 
* INPUT : wl1_46 
* INPUT : wl0_47 
* INPUT : wl1_47 
* INPUT : wl0_48 
* INPUT : wl1_48 
* INPUT : wl0_49 
* INPUT : wl1_49 
* INPUT : wl0_50 
* INPUT : wl1_50 
* INPUT : wl0_51 
* INPUT : wl1_51 
* INPUT : wl0_52 
* INPUT : wl1_52 
* INPUT : wl0_53 
* INPUT : wl1_53 
* INPUT : wl0_54 
* INPUT : wl1_54 
* INPUT : wl0_55 
* INPUT : wl1_55 
* INPUT : wl0_56 
* INPUT : wl1_56 
* INPUT : wl0_57 
* INPUT : wl1_57 
* INPUT : wl0_58 
* INPUT : wl1_58 
* INPUT : wl0_59 
* INPUT : wl1_59 
* INPUT : wl0_60 
* INPUT : wl1_60 
* INPUT : wl0_61 
* INPUT : wl1_61 
* INPUT : wl0_62 
* INPUT : wl1_62 
* INPUT : wl0_63 
* INPUT : wl1_63 
* INPUT : wl0_64 
* INPUT : wl1_64 
* INPUT : wl0_65 
* INPUT : wl1_65 
* INPUT : wl0_66 
* INPUT : wl1_66 
* INPUT : wl0_67 
* INPUT : wl1_67 
* INPUT : wl0_68 
* INPUT : wl1_68 
* INPUT : wl0_69 
* INPUT : wl1_69 
* INPUT : wl0_70 
* INPUT : wl1_70 
* INPUT : wl0_71 
* INPUT : wl1_71 
* INPUT : wl0_72 
* INPUT : wl1_72 
* INPUT : wl0_73 
* INPUT : wl1_73 
* INPUT : wl0_74 
* INPUT : wl1_74 
* INPUT : wl0_75 
* INPUT : wl1_75 
* INPUT : wl0_76 
* INPUT : wl1_76 
* INPUT : wl0_77 
* INPUT : wl1_77 
* INPUT : wl0_78 
* INPUT : wl1_78 
* INPUT : wl0_79 
* INPUT : wl1_79 
* INPUT : wl0_80 
* INPUT : wl1_80 
* INPUT : wl0_81 
* INPUT : wl1_81 
* INPUT : wl0_82 
* INPUT : wl1_82 
* INPUT : wl0_83 
* INPUT : wl1_83 
* INPUT : wl0_84 
* INPUT : wl1_84 
* INPUT : wl0_85 
* INPUT : wl1_85 
* INPUT : wl0_86 
* INPUT : wl1_86 
* INPUT : wl0_87 
* INPUT : wl1_87 
* INPUT : wl0_88 
* INPUT : wl1_88 
* INPUT : wl0_89 
* INPUT : wl1_89 
* INPUT : wl0_90 
* INPUT : wl1_90 
* INPUT : wl0_91 
* INPUT : wl1_91 
* INPUT : wl0_92 
* INPUT : wl1_92 
* INPUT : wl0_93 
* INPUT : wl1_93 
* INPUT : wl0_94 
* INPUT : wl1_94 
* INPUT : wl0_95 
* INPUT : wl1_95 
* INPUT : wl0_96 
* INPUT : wl1_96 
* INPUT : wl0_97 
* INPUT : wl1_97 
* INPUT : wl0_98 
* INPUT : wl1_98 
* INPUT : wl0_99 
* INPUT : wl1_99 
* INPUT : wl0_100 
* INPUT : wl1_100 
* INPUT : wl0_101 
* INPUT : wl1_101 
* INPUT : wl0_102 
* INPUT : wl1_102 
* INPUT : wl0_103 
* INPUT : wl1_103 
* INPUT : wl0_104 
* INPUT : wl1_104 
* INPUT : wl0_105 
* INPUT : wl1_105 
* INPUT : wl0_106 
* INPUT : wl1_106 
* INPUT : wl0_107 
* INPUT : wl1_107 
* INPUT : wl0_108 
* INPUT : wl1_108 
* INPUT : wl0_109 
* INPUT : wl1_109 
* INPUT : wl0_110 
* INPUT : wl1_110 
* INPUT : wl0_111 
* INPUT : wl1_111 
* INPUT : wl0_112 
* INPUT : wl1_112 
* INPUT : wl0_113 
* INPUT : wl1_113 
* INPUT : wl0_114 
* INPUT : wl1_114 
* INPUT : wl0_115 
* INPUT : wl1_115 
* INPUT : wl0_116 
* INPUT : wl1_116 
* INPUT : wl0_117 
* INPUT : wl1_117 
* INPUT : wl0_118 
* INPUT : wl1_118 
* INPUT : wl0_119 
* INPUT : wl1_119 
* INPUT : wl0_120 
* INPUT : wl1_120 
* INPUT : wl0_121 
* INPUT : wl1_121 
* INPUT : wl0_122 
* INPUT : wl1_122 
* INPUT : wl0_123 
* INPUT : wl1_123 
* INPUT : wl0_124 
* INPUT : wl1_124 
* INPUT : wl0_125 
* INPUT : wl1_125 
* INPUT : wl0_126 
* INPUT : wl1_126 
* INPUT : wl0_127 
* INPUT : wl1_127 
* INPUT : wl0_128 
* INPUT : wl1_128 
* INPUT : wl0_129 
* INPUT : wl1_129 
* INPUT : wl0_130 
* INPUT : wl1_130 
* INPUT : wl0_131 
* INPUT : wl1_131 
* POWER : vdd 
* GROUND: gnd 
Xrbc_1 bl0_0 br0_0 bl1_0 br1_0 wl0_1 wl1_1 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xrbc_2 bl0_0 br0_0 bl1_0 br1_0 wl0_2 wl1_2 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_3 bl0_0 br0_0 bl1_0 br1_0 wl0_3 wl1_3 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_4 bl0_0 br0_0 bl1_0 br1_0 wl0_4 wl1_4 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_5 bl0_0 br0_0 bl1_0 br1_0 wl0_5 wl1_5 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_6 bl0_0 br0_0 bl1_0 br1_0 wl0_6 wl1_6 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_7 bl0_0 br0_0 bl1_0 br1_0 wl0_7 wl1_7 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_8 bl0_0 br0_0 bl1_0 br1_0 wl0_8 wl1_8 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_9 bl0_0 br0_0 bl1_0 br1_0 wl0_9 wl1_9 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_10 bl0_0 br0_0 bl1_0 br1_0 wl0_10 wl1_10 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_11 bl0_0 br0_0 bl1_0 br1_0 wl0_11 wl1_11 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_12 bl0_0 br0_0 bl1_0 br1_0 wl0_12 wl1_12 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_13 bl0_0 br0_0 bl1_0 br1_0 wl0_13 wl1_13 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_14 bl0_0 br0_0 bl1_0 br1_0 wl0_14 wl1_14 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_15 bl0_0 br0_0 bl1_0 br1_0 wl0_15 wl1_15 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_16 bl0_0 br0_0 bl1_0 br1_0 wl0_16 wl1_16 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_17 bl0_0 br0_0 bl1_0 br1_0 wl0_17 wl1_17 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_18 bl0_0 br0_0 bl1_0 br1_0 wl0_18 wl1_18 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_19 bl0_0 br0_0 bl1_0 br1_0 wl0_19 wl1_19 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_20 bl0_0 br0_0 bl1_0 br1_0 wl0_20 wl1_20 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_21 bl0_0 br0_0 bl1_0 br1_0 wl0_21 wl1_21 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_22 bl0_0 br0_0 bl1_0 br1_0 wl0_22 wl1_22 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_23 bl0_0 br0_0 bl1_0 br1_0 wl0_23 wl1_23 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_24 bl0_0 br0_0 bl1_0 br1_0 wl0_24 wl1_24 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_25 bl0_0 br0_0 bl1_0 br1_0 wl0_25 wl1_25 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_26 bl0_0 br0_0 bl1_0 br1_0 wl0_26 wl1_26 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_27 bl0_0 br0_0 bl1_0 br1_0 wl0_27 wl1_27 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_28 bl0_0 br0_0 bl1_0 br1_0 wl0_28 wl1_28 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_29 bl0_0 br0_0 bl1_0 br1_0 wl0_29 wl1_29 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_30 bl0_0 br0_0 bl1_0 br1_0 wl0_30 wl1_30 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_31 bl0_0 br0_0 bl1_0 br1_0 wl0_31 wl1_31 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_32 bl0_0 br0_0 bl1_0 br1_0 wl0_32 wl1_32 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_33 bl0_0 br0_0 bl1_0 br1_0 wl0_33 wl1_33 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_34 bl0_0 br0_0 bl1_0 br1_0 wl0_34 wl1_34 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_35 bl0_0 br0_0 bl1_0 br1_0 wl0_35 wl1_35 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_36 bl0_0 br0_0 bl1_0 br1_0 wl0_36 wl1_36 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_37 bl0_0 br0_0 bl1_0 br1_0 wl0_37 wl1_37 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_38 bl0_0 br0_0 bl1_0 br1_0 wl0_38 wl1_38 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_39 bl0_0 br0_0 bl1_0 br1_0 wl0_39 wl1_39 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_40 bl0_0 br0_0 bl1_0 br1_0 wl0_40 wl1_40 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_41 bl0_0 br0_0 bl1_0 br1_0 wl0_41 wl1_41 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_42 bl0_0 br0_0 bl1_0 br1_0 wl0_42 wl1_42 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_43 bl0_0 br0_0 bl1_0 br1_0 wl0_43 wl1_43 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_44 bl0_0 br0_0 bl1_0 br1_0 wl0_44 wl1_44 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_45 bl0_0 br0_0 bl1_0 br1_0 wl0_45 wl1_45 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_46 bl0_0 br0_0 bl1_0 br1_0 wl0_46 wl1_46 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_47 bl0_0 br0_0 bl1_0 br1_0 wl0_47 wl1_47 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_48 bl0_0 br0_0 bl1_0 br1_0 wl0_48 wl1_48 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_49 bl0_0 br0_0 bl1_0 br1_0 wl0_49 wl1_49 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_50 bl0_0 br0_0 bl1_0 br1_0 wl0_50 wl1_50 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_51 bl0_0 br0_0 bl1_0 br1_0 wl0_51 wl1_51 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_52 bl0_0 br0_0 bl1_0 br1_0 wl0_52 wl1_52 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_53 bl0_0 br0_0 bl1_0 br1_0 wl0_53 wl1_53 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_54 bl0_0 br0_0 bl1_0 br1_0 wl0_54 wl1_54 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_55 bl0_0 br0_0 bl1_0 br1_0 wl0_55 wl1_55 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_56 bl0_0 br0_0 bl1_0 br1_0 wl0_56 wl1_56 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_57 bl0_0 br0_0 bl1_0 br1_0 wl0_57 wl1_57 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_58 bl0_0 br0_0 bl1_0 br1_0 wl0_58 wl1_58 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_59 bl0_0 br0_0 bl1_0 br1_0 wl0_59 wl1_59 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_60 bl0_0 br0_0 bl1_0 br1_0 wl0_60 wl1_60 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_61 bl0_0 br0_0 bl1_0 br1_0 wl0_61 wl1_61 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_62 bl0_0 br0_0 bl1_0 br1_0 wl0_62 wl1_62 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_63 bl0_0 br0_0 bl1_0 br1_0 wl0_63 wl1_63 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_64 bl0_0 br0_0 bl1_0 br1_0 wl0_64 wl1_64 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_65 bl0_0 br0_0 bl1_0 br1_0 wl0_65 wl1_65 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_66 bl0_0 br0_0 bl1_0 br1_0 wl0_66 wl1_66 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_67 bl0_0 br0_0 bl1_0 br1_0 wl0_67 wl1_67 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_68 bl0_0 br0_0 bl1_0 br1_0 wl0_68 wl1_68 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_69 bl0_0 br0_0 bl1_0 br1_0 wl0_69 wl1_69 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_70 bl0_0 br0_0 bl1_0 br1_0 wl0_70 wl1_70 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_71 bl0_0 br0_0 bl1_0 br1_0 wl0_71 wl1_71 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_72 bl0_0 br0_0 bl1_0 br1_0 wl0_72 wl1_72 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_73 bl0_0 br0_0 bl1_0 br1_0 wl0_73 wl1_73 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_74 bl0_0 br0_0 bl1_0 br1_0 wl0_74 wl1_74 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_75 bl0_0 br0_0 bl1_0 br1_0 wl0_75 wl1_75 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_76 bl0_0 br0_0 bl1_0 br1_0 wl0_76 wl1_76 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_77 bl0_0 br0_0 bl1_0 br1_0 wl0_77 wl1_77 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_78 bl0_0 br0_0 bl1_0 br1_0 wl0_78 wl1_78 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_79 bl0_0 br0_0 bl1_0 br1_0 wl0_79 wl1_79 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_80 bl0_0 br0_0 bl1_0 br1_0 wl0_80 wl1_80 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_81 bl0_0 br0_0 bl1_0 br1_0 wl0_81 wl1_81 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_82 bl0_0 br0_0 bl1_0 br1_0 wl0_82 wl1_82 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_83 bl0_0 br0_0 bl1_0 br1_0 wl0_83 wl1_83 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_84 bl0_0 br0_0 bl1_0 br1_0 wl0_84 wl1_84 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_85 bl0_0 br0_0 bl1_0 br1_0 wl0_85 wl1_85 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_86 bl0_0 br0_0 bl1_0 br1_0 wl0_86 wl1_86 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_87 bl0_0 br0_0 bl1_0 br1_0 wl0_87 wl1_87 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_88 bl0_0 br0_0 bl1_0 br1_0 wl0_88 wl1_88 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_89 bl0_0 br0_0 bl1_0 br1_0 wl0_89 wl1_89 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_90 bl0_0 br0_0 bl1_0 br1_0 wl0_90 wl1_90 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_91 bl0_0 br0_0 bl1_0 br1_0 wl0_91 wl1_91 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_92 bl0_0 br0_0 bl1_0 br1_0 wl0_92 wl1_92 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_93 bl0_0 br0_0 bl1_0 br1_0 wl0_93 wl1_93 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_94 bl0_0 br0_0 bl1_0 br1_0 wl0_94 wl1_94 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_95 bl0_0 br0_0 bl1_0 br1_0 wl0_95 wl1_95 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_96 bl0_0 br0_0 bl1_0 br1_0 wl0_96 wl1_96 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_97 bl0_0 br0_0 bl1_0 br1_0 wl0_97 wl1_97 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_98 bl0_0 br0_0 bl1_0 br1_0 wl0_98 wl1_98 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_99 bl0_0 br0_0 bl1_0 br1_0 wl0_99 wl1_99 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_100 bl0_0 br0_0 bl1_0 br1_0 wl0_100 wl1_100 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_101 bl0_0 br0_0 bl1_0 br1_0 wl0_101 wl1_101 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_102 bl0_0 br0_0 bl1_0 br1_0 wl0_102 wl1_102 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_103 bl0_0 br0_0 bl1_0 br1_0 wl0_103 wl1_103 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_104 bl0_0 br0_0 bl1_0 br1_0 wl0_104 wl1_104 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_105 bl0_0 br0_0 bl1_0 br1_0 wl0_105 wl1_105 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_106 bl0_0 br0_0 bl1_0 br1_0 wl0_106 wl1_106 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_107 bl0_0 br0_0 bl1_0 br1_0 wl0_107 wl1_107 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_108 bl0_0 br0_0 bl1_0 br1_0 wl0_108 wl1_108 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_109 bl0_0 br0_0 bl1_0 br1_0 wl0_109 wl1_109 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_110 bl0_0 br0_0 bl1_0 br1_0 wl0_110 wl1_110 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_111 bl0_0 br0_0 bl1_0 br1_0 wl0_111 wl1_111 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_112 bl0_0 br0_0 bl1_0 br1_0 wl0_112 wl1_112 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_113 bl0_0 br0_0 bl1_0 br1_0 wl0_113 wl1_113 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_114 bl0_0 br0_0 bl1_0 br1_0 wl0_114 wl1_114 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_115 bl0_0 br0_0 bl1_0 br1_0 wl0_115 wl1_115 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_116 bl0_0 br0_0 bl1_0 br1_0 wl0_116 wl1_116 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_117 bl0_0 br0_0 bl1_0 br1_0 wl0_117 wl1_117 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_118 bl0_0 br0_0 bl1_0 br1_0 wl0_118 wl1_118 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_119 bl0_0 br0_0 bl1_0 br1_0 wl0_119 wl1_119 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_120 bl0_0 br0_0 bl1_0 br1_0 wl0_120 wl1_120 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_121 bl0_0 br0_0 bl1_0 br1_0 wl0_121 wl1_121 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_122 bl0_0 br0_0 bl1_0 br1_0 wl0_122 wl1_122 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_123 bl0_0 br0_0 bl1_0 br1_0 wl0_123 wl1_123 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_124 bl0_0 br0_0 bl1_0 br1_0 wl0_124 wl1_124 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_125 bl0_0 br0_0 bl1_0 br1_0 wl0_125 wl1_125 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_126 bl0_0 br0_0 bl1_0 br1_0 wl0_126 wl1_126 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_127 bl0_0 br0_0 bl1_0 br1_0 wl0_127 wl1_127 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_128 bl0_0 br0_0 bl1_0 br1_0 wl0_128 wl1_128 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_129 bl0_0 br0_0 bl1_0 br1_0 wl0_129 wl1_129 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
Xrbc_130 bl0_0 br0_0 bl1_0 br1_0 wl0_130 wl1_130 vdd gnd sky130_fd_bd_sram__openram_dp_cell_replica
.ENDS replica_column_0

.SUBCKT dummy_array bl0_0 br0_0 bl1_0 br1_0 bl0_1 br0_1 bl1_1 br1_1 bl0_2 br0_2 bl1_2 br1_2 bl0_3 br0_3 bl1_3 br1_3 bl0_4 br0_4 bl1_4 br1_4 bl0_5 br0_5 bl1_5 br1_5 bl0_6 br0_6 bl1_6 br1_6 bl0_7 br0_7 bl1_7 br1_7 bl0_8 br0_8 bl1_8 br1_8 bl0_9 br0_9 bl1_9 br1_9 bl0_10 br0_10 bl1_10 br1_10 bl0_11 br0_11 bl1_11 br1_11 bl0_12 br0_12 bl1_12 br1_12 bl0_13 br0_13 bl1_13 br1_13 bl0_14 br0_14 bl1_14 br1_14 bl0_15 br0_15 bl1_15 br1_15 bl0_16 br0_16 bl1_16 br1_16 bl0_17 br0_17 bl1_17 br1_17 bl0_18 br0_18 bl1_18 br1_18 bl0_19 br0_19 bl1_19 br1_19 bl0_20 br0_20 bl1_20 br1_20 bl0_21 br0_21 bl1_21 br1_21 bl0_22 br0_22 bl1_22 br1_22 bl0_23 br0_23 bl1_23 br1_23 bl0_24 br0_24 bl1_24 br1_24 bl0_25 br0_25 bl1_25 br1_25 bl0_26 br0_26 bl1_26 br1_26 bl0_27 br0_27 bl1_27 br1_27 bl0_28 br0_28 bl1_28 br1_28 bl0_29 br0_29 bl1_29 br1_29 bl0_30 br0_30 bl1_30 br1_30 bl0_31 br0_31 bl1_31 br1_31 bl0_32 br0_32 bl1_32 br1_32 bl0_33 br0_33 bl1_33 br1_33 bl0_34 br0_34 bl1_34 br1_34 bl0_35 br0_35 bl1_35 br1_35 bl0_36 br0_36 bl1_36 br1_36 bl0_37 br0_37 bl1_37 br1_37 bl0_38 br0_38 bl1_38 br1_38 bl0_39 br0_39 bl1_39 br1_39 bl0_40 br0_40 bl1_40 br1_40 bl0_41 br0_41 bl1_41 br1_41 bl0_42 br0_42 bl1_42 br1_42 bl0_43 br0_43 bl1_43 br1_43 bl0_44 br0_44 bl1_44 br1_44 bl0_45 br0_45 bl1_45 br1_45 bl0_46 br0_46 bl1_46 br1_46 bl0_47 br0_47 bl1_47 br1_47 bl0_48 br0_48 bl1_48 br1_48 bl0_49 br0_49 bl1_49 br1_49 bl0_50 br0_50 bl1_50 br1_50 bl0_51 br0_51 bl1_51 br1_51 bl0_52 br0_52 bl1_52 br1_52 bl0_53 br0_53 bl1_53 br1_53 bl0_54 br0_54 bl1_54 br1_54 bl0_55 br0_55 bl1_55 br1_55 bl0_56 br0_56 bl1_56 br1_56 bl0_57 br0_57 bl1_57 br1_57 bl0_58 br0_58 bl1_58 br1_58 bl0_59 br0_59 bl1_59 br1_59 bl0_60 br0_60 bl1_60 br1_60 bl0_61 br0_61 bl1_61 br1_61 bl0_62 br0_62 bl1_62 br1_62 bl0_63 br0_63 bl1_63 br1_63 wl0_0 wl1_0 vdd gnd
* INOUT : bl0_0 
* INOUT : br0_0 
* INOUT : bl1_0 
* INOUT : br1_0 
* INOUT : bl0_1 
* INOUT : br0_1 
* INOUT : bl1_1 
* INOUT : br1_1 
* INOUT : bl0_2 
* INOUT : br0_2 
* INOUT : bl1_2 
* INOUT : br1_2 
* INOUT : bl0_3 
* INOUT : br0_3 
* INOUT : bl1_3 
* INOUT : br1_3 
* INOUT : bl0_4 
* INOUT : br0_4 
* INOUT : bl1_4 
* INOUT : br1_4 
* INOUT : bl0_5 
* INOUT : br0_5 
* INOUT : bl1_5 
* INOUT : br1_5 
* INOUT : bl0_6 
* INOUT : br0_6 
* INOUT : bl1_6 
* INOUT : br1_6 
* INOUT : bl0_7 
* INOUT : br0_7 
* INOUT : bl1_7 
* INOUT : br1_7 
* INOUT : bl0_8 
* INOUT : br0_8 
* INOUT : bl1_8 
* INOUT : br1_8 
* INOUT : bl0_9 
* INOUT : br0_9 
* INOUT : bl1_9 
* INOUT : br1_9 
* INOUT : bl0_10 
* INOUT : br0_10 
* INOUT : bl1_10 
* INOUT : br1_10 
* INOUT : bl0_11 
* INOUT : br0_11 
* INOUT : bl1_11 
* INOUT : br1_11 
* INOUT : bl0_12 
* INOUT : br0_12 
* INOUT : bl1_12 
* INOUT : br1_12 
* INOUT : bl0_13 
* INOUT : br0_13 
* INOUT : bl1_13 
* INOUT : br1_13 
* INOUT : bl0_14 
* INOUT : br0_14 
* INOUT : bl1_14 
* INOUT : br1_14 
* INOUT : bl0_15 
* INOUT : br0_15 
* INOUT : bl1_15 
* INOUT : br1_15 
* INOUT : bl0_16 
* INOUT : br0_16 
* INOUT : bl1_16 
* INOUT : br1_16 
* INOUT : bl0_17 
* INOUT : br0_17 
* INOUT : bl1_17 
* INOUT : br1_17 
* INOUT : bl0_18 
* INOUT : br0_18 
* INOUT : bl1_18 
* INOUT : br1_18 
* INOUT : bl0_19 
* INOUT : br0_19 
* INOUT : bl1_19 
* INOUT : br1_19 
* INOUT : bl0_20 
* INOUT : br0_20 
* INOUT : bl1_20 
* INOUT : br1_20 
* INOUT : bl0_21 
* INOUT : br0_21 
* INOUT : bl1_21 
* INOUT : br1_21 
* INOUT : bl0_22 
* INOUT : br0_22 
* INOUT : bl1_22 
* INOUT : br1_22 
* INOUT : bl0_23 
* INOUT : br0_23 
* INOUT : bl1_23 
* INOUT : br1_23 
* INOUT : bl0_24 
* INOUT : br0_24 
* INOUT : bl1_24 
* INOUT : br1_24 
* INOUT : bl0_25 
* INOUT : br0_25 
* INOUT : bl1_25 
* INOUT : br1_25 
* INOUT : bl0_26 
* INOUT : br0_26 
* INOUT : bl1_26 
* INOUT : br1_26 
* INOUT : bl0_27 
* INOUT : br0_27 
* INOUT : bl1_27 
* INOUT : br1_27 
* INOUT : bl0_28 
* INOUT : br0_28 
* INOUT : bl1_28 
* INOUT : br1_28 
* INOUT : bl0_29 
* INOUT : br0_29 
* INOUT : bl1_29 
* INOUT : br1_29 
* INOUT : bl0_30 
* INOUT : br0_30 
* INOUT : bl1_30 
* INOUT : br1_30 
* INOUT : bl0_31 
* INOUT : br0_31 
* INOUT : bl1_31 
* INOUT : br1_31 
* INOUT : bl0_32 
* INOUT : br0_32 
* INOUT : bl1_32 
* INOUT : br1_32 
* INOUT : bl0_33 
* INOUT : br0_33 
* INOUT : bl1_33 
* INOUT : br1_33 
* INOUT : bl0_34 
* INOUT : br0_34 
* INOUT : bl1_34 
* INOUT : br1_34 
* INOUT : bl0_35 
* INOUT : br0_35 
* INOUT : bl1_35 
* INOUT : br1_35 
* INOUT : bl0_36 
* INOUT : br0_36 
* INOUT : bl1_36 
* INOUT : br1_36 
* INOUT : bl0_37 
* INOUT : br0_37 
* INOUT : bl1_37 
* INOUT : br1_37 
* INOUT : bl0_38 
* INOUT : br0_38 
* INOUT : bl1_38 
* INOUT : br1_38 
* INOUT : bl0_39 
* INOUT : br0_39 
* INOUT : bl1_39 
* INOUT : br1_39 
* INOUT : bl0_40 
* INOUT : br0_40 
* INOUT : bl1_40 
* INOUT : br1_40 
* INOUT : bl0_41 
* INOUT : br0_41 
* INOUT : bl1_41 
* INOUT : br1_41 
* INOUT : bl0_42 
* INOUT : br0_42 
* INOUT : bl1_42 
* INOUT : br1_42 
* INOUT : bl0_43 
* INOUT : br0_43 
* INOUT : bl1_43 
* INOUT : br1_43 
* INOUT : bl0_44 
* INOUT : br0_44 
* INOUT : bl1_44 
* INOUT : br1_44 
* INOUT : bl0_45 
* INOUT : br0_45 
* INOUT : bl1_45 
* INOUT : br1_45 
* INOUT : bl0_46 
* INOUT : br0_46 
* INOUT : bl1_46 
* INOUT : br1_46 
* INOUT : bl0_47 
* INOUT : br0_47 
* INOUT : bl1_47 
* INOUT : br1_47 
* INOUT : bl0_48 
* INOUT : br0_48 
* INOUT : bl1_48 
* INOUT : br1_48 
* INOUT : bl0_49 
* INOUT : br0_49 
* INOUT : bl1_49 
* INOUT : br1_49 
* INOUT : bl0_50 
* INOUT : br0_50 
* INOUT : bl1_50 
* INOUT : br1_50 
* INOUT : bl0_51 
* INOUT : br0_51 
* INOUT : bl1_51 
* INOUT : br1_51 
* INOUT : bl0_52 
* INOUT : br0_52 
* INOUT : bl1_52 
* INOUT : br1_52 
* INOUT : bl0_53 
* INOUT : br0_53 
* INOUT : bl1_53 
* INOUT : br1_53 
* INOUT : bl0_54 
* INOUT : br0_54 
* INOUT : bl1_54 
* INOUT : br1_54 
* INOUT : bl0_55 
* INOUT : br0_55 
* INOUT : bl1_55 
* INOUT : br1_55 
* INOUT : bl0_56 
* INOUT : br0_56 
* INOUT : bl1_56 
* INOUT : br1_56 
* INOUT : bl0_57 
* INOUT : br0_57 
* INOUT : bl1_57 
* INOUT : br1_57 
* INOUT : bl0_58 
* INOUT : br0_58 
* INOUT : bl1_58 
* INOUT : br1_58 
* INOUT : bl0_59 
* INOUT : br0_59 
* INOUT : bl1_59 
* INOUT : br1_59 
* INOUT : bl0_60 
* INOUT : br0_60 
* INOUT : bl1_60 
* INOUT : br1_60 
* INOUT : bl0_61 
* INOUT : br0_61 
* INOUT : bl1_61 
* INOUT : br1_61 
* INOUT : bl0_62 
* INOUT : br0_62 
* INOUT : bl1_62 
* INOUT : br1_62 
* INOUT : bl0_63 
* INOUT : br0_63 
* INOUT : bl1_63 
* INOUT : br1_63 
* INPUT : wl0_0 
* INPUT : wl1_0 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 64
Xbit_r0_c0 bl0_0 br0_0 bl1_0 br1_0 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c1 bl0_1 br0_1 bl1_1 br1_1 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c2 bl0_2 br0_2 bl1_2 br1_2 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c3 bl0_3 br0_3 bl1_3 br1_3 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c4 bl0_4 br0_4 bl1_4 br1_4 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c5 bl0_5 br0_5 bl1_5 br1_5 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c6 bl0_6 br0_6 bl1_6 br1_6 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c7 bl0_7 br0_7 bl1_7 br1_7 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c8 bl0_8 br0_8 bl1_8 br1_8 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c9 bl0_9 br0_9 bl1_9 br1_9 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c10 bl0_10 br0_10 bl1_10 br1_10 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c11 bl0_11 br0_11 bl1_11 br1_11 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c12 bl0_12 br0_12 bl1_12 br1_12 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c13 bl0_13 br0_13 bl1_13 br1_13 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c14 bl0_14 br0_14 bl1_14 br1_14 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c15 bl0_15 br0_15 bl1_15 br1_15 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c16 bl0_16 br0_16 bl1_16 br1_16 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c17 bl0_17 br0_17 bl1_17 br1_17 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c18 bl0_18 br0_18 bl1_18 br1_18 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c19 bl0_19 br0_19 bl1_19 br1_19 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c20 bl0_20 br0_20 bl1_20 br1_20 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c21 bl0_21 br0_21 bl1_21 br1_21 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c22 bl0_22 br0_22 bl1_22 br1_22 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c23 bl0_23 br0_23 bl1_23 br1_23 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c24 bl0_24 br0_24 bl1_24 br1_24 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c25 bl0_25 br0_25 bl1_25 br1_25 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c26 bl0_26 br0_26 bl1_26 br1_26 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c27 bl0_27 br0_27 bl1_27 br1_27 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c28 bl0_28 br0_28 bl1_28 br1_28 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c29 bl0_29 br0_29 bl1_29 br1_29 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c30 bl0_30 br0_30 bl1_30 br1_30 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c31 bl0_31 br0_31 bl1_31 br1_31 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c32 bl0_32 br0_32 bl1_32 br1_32 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c33 bl0_33 br0_33 bl1_33 br1_33 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c34 bl0_34 br0_34 bl1_34 br1_34 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c35 bl0_35 br0_35 bl1_35 br1_35 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c36 bl0_36 br0_36 bl1_36 br1_36 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c37 bl0_37 br0_37 bl1_37 br1_37 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c38 bl0_38 br0_38 bl1_38 br1_38 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c39 bl0_39 br0_39 bl1_39 br1_39 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c40 bl0_40 br0_40 bl1_40 br1_40 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c41 bl0_41 br0_41 bl1_41 br1_41 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c42 bl0_42 br0_42 bl1_42 br1_42 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c43 bl0_43 br0_43 bl1_43 br1_43 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c44 bl0_44 br0_44 bl1_44 br1_44 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c45 bl0_45 br0_45 bl1_45 br1_45 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c46 bl0_46 br0_46 bl1_46 br1_46 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c47 bl0_47 br0_47 bl1_47 br1_47 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c48 bl0_48 br0_48 bl1_48 br1_48 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c49 bl0_49 br0_49 bl1_49 br1_49 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c50 bl0_50 br0_50 bl1_50 br1_50 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c51 bl0_51 br0_51 bl1_51 br1_51 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c52 bl0_52 br0_52 bl1_52 br1_52 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c53 bl0_53 br0_53 bl1_53 br1_53 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c54 bl0_54 br0_54 bl1_54 br1_54 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c55 bl0_55 br0_55 bl1_55 br1_55 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c56 bl0_56 br0_56 bl1_56 br1_56 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c57 bl0_57 br0_57 bl1_57 br1_57 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c58 bl0_58 br0_58 bl1_58 br1_58 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c59 bl0_59 br0_59 bl1_59 br1_59 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c60 bl0_60 br0_60 bl1_60 br1_60 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c61 bl0_61 br0_61 bl1_61 br1_61 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c62 bl0_62 br0_62 bl1_62 br1_62 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xbit_r0_c63 bl0_63 br0_63 bl1_63 br1_63 wl0_0 wl1_0 vdd gnd sky130_fd_bd_sram__openram_dp_cell_dummy
.ENDS dummy_array

.SUBCKT replica_bitcell_array bl0_0 br0_0 bl1_0 br1_0 bl0_1 br0_1 bl1_1 br1_1 bl0_2 br0_2 bl1_2 br1_2 bl0_3 br0_3 bl1_3 br1_3 bl0_4 br0_4 bl1_4 br1_4 bl0_5 br0_5 bl1_5 br1_5 bl0_6 br0_6 bl1_6 br1_6 bl0_7 br0_7 bl1_7 br1_7 bl0_8 br0_8 bl1_8 br1_8 bl0_9 br0_9 bl1_9 br1_9 bl0_10 br0_10 bl1_10 br1_10 bl0_11 br0_11 bl1_11 br1_11 bl0_12 br0_12 bl1_12 br1_12 bl0_13 br0_13 bl1_13 br1_13 bl0_14 br0_14 bl1_14 br1_14 bl0_15 br0_15 bl1_15 br1_15 bl0_16 br0_16 bl1_16 br1_16 bl0_17 br0_17 bl1_17 br1_17 bl0_18 br0_18 bl1_18 br1_18 bl0_19 br0_19 bl1_19 br1_19 bl0_20 br0_20 bl1_20 br1_20 bl0_21 br0_21 bl1_21 br1_21 bl0_22 br0_22 bl1_22 br1_22 bl0_23 br0_23 bl1_23 br1_23 bl0_24 br0_24 bl1_24 br1_24 bl0_25 br0_25 bl1_25 br1_25 bl0_26 br0_26 bl1_26 br1_26 bl0_27 br0_27 bl1_27 br1_27 bl0_28 br0_28 bl1_28 br1_28 bl0_29 br0_29 bl1_29 br1_29 bl0_30 br0_30 bl1_30 br1_30 bl0_31 br0_31 bl1_31 br1_31 bl0_32 br0_32 bl1_32 br1_32 bl0_33 br0_33 bl1_33 br1_33 bl0_34 br0_34 bl1_34 br1_34 bl0_35 br0_35 bl1_35 br1_35 bl0_36 br0_36 bl1_36 br1_36 bl0_37 br0_37 bl1_37 br1_37 bl0_38 br0_38 bl1_38 br1_38 bl0_39 br0_39 bl1_39 br1_39 bl0_40 br0_40 bl1_40 br1_40 bl0_41 br0_41 bl1_41 br1_41 bl0_42 br0_42 bl1_42 br1_42 bl0_43 br0_43 bl1_43 br1_43 bl0_44 br0_44 bl1_44 br1_44 bl0_45 br0_45 bl1_45 br1_45 bl0_46 br0_46 bl1_46 br1_46 bl0_47 br0_47 bl1_47 br1_47 bl0_48 br0_48 bl1_48 br1_48 bl0_49 br0_49 bl1_49 br1_49 bl0_50 br0_50 bl1_50 br1_50 bl0_51 br0_51 bl1_51 br1_51 bl0_52 br0_52 bl1_52 br1_52 bl0_53 br0_53 bl1_53 br1_53 bl0_54 br0_54 bl1_54 br1_54 bl0_55 br0_55 bl1_55 br1_55 bl0_56 br0_56 bl1_56 br1_56 bl0_57 br0_57 bl1_57 br1_57 bl0_58 br0_58 bl1_58 br1_58 bl0_59 br0_59 bl1_59 br1_59 bl0_60 br0_60 bl1_60 br1_60 bl0_61 br0_61 bl1_61 br1_61 bl0_62 br0_62 bl1_62 br1_62 bl0_63 br0_63 bl1_63 br1_63 rbl_bl0_0 rbl_br0_0 rbl_bl1_1 rbl_br1_1 wl0_0 wl1_0 wl0_1 wl1_1 wl0_2 wl1_2 wl0_3 wl1_3 wl0_4 wl1_4 wl0_5 wl1_5 wl0_6 wl1_6 wl0_7 wl1_7 wl0_8 wl1_8 wl0_9 wl1_9 wl0_10 wl1_10 wl0_11 wl1_11 wl0_12 wl1_12 wl0_13 wl1_13 wl0_14 wl1_14 wl0_15 wl1_15 wl0_16 wl1_16 wl0_17 wl1_17 wl0_18 wl1_18 wl0_19 wl1_19 wl0_20 wl1_20 wl0_21 wl1_21 wl0_22 wl1_22 wl0_23 wl1_23 wl0_24 wl1_24 wl0_25 wl1_25 wl0_26 wl1_26 wl0_27 wl1_27 wl0_28 wl1_28 wl0_29 wl1_29 wl0_30 wl1_30 wl0_31 wl1_31 wl0_32 wl1_32 wl0_33 wl1_33 wl0_34 wl1_34 wl0_35 wl1_35 wl0_36 wl1_36 wl0_37 wl1_37 wl0_38 wl1_38 wl0_39 wl1_39 wl0_40 wl1_40 wl0_41 wl1_41 wl0_42 wl1_42 wl0_43 wl1_43 wl0_44 wl1_44 wl0_45 wl1_45 wl0_46 wl1_46 wl0_47 wl1_47 wl0_48 wl1_48 wl0_49 wl1_49 wl0_50 wl1_50 wl0_51 wl1_51 wl0_52 wl1_52 wl0_53 wl1_53 wl0_54 wl1_54 wl0_55 wl1_55 wl0_56 wl1_56 wl0_57 wl1_57 wl0_58 wl1_58 wl0_59 wl1_59 wl0_60 wl1_60 wl0_61 wl1_61 wl0_62 wl1_62 wl0_63 wl1_63 wl0_64 wl1_64 wl0_65 wl1_65 wl0_66 wl1_66 wl0_67 wl1_67 wl0_68 wl1_68 wl0_69 wl1_69 wl0_70 wl1_70 wl0_71 wl1_71 wl0_72 wl1_72 wl0_73 wl1_73 wl0_74 wl1_74 wl0_75 wl1_75 wl0_76 wl1_76 wl0_77 wl1_77 wl0_78 wl1_78 wl0_79 wl1_79 wl0_80 wl1_80 wl0_81 wl1_81 wl0_82 wl1_82 wl0_83 wl1_83 wl0_84 wl1_84 wl0_85 wl1_85 wl0_86 wl1_86 wl0_87 wl1_87 wl0_88 wl1_88 wl0_89 wl1_89 wl0_90 wl1_90 wl0_91 wl1_91 wl0_92 wl1_92 wl0_93 wl1_93 wl0_94 wl1_94 wl0_95 wl1_95 wl0_96 wl1_96 wl0_97 wl1_97 wl0_98 wl1_98 wl0_99 wl1_99 wl0_100 wl1_100 wl0_101 wl1_101 wl0_102 wl1_102 wl0_103 wl1_103 wl0_104 wl1_104 wl0_105 wl1_105 wl0_106 wl1_106 wl0_107 wl1_107 wl0_108 wl1_108 wl0_109 wl1_109 wl0_110 wl1_110 wl0_111 wl1_111 wl0_112 wl1_112 wl0_113 wl1_113 wl0_114 wl1_114 wl0_115 wl1_115 wl0_116 wl1_116 wl0_117 wl1_117 wl0_118 wl1_118 wl0_119 wl1_119 wl0_120 wl1_120 wl0_121 wl1_121 wl0_122 wl1_122 wl0_123 wl1_123 wl0_124 wl1_124 wl0_125 wl1_125 wl0_126 wl1_126 wl0_127 wl1_127 rbl_wl0_0 rbl_wl1_1 vdd gnd
* INOUT : bl0_0 
* INOUT : br0_0 
* INOUT : bl1_0 
* INOUT : br1_0 
* INOUT : bl0_1 
* INOUT : br0_1 
* INOUT : bl1_1 
* INOUT : br1_1 
* INOUT : bl0_2 
* INOUT : br0_2 
* INOUT : bl1_2 
* INOUT : br1_2 
* INOUT : bl0_3 
* INOUT : br0_3 
* INOUT : bl1_3 
* INOUT : br1_3 
* INOUT : bl0_4 
* INOUT : br0_4 
* INOUT : bl1_4 
* INOUT : br1_4 
* INOUT : bl0_5 
* INOUT : br0_5 
* INOUT : bl1_5 
* INOUT : br1_5 
* INOUT : bl0_6 
* INOUT : br0_6 
* INOUT : bl1_6 
* INOUT : br1_6 
* INOUT : bl0_7 
* INOUT : br0_7 
* INOUT : bl1_7 
* INOUT : br1_7 
* INOUT : bl0_8 
* INOUT : br0_8 
* INOUT : bl1_8 
* INOUT : br1_8 
* INOUT : bl0_9 
* INOUT : br0_9 
* INOUT : bl1_9 
* INOUT : br1_9 
* INOUT : bl0_10 
* INOUT : br0_10 
* INOUT : bl1_10 
* INOUT : br1_10 
* INOUT : bl0_11 
* INOUT : br0_11 
* INOUT : bl1_11 
* INOUT : br1_11 
* INOUT : bl0_12 
* INOUT : br0_12 
* INOUT : bl1_12 
* INOUT : br1_12 
* INOUT : bl0_13 
* INOUT : br0_13 
* INOUT : bl1_13 
* INOUT : br1_13 
* INOUT : bl0_14 
* INOUT : br0_14 
* INOUT : bl1_14 
* INOUT : br1_14 
* INOUT : bl0_15 
* INOUT : br0_15 
* INOUT : bl1_15 
* INOUT : br1_15 
* INOUT : bl0_16 
* INOUT : br0_16 
* INOUT : bl1_16 
* INOUT : br1_16 
* INOUT : bl0_17 
* INOUT : br0_17 
* INOUT : bl1_17 
* INOUT : br1_17 
* INOUT : bl0_18 
* INOUT : br0_18 
* INOUT : bl1_18 
* INOUT : br1_18 
* INOUT : bl0_19 
* INOUT : br0_19 
* INOUT : bl1_19 
* INOUT : br1_19 
* INOUT : bl0_20 
* INOUT : br0_20 
* INOUT : bl1_20 
* INOUT : br1_20 
* INOUT : bl0_21 
* INOUT : br0_21 
* INOUT : bl1_21 
* INOUT : br1_21 
* INOUT : bl0_22 
* INOUT : br0_22 
* INOUT : bl1_22 
* INOUT : br1_22 
* INOUT : bl0_23 
* INOUT : br0_23 
* INOUT : bl1_23 
* INOUT : br1_23 
* INOUT : bl0_24 
* INOUT : br0_24 
* INOUT : bl1_24 
* INOUT : br1_24 
* INOUT : bl0_25 
* INOUT : br0_25 
* INOUT : bl1_25 
* INOUT : br1_25 
* INOUT : bl0_26 
* INOUT : br0_26 
* INOUT : bl1_26 
* INOUT : br1_26 
* INOUT : bl0_27 
* INOUT : br0_27 
* INOUT : bl1_27 
* INOUT : br1_27 
* INOUT : bl0_28 
* INOUT : br0_28 
* INOUT : bl1_28 
* INOUT : br1_28 
* INOUT : bl0_29 
* INOUT : br0_29 
* INOUT : bl1_29 
* INOUT : br1_29 
* INOUT : bl0_30 
* INOUT : br0_30 
* INOUT : bl1_30 
* INOUT : br1_30 
* INOUT : bl0_31 
* INOUT : br0_31 
* INOUT : bl1_31 
* INOUT : br1_31 
* INOUT : bl0_32 
* INOUT : br0_32 
* INOUT : bl1_32 
* INOUT : br1_32 
* INOUT : bl0_33 
* INOUT : br0_33 
* INOUT : bl1_33 
* INOUT : br1_33 
* INOUT : bl0_34 
* INOUT : br0_34 
* INOUT : bl1_34 
* INOUT : br1_34 
* INOUT : bl0_35 
* INOUT : br0_35 
* INOUT : bl1_35 
* INOUT : br1_35 
* INOUT : bl0_36 
* INOUT : br0_36 
* INOUT : bl1_36 
* INOUT : br1_36 
* INOUT : bl0_37 
* INOUT : br0_37 
* INOUT : bl1_37 
* INOUT : br1_37 
* INOUT : bl0_38 
* INOUT : br0_38 
* INOUT : bl1_38 
* INOUT : br1_38 
* INOUT : bl0_39 
* INOUT : br0_39 
* INOUT : bl1_39 
* INOUT : br1_39 
* INOUT : bl0_40 
* INOUT : br0_40 
* INOUT : bl1_40 
* INOUT : br1_40 
* INOUT : bl0_41 
* INOUT : br0_41 
* INOUT : bl1_41 
* INOUT : br1_41 
* INOUT : bl0_42 
* INOUT : br0_42 
* INOUT : bl1_42 
* INOUT : br1_42 
* INOUT : bl0_43 
* INOUT : br0_43 
* INOUT : bl1_43 
* INOUT : br1_43 
* INOUT : bl0_44 
* INOUT : br0_44 
* INOUT : bl1_44 
* INOUT : br1_44 
* INOUT : bl0_45 
* INOUT : br0_45 
* INOUT : bl1_45 
* INOUT : br1_45 
* INOUT : bl0_46 
* INOUT : br0_46 
* INOUT : bl1_46 
* INOUT : br1_46 
* INOUT : bl0_47 
* INOUT : br0_47 
* INOUT : bl1_47 
* INOUT : br1_47 
* INOUT : bl0_48 
* INOUT : br0_48 
* INOUT : bl1_48 
* INOUT : br1_48 
* INOUT : bl0_49 
* INOUT : br0_49 
* INOUT : bl1_49 
* INOUT : br1_49 
* INOUT : bl0_50 
* INOUT : br0_50 
* INOUT : bl1_50 
* INOUT : br1_50 
* INOUT : bl0_51 
* INOUT : br0_51 
* INOUT : bl1_51 
* INOUT : br1_51 
* INOUT : bl0_52 
* INOUT : br0_52 
* INOUT : bl1_52 
* INOUT : br1_52 
* INOUT : bl0_53 
* INOUT : br0_53 
* INOUT : bl1_53 
* INOUT : br1_53 
* INOUT : bl0_54 
* INOUT : br0_54 
* INOUT : bl1_54 
* INOUT : br1_54 
* INOUT : bl0_55 
* INOUT : br0_55 
* INOUT : bl1_55 
* INOUT : br1_55 
* INOUT : bl0_56 
* INOUT : br0_56 
* INOUT : bl1_56 
* INOUT : br1_56 
* INOUT : bl0_57 
* INOUT : br0_57 
* INOUT : bl1_57 
* INOUT : br1_57 
* INOUT : bl0_58 
* INOUT : br0_58 
* INOUT : bl1_58 
* INOUT : br1_58 
* INOUT : bl0_59 
* INOUT : br0_59 
* INOUT : bl1_59 
* INOUT : br1_59 
* INOUT : bl0_60 
* INOUT : br0_60 
* INOUT : bl1_60 
* INOUT : br1_60 
* INOUT : bl0_61 
* INOUT : br0_61 
* INOUT : bl1_61 
* INOUT : br1_61 
* INOUT : bl0_62 
* INOUT : br0_62 
* INOUT : bl1_62 
* INOUT : br1_62 
* INOUT : bl0_63 
* INOUT : br0_63 
* INOUT : bl1_63 
* INOUT : br1_63 
* OUTPUT: rbl_bl0_0 
* OUTPUT: rbl_br0_0 
* OUTPUT: rbl_bl1_1 
* OUTPUT: rbl_br1_1 
* INPUT : wl0_0 
* INPUT : wl1_0 
* INPUT : wl0_1 
* INPUT : wl1_1 
* INPUT : wl0_2 
* INPUT : wl1_2 
* INPUT : wl0_3 
* INPUT : wl1_3 
* INPUT : wl0_4 
* INPUT : wl1_4 
* INPUT : wl0_5 
* INPUT : wl1_5 
* INPUT : wl0_6 
* INPUT : wl1_6 
* INPUT : wl0_7 
* INPUT : wl1_7 
* INPUT : wl0_8 
* INPUT : wl1_8 
* INPUT : wl0_9 
* INPUT : wl1_9 
* INPUT : wl0_10 
* INPUT : wl1_10 
* INPUT : wl0_11 
* INPUT : wl1_11 
* INPUT : wl0_12 
* INPUT : wl1_12 
* INPUT : wl0_13 
* INPUT : wl1_13 
* INPUT : wl0_14 
* INPUT : wl1_14 
* INPUT : wl0_15 
* INPUT : wl1_15 
* INPUT : wl0_16 
* INPUT : wl1_16 
* INPUT : wl0_17 
* INPUT : wl1_17 
* INPUT : wl0_18 
* INPUT : wl1_18 
* INPUT : wl0_19 
* INPUT : wl1_19 
* INPUT : wl0_20 
* INPUT : wl1_20 
* INPUT : wl0_21 
* INPUT : wl1_21 
* INPUT : wl0_22 
* INPUT : wl1_22 
* INPUT : wl0_23 
* INPUT : wl1_23 
* INPUT : wl0_24 
* INPUT : wl1_24 
* INPUT : wl0_25 
* INPUT : wl1_25 
* INPUT : wl0_26 
* INPUT : wl1_26 
* INPUT : wl0_27 
* INPUT : wl1_27 
* INPUT : wl0_28 
* INPUT : wl1_28 
* INPUT : wl0_29 
* INPUT : wl1_29 
* INPUT : wl0_30 
* INPUT : wl1_30 
* INPUT : wl0_31 
* INPUT : wl1_31 
* INPUT : wl0_32 
* INPUT : wl1_32 
* INPUT : wl0_33 
* INPUT : wl1_33 
* INPUT : wl0_34 
* INPUT : wl1_34 
* INPUT : wl0_35 
* INPUT : wl1_35 
* INPUT : wl0_36 
* INPUT : wl1_36 
* INPUT : wl0_37 
* INPUT : wl1_37 
* INPUT : wl0_38 
* INPUT : wl1_38 
* INPUT : wl0_39 
* INPUT : wl1_39 
* INPUT : wl0_40 
* INPUT : wl1_40 
* INPUT : wl0_41 
* INPUT : wl1_41 
* INPUT : wl0_42 
* INPUT : wl1_42 
* INPUT : wl0_43 
* INPUT : wl1_43 
* INPUT : wl0_44 
* INPUT : wl1_44 
* INPUT : wl0_45 
* INPUT : wl1_45 
* INPUT : wl0_46 
* INPUT : wl1_46 
* INPUT : wl0_47 
* INPUT : wl1_47 
* INPUT : wl0_48 
* INPUT : wl1_48 
* INPUT : wl0_49 
* INPUT : wl1_49 
* INPUT : wl0_50 
* INPUT : wl1_50 
* INPUT : wl0_51 
* INPUT : wl1_51 
* INPUT : wl0_52 
* INPUT : wl1_52 
* INPUT : wl0_53 
* INPUT : wl1_53 
* INPUT : wl0_54 
* INPUT : wl1_54 
* INPUT : wl0_55 
* INPUT : wl1_55 
* INPUT : wl0_56 
* INPUT : wl1_56 
* INPUT : wl0_57 
* INPUT : wl1_57 
* INPUT : wl0_58 
* INPUT : wl1_58 
* INPUT : wl0_59 
* INPUT : wl1_59 
* INPUT : wl0_60 
* INPUT : wl1_60 
* INPUT : wl0_61 
* INPUT : wl1_61 
* INPUT : wl0_62 
* INPUT : wl1_62 
* INPUT : wl0_63 
* INPUT : wl1_63 
* INPUT : wl0_64 
* INPUT : wl1_64 
* INPUT : wl0_65 
* INPUT : wl1_65 
* INPUT : wl0_66 
* INPUT : wl1_66 
* INPUT : wl0_67 
* INPUT : wl1_67 
* INPUT : wl0_68 
* INPUT : wl1_68 
* INPUT : wl0_69 
* INPUT : wl1_69 
* INPUT : wl0_70 
* INPUT : wl1_70 
* INPUT : wl0_71 
* INPUT : wl1_71 
* INPUT : wl0_72 
* INPUT : wl1_72 
* INPUT : wl0_73 
* INPUT : wl1_73 
* INPUT : wl0_74 
* INPUT : wl1_74 
* INPUT : wl0_75 
* INPUT : wl1_75 
* INPUT : wl0_76 
* INPUT : wl1_76 
* INPUT : wl0_77 
* INPUT : wl1_77 
* INPUT : wl0_78 
* INPUT : wl1_78 
* INPUT : wl0_79 
* INPUT : wl1_79 
* INPUT : wl0_80 
* INPUT : wl1_80 
* INPUT : wl0_81 
* INPUT : wl1_81 
* INPUT : wl0_82 
* INPUT : wl1_82 
* INPUT : wl0_83 
* INPUT : wl1_83 
* INPUT : wl0_84 
* INPUT : wl1_84 
* INPUT : wl0_85 
* INPUT : wl1_85 
* INPUT : wl0_86 
* INPUT : wl1_86 
* INPUT : wl0_87 
* INPUT : wl1_87 
* INPUT : wl0_88 
* INPUT : wl1_88 
* INPUT : wl0_89 
* INPUT : wl1_89 
* INPUT : wl0_90 
* INPUT : wl1_90 
* INPUT : wl0_91 
* INPUT : wl1_91 
* INPUT : wl0_92 
* INPUT : wl1_92 
* INPUT : wl0_93 
* INPUT : wl1_93 
* INPUT : wl0_94 
* INPUT : wl1_94 
* INPUT : wl0_95 
* INPUT : wl1_95 
* INPUT : wl0_96 
* INPUT : wl1_96 
* INPUT : wl0_97 
* INPUT : wl1_97 
* INPUT : wl0_98 
* INPUT : wl1_98 
* INPUT : wl0_99 
* INPUT : wl1_99 
* INPUT : wl0_100 
* INPUT : wl1_100 
* INPUT : wl0_101 
* INPUT : wl1_101 
* INPUT : wl0_102 
* INPUT : wl1_102 
* INPUT : wl0_103 
* INPUT : wl1_103 
* INPUT : wl0_104 
* INPUT : wl1_104 
* INPUT : wl0_105 
* INPUT : wl1_105 
* INPUT : wl0_106 
* INPUT : wl1_106 
* INPUT : wl0_107 
* INPUT : wl1_107 
* INPUT : wl0_108 
* INPUT : wl1_108 
* INPUT : wl0_109 
* INPUT : wl1_109 
* INPUT : wl0_110 
* INPUT : wl1_110 
* INPUT : wl0_111 
* INPUT : wl1_111 
* INPUT : wl0_112 
* INPUT : wl1_112 
* INPUT : wl0_113 
* INPUT : wl1_113 
* INPUT : wl0_114 
* INPUT : wl1_114 
* INPUT : wl0_115 
* INPUT : wl1_115 
* INPUT : wl0_116 
* INPUT : wl1_116 
* INPUT : wl0_117 
* INPUT : wl1_117 
* INPUT : wl0_118 
* INPUT : wl1_118 
* INPUT : wl0_119 
* INPUT : wl1_119 
* INPUT : wl0_120 
* INPUT : wl1_120 
* INPUT : wl0_121 
* INPUT : wl1_121 
* INPUT : wl0_122 
* INPUT : wl1_122 
* INPUT : wl0_123 
* INPUT : wl1_123 
* INPUT : wl0_124 
* INPUT : wl1_124 
* INPUT : wl0_125 
* INPUT : wl1_125 
* INPUT : wl0_126 
* INPUT : wl1_126 
* INPUT : wl0_127 
* INPUT : wl1_127 
* INPUT : rbl_wl0_0 
* INPUT : rbl_wl1_1 
* POWER : vdd 
* GROUND: gnd 
* rows: 128 cols: 64
Xbitcell_array bl0_0 br0_0 bl1_0 br1_0 bl0_1 br0_1 bl1_1 br1_1 bl0_2 br0_2 bl1_2 br1_2 bl0_3 br0_3 bl1_3 br1_3 bl0_4 br0_4 bl1_4 br1_4 bl0_5 br0_5 bl1_5 br1_5 bl0_6 br0_6 bl1_6 br1_6 bl0_7 br0_7 bl1_7 br1_7 bl0_8 br0_8 bl1_8 br1_8 bl0_9 br0_9 bl1_9 br1_9 bl0_10 br0_10 bl1_10 br1_10 bl0_11 br0_11 bl1_11 br1_11 bl0_12 br0_12 bl1_12 br1_12 bl0_13 br0_13 bl1_13 br1_13 bl0_14 br0_14 bl1_14 br1_14 bl0_15 br0_15 bl1_15 br1_15 bl0_16 br0_16 bl1_16 br1_16 bl0_17 br0_17 bl1_17 br1_17 bl0_18 br0_18 bl1_18 br1_18 bl0_19 br0_19 bl1_19 br1_19 bl0_20 br0_20 bl1_20 br1_20 bl0_21 br0_21 bl1_21 br1_21 bl0_22 br0_22 bl1_22 br1_22 bl0_23 br0_23 bl1_23 br1_23 bl0_24 br0_24 bl1_24 br1_24 bl0_25 br0_25 bl1_25 br1_25 bl0_26 br0_26 bl1_26 br1_26 bl0_27 br0_27 bl1_27 br1_27 bl0_28 br0_28 bl1_28 br1_28 bl0_29 br0_29 bl1_29 br1_29 bl0_30 br0_30 bl1_30 br1_30 bl0_31 br0_31 bl1_31 br1_31 bl0_32 br0_32 bl1_32 br1_32 bl0_33 br0_33 bl1_33 br1_33 bl0_34 br0_34 bl1_34 br1_34 bl0_35 br0_35 bl1_35 br1_35 bl0_36 br0_36 bl1_36 br1_36 bl0_37 br0_37 bl1_37 br1_37 bl0_38 br0_38 bl1_38 br1_38 bl0_39 br0_39 bl1_39 br1_39 bl0_40 br0_40 bl1_40 br1_40 bl0_41 br0_41 bl1_41 br1_41 bl0_42 br0_42 bl1_42 br1_42 bl0_43 br0_43 bl1_43 br1_43 bl0_44 br0_44 bl1_44 br1_44 bl0_45 br0_45 bl1_45 br1_45 bl0_46 br0_46 bl1_46 br1_46 bl0_47 br0_47 bl1_47 br1_47 bl0_48 br0_48 bl1_48 br1_48 bl0_49 br0_49 bl1_49 br1_49 bl0_50 br0_50 bl1_50 br1_50 bl0_51 br0_51 bl1_51 br1_51 bl0_52 br0_52 bl1_52 br1_52 bl0_53 br0_53 bl1_53 br1_53 bl0_54 br0_54 bl1_54 br1_54 bl0_55 br0_55 bl1_55 br1_55 bl0_56 br0_56 bl1_56 br1_56 bl0_57 br0_57 bl1_57 br1_57 bl0_58 br0_58 bl1_58 br1_58 bl0_59 br0_59 bl1_59 br1_59 bl0_60 br0_60 bl1_60 br1_60 bl0_61 br0_61 bl1_61 br1_61 bl0_62 br0_62 bl1_62 br1_62 bl0_63 br0_63 bl1_63 br1_63 wl0_0 wl1_0 wl0_1 wl1_1 wl0_2 wl1_2 wl0_3 wl1_3 wl0_4 wl1_4 wl0_5 wl1_5 wl0_6 wl1_6 wl0_7 wl1_7 wl0_8 wl1_8 wl0_9 wl1_9 wl0_10 wl1_10 wl0_11 wl1_11 wl0_12 wl1_12 wl0_13 wl1_13 wl0_14 wl1_14 wl0_15 wl1_15 wl0_16 wl1_16 wl0_17 wl1_17 wl0_18 wl1_18 wl0_19 wl1_19 wl0_20 wl1_20 wl0_21 wl1_21 wl0_22 wl1_22 wl0_23 wl1_23 wl0_24 wl1_24 wl0_25 wl1_25 wl0_26 wl1_26 wl0_27 wl1_27 wl0_28 wl1_28 wl0_29 wl1_29 wl0_30 wl1_30 wl0_31 wl1_31 wl0_32 wl1_32 wl0_33 wl1_33 wl0_34 wl1_34 wl0_35 wl1_35 wl0_36 wl1_36 wl0_37 wl1_37 wl0_38 wl1_38 wl0_39 wl1_39 wl0_40 wl1_40 wl0_41 wl1_41 wl0_42 wl1_42 wl0_43 wl1_43 wl0_44 wl1_44 wl0_45 wl1_45 wl0_46 wl1_46 wl0_47 wl1_47 wl0_48 wl1_48 wl0_49 wl1_49 wl0_50 wl1_50 wl0_51 wl1_51 wl0_52 wl1_52 wl0_53 wl1_53 wl0_54 wl1_54 wl0_55 wl1_55 wl0_56 wl1_56 wl0_57 wl1_57 wl0_58 wl1_58 wl0_59 wl1_59 wl0_60 wl1_60 wl0_61 wl1_61 wl0_62 wl1_62 wl0_63 wl1_63 wl0_64 wl1_64 wl0_65 wl1_65 wl0_66 wl1_66 wl0_67 wl1_67 wl0_68 wl1_68 wl0_69 wl1_69 wl0_70 wl1_70 wl0_71 wl1_71 wl0_72 wl1_72 wl0_73 wl1_73 wl0_74 wl1_74 wl0_75 wl1_75 wl0_76 wl1_76 wl0_77 wl1_77 wl0_78 wl1_78 wl0_79 wl1_79 wl0_80 wl1_80 wl0_81 wl1_81 wl0_82 wl1_82 wl0_83 wl1_83 wl0_84 wl1_84 wl0_85 wl1_85 wl0_86 wl1_86 wl0_87 wl1_87 wl0_88 wl1_88 wl0_89 wl1_89 wl0_90 wl1_90 wl0_91 wl1_91 wl0_92 wl1_92 wl0_93 wl1_93 wl0_94 wl1_94 wl0_95 wl1_95 wl0_96 wl1_96 wl0_97 wl1_97 wl0_98 wl1_98 wl0_99 wl1_99 wl0_100 wl1_100 wl0_101 wl1_101 wl0_102 wl1_102 wl0_103 wl1_103 wl0_104 wl1_104 wl0_105 wl1_105 wl0_106 wl1_106 wl0_107 wl1_107 wl0_108 wl1_108 wl0_109 wl1_109 wl0_110 wl1_110 wl0_111 wl1_111 wl0_112 wl1_112 wl0_113 wl1_113 wl0_114 wl1_114 wl0_115 wl1_115 wl0_116 wl1_116 wl0_117 wl1_117 wl0_118 wl1_118 wl0_119 wl1_119 wl0_120 wl1_120 wl0_121 wl1_121 wl0_122 wl1_122 wl0_123 wl1_123 wl0_124 wl1_124 wl0_125 wl1_125 wl0_126 wl1_126 wl0_127 wl1_127 vdd gnd bitcell_array
Xreplica_col_0 rbl_bl0_0 rbl_br0_0 rbl_bl1_0 rbl_br1_0 dummy_wl0_bot dummy_wl1_bot rbl_wl0_0 gnd wl0_0 wl1_0 wl0_1 wl1_1 wl0_2 wl1_2 wl0_3 wl1_3 wl0_4 wl1_4 wl0_5 wl1_5 wl0_6 wl1_6 wl0_7 wl1_7 wl0_8 wl1_8 wl0_9 wl1_9 wl0_10 wl1_10 wl0_11 wl1_11 wl0_12 wl1_12 wl0_13 wl1_13 wl0_14 wl1_14 wl0_15 wl1_15 wl0_16 wl1_16 wl0_17 wl1_17 wl0_18 wl1_18 wl0_19 wl1_19 wl0_20 wl1_20 wl0_21 wl1_21 wl0_22 wl1_22 wl0_23 wl1_23 wl0_24 wl1_24 wl0_25 wl1_25 wl0_26 wl1_26 wl0_27 wl1_27 wl0_28 wl1_28 wl0_29 wl1_29 wl0_30 wl1_30 wl0_31 wl1_31 wl0_32 wl1_32 wl0_33 wl1_33 wl0_34 wl1_34 wl0_35 wl1_35 wl0_36 wl1_36 wl0_37 wl1_37 wl0_38 wl1_38 wl0_39 wl1_39 wl0_40 wl1_40 wl0_41 wl1_41 wl0_42 wl1_42 wl0_43 wl1_43 wl0_44 wl1_44 wl0_45 wl1_45 wl0_46 wl1_46 wl0_47 wl1_47 wl0_48 wl1_48 wl0_49 wl1_49 wl0_50 wl1_50 wl0_51 wl1_51 wl0_52 wl1_52 wl0_53 wl1_53 wl0_54 wl1_54 wl0_55 wl1_55 wl0_56 wl1_56 wl0_57 wl1_57 wl0_58 wl1_58 wl0_59 wl1_59 wl0_60 wl1_60 wl0_61 wl1_61 wl0_62 wl1_62 wl0_63 wl1_63 wl0_64 wl1_64 wl0_65 wl1_65 wl0_66 wl1_66 wl0_67 wl1_67 wl0_68 wl1_68 wl0_69 wl1_69 wl0_70 wl1_70 wl0_71 wl1_71 wl0_72 wl1_72 wl0_73 wl1_73 wl0_74 wl1_74 wl0_75 wl1_75 wl0_76 wl1_76 wl0_77 wl1_77 wl0_78 wl1_78 wl0_79 wl1_79 wl0_80 wl1_80 wl0_81 wl1_81 wl0_82 wl1_82 wl0_83 wl1_83 wl0_84 wl1_84 wl0_85 wl1_85 wl0_86 wl1_86 wl0_87 wl1_87 wl0_88 wl1_88 wl0_89 wl1_89 wl0_90 wl1_90 wl0_91 wl1_91 wl0_92 wl1_92 wl0_93 wl1_93 wl0_94 wl1_94 wl0_95 wl1_95 wl0_96 wl1_96 wl0_97 wl1_97 wl0_98 wl1_98 wl0_99 wl1_99 wl0_100 wl1_100 wl0_101 wl1_101 wl0_102 wl1_102 wl0_103 wl1_103 wl0_104 wl1_104 wl0_105 wl1_105 wl0_106 wl1_106 wl0_107 wl1_107 wl0_108 wl1_108 wl0_109 wl1_109 wl0_110 wl1_110 wl0_111 wl1_111 wl0_112 wl1_112 wl0_113 wl1_113 wl0_114 wl1_114 wl0_115 wl1_115 wl0_116 wl1_116 wl0_117 wl1_117 wl0_118 wl1_118 wl0_119 wl1_119 wl0_120 wl1_120 wl0_121 wl1_121 wl0_122 wl1_122 wl0_123 wl1_123 wl0_124 wl1_124 wl0_125 wl1_125 wl0_126 wl1_126 wl0_127 wl1_127 gnd rbl_wl1_1 dummy_wl0_top dummy_wl1_top vdd gnd replica_column
Xreplica_col_1 rbl_bl0_1 rbl_br0_1 rbl_bl1_1 rbl_br1_1 dummy_wl0_bot dummy_wl1_bot rbl_wl0_0 gnd wl0_0 wl1_0 wl0_1 wl1_1 wl0_2 wl1_2 wl0_3 wl1_3 wl0_4 wl1_4 wl0_5 wl1_5 wl0_6 wl1_6 wl0_7 wl1_7 wl0_8 wl1_8 wl0_9 wl1_9 wl0_10 wl1_10 wl0_11 wl1_11 wl0_12 wl1_12 wl0_13 wl1_13 wl0_14 wl1_14 wl0_15 wl1_15 wl0_16 wl1_16 wl0_17 wl1_17 wl0_18 wl1_18 wl0_19 wl1_19 wl0_20 wl1_20 wl0_21 wl1_21 wl0_22 wl1_22 wl0_23 wl1_23 wl0_24 wl1_24 wl0_25 wl1_25 wl0_26 wl1_26 wl0_27 wl1_27 wl0_28 wl1_28 wl0_29 wl1_29 wl0_30 wl1_30 wl0_31 wl1_31 wl0_32 wl1_32 wl0_33 wl1_33 wl0_34 wl1_34 wl0_35 wl1_35 wl0_36 wl1_36 wl0_37 wl1_37 wl0_38 wl1_38 wl0_39 wl1_39 wl0_40 wl1_40 wl0_41 wl1_41 wl0_42 wl1_42 wl0_43 wl1_43 wl0_44 wl1_44 wl0_45 wl1_45 wl0_46 wl1_46 wl0_47 wl1_47 wl0_48 wl1_48 wl0_49 wl1_49 wl0_50 wl1_50 wl0_51 wl1_51 wl0_52 wl1_52 wl0_53 wl1_53 wl0_54 wl1_54 wl0_55 wl1_55 wl0_56 wl1_56 wl0_57 wl1_57 wl0_58 wl1_58 wl0_59 wl1_59 wl0_60 wl1_60 wl0_61 wl1_61 wl0_62 wl1_62 wl0_63 wl1_63 wl0_64 wl1_64 wl0_65 wl1_65 wl0_66 wl1_66 wl0_67 wl1_67 wl0_68 wl1_68 wl0_69 wl1_69 wl0_70 wl1_70 wl0_71 wl1_71 wl0_72 wl1_72 wl0_73 wl1_73 wl0_74 wl1_74 wl0_75 wl1_75 wl0_76 wl1_76 wl0_77 wl1_77 wl0_78 wl1_78 wl0_79 wl1_79 wl0_80 wl1_80 wl0_81 wl1_81 wl0_82 wl1_82 wl0_83 wl1_83 wl0_84 wl1_84 wl0_85 wl1_85 wl0_86 wl1_86 wl0_87 wl1_87 wl0_88 wl1_88 wl0_89 wl1_89 wl0_90 wl1_90 wl0_91 wl1_91 wl0_92 wl1_92 wl0_93 wl1_93 wl0_94 wl1_94 wl0_95 wl1_95 wl0_96 wl1_96 wl0_97 wl1_97 wl0_98 wl1_98 wl0_99 wl1_99 wl0_100 wl1_100 wl0_101 wl1_101 wl0_102 wl1_102 wl0_103 wl1_103 wl0_104 wl1_104 wl0_105 wl1_105 wl0_106 wl1_106 wl0_107 wl1_107 wl0_108 wl1_108 wl0_109 wl1_109 wl0_110 wl1_110 wl0_111 wl1_111 wl0_112 wl1_112 wl0_113 wl1_113 wl0_114 wl1_114 wl0_115 wl1_115 wl0_116 wl1_116 wl0_117 wl1_117 wl0_118 wl1_118 wl0_119 wl1_119 wl0_120 wl1_120 wl0_121 wl1_121 wl0_122 wl1_122 wl0_123 wl1_123 wl0_124 wl1_124 wl0_125 wl1_125 wl0_126 wl1_126 wl0_127 wl1_127 gnd rbl_wl1_1 dummy_wl0_top dummy_wl1_top vdd gnd replica_column_0
Xdummy_row_0 bl0_0 br0_0 bl1_0 br1_0 bl0_1 br0_1 bl1_1 br1_1 bl0_2 br0_2 bl1_2 br1_2 bl0_3 br0_3 bl1_3 br1_3 bl0_4 br0_4 bl1_4 br1_4 bl0_5 br0_5 bl1_5 br1_5 bl0_6 br0_6 bl1_6 br1_6 bl0_7 br0_7 bl1_7 br1_7 bl0_8 br0_8 bl1_8 br1_8 bl0_9 br0_9 bl1_9 br1_9 bl0_10 br0_10 bl1_10 br1_10 bl0_11 br0_11 bl1_11 br1_11 bl0_12 br0_12 bl1_12 br1_12 bl0_13 br0_13 bl1_13 br1_13 bl0_14 br0_14 bl1_14 br1_14 bl0_15 br0_15 bl1_15 br1_15 bl0_16 br0_16 bl1_16 br1_16 bl0_17 br0_17 bl1_17 br1_17 bl0_18 br0_18 bl1_18 br1_18 bl0_19 br0_19 bl1_19 br1_19 bl0_20 br0_20 bl1_20 br1_20 bl0_21 br0_21 bl1_21 br1_21 bl0_22 br0_22 bl1_22 br1_22 bl0_23 br0_23 bl1_23 br1_23 bl0_24 br0_24 bl1_24 br1_24 bl0_25 br0_25 bl1_25 br1_25 bl0_26 br0_26 bl1_26 br1_26 bl0_27 br0_27 bl1_27 br1_27 bl0_28 br0_28 bl1_28 br1_28 bl0_29 br0_29 bl1_29 br1_29 bl0_30 br0_30 bl1_30 br1_30 bl0_31 br0_31 bl1_31 br1_31 bl0_32 br0_32 bl1_32 br1_32 bl0_33 br0_33 bl1_33 br1_33 bl0_34 br0_34 bl1_34 br1_34 bl0_35 br0_35 bl1_35 br1_35 bl0_36 br0_36 bl1_36 br1_36 bl0_37 br0_37 bl1_37 br1_37 bl0_38 br0_38 bl1_38 br1_38 bl0_39 br0_39 bl1_39 br1_39 bl0_40 br0_40 bl1_40 br1_40 bl0_41 br0_41 bl1_41 br1_41 bl0_42 br0_42 bl1_42 br1_42 bl0_43 br0_43 bl1_43 br1_43 bl0_44 br0_44 bl1_44 br1_44 bl0_45 br0_45 bl1_45 br1_45 bl0_46 br0_46 bl1_46 br1_46 bl0_47 br0_47 bl1_47 br1_47 bl0_48 br0_48 bl1_48 br1_48 bl0_49 br0_49 bl1_49 br1_49 bl0_50 br0_50 bl1_50 br1_50 bl0_51 br0_51 bl1_51 br1_51 bl0_52 br0_52 bl1_52 br1_52 bl0_53 br0_53 bl1_53 br1_53 bl0_54 br0_54 bl1_54 br1_54 bl0_55 br0_55 bl1_55 br1_55 bl0_56 br0_56 bl1_56 br1_56 bl0_57 br0_57 bl1_57 br1_57 bl0_58 br0_58 bl1_58 br1_58 bl0_59 br0_59 bl1_59 br1_59 bl0_60 br0_60 bl1_60 br1_60 bl0_61 br0_61 bl1_61 br1_61 bl0_62 br0_62 bl1_62 br1_62 bl0_63 br0_63 bl1_63 br1_63 rbl_wl0_0 gnd vdd gnd dummy_array
Xdummy_row_1 bl0_0 br0_0 bl1_0 br1_0 bl0_1 br0_1 bl1_1 br1_1 bl0_2 br0_2 bl1_2 br1_2 bl0_3 br0_3 bl1_3 br1_3 bl0_4 br0_4 bl1_4 br1_4 bl0_5 br0_5 bl1_5 br1_5 bl0_6 br0_6 bl1_6 br1_6 bl0_7 br0_7 bl1_7 br1_7 bl0_8 br0_8 bl1_8 br1_8 bl0_9 br0_9 bl1_9 br1_9 bl0_10 br0_10 bl1_10 br1_10 bl0_11 br0_11 bl1_11 br1_11 bl0_12 br0_12 bl1_12 br1_12 bl0_13 br0_13 bl1_13 br1_13 bl0_14 br0_14 bl1_14 br1_14 bl0_15 br0_15 bl1_15 br1_15 bl0_16 br0_16 bl1_16 br1_16 bl0_17 br0_17 bl1_17 br1_17 bl0_18 br0_18 bl1_18 br1_18 bl0_19 br0_19 bl1_19 br1_19 bl0_20 br0_20 bl1_20 br1_20 bl0_21 br0_21 bl1_21 br1_21 bl0_22 br0_22 bl1_22 br1_22 bl0_23 br0_23 bl1_23 br1_23 bl0_24 br0_24 bl1_24 br1_24 bl0_25 br0_25 bl1_25 br1_25 bl0_26 br0_26 bl1_26 br1_26 bl0_27 br0_27 bl1_27 br1_27 bl0_28 br0_28 bl1_28 br1_28 bl0_29 br0_29 bl1_29 br1_29 bl0_30 br0_30 bl1_30 br1_30 bl0_31 br0_31 bl1_31 br1_31 bl0_32 br0_32 bl1_32 br1_32 bl0_33 br0_33 bl1_33 br1_33 bl0_34 br0_34 bl1_34 br1_34 bl0_35 br0_35 bl1_35 br1_35 bl0_36 br0_36 bl1_36 br1_36 bl0_37 br0_37 bl1_37 br1_37 bl0_38 br0_38 bl1_38 br1_38 bl0_39 br0_39 bl1_39 br1_39 bl0_40 br0_40 bl1_40 br1_40 bl0_41 br0_41 bl1_41 br1_41 bl0_42 br0_42 bl1_42 br1_42 bl0_43 br0_43 bl1_43 br1_43 bl0_44 br0_44 bl1_44 br1_44 bl0_45 br0_45 bl1_45 br1_45 bl0_46 br0_46 bl1_46 br1_46 bl0_47 br0_47 bl1_47 br1_47 bl0_48 br0_48 bl1_48 br1_48 bl0_49 br0_49 bl1_49 br1_49 bl0_50 br0_50 bl1_50 br1_50 bl0_51 br0_51 bl1_51 br1_51 bl0_52 br0_52 bl1_52 br1_52 bl0_53 br0_53 bl1_53 br1_53 bl0_54 br0_54 bl1_54 br1_54 bl0_55 br0_55 bl1_55 br1_55 bl0_56 br0_56 bl1_56 br1_56 bl0_57 br0_57 bl1_57 br1_57 bl0_58 br0_58 bl1_58 br1_58 bl0_59 br0_59 bl1_59 br1_59 bl0_60 br0_60 bl1_60 br1_60 bl0_61 br0_61 bl1_61 br1_61 bl0_62 br0_62 bl1_62 br1_62 bl0_63 br0_63 bl1_63 br1_63 gnd rbl_wl1_1 vdd gnd dummy_array
.ENDS replica_bitcell_array

.SUBCKT pinv_0 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u
.ENDS pinv_0

.SUBCKT pinv_1 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS pinv_1

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=1.68 l=0.15 pd=3.66 ps=3.66 as=0.63u ad=0.63u

* ptx M{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=1.65 l=0.15 pd=3.60 ps=3.60 as=0.62u ad=0.62u

.SUBCKT pinv_2 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.65 l=0.15 pd=3.60 ps=3.60 as=0.62u ad=0.62u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=1.68 l=0.15 pd=3.66 ps=3.66 as=0.63u ad=0.63u
.ENDS pinv_2

.SUBCKT pinvbuf A Zb Z vdd gnd
* INOUT : A 
* INOUT : Zb 
* INOUT : Z 
* INOUT : vdd 
* INOUT : gnd 
Xbuf_inv1 A zb_int vdd gnd pinv_0
Xbuf_inv2 zb_int z_int vdd gnd pinv_1
Xbuf_inv3 z_int Zb vdd gnd pinv_2
Xbuf_inv4 zb_int Z vdd gnd pinv_2
.ENDS pinvbuf

.SUBCKT bank dout0_0 dout0_1 dout0_2 dout0_3 dout0_4 dout0_5 dout0_6 dout0_7 dout0_8 dout0_9 dout0_10 dout0_11 dout0_12 dout0_13 dout0_14 dout0_15 dout0_16 dout0_17 dout0_18 dout0_19 dout0_20 dout0_21 dout0_22 dout0_23 dout0_24 dout0_25 dout0_26 dout0_27 dout0_28 dout0_29 dout0_30 dout0_31 dout1_0 dout1_1 dout1_2 dout1_3 dout1_4 dout1_5 dout1_6 dout1_7 dout1_8 dout1_9 dout1_10 dout1_11 dout1_12 dout1_13 dout1_14 dout1_15 dout1_16 dout1_17 dout1_18 dout1_19 dout1_20 dout1_21 dout1_22 dout1_23 dout1_24 dout1_25 dout1_26 dout1_27 dout1_28 dout1_29 dout1_30 dout1_31 rbl_bl0_0 rbl_bl1_1 din0_0 din0_1 din0_2 din0_3 din0_4 din0_5 din0_6 din0_7 din0_8 din0_9 din0_10 din0_11 din0_12 din0_13 din0_14 din0_15 din0_16 din0_17 din0_18 din0_19 din0_20 din0_21 din0_22 din0_23 din0_24 din0_25 din0_26 din0_27 din0_28 din0_29 din0_30 din0_31 addr0_0 addr0_1 addr0_2 addr0_3 addr0_4 addr0_5 addr0_6 addr0_7 addr1_0 addr1_1 addr1_2 addr1_3 addr1_4 addr1_5 addr1_6 addr1_7 s_en0 s_en1 p_en_bar0 p_en_bar1 w_en0 bank_wmask0_0 bank_wmask0_1 bank_wmask0_2 bank_wmask0_3 wl_en0 wl_en1 vdd gnd
* OUTPUT: dout0_0 
* OUTPUT: dout0_1 
* OUTPUT: dout0_2 
* OUTPUT: dout0_3 
* OUTPUT: dout0_4 
* OUTPUT: dout0_5 
* OUTPUT: dout0_6 
* OUTPUT: dout0_7 
* OUTPUT: dout0_8 
* OUTPUT: dout0_9 
* OUTPUT: dout0_10 
* OUTPUT: dout0_11 
* OUTPUT: dout0_12 
* OUTPUT: dout0_13 
* OUTPUT: dout0_14 
* OUTPUT: dout0_15 
* OUTPUT: dout0_16 
* OUTPUT: dout0_17 
* OUTPUT: dout0_18 
* OUTPUT: dout0_19 
* OUTPUT: dout0_20 
* OUTPUT: dout0_21 
* OUTPUT: dout0_22 
* OUTPUT: dout0_23 
* OUTPUT: dout0_24 
* OUTPUT: dout0_25 
* OUTPUT: dout0_26 
* OUTPUT: dout0_27 
* OUTPUT: dout0_28 
* OUTPUT: dout0_29 
* OUTPUT: dout0_30 
* OUTPUT: dout0_31 
* OUTPUT: dout1_0 
* OUTPUT: dout1_1 
* OUTPUT: dout1_2 
* OUTPUT: dout1_3 
* OUTPUT: dout1_4 
* OUTPUT: dout1_5 
* OUTPUT: dout1_6 
* OUTPUT: dout1_7 
* OUTPUT: dout1_8 
* OUTPUT: dout1_9 
* OUTPUT: dout1_10 
* OUTPUT: dout1_11 
* OUTPUT: dout1_12 
* OUTPUT: dout1_13 
* OUTPUT: dout1_14 
* OUTPUT: dout1_15 
* OUTPUT: dout1_16 
* OUTPUT: dout1_17 
* OUTPUT: dout1_18 
* OUTPUT: dout1_19 
* OUTPUT: dout1_20 
* OUTPUT: dout1_21 
* OUTPUT: dout1_22 
* OUTPUT: dout1_23 
* OUTPUT: dout1_24 
* OUTPUT: dout1_25 
* OUTPUT: dout1_26 
* OUTPUT: dout1_27 
* OUTPUT: dout1_28 
* OUTPUT: dout1_29 
* OUTPUT: dout1_30 
* OUTPUT: dout1_31 
* OUTPUT: rbl_bl0_0 
* OUTPUT: rbl_bl1_1 
* INPUT : din0_0 
* INPUT : din0_1 
* INPUT : din0_2 
* INPUT : din0_3 
* INPUT : din0_4 
* INPUT : din0_5 
* INPUT : din0_6 
* INPUT : din0_7 
* INPUT : din0_8 
* INPUT : din0_9 
* INPUT : din0_10 
* INPUT : din0_11 
* INPUT : din0_12 
* INPUT : din0_13 
* INPUT : din0_14 
* INPUT : din0_15 
* INPUT : din0_16 
* INPUT : din0_17 
* INPUT : din0_18 
* INPUT : din0_19 
* INPUT : din0_20 
* INPUT : din0_21 
* INPUT : din0_22 
* INPUT : din0_23 
* INPUT : din0_24 
* INPUT : din0_25 
* INPUT : din0_26 
* INPUT : din0_27 
* INPUT : din0_28 
* INPUT : din0_29 
* INPUT : din0_30 
* INPUT : din0_31 
* INPUT : addr0_0 
* INPUT : addr0_1 
* INPUT : addr0_2 
* INPUT : addr0_3 
* INPUT : addr0_4 
* INPUT : addr0_5 
* INPUT : addr0_6 
* INPUT : addr0_7 
* INPUT : addr1_0 
* INPUT : addr1_1 
* INPUT : addr1_2 
* INPUT : addr1_3 
* INPUT : addr1_4 
* INPUT : addr1_5 
* INPUT : addr1_6 
* INPUT : addr1_7 
* INPUT : s_en0 
* INPUT : s_en1 
* INPUT : p_en_bar0 
* INPUT : p_en_bar1 
* INPUT : w_en0 
* INPUT : bank_wmask0_0 
* INPUT : bank_wmask0_1 
* INPUT : bank_wmask0_2 
* INPUT : bank_wmask0_3 
* INPUT : wl_en0 
* INPUT : wl_en1 
* POWER : vdd 
* GROUND: gnd 
Xreplica_bitcell_array bl0_0 br0_0 bl1_0 br1_0 bl0_1 br0_1 bl1_1 br1_1 bl0_2 br0_2 bl1_2 br1_2 bl0_3 br0_3 bl1_3 br1_3 bl0_4 br0_4 bl1_4 br1_4 bl0_5 br0_5 bl1_5 br1_5 bl0_6 br0_6 bl1_6 br1_6 bl0_7 br0_7 bl1_7 br1_7 bl0_8 br0_8 bl1_8 br1_8 bl0_9 br0_9 bl1_9 br1_9 bl0_10 br0_10 bl1_10 br1_10 bl0_11 br0_11 bl1_11 br1_11 bl0_12 br0_12 bl1_12 br1_12 bl0_13 br0_13 bl1_13 br1_13 bl0_14 br0_14 bl1_14 br1_14 bl0_15 br0_15 bl1_15 br1_15 bl0_16 br0_16 bl1_16 br1_16 bl0_17 br0_17 bl1_17 br1_17 bl0_18 br0_18 bl1_18 br1_18 bl0_19 br0_19 bl1_19 br1_19 bl0_20 br0_20 bl1_20 br1_20 bl0_21 br0_21 bl1_21 br1_21 bl0_22 br0_22 bl1_22 br1_22 bl0_23 br0_23 bl1_23 br1_23 bl0_24 br0_24 bl1_24 br1_24 bl0_25 br0_25 bl1_25 br1_25 bl0_26 br0_26 bl1_26 br1_26 bl0_27 br0_27 bl1_27 br1_27 bl0_28 br0_28 bl1_28 br1_28 bl0_29 br0_29 bl1_29 br1_29 bl0_30 br0_30 bl1_30 br1_30 bl0_31 br0_31 bl1_31 br1_31 bl0_32 br0_32 bl1_32 br1_32 bl0_33 br0_33 bl1_33 br1_33 bl0_34 br0_34 bl1_34 br1_34 bl0_35 br0_35 bl1_35 br1_35 bl0_36 br0_36 bl1_36 br1_36 bl0_37 br0_37 bl1_37 br1_37 bl0_38 br0_38 bl1_38 br1_38 bl0_39 br0_39 bl1_39 br1_39 bl0_40 br0_40 bl1_40 br1_40 bl0_41 br0_41 bl1_41 br1_41 bl0_42 br0_42 bl1_42 br1_42 bl0_43 br0_43 bl1_43 br1_43 bl0_44 br0_44 bl1_44 br1_44 bl0_45 br0_45 bl1_45 br1_45 bl0_46 br0_46 bl1_46 br1_46 bl0_47 br0_47 bl1_47 br1_47 bl0_48 br0_48 bl1_48 br1_48 bl0_49 br0_49 bl1_49 br1_49 bl0_50 br0_50 bl1_50 br1_50 bl0_51 br0_51 bl1_51 br1_51 bl0_52 br0_52 bl1_52 br1_52 bl0_53 br0_53 bl1_53 br1_53 bl0_54 br0_54 bl1_54 br1_54 bl0_55 br0_55 bl1_55 br1_55 bl0_56 br0_56 bl1_56 br1_56 bl0_57 br0_57 bl1_57 br1_57 bl0_58 br0_58 bl1_58 br1_58 bl0_59 br0_59 bl1_59 br1_59 bl0_60 br0_60 bl1_60 br1_60 bl0_61 br0_61 bl1_61 br1_61 bl0_62 br0_62 bl1_62 br1_62 bl0_63 br0_63 bl1_63 br1_63 rbl_bl0_0 rbl_br0_0 rbl_bl1_1 rbl_br1_1 wl0_0 wl1_0 wl0_1 wl1_1 wl0_2 wl1_2 wl0_3 wl1_3 wl0_4 wl1_4 wl0_5 wl1_5 wl0_6 wl1_6 wl0_7 wl1_7 wl0_8 wl1_8 wl0_9 wl1_9 wl0_10 wl1_10 wl0_11 wl1_11 wl0_12 wl1_12 wl0_13 wl1_13 wl0_14 wl1_14 wl0_15 wl1_15 wl0_16 wl1_16 wl0_17 wl1_17 wl0_18 wl1_18 wl0_19 wl1_19 wl0_20 wl1_20 wl0_21 wl1_21 wl0_22 wl1_22 wl0_23 wl1_23 wl0_24 wl1_24 wl0_25 wl1_25 wl0_26 wl1_26 wl0_27 wl1_27 wl0_28 wl1_28 wl0_29 wl1_29 wl0_30 wl1_30 wl0_31 wl1_31 wl0_32 wl1_32 wl0_33 wl1_33 wl0_34 wl1_34 wl0_35 wl1_35 wl0_36 wl1_36 wl0_37 wl1_37 wl0_38 wl1_38 wl0_39 wl1_39 wl0_40 wl1_40 wl0_41 wl1_41 wl0_42 wl1_42 wl0_43 wl1_43 wl0_44 wl1_44 wl0_45 wl1_45 wl0_46 wl1_46 wl0_47 wl1_47 wl0_48 wl1_48 wl0_49 wl1_49 wl0_50 wl1_50 wl0_51 wl1_51 wl0_52 wl1_52 wl0_53 wl1_53 wl0_54 wl1_54 wl0_55 wl1_55 wl0_56 wl1_56 wl0_57 wl1_57 wl0_58 wl1_58 wl0_59 wl1_59 wl0_60 wl1_60 wl0_61 wl1_61 wl0_62 wl1_62 wl0_63 wl1_63 wl0_64 wl1_64 wl0_65 wl1_65 wl0_66 wl1_66 wl0_67 wl1_67 wl0_68 wl1_68 wl0_69 wl1_69 wl0_70 wl1_70 wl0_71 wl1_71 wl0_72 wl1_72 wl0_73 wl1_73 wl0_74 wl1_74 wl0_75 wl1_75 wl0_76 wl1_76 wl0_77 wl1_77 wl0_78 wl1_78 wl0_79 wl1_79 wl0_80 wl1_80 wl0_81 wl1_81 wl0_82 wl1_82 wl0_83 wl1_83 wl0_84 wl1_84 wl0_85 wl1_85 wl0_86 wl1_86 wl0_87 wl1_87 wl0_88 wl1_88 wl0_89 wl1_89 wl0_90 wl1_90 wl0_91 wl1_91 wl0_92 wl1_92 wl0_93 wl1_93 wl0_94 wl1_94 wl0_95 wl1_95 wl0_96 wl1_96 wl0_97 wl1_97 wl0_98 wl1_98 wl0_99 wl1_99 wl0_100 wl1_100 wl0_101 wl1_101 wl0_102 wl1_102 wl0_103 wl1_103 wl0_104 wl1_104 wl0_105 wl1_105 wl0_106 wl1_106 wl0_107 wl1_107 wl0_108 wl1_108 wl0_109 wl1_109 wl0_110 wl1_110 wl0_111 wl1_111 wl0_112 wl1_112 wl0_113 wl1_113 wl0_114 wl1_114 wl0_115 wl1_115 wl0_116 wl1_116 wl0_117 wl1_117 wl0_118 wl1_118 wl0_119 wl1_119 wl0_120 wl1_120 wl0_121 wl1_121 wl0_122 wl1_122 wl0_123 wl1_123 wl0_124 wl1_124 wl0_125 wl1_125 wl0_126 wl1_126 wl0_127 wl1_127 wl_en0 wl_en1 vdd gnd replica_bitcell_array
Xport_data0 rbl_bl0_0 rbl_br0_0 bl0_0 br0_0 bl0_1 br0_1 bl0_2 br0_2 bl0_3 br0_3 bl0_4 br0_4 bl0_5 br0_5 bl0_6 br0_6 bl0_7 br0_7 bl0_8 br0_8 bl0_9 br0_9 bl0_10 br0_10 bl0_11 br0_11 bl0_12 br0_12 bl0_13 br0_13 bl0_14 br0_14 bl0_15 br0_15 bl0_16 br0_16 bl0_17 br0_17 bl0_18 br0_18 bl0_19 br0_19 bl0_20 br0_20 bl0_21 br0_21 bl0_22 br0_22 bl0_23 br0_23 bl0_24 br0_24 bl0_25 br0_25 bl0_26 br0_26 bl0_27 br0_27 bl0_28 br0_28 bl0_29 br0_29 bl0_30 br0_30 bl0_31 br0_31 bl0_32 br0_32 bl0_33 br0_33 bl0_34 br0_34 bl0_35 br0_35 bl0_36 br0_36 bl0_37 br0_37 bl0_38 br0_38 bl0_39 br0_39 bl0_40 br0_40 bl0_41 br0_41 bl0_42 br0_42 bl0_43 br0_43 bl0_44 br0_44 bl0_45 br0_45 bl0_46 br0_46 bl0_47 br0_47 bl0_48 br0_48 bl0_49 br0_49 bl0_50 br0_50 bl0_51 br0_51 bl0_52 br0_52 bl0_53 br0_53 bl0_54 br0_54 bl0_55 br0_55 bl0_56 br0_56 bl0_57 br0_57 bl0_58 br0_58 bl0_59 br0_59 bl0_60 br0_60 bl0_61 br0_61 bl0_62 br0_62 bl0_63 br0_63 dout0_0 dout0_1 dout0_2 dout0_3 dout0_4 dout0_5 dout0_6 dout0_7 dout0_8 dout0_9 dout0_10 dout0_11 dout0_12 dout0_13 dout0_14 dout0_15 dout0_16 dout0_17 dout0_18 dout0_19 dout0_20 dout0_21 dout0_22 dout0_23 dout0_24 dout0_25 dout0_26 dout0_27 dout0_28 dout0_29 dout0_30 dout0_31 din0_0 din0_1 din0_2 din0_3 din0_4 din0_5 din0_6 din0_7 din0_8 din0_9 din0_10 din0_11 din0_12 din0_13 din0_14 din0_15 din0_16 din0_17 din0_18 din0_19 din0_20 din0_21 din0_22 din0_23 din0_24 din0_25 din0_26 din0_27 din0_28 din0_29 din0_30 din0_31 sel0_0 sel0_1 s_en0 p_en_bar0 w_en0 bank_wmask0_0 bank_wmask0_1 bank_wmask0_2 bank_wmask0_3 vdd gnd port_data
Xport_data1 rbl_bl1_1 rbl_br1_1 bl1_0 br1_0 bl1_1 br1_1 bl1_2 br1_2 bl1_3 br1_3 bl1_4 br1_4 bl1_5 br1_5 bl1_6 br1_6 bl1_7 br1_7 bl1_8 br1_8 bl1_9 br1_9 bl1_10 br1_10 bl1_11 br1_11 bl1_12 br1_12 bl1_13 br1_13 bl1_14 br1_14 bl1_15 br1_15 bl1_16 br1_16 bl1_17 br1_17 bl1_18 br1_18 bl1_19 br1_19 bl1_20 br1_20 bl1_21 br1_21 bl1_22 br1_22 bl1_23 br1_23 bl1_24 br1_24 bl1_25 br1_25 bl1_26 br1_26 bl1_27 br1_27 bl1_28 br1_28 bl1_29 br1_29 bl1_30 br1_30 bl1_31 br1_31 bl1_32 br1_32 bl1_33 br1_33 bl1_34 br1_34 bl1_35 br1_35 bl1_36 br1_36 bl1_37 br1_37 bl1_38 br1_38 bl1_39 br1_39 bl1_40 br1_40 bl1_41 br1_41 bl1_42 br1_42 bl1_43 br1_43 bl1_44 br1_44 bl1_45 br1_45 bl1_46 br1_46 bl1_47 br1_47 bl1_48 br1_48 bl1_49 br1_49 bl1_50 br1_50 bl1_51 br1_51 bl1_52 br1_52 bl1_53 br1_53 bl1_54 br1_54 bl1_55 br1_55 bl1_56 br1_56 bl1_57 br1_57 bl1_58 br1_58 bl1_59 br1_59 bl1_60 br1_60 bl1_61 br1_61 bl1_62 br1_62 bl1_63 br1_63 dout1_0 dout1_1 dout1_2 dout1_3 dout1_4 dout1_5 dout1_6 dout1_7 dout1_8 dout1_9 dout1_10 dout1_11 dout1_12 dout1_13 dout1_14 dout1_15 dout1_16 dout1_17 dout1_18 dout1_19 dout1_20 dout1_21 dout1_22 dout1_23 dout1_24 dout1_25 dout1_26 dout1_27 dout1_28 dout1_29 dout1_30 dout1_31 sel1_0 sel1_1 s_en1 p_en_bar1 vdd gnd port_data_0
Xport_address0 addr0_1 addr0_2 addr0_3 addr0_4 addr0_5 addr0_6 addr0_7 wl_en0 wl0_0 wl0_1 wl0_2 wl0_3 wl0_4 wl0_5 wl0_6 wl0_7 wl0_8 wl0_9 wl0_10 wl0_11 wl0_12 wl0_13 wl0_14 wl0_15 wl0_16 wl0_17 wl0_18 wl0_19 wl0_20 wl0_21 wl0_22 wl0_23 wl0_24 wl0_25 wl0_26 wl0_27 wl0_28 wl0_29 wl0_30 wl0_31 wl0_32 wl0_33 wl0_34 wl0_35 wl0_36 wl0_37 wl0_38 wl0_39 wl0_40 wl0_41 wl0_42 wl0_43 wl0_44 wl0_45 wl0_46 wl0_47 wl0_48 wl0_49 wl0_50 wl0_51 wl0_52 wl0_53 wl0_54 wl0_55 wl0_56 wl0_57 wl0_58 wl0_59 wl0_60 wl0_61 wl0_62 wl0_63 wl0_64 wl0_65 wl0_66 wl0_67 wl0_68 wl0_69 wl0_70 wl0_71 wl0_72 wl0_73 wl0_74 wl0_75 wl0_76 wl0_77 wl0_78 wl0_79 wl0_80 wl0_81 wl0_82 wl0_83 wl0_84 wl0_85 wl0_86 wl0_87 wl0_88 wl0_89 wl0_90 wl0_91 wl0_92 wl0_93 wl0_94 wl0_95 wl0_96 wl0_97 wl0_98 wl0_99 wl0_100 wl0_101 wl0_102 wl0_103 wl0_104 wl0_105 wl0_106 wl0_107 wl0_108 wl0_109 wl0_110 wl0_111 wl0_112 wl0_113 wl0_114 wl0_115 wl0_116 wl0_117 wl0_118 wl0_119 wl0_120 wl0_121 wl0_122 wl0_123 wl0_124 wl0_125 wl0_126 wl0_127 vdd gnd port_address
Xport_address1 addr1_1 addr1_2 addr1_3 addr1_4 addr1_5 addr1_6 addr1_7 wl_en1 wl1_0 wl1_1 wl1_2 wl1_3 wl1_4 wl1_5 wl1_6 wl1_7 wl1_8 wl1_9 wl1_10 wl1_11 wl1_12 wl1_13 wl1_14 wl1_15 wl1_16 wl1_17 wl1_18 wl1_19 wl1_20 wl1_21 wl1_22 wl1_23 wl1_24 wl1_25 wl1_26 wl1_27 wl1_28 wl1_29 wl1_30 wl1_31 wl1_32 wl1_33 wl1_34 wl1_35 wl1_36 wl1_37 wl1_38 wl1_39 wl1_40 wl1_41 wl1_42 wl1_43 wl1_44 wl1_45 wl1_46 wl1_47 wl1_48 wl1_49 wl1_50 wl1_51 wl1_52 wl1_53 wl1_54 wl1_55 wl1_56 wl1_57 wl1_58 wl1_59 wl1_60 wl1_61 wl1_62 wl1_63 wl1_64 wl1_65 wl1_66 wl1_67 wl1_68 wl1_69 wl1_70 wl1_71 wl1_72 wl1_73 wl1_74 wl1_75 wl1_76 wl1_77 wl1_78 wl1_79 wl1_80 wl1_81 wl1_82 wl1_83 wl1_84 wl1_85 wl1_86 wl1_87 wl1_88 wl1_89 wl1_90 wl1_91 wl1_92 wl1_93 wl1_94 wl1_95 wl1_96 wl1_97 wl1_98 wl1_99 wl1_100 wl1_101 wl1_102 wl1_103 wl1_104 wl1_105 wl1_106 wl1_107 wl1_108 wl1_109 wl1_110 wl1_111 wl1_112 wl1_113 wl1_114 wl1_115 wl1_116 wl1_117 wl1_118 wl1_119 wl1_120 wl1_121 wl1_122 wl1_123 wl1_124 wl1_125 wl1_126 wl1_127 vdd gnd port_address
Xcol_address_decoder0 addr0_0 sel0_0 sel0_1 vdd gnd pinvbuf
Xcol_address_decoder1 addr1_0 sel1_0 sel1_1 vdd gnd pinvbuf
.ENDS bank

.SUBCKT dff_buf_0 D Q Qb clk vdd gnd
* INPUT : D 
* OUTPUT: Q 
* OUTPUT: Qb 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* inv1: 2 inv2: 4
Xdff_buf_dff D qint clk vdd gnd dff
Xdff_buf_inv1 qint Qb vdd gnd pinv_1
Xdff_buf_inv2 Qb Q vdd gnd pinv_2
.ENDS dff_buf_0

.SUBCKT dff_buf_array din_0 din_1 dout_0 dout_bar_0 dout_1 dout_bar_1 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* OUTPUT: dout_0 
* OUTPUT: dout_bar_0 
* OUTPUT: dout_1 
* OUTPUT: dout_bar_1 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* inv1: 2 inv2: 4
Xdff_r0_c0 din_0 dout_0 dout_bar_0 clk vdd gnd dff_buf_0
Xdff_r1_c0 din_1 dout_1 dout_bar_1 clk vdd gnd dff_buf_0
.ENDS dff_buf_array

.SUBCKT pnand2_0 A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpnand2_pmos1 vdd A Z vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
XMpnand2_pmos2 Z B vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
XMpnand2_nmos1 Z B net1 gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
XMpnand2_nmos2 net1 A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS pnand2_0

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=1.68 l=0.15 pd=3.66 ps=3.66 as=0.63u ad=0.63u

* ptx M{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_3 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=1.68 l=0.15 pd=3.66 ps=3.66 as=0.63u ad=0.63u
.ENDS pinv_3

.SUBCKT pdriver_0 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [12]
Xbuf_inv1 A Z vdd gnd pinv_3
.ENDS pdriver_0

.SUBCKT pand2_0 A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpand2_nand A B zb_int vdd gnd pnand2_0
Xpand2_inv zb_int Z vdd gnd pdriver_0
.ENDS pand2_0

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

* ptx M{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_4 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS pinv_4

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

* ptx M{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_5 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS pinv_5

.SUBCKT pbuf A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xbuf_inv1 A zb_int vdd gnd pinv_4
Xbuf_inv2 zb_int Z vdd gnd pinv_5
.ENDS pbuf

.SUBCKT pinv_6 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u
.ENDS pinv_6

.SUBCKT pinv_7 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u
.ENDS pinv_7

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=1.26 l=0.15 pd=2.82 ps=2.82 as=0.47u ad=0.47u

* ptx M{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=1.65 l=0.15 pd=3.60 ps=3.60 as=0.62u ad=0.62u

.SUBCKT pinv_8 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.65 l=0.15 pd=3.60 ps=3.60 as=0.62u ad=0.62u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=1.26 l=0.15 pd=2.82 ps=2.82 as=0.47u ad=0.47u
.ENDS pinv_8

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=1.68 l=0.15 pd=3.66 ps=3.66 as=0.63u ad=0.63u

* ptx M{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_9 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=1.68 l=0.15 pd=3.66 ps=3.66 as=0.63u ad=0.63u
.ENDS pinv_9

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

* ptx M{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_10 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS pinv_10

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

* ptx M{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_11 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS pinv_11

.SUBCKT pdriver_1 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 3, 8, 24, 73]
Xbuf_inv1 A Zb1_int vdd gnd pinv_6
Xbuf_inv2 Zb1_int Zb2_int vdd gnd pinv_7
Xbuf_inv3 Zb2_int Zb3_int vdd gnd pinv_8
Xbuf_inv4 Zb3_int Zb4_int vdd gnd pinv_9
Xbuf_inv5 Zb4_int Zb5_int vdd gnd pinv_10
Xbuf_inv6 Zb5_int Z vdd gnd pinv_11
.ENDS pdriver_1

.SUBCKT pinv_12 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS pinv_12

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

* ptx M{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_13 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS pinv_13

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=1.68 l=0.15 pd=3.66 ps=3.66 as=0.63u ad=0.63u

* ptx M{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_14 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=1.68 l=0.15 pd=3.66 ps=3.66 as=0.63u ad=0.63u
.ENDS pinv_14

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

* ptx M{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_15 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS pinv_15

.SUBCKT pdriver_2 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 2, 5, 14, 43]
Xbuf_inv1 A Zb1_int vdd gnd pinv_6
Xbuf_inv2 Zb1_int Zb2_int vdd gnd pinv_7
Xbuf_inv3 Zb2_int Zb3_int vdd gnd pinv_12
Xbuf_inv4 Zb3_int Zb4_int vdd gnd pinv_13
Xbuf_inv5 Zb4_int Zb5_int vdd gnd pinv_14
Xbuf_inv6 Zb5_int Z vdd gnd pinv_15
.ENDS pdriver_2

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u

.SUBCKT pnand3 A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpnand3_pmos1 vdd A Z vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
XMpnand3_pmos2 Z B vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
XMpnand3_pmos3 Z C vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
XMpnand3_nmos1 Z C net1 gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
XMpnand3_nmos2 net1 B net2 gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
XMpnand3_nmos3 net2 A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS pnand3

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

* ptx M{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_16 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS pinv_16

.SUBCKT pdriver_3 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [40]
Xbuf_inv1 A Z vdd gnd pinv_16
.ENDS pdriver_3

.SUBCKT pand3 A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpand3_nand A B C zb_int vdd gnd pnand3
Xpand3_inv zb_int Z vdd gnd pdriver_3
.ENDS pand3

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

* ptx M{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_17 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS pinv_17

.SUBCKT pdriver_4 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [32]
Xbuf_inv1 A Z vdd gnd pinv_17
.ENDS pdriver_4

.SUBCKT pand3_0 A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpand3_nand A B C zb_int vdd gnd pnand3
Xpand3_inv zb_int Z vdd gnd pdriver_4
.ENDS pand3_0

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=1.26 l=0.15 pd=2.82 ps=2.82 as=0.47u ad=0.47u

* ptx M{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_18 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=1.26 l=0.15 pd=2.82 ps=2.82 as=0.47u ad=0.47u
.ENDS pinv_18

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

* ptx M{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_19 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS pinv_19

.SUBCKT pdriver_5 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 2, 7, 21]
Xbuf_inv1 A Zb1_int vdd gnd pinv_6
Xbuf_inv2 Zb1_int Zb2_int vdd gnd pinv_12
Xbuf_inv3 Zb2_int Zb3_int vdd gnd pinv_18
Xbuf_inv4 Zb3_int Z vdd gnd pinv_19
.ENDS pdriver_5

.SUBCKT pnand2_1 A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpnand2_pmos1 vdd A Z vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
XMpnand2_pmos2 Z B vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
XMpnand2_nmos1 Z B net1 gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
XMpnand2_nmos2 net1 A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS pnand2_1

.SUBCKT pinv_20 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u
.ENDS pinv_20

.SUBCKT delay_chain in out vdd gnd
* INPUT : in 
* OUTPUT: out 
* POWER : vdd 
* GROUND: gnd 
* fanouts: [4, 4, 4, 4, 4, 4, 4, 4, 4]
Xdinv0 in dout_1 vdd gnd pinv_20
Xdload_0_0 dout_1 n_0_0 vdd gnd pinv_20
Xdload_0_1 dout_1 n_0_1 vdd gnd pinv_20
Xdload_0_2 dout_1 n_0_2 vdd gnd pinv_20
Xdload_0_3 dout_1 n_0_3 vdd gnd pinv_20
Xdinv1 dout_1 dout_2 vdd gnd pinv_20
Xdload_1_0 dout_2 n_1_0 vdd gnd pinv_20
Xdload_1_1 dout_2 n_1_1 vdd gnd pinv_20
Xdload_1_2 dout_2 n_1_2 vdd gnd pinv_20
Xdload_1_3 dout_2 n_1_3 vdd gnd pinv_20
Xdinv2 dout_2 dout_3 vdd gnd pinv_20
Xdload_2_0 dout_3 n_2_0 vdd gnd pinv_20
Xdload_2_1 dout_3 n_2_1 vdd gnd pinv_20
Xdload_2_2 dout_3 n_2_2 vdd gnd pinv_20
Xdload_2_3 dout_3 n_2_3 vdd gnd pinv_20
Xdinv3 dout_3 dout_4 vdd gnd pinv_20
Xdload_3_0 dout_4 n_3_0 vdd gnd pinv_20
Xdload_3_1 dout_4 n_3_1 vdd gnd pinv_20
Xdload_3_2 dout_4 n_3_2 vdd gnd pinv_20
Xdload_3_3 dout_4 n_3_3 vdd gnd pinv_20
Xdinv4 dout_4 dout_5 vdd gnd pinv_20
Xdload_4_0 dout_5 n_4_0 vdd gnd pinv_20
Xdload_4_1 dout_5 n_4_1 vdd gnd pinv_20
Xdload_4_2 dout_5 n_4_2 vdd gnd pinv_20
Xdload_4_3 dout_5 n_4_3 vdd gnd pinv_20
Xdinv5 dout_5 dout_6 vdd gnd pinv_20
Xdload_5_0 dout_6 n_5_0 vdd gnd pinv_20
Xdload_5_1 dout_6 n_5_1 vdd gnd pinv_20
Xdload_5_2 dout_6 n_5_2 vdd gnd pinv_20
Xdload_5_3 dout_6 n_5_3 vdd gnd pinv_20
Xdinv6 dout_6 dout_7 vdd gnd pinv_20
Xdload_6_0 dout_7 n_6_0 vdd gnd pinv_20
Xdload_6_1 dout_7 n_6_1 vdd gnd pinv_20
Xdload_6_2 dout_7 n_6_2 vdd gnd pinv_20
Xdload_6_3 dout_7 n_6_3 vdd gnd pinv_20
Xdinv7 dout_7 dout_8 vdd gnd pinv_20
Xdload_7_0 dout_8 n_7_0 vdd gnd pinv_20
Xdload_7_1 dout_8 n_7_1 vdd gnd pinv_20
Xdload_7_2 dout_8 n_7_2 vdd gnd pinv_20
Xdload_7_3 dout_8 n_7_3 vdd gnd pinv_20
Xdinv8 dout_8 out vdd gnd pinv_20
Xdload_8_0 out n_8_0 vdd gnd pinv_20
Xdload_8_1 out n_8_1 vdd gnd pinv_20
Xdload_8_2 out n_8_2 vdd gnd pinv_20
Xdload_8_3 out n_8_3 vdd gnd pinv_20
.ENDS delay_chain

.SUBCKT control_logic_rw csb web clk rbl_bl s_en w_en p_en_bar wl_en clk_buf vdd gnd
* INPUT : csb 
* INPUT : web 
* INPUT : clk 
* INPUT : rbl_bl 
* OUTPUT: s_en 
* OUTPUT: w_en 
* OUTPUT: p_en_bar 
* OUTPUT: wl_en 
* OUTPUT: clk_buf 
* POWER : vdd 
* GROUND: gnd 
* word_size 32
Xctrl_dffs csb web cs_bar cs we_bar we clk_buf vdd gnd dff_buf_array
Xclkbuf clk clk_buf vdd gnd pdriver_1
Xinv_clk_bar clk_buf clk_bar vdd gnd pinv_0
Xand2_gated_clk_bar clk_bar cs gated_clk_bar vdd gnd pand2_0
Xand2_gated_clk_buf clk_buf cs gated_clk_buf vdd gnd pand2_0
Xbuf_wl_en gated_clk_bar wl_en vdd gnd pdriver_2
Xrbl_bl_delay_inv rbl_bl_delay rbl_bl_delay_bar vdd gnd pinv_0
Xw_en_and we rbl_bl_delay_bar gated_clk_bar w_en vdd gnd pand3
Xbuf_s_en_and rbl_bl_delay gated_clk_bar we_bar s_en vdd gnd pand3_0
Xdelay_chain rbl_bl rbl_bl_delay vdd gnd delay_chain
Xnand_p_en_bar gated_clk_buf rbl_bl_delay p_en_bar_unbuf vdd gnd pnand2_1
Xbuf_p_en_bar p_en_bar_unbuf p_en_bar vdd gnd pdriver_5
.ENDS control_logic_rw

.SUBCKT dff_buf_array_0 din_0 dout_0 dout_bar_0 clk vdd gnd
* INPUT : din_0 
* OUTPUT: dout_0 
* OUTPUT: dout_bar_0 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* inv1: 2 inv2: 4
Xdff_r0_c0 din_0 dout_0 dout_bar_0 clk vdd gnd dff_buf_0
.ENDS dff_buf_array_0

* ptx M{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

* ptx M{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT pinv_21 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
XMpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
XMpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS pinv_21

.SUBCKT pdriver_6 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 3, 8, 24, 72]
Xbuf_inv1 A Zb1_int vdd gnd pinv_6
Xbuf_inv2 Zb1_int Zb2_int vdd gnd pinv_7
Xbuf_inv3 Zb2_int Zb3_int vdd gnd pinv_8
Xbuf_inv4 Zb3_int Zb4_int vdd gnd pinv_9
Xbuf_inv5 Zb4_int Zb5_int vdd gnd pinv_10
Xbuf_inv6 Zb5_int Z vdd gnd pinv_21
.ENDS pdriver_6

.SUBCKT control_logic_r csb clk rbl_bl s_en p_en_bar wl_en clk_buf vdd gnd
* INPUT : csb 
* INPUT : clk 
* INPUT : rbl_bl 
* OUTPUT: s_en 
* OUTPUT: p_en_bar 
* OUTPUT: wl_en 
* OUTPUT: clk_buf 
* POWER : vdd 
* GROUND: gnd 
* word_size 32
Xctrl_dffs csb cs_bar cs clk_buf vdd gnd dff_buf_array_0
Xclkbuf clk clk_buf vdd gnd pdriver_6
Xinv_clk_bar clk_buf clk_bar vdd gnd pinv_0
Xand2_gated_clk_bar clk_bar cs gated_clk_bar vdd gnd pand2_0
Xand2_gated_clk_buf clk_buf cs gated_clk_buf vdd gnd pand2_0
Xbuf_wl_en gated_clk_bar wl_en vdd gnd pdriver_2
Xbuf_s_en_and rbl_bl_delay gated_clk_bar cs s_en vdd gnd pand3_0
Xdelay_chain rbl_bl rbl_bl_delay vdd gnd delay_chain
Xnand_p_en_bar gated_clk_buf rbl_bl_delay p_en_bar_unbuf vdd gnd pnand2_1
Xbuf_p_en_bar p_en_bar_unbuf p_en_bar vdd gnd pdriver_5
.ENDS control_logic_r

.SUBCKT sram_1rw1r_32_256_8_sky130  din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6] din0[7] din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15] din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22] din0[23] din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[30] din0[31] addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] addr1[0] addr1[1] addr1[2] addr1[3] addr1[4] addr1[5] addr1[6] addr1[7] csb0 csb1 web0 clk0 clk1 wmask0[0] wmask0[1] wmask0[2] wmask0[3] dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19] dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[30] dout0[31] dout1[0] dout1[1] dout1[2] dout1[3] dout1[4] dout1[5] dout1[6] dout1[7] dout1[8] dout1[9] dout1[10] dout1[11] dout1[12] dout1[13] dout1[14] dout1[15] dout1[16] dout1[17] dout1[18] dout1[19] dout1[20] dout1[21] dout1[22] dout1[23] dout1[24] dout1[25] dout1[26] dout1[27] dout1[28] dout1[29] dout1[30] dout1[31] vdd gnd
* INPUT : din0[0] 
* INPUT : din0[1] 
* INPUT : din0[2] 
* INPUT : din0[3] 
* INPUT : din0[4] 
* INPUT : din0[5] 
* INPUT : din0[6] 
* INPUT : din0[7] 
* INPUT : din0[8] 
* INPUT : din0[9] 
* INPUT : din0[10] 
* INPUT : din0[11] 
* INPUT : din0[12] 
* INPUT : din0[13] 
* INPUT : din0[14] 
* INPUT : din0[15] 
* INPUT : din0[16] 
* INPUT : din0[17] 
* INPUT : din0[18] 
* INPUT : din0[19] 
* INPUT : din0[20] 
* INPUT : din0[21] 
* INPUT : din0[22] 
* INPUT : din0[23] 
* INPUT : din0[24] 
* INPUT : din0[25] 
* INPUT : din0[26] 
* INPUT : din0[27] 
* INPUT : din0[28] 
* INPUT : din0[29] 
* INPUT : din0[30] 
* INPUT : din0[31] 
* INPUT : addr0[0] 
* INPUT : addr0[1] 
* INPUT : addr0[2] 
* INPUT : addr0[3] 
* INPUT : addr0[4] 
* INPUT : addr0[5] 
* INPUT : addr0[6] 
* INPUT : addr0[7] 
* INPUT : addr1[0] 
* INPUT : addr1[1] 
* INPUT : addr1[2] 
* INPUT : addr1[3] 
* INPUT : addr1[4] 
* INPUT : addr1[5] 
* INPUT : addr1[6] 
* INPUT : addr1[7] 
* INPUT : csb0 
* INPUT : csb1 
* INPUT : web0 
* INPUT : clk0 
* INPUT : clk1 
* INPUT : wmask0[0] 
* INPUT : wmask0[1] 
* INPUT : wmask0[2] 
* INPUT : wmask0[3] 
* OUTPUT: dout0[0] 
* OUTPUT: dout0[1] 
* OUTPUT: dout0[2] 
* OUTPUT: dout0[3] 
* OUTPUT: dout0[4] 
* OUTPUT: dout0[5] 
* OUTPUT: dout0[6] 
* OUTPUT: dout0[7] 
* OUTPUT: dout0[8] 
* OUTPUT: dout0[9] 
* OUTPUT: dout0[10] 
* OUTPUT: dout0[11] 
* OUTPUT: dout0[12] 
* OUTPUT: dout0[13] 
* OUTPUT: dout0[14] 
* OUTPUT: dout0[15] 
* OUTPUT: dout0[16] 
* OUTPUT: dout0[17] 
* OUTPUT: dout0[18] 
* OUTPUT: dout0[19] 
* OUTPUT: dout0[20] 
* OUTPUT: dout0[21] 
* OUTPUT: dout0[22] 
* OUTPUT: dout0[23] 
* OUTPUT: dout0[24] 
* OUTPUT: dout0[25] 
* OUTPUT: dout0[26] 
* OUTPUT: dout0[27] 
* OUTPUT: dout0[28] 
* OUTPUT: dout0[29] 
* OUTPUT: dout0[30] 
* OUTPUT: dout0[31] 
* OUTPUT: dout1[0] 
* OUTPUT: dout1[1] 
* OUTPUT: dout1[2] 
* OUTPUT: dout1[3] 
* OUTPUT: dout1[4] 
* OUTPUT: dout1[5] 
* OUTPUT: dout1[6] 
* OUTPUT: dout1[7] 
* OUTPUT: dout1[8] 
* OUTPUT: dout1[9] 
* OUTPUT: dout1[10] 
* OUTPUT: dout1[11] 
* OUTPUT: dout1[12] 
* OUTPUT: dout1[13] 
* OUTPUT: dout1[14] 
* OUTPUT: dout1[15] 
* OUTPUT: dout1[16] 
* OUTPUT: dout1[17] 
* OUTPUT: dout1[18] 
* OUTPUT: dout1[19] 
* OUTPUT: dout1[20] 
* OUTPUT: dout1[21] 
* OUTPUT: dout1[22] 
* OUTPUT: dout1[23] 
* OUTPUT: dout1[24] 
* OUTPUT: dout1[25] 
* OUTPUT: dout1[26] 
* OUTPUT: dout1[27] 
* OUTPUT: dout1[28] 
* OUTPUT: dout1[29] 
* OUTPUT: dout1[30] 
* OUTPUT: dout1[31] 
* POWER : vdd 
* GROUND: gnd 
Xbank0 dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19] dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[30] dout0[31] dout1[0] dout1[1] dout1[2] dout1[3] dout1[4] dout1[5] dout1[6] dout1[7] dout1[8] dout1[9] dout1[10] dout1[11] dout1[12] dout1[13] dout1[14] dout1[15] dout1[16] dout1[17] dout1[18] dout1[19] dout1[20] dout1[21] dout1[22] dout1[23] dout1[24] dout1[25] dout1[26] dout1[27] dout1[28] dout1[29] dout1[30] dout1[31] rbl_bl0 rbl_bl1 bank_din0[0] bank_din0[1] bank_din0[2] bank_din0[3] bank_din0[4] bank_din0[5] bank_din0[6] bank_din0[7] bank_din0[8] bank_din0[9] bank_din0[10] bank_din0[11] bank_din0[12] bank_din0[13] bank_din0[14] bank_din0[15] bank_din0[16] bank_din0[17] bank_din0[18] bank_din0[19] bank_din0[20] bank_din0[21] bank_din0[22] bank_din0[23] bank_din0[24] bank_din0[25] bank_din0[26] bank_din0[27] bank_din0[28] bank_din0[29] bank_din0[30] bank_din0[31] a0[0] a0[1] a0[2] a0[3] a0[4] a0[5] a0[6] a0[7] a1[0] a1[1] a1[2] a1[3] a1[4] a1[5] a1[6] a1[7] s_en0 s_en1 p_en_bar0 p_en_bar1 w_en0 bank_wmask0[0] bank_wmask0[1] bank_wmask0[2] bank_wmask0[3] wl_en0 wl_en1 vdd gnd bank
Xcontrol0 csb0 web0 clk0 rbl_bl0 s_en0 w_en0 p_en_bar0 wl_en0 clk_buf0 vdd gnd control_logic_rw
Xcontrol1 csb1 clk1 rbl_bl1 s_en1 p_en_bar1 wl_en1 clk_buf1 vdd gnd control_logic_r
Xrow_address0 addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] a0[1] a0[2] a0[3] a0[4] a0[5] a0[6] a0[7] clk_buf0 vdd gnd row_addr_dff
Xrow_address1 addr1[1] addr1[2] addr1[3] addr1[4] addr1[5] addr1[6] addr1[7] a1[1] a1[2] a1[3] a1[4] a1[5] a1[6] a1[7] clk_buf1 vdd gnd row_addr_dff
Xcol_address0 addr0[0] a0[0] clk_buf0 vdd gnd col_addr_dff
Xcol_address1 addr1[0] a1[0] clk_buf1 vdd gnd col_addr_dff
Xwmask_dff0 wmask0[0] wmask0[1] wmask0[2] wmask0[3] bank_wmask0[0] bank_wmask0[1] bank_wmask0[2] bank_wmask0[3] clk_buf0 vdd gnd wmask_dff
Xdata_dff0 din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6] din0[7] din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15] din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22] din0[23] din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[30] din0[31] bank_din0[0] bank_din0[1] bank_din0[2] bank_din0[3] bank_din0[4] bank_din0[5] bank_din0[6] bank_din0[7] bank_din0[8] bank_din0[9] bank_din0[10] bank_din0[11] bank_din0[12] bank_din0[13] bank_din0[14] bank_din0[15] bank_din0[16] bank_din0[17] bank_din0[18] bank_din0[19] bank_din0[20] bank_din0[21] bank_din0[22] bank_din0[23] bank_din0[24] bank_din0[25] bank_din0[26] bank_din0[27] bank_din0[28] bank_din0[29] bank_din0[30] bank_din0[31] clk_buf0 vdd gnd data_dff
.ENDS sram_1rw1r_32_256_8_sky130
