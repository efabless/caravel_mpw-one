* NGSPICE file created from (UNNAMED).ext - technology: sky130A

.subckt x(UNNAMED)
.ends

