magic
tech sky130A
magscale 1 2
timestamp 1608935505
<< obsli1 >>
rect 1104 2159 428812 179231
<< obsm1 >>
rect 566 892 429166 179716
<< metal2 >>
rect 754 179200 810 180000
rect 1122 179200 1178 180000
rect 1490 179200 1546 180000
rect 1858 179200 1914 180000
rect 2226 179200 2282 180000
rect 2594 179200 2650 180000
rect 2962 179200 3018 180000
rect 3330 179200 3386 180000
rect 3698 179200 3754 180000
rect 4066 179200 4122 180000
rect 4434 179200 4490 180000
rect 4802 179200 4858 180000
rect 5170 179200 5226 180000
rect 5538 179200 5594 180000
rect 5906 179200 5962 180000
rect 6274 179200 6330 180000
rect 6642 179200 6698 180000
rect 7010 179200 7066 180000
rect 7378 179200 7434 180000
rect 7746 179200 7802 180000
rect 8114 179200 8170 180000
rect 8482 179200 8538 180000
rect 8850 179200 8906 180000
rect 9218 179200 9274 180000
rect 9586 179200 9642 180000
rect 9954 179200 10010 180000
rect 10322 179200 10378 180000
rect 10690 179200 10746 180000
rect 11058 179200 11114 180000
rect 11426 179200 11482 180000
rect 11794 179200 11850 180000
rect 12162 179200 12218 180000
rect 12530 179200 12586 180000
rect 12898 179200 12954 180000
rect 13266 179200 13322 180000
rect 13634 179200 13690 180000
rect 14002 179200 14058 180000
rect 14370 179200 14426 180000
rect 14738 179200 14794 180000
rect 15106 179200 15162 180000
rect 15474 179200 15530 180000
rect 15842 179200 15898 180000
rect 16210 179200 16266 180000
rect 16578 179200 16634 180000
rect 16946 179200 17002 180000
rect 17314 179200 17370 180000
rect 17682 179200 17738 180000
rect 18050 179200 18106 180000
rect 18418 179200 18474 180000
rect 18786 179200 18842 180000
rect 19154 179200 19210 180000
rect 19522 179200 19578 180000
rect 19890 179200 19946 180000
rect 20258 179200 20314 180000
rect 20626 179200 20682 180000
rect 20994 179200 21050 180000
rect 21362 179200 21418 180000
rect 21730 179200 21786 180000
rect 22098 179200 22154 180000
rect 22466 179200 22522 180000
rect 22834 179200 22890 180000
rect 23202 179200 23258 180000
rect 23570 179200 23626 180000
rect 23938 179200 23994 180000
rect 24306 179200 24362 180000
rect 24674 179200 24730 180000
rect 25042 179200 25098 180000
rect 25410 179200 25466 180000
rect 25778 179200 25834 180000
rect 26146 179200 26202 180000
rect 26514 179200 26570 180000
rect 26882 179200 26938 180000
rect 27250 179200 27306 180000
rect 27618 179200 27674 180000
rect 27986 179200 28042 180000
rect 28354 179200 28410 180000
rect 28722 179200 28778 180000
rect 29090 179200 29146 180000
rect 29458 179200 29514 180000
rect 29826 179200 29882 180000
rect 30194 179200 30250 180000
rect 30562 179200 30618 180000
rect 30930 179200 30986 180000
rect 31298 179200 31354 180000
rect 31666 179200 31722 180000
rect 32034 179200 32090 180000
rect 32402 179200 32458 180000
rect 32770 179200 32826 180000
rect 33138 179200 33194 180000
rect 33506 179200 33562 180000
rect 33874 179200 33930 180000
rect 34242 179200 34298 180000
rect 34610 179200 34666 180000
rect 34978 179200 35034 180000
rect 35346 179200 35402 180000
rect 35714 179200 35770 180000
rect 36082 179200 36138 180000
rect 36450 179200 36506 180000
rect 36818 179200 36874 180000
rect 37186 179200 37242 180000
rect 37554 179200 37610 180000
rect 37922 179200 37978 180000
rect 38290 179200 38346 180000
rect 38658 179200 38714 180000
rect 39026 179200 39082 180000
rect 39394 179200 39450 180000
rect 39762 179200 39818 180000
rect 40130 179200 40186 180000
rect 40498 179200 40554 180000
rect 40866 179200 40922 180000
rect 41234 179200 41290 180000
rect 41602 179200 41658 180000
rect 41970 179200 42026 180000
rect 42338 179200 42394 180000
rect 42706 179200 42762 180000
rect 43074 179200 43130 180000
rect 43442 179200 43498 180000
rect 43810 179200 43866 180000
rect 44178 179200 44234 180000
rect 44546 179200 44602 180000
rect 44914 179200 44970 180000
rect 45282 179200 45338 180000
rect 45650 179200 45706 180000
rect 46018 179200 46074 180000
rect 46386 179200 46442 180000
rect 46754 179200 46810 180000
rect 47122 179200 47178 180000
rect 47490 179200 47546 180000
rect 47858 179200 47914 180000
rect 48226 179200 48282 180000
rect 48594 179200 48650 180000
rect 48962 179200 49018 180000
rect 49330 179200 49386 180000
rect 49698 179200 49754 180000
rect 50066 179200 50122 180000
rect 50434 179200 50490 180000
rect 50802 179200 50858 180000
rect 51170 179200 51226 180000
rect 51538 179200 51594 180000
rect 51906 179200 51962 180000
rect 52274 179200 52330 180000
rect 52642 179200 52698 180000
rect 53010 179200 53066 180000
rect 53378 179200 53434 180000
rect 53746 179200 53802 180000
rect 54114 179200 54170 180000
rect 54482 179200 54538 180000
rect 54850 179200 54906 180000
rect 55218 179200 55274 180000
rect 55586 179200 55642 180000
rect 55954 179200 56010 180000
rect 56322 179200 56378 180000
rect 56690 179200 56746 180000
rect 57058 179200 57114 180000
rect 57426 179200 57482 180000
rect 57794 179200 57850 180000
rect 58162 179200 58218 180000
rect 58530 179200 58586 180000
rect 58898 179200 58954 180000
rect 59266 179200 59322 180000
rect 59634 179200 59690 180000
rect 60002 179200 60058 180000
rect 60370 179200 60426 180000
rect 60738 179200 60794 180000
rect 61106 179200 61162 180000
rect 61474 179200 61530 180000
rect 61842 179200 61898 180000
rect 62210 179200 62266 180000
rect 62578 179200 62634 180000
rect 62946 179200 63002 180000
rect 63314 179200 63370 180000
rect 63682 179200 63738 180000
rect 64050 179200 64106 180000
rect 64418 179200 64474 180000
rect 64786 179200 64842 180000
rect 65154 179200 65210 180000
rect 65522 179200 65578 180000
rect 65890 179200 65946 180000
rect 66258 179200 66314 180000
rect 66626 179200 66682 180000
rect 66994 179200 67050 180000
rect 67362 179200 67418 180000
rect 67730 179200 67786 180000
rect 68098 179200 68154 180000
rect 68466 179200 68522 180000
rect 68834 179200 68890 180000
rect 69202 179200 69258 180000
rect 69570 179200 69626 180000
rect 69938 179200 69994 180000
rect 70306 179200 70362 180000
rect 70674 179200 70730 180000
rect 71042 179200 71098 180000
rect 71410 179200 71466 180000
rect 71778 179200 71834 180000
rect 72146 179200 72202 180000
rect 72514 179200 72570 180000
rect 72882 179200 72938 180000
rect 73250 179200 73306 180000
rect 73618 179200 73674 180000
rect 73986 179200 74042 180000
rect 74354 179200 74410 180000
rect 74722 179200 74778 180000
rect 75090 179200 75146 180000
rect 75458 179200 75514 180000
rect 75826 179200 75882 180000
rect 76194 179200 76250 180000
rect 76562 179200 76618 180000
rect 76930 179200 76986 180000
rect 77298 179200 77354 180000
rect 77666 179200 77722 180000
rect 78034 179200 78090 180000
rect 78402 179200 78458 180000
rect 78770 179200 78826 180000
rect 79138 179200 79194 180000
rect 79506 179200 79562 180000
rect 79874 179200 79930 180000
rect 80242 179200 80298 180000
rect 80610 179200 80666 180000
rect 80978 179200 81034 180000
rect 81346 179200 81402 180000
rect 81714 179200 81770 180000
rect 82082 179200 82138 180000
rect 82450 179200 82506 180000
rect 82818 179200 82874 180000
rect 83186 179200 83242 180000
rect 83554 179200 83610 180000
rect 83922 179200 83978 180000
rect 84290 179200 84346 180000
rect 84658 179200 84714 180000
rect 85026 179200 85082 180000
rect 85394 179200 85450 180000
rect 85762 179200 85818 180000
rect 86130 179200 86186 180000
rect 86498 179200 86554 180000
rect 86866 179200 86922 180000
rect 87234 179200 87290 180000
rect 87602 179200 87658 180000
rect 87970 179200 88026 180000
rect 88338 179200 88394 180000
rect 88706 179200 88762 180000
rect 89074 179200 89130 180000
rect 89442 179200 89498 180000
rect 89810 179200 89866 180000
rect 90178 179200 90234 180000
rect 90546 179200 90602 180000
rect 90914 179200 90970 180000
rect 91282 179200 91338 180000
rect 91650 179200 91706 180000
rect 92018 179200 92074 180000
rect 92386 179200 92442 180000
rect 92754 179200 92810 180000
rect 93122 179200 93178 180000
rect 93490 179200 93546 180000
rect 93858 179200 93914 180000
rect 94226 179200 94282 180000
rect 94594 179200 94650 180000
rect 94962 179200 95018 180000
rect 95330 179200 95386 180000
rect 95698 179200 95754 180000
rect 96066 179200 96122 180000
rect 96434 179200 96490 180000
rect 96802 179200 96858 180000
rect 97170 179200 97226 180000
rect 97538 179200 97594 180000
rect 97906 179200 97962 180000
rect 98274 179200 98330 180000
rect 98642 179200 98698 180000
rect 99010 179200 99066 180000
rect 99378 179200 99434 180000
rect 99746 179200 99802 180000
rect 100114 179200 100170 180000
rect 100482 179200 100538 180000
rect 100850 179200 100906 180000
rect 101218 179200 101274 180000
rect 101586 179200 101642 180000
rect 101954 179200 102010 180000
rect 102322 179200 102378 180000
rect 102690 179200 102746 180000
rect 103058 179200 103114 180000
rect 103426 179200 103482 180000
rect 103794 179200 103850 180000
rect 104162 179200 104218 180000
rect 104530 179200 104586 180000
rect 104898 179200 104954 180000
rect 105266 179200 105322 180000
rect 105634 179200 105690 180000
rect 106002 179200 106058 180000
rect 106370 179200 106426 180000
rect 106738 179200 106794 180000
rect 107106 179200 107162 180000
rect 107474 179200 107530 180000
rect 107842 179200 107898 180000
rect 108210 179200 108266 180000
rect 108578 179200 108634 180000
rect 108946 179200 109002 180000
rect 109314 179200 109370 180000
rect 109682 179200 109738 180000
rect 110050 179200 110106 180000
rect 110418 179200 110474 180000
rect 110786 179200 110842 180000
rect 111154 179200 111210 180000
rect 111522 179200 111578 180000
rect 111890 179200 111946 180000
rect 112258 179200 112314 180000
rect 112626 179200 112682 180000
rect 112994 179200 113050 180000
rect 113362 179200 113418 180000
rect 113730 179200 113786 180000
rect 114098 179200 114154 180000
rect 114466 179200 114522 180000
rect 114834 179200 114890 180000
rect 115202 179200 115258 180000
rect 115570 179200 115626 180000
rect 115938 179200 115994 180000
rect 116306 179200 116362 180000
rect 116674 179200 116730 180000
rect 117042 179200 117098 180000
rect 117410 179200 117466 180000
rect 117778 179200 117834 180000
rect 118146 179200 118202 180000
rect 118514 179200 118570 180000
rect 118882 179200 118938 180000
rect 119250 179200 119306 180000
rect 119618 179200 119674 180000
rect 119986 179200 120042 180000
rect 120354 179200 120410 180000
rect 120722 179200 120778 180000
rect 121090 179200 121146 180000
rect 121458 179200 121514 180000
rect 121826 179200 121882 180000
rect 122194 179200 122250 180000
rect 122562 179200 122618 180000
rect 122930 179200 122986 180000
rect 123298 179200 123354 180000
rect 123666 179200 123722 180000
rect 124034 179200 124090 180000
rect 124402 179200 124458 180000
rect 124770 179200 124826 180000
rect 125138 179200 125194 180000
rect 125506 179200 125562 180000
rect 125874 179200 125930 180000
rect 126242 179200 126298 180000
rect 126610 179200 126666 180000
rect 126978 179200 127034 180000
rect 127346 179200 127402 180000
rect 127714 179200 127770 180000
rect 128082 179200 128138 180000
rect 128450 179200 128506 180000
rect 128818 179200 128874 180000
rect 129186 179200 129242 180000
rect 129554 179200 129610 180000
rect 129922 179200 129978 180000
rect 130290 179200 130346 180000
rect 130658 179200 130714 180000
rect 131026 179200 131082 180000
rect 131394 179200 131450 180000
rect 131762 179200 131818 180000
rect 132130 179200 132186 180000
rect 132498 179200 132554 180000
rect 132866 179200 132922 180000
rect 133234 179200 133290 180000
rect 133602 179200 133658 180000
rect 133970 179200 134026 180000
rect 134338 179200 134394 180000
rect 134706 179200 134762 180000
rect 135074 179200 135130 180000
rect 135442 179200 135498 180000
rect 135810 179200 135866 180000
rect 136178 179200 136234 180000
rect 136546 179200 136602 180000
rect 136914 179200 136970 180000
rect 137282 179200 137338 180000
rect 137650 179200 137706 180000
rect 138018 179200 138074 180000
rect 138386 179200 138442 180000
rect 138754 179200 138810 180000
rect 139122 179200 139178 180000
rect 139490 179200 139546 180000
rect 139858 179200 139914 180000
rect 140226 179200 140282 180000
rect 140594 179200 140650 180000
rect 140962 179200 141018 180000
rect 141330 179200 141386 180000
rect 141698 179200 141754 180000
rect 142066 179200 142122 180000
rect 142434 179200 142490 180000
rect 142802 179200 142858 180000
rect 143170 179200 143226 180000
rect 143538 179200 143594 180000
rect 143906 179200 143962 180000
rect 144274 179200 144330 180000
rect 144642 179200 144698 180000
rect 145010 179200 145066 180000
rect 145378 179200 145434 180000
rect 145746 179200 145802 180000
rect 146114 179200 146170 180000
rect 146482 179200 146538 180000
rect 146850 179200 146906 180000
rect 147218 179200 147274 180000
rect 147586 179200 147642 180000
rect 147954 179200 148010 180000
rect 148322 179200 148378 180000
rect 148690 179200 148746 180000
rect 149058 179200 149114 180000
rect 149426 179200 149482 180000
rect 149794 179200 149850 180000
rect 150162 179200 150218 180000
rect 150530 179200 150586 180000
rect 150898 179200 150954 180000
rect 151266 179200 151322 180000
rect 151634 179200 151690 180000
rect 152002 179200 152058 180000
rect 152370 179200 152426 180000
rect 152738 179200 152794 180000
rect 153106 179200 153162 180000
rect 153474 179200 153530 180000
rect 153842 179200 153898 180000
rect 154210 179200 154266 180000
rect 154578 179200 154634 180000
rect 154946 179200 155002 180000
rect 155314 179200 155370 180000
rect 155682 179200 155738 180000
rect 156050 179200 156106 180000
rect 156418 179200 156474 180000
rect 156786 179200 156842 180000
rect 157154 179200 157210 180000
rect 157522 179200 157578 180000
rect 157890 179200 157946 180000
rect 158258 179200 158314 180000
rect 158626 179200 158682 180000
rect 158994 179200 159050 180000
rect 159362 179200 159418 180000
rect 159730 179200 159786 180000
rect 160098 179200 160154 180000
rect 160466 179200 160522 180000
rect 160834 179200 160890 180000
rect 161202 179200 161258 180000
rect 161570 179200 161626 180000
rect 161938 179200 161994 180000
rect 162306 179200 162362 180000
rect 162674 179200 162730 180000
rect 163042 179200 163098 180000
rect 163410 179200 163466 180000
rect 163778 179200 163834 180000
rect 164146 179200 164202 180000
rect 164514 179200 164570 180000
rect 164882 179200 164938 180000
rect 165250 179200 165306 180000
rect 165618 179200 165674 180000
rect 165986 179200 166042 180000
rect 166354 179200 166410 180000
rect 166722 179200 166778 180000
rect 167090 179200 167146 180000
rect 167458 179200 167514 180000
rect 167826 179200 167882 180000
rect 168194 179200 168250 180000
rect 168562 179200 168618 180000
rect 168930 179200 168986 180000
rect 169298 179200 169354 180000
rect 169666 179200 169722 180000
rect 170034 179200 170090 180000
rect 170402 179200 170458 180000
rect 170770 179200 170826 180000
rect 171138 179200 171194 180000
rect 171506 179200 171562 180000
rect 171874 179200 171930 180000
rect 172242 179200 172298 180000
rect 172610 179200 172666 180000
rect 172978 179200 173034 180000
rect 173346 179200 173402 180000
rect 173714 179200 173770 180000
rect 174082 179200 174138 180000
rect 174450 179200 174506 180000
rect 174818 179200 174874 180000
rect 210146 179200 210202 180000
rect 287058 179200 287114 180000
rect 295154 179200 295210 180000
rect 299938 179200 299994 180000
rect 338578 179200 338634 180000
rect 426898 179200 426954 180000
rect 427266 179200 427322 180000
rect 427634 179200 427690 180000
rect 428002 179200 428058 180000
rect 428370 179200 428426 180000
rect 428738 179200 428794 180000
rect 429106 179200 429162 180000
rect 570 0 626 800
rect 754 0 810 800
rect 938 0 994 800
rect 1122 0 1178 800
rect 1306 0 1362 800
rect 1490 0 1546 800
rect 1674 0 1730 800
rect 1858 0 1914 800
rect 2042 0 2098 800
rect 2226 0 2282 800
rect 2410 0 2466 800
rect 2594 0 2650 800
rect 2778 0 2834 800
rect 2962 0 3018 800
rect 3146 0 3202 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3882 0 3938 800
rect 4066 0 4122 800
rect 4250 0 4306 800
rect 4434 0 4490 800
rect 4618 0 4674 800
rect 4802 0 4858 800
rect 4986 0 5042 800
rect 5170 0 5226 800
rect 5354 0 5410 800
rect 5538 0 5594 800
rect 5722 0 5778 800
rect 5906 0 5962 800
rect 6090 0 6146 800
rect 6274 0 6330 800
rect 6458 0 6514 800
rect 6642 0 6698 800
rect 6826 0 6882 800
rect 7010 0 7066 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7562 0 7618 800
rect 7746 0 7802 800
rect 7930 0 7986 800
rect 8114 0 8170 800
rect 8298 0 8354 800
rect 8482 0 8538 800
rect 8666 0 8722 800
rect 8850 0 8906 800
rect 9034 0 9090 800
rect 9218 0 9274 800
rect 9402 0 9458 800
rect 9586 0 9642 800
rect 9770 0 9826 800
rect 9954 0 10010 800
rect 10138 0 10194 800
rect 10322 0 10378 800
rect 10506 0 10562 800
rect 10690 0 10746 800
rect 10874 0 10930 800
rect 11058 0 11114 800
rect 11242 0 11298 800
rect 11426 0 11482 800
rect 11610 0 11666 800
rect 11794 0 11850 800
rect 11978 0 12034 800
rect 12162 0 12218 800
rect 12346 0 12402 800
rect 12530 0 12586 800
rect 12714 0 12770 800
rect 12898 0 12954 800
rect 13082 0 13138 800
rect 13266 0 13322 800
rect 13450 0 13506 800
rect 13634 0 13690 800
rect 13818 0 13874 800
rect 14002 0 14058 800
rect 14186 0 14242 800
rect 14370 0 14426 800
rect 14554 0 14610 800
rect 14738 0 14794 800
rect 14922 0 14978 800
rect 15106 0 15162 800
rect 15290 0 15346 800
rect 15474 0 15530 800
rect 15658 0 15714 800
rect 15842 0 15898 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20810 0 20866 800
rect 21178 0 21234 800
rect 21546 0 21602 800
rect 21914 0 21970 800
rect 22282 0 22338 800
rect 22650 0 22706 800
rect 23018 0 23074 800
rect 23386 0 23442 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24858 0 24914 800
rect 25226 0 25282 800
rect 25594 0 25650 800
rect 25962 0 26018 800
rect 26330 0 26386 800
rect 26698 0 26754 800
rect 27066 0 27122 800
rect 27434 0 27490 800
rect 27802 0 27858 800
rect 28170 0 28226 800
rect 28538 0 28594 800
rect 28906 0 28962 800
rect 29274 0 29330 800
rect 29642 0 29698 800
rect 30010 0 30066 800
rect 30378 0 30434 800
rect 30746 0 30802 800
rect 31114 0 31170 800
rect 31482 0 31538 800
rect 31850 0 31906 800
rect 32218 0 32274 800
rect 32586 0 32642 800
rect 32954 0 33010 800
rect 33322 0 33378 800
rect 33690 0 33746 800
<< obsm2 >>
rect 572 179144 698 179722
rect 866 179144 1066 179722
rect 1234 179144 1434 179722
rect 1602 179144 1802 179722
rect 1970 179144 2170 179722
rect 2338 179144 2538 179722
rect 2706 179144 2906 179722
rect 3074 179144 3274 179722
rect 3442 179144 3642 179722
rect 3810 179144 4010 179722
rect 4178 179144 4378 179722
rect 4546 179144 4746 179722
rect 4914 179144 5114 179722
rect 5282 179144 5482 179722
rect 5650 179144 5850 179722
rect 6018 179144 6218 179722
rect 6386 179144 6586 179722
rect 6754 179144 6954 179722
rect 7122 179144 7322 179722
rect 7490 179144 7690 179722
rect 7858 179144 8058 179722
rect 8226 179144 8426 179722
rect 8594 179144 8794 179722
rect 8962 179144 9162 179722
rect 9330 179144 9530 179722
rect 9698 179144 9898 179722
rect 10066 179144 10266 179722
rect 10434 179144 10634 179722
rect 10802 179144 11002 179722
rect 11170 179144 11370 179722
rect 11538 179144 11738 179722
rect 11906 179144 12106 179722
rect 12274 179144 12474 179722
rect 12642 179144 12842 179722
rect 13010 179144 13210 179722
rect 13378 179144 13578 179722
rect 13746 179144 13946 179722
rect 14114 179144 14314 179722
rect 14482 179144 14682 179722
rect 14850 179144 15050 179722
rect 15218 179144 15418 179722
rect 15586 179144 15786 179722
rect 15954 179144 16154 179722
rect 16322 179144 16522 179722
rect 16690 179144 16890 179722
rect 17058 179144 17258 179722
rect 17426 179144 17626 179722
rect 17794 179144 17994 179722
rect 18162 179144 18362 179722
rect 18530 179144 18730 179722
rect 18898 179144 19098 179722
rect 19266 179144 19466 179722
rect 19634 179144 19834 179722
rect 20002 179144 20202 179722
rect 20370 179144 20570 179722
rect 20738 179144 20938 179722
rect 21106 179144 21306 179722
rect 21474 179144 21674 179722
rect 21842 179144 22042 179722
rect 22210 179144 22410 179722
rect 22578 179144 22778 179722
rect 22946 179144 23146 179722
rect 23314 179144 23514 179722
rect 23682 179144 23882 179722
rect 24050 179144 24250 179722
rect 24418 179144 24618 179722
rect 24786 179144 24986 179722
rect 25154 179144 25354 179722
rect 25522 179144 25722 179722
rect 25890 179144 26090 179722
rect 26258 179144 26458 179722
rect 26626 179144 26826 179722
rect 26994 179144 27194 179722
rect 27362 179144 27562 179722
rect 27730 179144 27930 179722
rect 28098 179144 28298 179722
rect 28466 179144 28666 179722
rect 28834 179144 29034 179722
rect 29202 179144 29402 179722
rect 29570 179144 29770 179722
rect 29938 179144 30138 179722
rect 30306 179144 30506 179722
rect 30674 179144 30874 179722
rect 31042 179144 31242 179722
rect 31410 179144 31610 179722
rect 31778 179144 31978 179722
rect 32146 179144 32346 179722
rect 32514 179144 32714 179722
rect 32882 179144 33082 179722
rect 33250 179144 33450 179722
rect 33618 179144 33818 179722
rect 33986 179144 34186 179722
rect 34354 179144 34554 179722
rect 34722 179144 34922 179722
rect 35090 179144 35290 179722
rect 35458 179144 35658 179722
rect 35826 179144 36026 179722
rect 36194 179144 36394 179722
rect 36562 179144 36762 179722
rect 36930 179144 37130 179722
rect 37298 179144 37498 179722
rect 37666 179144 37866 179722
rect 38034 179144 38234 179722
rect 38402 179144 38602 179722
rect 38770 179144 38970 179722
rect 39138 179144 39338 179722
rect 39506 179144 39706 179722
rect 39874 179144 40074 179722
rect 40242 179144 40442 179722
rect 40610 179144 40810 179722
rect 40978 179144 41178 179722
rect 41346 179144 41546 179722
rect 41714 179144 41914 179722
rect 42082 179144 42282 179722
rect 42450 179144 42650 179722
rect 42818 179144 43018 179722
rect 43186 179144 43386 179722
rect 43554 179144 43754 179722
rect 43922 179144 44122 179722
rect 44290 179144 44490 179722
rect 44658 179144 44858 179722
rect 45026 179144 45226 179722
rect 45394 179144 45594 179722
rect 45762 179144 45962 179722
rect 46130 179144 46330 179722
rect 46498 179144 46698 179722
rect 46866 179144 47066 179722
rect 47234 179144 47434 179722
rect 47602 179144 47802 179722
rect 47970 179144 48170 179722
rect 48338 179144 48538 179722
rect 48706 179144 48906 179722
rect 49074 179144 49274 179722
rect 49442 179144 49642 179722
rect 49810 179144 50010 179722
rect 50178 179144 50378 179722
rect 50546 179144 50746 179722
rect 50914 179144 51114 179722
rect 51282 179144 51482 179722
rect 51650 179144 51850 179722
rect 52018 179144 52218 179722
rect 52386 179144 52586 179722
rect 52754 179144 52954 179722
rect 53122 179144 53322 179722
rect 53490 179144 53690 179722
rect 53858 179144 54058 179722
rect 54226 179144 54426 179722
rect 54594 179144 54794 179722
rect 54962 179144 55162 179722
rect 55330 179144 55530 179722
rect 55698 179144 55898 179722
rect 56066 179144 56266 179722
rect 56434 179144 56634 179722
rect 56802 179144 57002 179722
rect 57170 179144 57370 179722
rect 57538 179144 57738 179722
rect 57906 179144 58106 179722
rect 58274 179144 58474 179722
rect 58642 179144 58842 179722
rect 59010 179144 59210 179722
rect 59378 179144 59578 179722
rect 59746 179144 59946 179722
rect 60114 179144 60314 179722
rect 60482 179144 60682 179722
rect 60850 179144 61050 179722
rect 61218 179144 61418 179722
rect 61586 179144 61786 179722
rect 61954 179144 62154 179722
rect 62322 179144 62522 179722
rect 62690 179144 62890 179722
rect 63058 179144 63258 179722
rect 63426 179144 63626 179722
rect 63794 179144 63994 179722
rect 64162 179144 64362 179722
rect 64530 179144 64730 179722
rect 64898 179144 65098 179722
rect 65266 179144 65466 179722
rect 65634 179144 65834 179722
rect 66002 179144 66202 179722
rect 66370 179144 66570 179722
rect 66738 179144 66938 179722
rect 67106 179144 67306 179722
rect 67474 179144 67674 179722
rect 67842 179144 68042 179722
rect 68210 179144 68410 179722
rect 68578 179144 68778 179722
rect 68946 179144 69146 179722
rect 69314 179144 69514 179722
rect 69682 179144 69882 179722
rect 70050 179144 70250 179722
rect 70418 179144 70618 179722
rect 70786 179144 70986 179722
rect 71154 179144 71354 179722
rect 71522 179144 71722 179722
rect 71890 179144 72090 179722
rect 72258 179144 72458 179722
rect 72626 179144 72826 179722
rect 72994 179144 73194 179722
rect 73362 179144 73562 179722
rect 73730 179144 73930 179722
rect 74098 179144 74298 179722
rect 74466 179144 74666 179722
rect 74834 179144 75034 179722
rect 75202 179144 75402 179722
rect 75570 179144 75770 179722
rect 75938 179144 76138 179722
rect 76306 179144 76506 179722
rect 76674 179144 76874 179722
rect 77042 179144 77242 179722
rect 77410 179144 77610 179722
rect 77778 179144 77978 179722
rect 78146 179144 78346 179722
rect 78514 179144 78714 179722
rect 78882 179144 79082 179722
rect 79250 179144 79450 179722
rect 79618 179144 79818 179722
rect 79986 179144 80186 179722
rect 80354 179144 80554 179722
rect 80722 179144 80922 179722
rect 81090 179144 81290 179722
rect 81458 179144 81658 179722
rect 81826 179144 82026 179722
rect 82194 179144 82394 179722
rect 82562 179144 82762 179722
rect 82930 179144 83130 179722
rect 83298 179144 83498 179722
rect 83666 179144 83866 179722
rect 84034 179144 84234 179722
rect 84402 179144 84602 179722
rect 84770 179144 84970 179722
rect 85138 179144 85338 179722
rect 85506 179144 85706 179722
rect 85874 179144 86074 179722
rect 86242 179144 86442 179722
rect 86610 179144 86810 179722
rect 86978 179144 87178 179722
rect 87346 179144 87546 179722
rect 87714 179144 87914 179722
rect 88082 179144 88282 179722
rect 88450 179144 88650 179722
rect 88818 179144 89018 179722
rect 89186 179144 89386 179722
rect 89554 179144 89754 179722
rect 89922 179144 90122 179722
rect 90290 179144 90490 179722
rect 90658 179144 90858 179722
rect 91026 179144 91226 179722
rect 91394 179144 91594 179722
rect 91762 179144 91962 179722
rect 92130 179144 92330 179722
rect 92498 179144 92698 179722
rect 92866 179144 93066 179722
rect 93234 179144 93434 179722
rect 93602 179144 93802 179722
rect 93970 179144 94170 179722
rect 94338 179144 94538 179722
rect 94706 179144 94906 179722
rect 95074 179144 95274 179722
rect 95442 179144 95642 179722
rect 95810 179144 96010 179722
rect 96178 179144 96378 179722
rect 96546 179144 96746 179722
rect 96914 179144 97114 179722
rect 97282 179144 97482 179722
rect 97650 179144 97850 179722
rect 98018 179144 98218 179722
rect 98386 179144 98586 179722
rect 98754 179144 98954 179722
rect 99122 179144 99322 179722
rect 99490 179144 99690 179722
rect 99858 179144 100058 179722
rect 100226 179144 100426 179722
rect 100594 179144 100794 179722
rect 100962 179144 101162 179722
rect 101330 179144 101530 179722
rect 101698 179144 101898 179722
rect 102066 179144 102266 179722
rect 102434 179144 102634 179722
rect 102802 179144 103002 179722
rect 103170 179144 103370 179722
rect 103538 179144 103738 179722
rect 103906 179144 104106 179722
rect 104274 179144 104474 179722
rect 104642 179144 104842 179722
rect 105010 179144 105210 179722
rect 105378 179144 105578 179722
rect 105746 179144 105946 179722
rect 106114 179144 106314 179722
rect 106482 179144 106682 179722
rect 106850 179144 107050 179722
rect 107218 179144 107418 179722
rect 107586 179144 107786 179722
rect 107954 179144 108154 179722
rect 108322 179144 108522 179722
rect 108690 179144 108890 179722
rect 109058 179144 109258 179722
rect 109426 179144 109626 179722
rect 109794 179144 109994 179722
rect 110162 179144 110362 179722
rect 110530 179144 110730 179722
rect 110898 179144 111098 179722
rect 111266 179144 111466 179722
rect 111634 179144 111834 179722
rect 112002 179144 112202 179722
rect 112370 179144 112570 179722
rect 112738 179144 112938 179722
rect 113106 179144 113306 179722
rect 113474 179144 113674 179722
rect 113842 179144 114042 179722
rect 114210 179144 114410 179722
rect 114578 179144 114778 179722
rect 114946 179144 115146 179722
rect 115314 179144 115514 179722
rect 115682 179144 115882 179722
rect 116050 179144 116250 179722
rect 116418 179144 116618 179722
rect 116786 179144 116986 179722
rect 117154 179144 117354 179722
rect 117522 179144 117722 179722
rect 117890 179144 118090 179722
rect 118258 179144 118458 179722
rect 118626 179144 118826 179722
rect 118994 179144 119194 179722
rect 119362 179144 119562 179722
rect 119730 179144 119930 179722
rect 120098 179144 120298 179722
rect 120466 179144 120666 179722
rect 120834 179144 121034 179722
rect 121202 179144 121402 179722
rect 121570 179144 121770 179722
rect 121938 179144 122138 179722
rect 122306 179144 122506 179722
rect 122674 179144 122874 179722
rect 123042 179144 123242 179722
rect 123410 179144 123610 179722
rect 123778 179144 123978 179722
rect 124146 179144 124346 179722
rect 124514 179144 124714 179722
rect 124882 179144 125082 179722
rect 125250 179144 125450 179722
rect 125618 179144 125818 179722
rect 125986 179144 126186 179722
rect 126354 179144 126554 179722
rect 126722 179144 126922 179722
rect 127090 179144 127290 179722
rect 127458 179144 127658 179722
rect 127826 179144 128026 179722
rect 128194 179144 128394 179722
rect 128562 179144 128762 179722
rect 128930 179144 129130 179722
rect 129298 179144 129498 179722
rect 129666 179144 129866 179722
rect 130034 179144 130234 179722
rect 130402 179144 130602 179722
rect 130770 179144 130970 179722
rect 131138 179144 131338 179722
rect 131506 179144 131706 179722
rect 131874 179144 132074 179722
rect 132242 179144 132442 179722
rect 132610 179144 132810 179722
rect 132978 179144 133178 179722
rect 133346 179144 133546 179722
rect 133714 179144 133914 179722
rect 134082 179144 134282 179722
rect 134450 179144 134650 179722
rect 134818 179144 135018 179722
rect 135186 179144 135386 179722
rect 135554 179144 135754 179722
rect 135922 179144 136122 179722
rect 136290 179144 136490 179722
rect 136658 179144 136858 179722
rect 137026 179144 137226 179722
rect 137394 179144 137594 179722
rect 137762 179144 137962 179722
rect 138130 179144 138330 179722
rect 138498 179144 138698 179722
rect 138866 179144 139066 179722
rect 139234 179144 139434 179722
rect 139602 179144 139802 179722
rect 139970 179144 140170 179722
rect 140338 179144 140538 179722
rect 140706 179144 140906 179722
rect 141074 179144 141274 179722
rect 141442 179144 141642 179722
rect 141810 179144 142010 179722
rect 142178 179144 142378 179722
rect 142546 179144 142746 179722
rect 142914 179144 143114 179722
rect 143282 179144 143482 179722
rect 143650 179144 143850 179722
rect 144018 179144 144218 179722
rect 144386 179144 144586 179722
rect 144754 179144 144954 179722
rect 145122 179144 145322 179722
rect 145490 179144 145690 179722
rect 145858 179144 146058 179722
rect 146226 179144 146426 179722
rect 146594 179144 146794 179722
rect 146962 179144 147162 179722
rect 147330 179144 147530 179722
rect 147698 179144 147898 179722
rect 148066 179144 148266 179722
rect 148434 179144 148634 179722
rect 148802 179144 149002 179722
rect 149170 179144 149370 179722
rect 149538 179144 149738 179722
rect 149906 179144 150106 179722
rect 150274 179144 150474 179722
rect 150642 179144 150842 179722
rect 151010 179144 151210 179722
rect 151378 179144 151578 179722
rect 151746 179144 151946 179722
rect 152114 179144 152314 179722
rect 152482 179144 152682 179722
rect 152850 179144 153050 179722
rect 153218 179144 153418 179722
rect 153586 179144 153786 179722
rect 153954 179144 154154 179722
rect 154322 179144 154522 179722
rect 154690 179144 154890 179722
rect 155058 179144 155258 179722
rect 155426 179144 155626 179722
rect 155794 179144 155994 179722
rect 156162 179144 156362 179722
rect 156530 179144 156730 179722
rect 156898 179144 157098 179722
rect 157266 179144 157466 179722
rect 157634 179144 157834 179722
rect 158002 179144 158202 179722
rect 158370 179144 158570 179722
rect 158738 179144 158938 179722
rect 159106 179144 159306 179722
rect 159474 179144 159674 179722
rect 159842 179144 160042 179722
rect 160210 179144 160410 179722
rect 160578 179144 160778 179722
rect 160946 179144 161146 179722
rect 161314 179144 161514 179722
rect 161682 179144 161882 179722
rect 162050 179144 162250 179722
rect 162418 179144 162618 179722
rect 162786 179144 162986 179722
rect 163154 179144 163354 179722
rect 163522 179144 163722 179722
rect 163890 179144 164090 179722
rect 164258 179144 164458 179722
rect 164626 179144 164826 179722
rect 164994 179144 165194 179722
rect 165362 179144 165562 179722
rect 165730 179144 165930 179722
rect 166098 179144 166298 179722
rect 166466 179144 166666 179722
rect 166834 179144 167034 179722
rect 167202 179144 167402 179722
rect 167570 179144 167770 179722
rect 167938 179144 168138 179722
rect 168306 179144 168506 179722
rect 168674 179144 168874 179722
rect 169042 179144 169242 179722
rect 169410 179144 169610 179722
rect 169778 179144 169978 179722
rect 170146 179144 170346 179722
rect 170514 179144 170714 179722
rect 170882 179144 171082 179722
rect 171250 179144 171450 179722
rect 171618 179144 171818 179722
rect 171986 179144 172186 179722
rect 172354 179144 172554 179722
rect 172722 179144 172922 179722
rect 173090 179144 173290 179722
rect 173458 179144 173658 179722
rect 173826 179144 174026 179722
rect 174194 179144 174394 179722
rect 174562 179144 174762 179722
rect 174930 179144 210090 179722
rect 210258 179144 287002 179722
rect 287170 179144 295098 179722
rect 295266 179144 299882 179722
rect 300050 179144 338522 179722
rect 338690 179144 426842 179722
rect 427010 179144 427210 179722
rect 427378 179144 427578 179722
rect 427746 179144 427946 179722
rect 428114 179144 428314 179722
rect 428482 179144 428682 179722
rect 428850 179144 429050 179722
rect 572 856 429160 179144
rect 682 800 698 856
rect 866 800 882 856
rect 1050 800 1066 856
rect 1234 800 1250 856
rect 1418 800 1434 856
rect 1602 800 1618 856
rect 1786 800 1802 856
rect 1970 800 1986 856
rect 2154 800 2170 856
rect 2338 800 2354 856
rect 2522 800 2538 856
rect 2706 800 2722 856
rect 2890 800 2906 856
rect 3074 800 3090 856
rect 3258 800 3274 856
rect 3442 800 3458 856
rect 3626 800 3642 856
rect 3810 800 3826 856
rect 3994 800 4010 856
rect 4178 800 4194 856
rect 4362 800 4378 856
rect 4546 800 4562 856
rect 4730 800 4746 856
rect 4914 800 4930 856
rect 5098 800 5114 856
rect 5282 800 5298 856
rect 5466 800 5482 856
rect 5650 800 5666 856
rect 5834 800 5850 856
rect 6018 800 6034 856
rect 6202 800 6218 856
rect 6386 800 6402 856
rect 6570 800 6586 856
rect 6754 800 6770 856
rect 6938 800 6954 856
rect 7122 800 7138 856
rect 7306 800 7322 856
rect 7490 800 7506 856
rect 7674 800 7690 856
rect 7858 800 7874 856
rect 8042 800 8058 856
rect 8226 800 8242 856
rect 8410 800 8426 856
rect 8594 800 8610 856
rect 8778 800 8794 856
rect 8962 800 8978 856
rect 9146 800 9162 856
rect 9330 800 9346 856
rect 9514 800 9530 856
rect 9698 800 9714 856
rect 9882 800 9898 856
rect 10066 800 10082 856
rect 10250 800 10266 856
rect 10434 800 10450 856
rect 10618 800 10634 856
rect 10802 800 10818 856
rect 10986 800 11002 856
rect 11170 800 11186 856
rect 11354 800 11370 856
rect 11538 800 11554 856
rect 11722 800 11738 856
rect 11906 800 11922 856
rect 12090 800 12106 856
rect 12274 800 12290 856
rect 12458 800 12474 856
rect 12642 800 12658 856
rect 12826 800 12842 856
rect 13010 800 13026 856
rect 13194 800 13210 856
rect 13378 800 13394 856
rect 13562 800 13578 856
rect 13746 800 13762 856
rect 13930 800 13946 856
rect 14114 800 14130 856
rect 14298 800 14314 856
rect 14482 800 14498 856
rect 14666 800 14682 856
rect 14850 800 14866 856
rect 15034 800 15050 856
rect 15218 800 15234 856
rect 15402 800 15418 856
rect 15586 800 15602 856
rect 15770 800 15786 856
rect 15954 800 15970 856
rect 16138 800 16338 856
rect 16506 800 16706 856
rect 16874 800 17074 856
rect 17242 800 17442 856
rect 17610 800 17810 856
rect 17978 800 18178 856
rect 18346 800 18546 856
rect 18714 800 18914 856
rect 19082 800 19282 856
rect 19450 800 19650 856
rect 19818 800 20018 856
rect 20186 800 20386 856
rect 20554 800 20754 856
rect 20922 800 21122 856
rect 21290 800 21490 856
rect 21658 800 21858 856
rect 22026 800 22226 856
rect 22394 800 22594 856
rect 22762 800 22962 856
rect 23130 800 23330 856
rect 23498 800 23698 856
rect 23866 800 24066 856
rect 24234 800 24434 856
rect 24602 800 24802 856
rect 24970 800 25170 856
rect 25338 800 25538 856
rect 25706 800 25906 856
rect 26074 800 26274 856
rect 26442 800 26642 856
rect 26810 800 27010 856
rect 27178 800 27378 856
rect 27546 800 27746 856
rect 27914 800 28114 856
rect 28282 800 28482 856
rect 28650 800 28850 856
rect 29018 800 29218 856
rect 29386 800 29586 856
rect 29754 800 29954 856
rect 30122 800 30322 856
rect 30490 800 30690 856
rect 30858 800 31058 856
rect 31226 800 31426 856
rect 31594 800 31794 856
rect 31962 800 32162 856
rect 32330 800 32530 856
rect 32698 800 32898 856
rect 33066 800 33266 856
rect 33434 800 33634 856
rect 33802 800 429160 856
<< metal3 >>
rect 0 178984 800 179104
rect 429200 178984 430000 179104
rect 0 178440 800 178560
rect 429200 178440 430000 178560
rect 0 177896 800 178016
rect 429200 177896 430000 178016
rect 0 177352 800 177472
rect 429200 177352 430000 177472
rect 0 176808 800 176928
rect 429200 176808 430000 176928
rect 0 176264 800 176384
rect 0 175720 800 175840
rect 0 175176 800 175296
rect 0 174632 800 174752
rect 0 174088 800 174208
rect 0 173544 800 173664
rect 0 173000 800 173120
rect 0 172456 800 172576
rect 0 171912 800 172032
rect 0 171368 800 171488
rect 0 170824 800 170944
rect 0 170280 800 170400
rect 0 169736 800 169856
rect 0 169192 800 169312
rect 0 168648 800 168768
rect 0 168104 800 168224
rect 0 167560 800 167680
rect 0 167016 800 167136
rect 0 166472 800 166592
rect 0 165928 800 166048
rect 0 165384 800 165504
rect 0 164840 800 164960
rect 0 164296 800 164416
rect 0 163752 800 163872
rect 0 163208 800 163328
rect 0 162664 800 162784
rect 0 162120 800 162240
rect 0 161576 800 161696
rect 0 161032 800 161152
rect 0 160488 800 160608
rect 0 159944 800 160064
rect 0 159400 800 159520
rect 0 158856 800 158976
rect 0 158312 800 158432
rect 0 157768 800 157888
rect 429200 157224 430000 157344
rect 0 149064 800 149184
rect 429200 113160 430000 113280
rect 429200 112616 430000 112736
rect 429200 112072 430000 112192
rect 429200 68008 430000 68128
rect 429200 67464 430000 67584
rect 429200 66920 430000 67040
rect 429200 66376 430000 66496
rect 429200 50600 430000 50720
rect 0 48424 800 48544
rect 0 47880 800 48000
rect 0 47336 800 47456
rect 0 46792 800 46912
rect 0 46248 800 46368
rect 0 45704 800 45824
rect 0 45160 800 45280
rect 0 44616 800 44736
rect 0 44072 800 44192
rect 0 43528 800 43648
rect 0 42984 800 43104
rect 0 42440 800 42560
rect 0 41896 800 42016
rect 0 41352 800 41472
rect 0 40808 800 40928
rect 0 40264 800 40384
rect 0 39720 800 39840
rect 0 39176 800 39296
rect 0 38632 800 38752
rect 0 38088 800 38208
rect 0 37544 800 37664
rect 0 37000 800 37120
rect 0 36456 800 36576
rect 0 35912 800 36032
rect 0 35368 800 35488
rect 429200 35368 430000 35488
rect 0 34824 800 34944
rect 429200 34824 430000 34944
rect 0 34280 800 34400
rect 429200 34280 430000 34400
rect 0 33736 800 33856
rect 429200 33736 430000 33856
rect 0 33192 800 33312
rect 429200 33192 430000 33312
rect 0 32648 800 32768
rect 429200 32648 430000 32768
rect 0 32104 800 32224
rect 429200 32104 430000 32224
rect 0 31560 800 31680
rect 429200 31560 430000 31680
rect 0 31016 800 31136
rect 429200 31016 430000 31136
rect 0 30472 800 30592
rect 429200 30472 430000 30592
rect 0 29928 800 30048
rect 429200 29928 430000 30048
rect 0 29384 800 29504
rect 429200 29384 430000 29504
rect 0 28840 800 28960
rect 429200 28840 430000 28960
rect 0 28296 800 28416
rect 429200 28296 430000 28416
rect 0 27752 800 27872
rect 429200 27752 430000 27872
rect 0 27208 800 27328
rect 429200 27208 430000 27328
rect 0 26664 800 26784
rect 429200 26664 430000 26784
rect 0 26120 800 26240
rect 429200 26120 430000 26240
rect 0 25576 800 25696
rect 429200 25576 430000 25696
rect 0 25032 800 25152
rect 429200 25032 430000 25152
rect 0 24488 800 24608
rect 429200 24488 430000 24608
rect 0 23944 800 24064
rect 429200 23944 430000 24064
rect 0 23400 800 23520
rect 429200 23400 430000 23520
rect 0 22856 800 22976
rect 429200 22856 430000 22976
rect 0 22312 800 22432
rect 429200 22312 430000 22432
rect 0 21768 800 21888
rect 429200 21768 430000 21888
rect 0 21224 800 21344
rect 429200 21224 430000 21344
rect 0 20680 800 20800
rect 429200 20680 430000 20800
rect 0 20136 800 20256
rect 429200 20136 430000 20256
rect 0 19592 800 19712
rect 429200 19592 430000 19712
rect 0 19048 800 19168
rect 429200 19048 430000 19168
rect 0 18504 800 18624
rect 429200 18504 430000 18624
rect 0 17960 800 18080
rect 0 17416 800 17536
rect 0 16872 800 16992
rect 0 16328 800 16448
rect 0 15784 800 15904
rect 0 15240 800 15360
rect 0 14696 800 14816
rect 0 14152 800 14272
rect 0 13608 800 13728
rect 0 13064 800 13184
rect 0 12520 800 12640
rect 0 11976 800 12096
rect 0 11432 800 11552
rect 0 10888 800 11008
rect 0 10344 800 10464
rect 0 9800 800 9920
rect 0 9256 800 9376
rect 0 8712 800 8832
rect 0 8168 800 8288
rect 0 7624 800 7744
rect 0 7080 800 7200
rect 0 6536 800 6656
rect 0 5992 800 6112
rect 0 5448 800 5568
rect 0 4904 800 5024
rect 0 4360 800 4480
rect 0 3816 800 3936
rect 0 3272 800 3392
rect 0 2728 800 2848
rect 0 2184 800 2304
rect 0 1640 800 1760
rect 0 1096 800 1216
<< obsm3 >>
rect 880 178904 429120 179077
rect 798 178640 429210 178904
rect 880 178360 429120 178640
rect 798 178096 429210 178360
rect 880 177816 429120 178096
rect 798 177552 429210 177816
rect 880 177272 429120 177552
rect 798 177008 429210 177272
rect 880 176728 429120 177008
rect 798 176464 429210 176728
rect 880 176184 429210 176464
rect 798 175920 429210 176184
rect 880 175640 429210 175920
rect 798 175376 429210 175640
rect 880 175096 429210 175376
rect 798 174832 429210 175096
rect 880 174552 429210 174832
rect 798 174288 429210 174552
rect 880 174008 429210 174288
rect 798 173744 429210 174008
rect 880 173464 429210 173744
rect 798 173200 429210 173464
rect 880 172920 429210 173200
rect 798 172656 429210 172920
rect 880 172376 429210 172656
rect 798 172112 429210 172376
rect 880 171832 429210 172112
rect 798 171568 429210 171832
rect 880 171288 429210 171568
rect 798 171024 429210 171288
rect 880 170744 429210 171024
rect 798 170480 429210 170744
rect 880 170200 429210 170480
rect 798 169936 429210 170200
rect 880 169656 429210 169936
rect 798 169392 429210 169656
rect 880 169112 429210 169392
rect 798 168848 429210 169112
rect 880 168568 429210 168848
rect 798 168304 429210 168568
rect 880 168024 429210 168304
rect 798 167760 429210 168024
rect 880 167480 429210 167760
rect 798 167216 429210 167480
rect 880 166936 429210 167216
rect 798 166672 429210 166936
rect 880 166392 429210 166672
rect 798 166128 429210 166392
rect 880 165848 429210 166128
rect 798 165584 429210 165848
rect 880 165304 429210 165584
rect 798 165040 429210 165304
rect 880 164760 429210 165040
rect 798 164496 429210 164760
rect 880 164216 429210 164496
rect 798 163952 429210 164216
rect 880 163672 429210 163952
rect 798 163408 429210 163672
rect 880 163128 429210 163408
rect 798 162864 429210 163128
rect 880 162584 429210 162864
rect 798 162320 429210 162584
rect 880 162040 429210 162320
rect 798 161776 429210 162040
rect 880 161496 429210 161776
rect 798 161232 429210 161496
rect 880 160952 429210 161232
rect 798 160688 429210 160952
rect 880 160408 429210 160688
rect 798 160144 429210 160408
rect 880 159864 429210 160144
rect 798 159600 429210 159864
rect 880 159320 429210 159600
rect 798 159056 429210 159320
rect 880 158776 429210 159056
rect 798 158512 429210 158776
rect 880 158232 429210 158512
rect 798 157968 429210 158232
rect 880 157688 429210 157968
rect 798 157424 429210 157688
rect 798 157144 429120 157424
rect 798 149264 429210 157144
rect 880 148984 429210 149264
rect 798 113360 429210 148984
rect 798 113080 429120 113360
rect 798 112816 429210 113080
rect 798 112536 429120 112816
rect 798 112272 429210 112536
rect 798 111992 429120 112272
rect 798 68208 429210 111992
rect 798 67928 429120 68208
rect 798 67664 429210 67928
rect 798 67384 429120 67664
rect 798 67120 429210 67384
rect 798 66840 429120 67120
rect 798 66576 429210 66840
rect 798 66296 429120 66576
rect 798 50800 429210 66296
rect 798 50520 429120 50800
rect 798 48624 429210 50520
rect 880 48344 429210 48624
rect 798 48080 429210 48344
rect 880 47800 429210 48080
rect 798 47536 429210 47800
rect 880 47256 429210 47536
rect 798 46992 429210 47256
rect 880 46712 429210 46992
rect 798 46448 429210 46712
rect 880 46168 429210 46448
rect 798 45904 429210 46168
rect 880 45624 429210 45904
rect 798 45360 429210 45624
rect 880 45080 429210 45360
rect 798 44816 429210 45080
rect 880 44536 429210 44816
rect 798 44272 429210 44536
rect 880 43992 429210 44272
rect 798 43728 429210 43992
rect 880 43448 429210 43728
rect 798 43184 429210 43448
rect 880 42904 429210 43184
rect 798 42640 429210 42904
rect 880 42360 429210 42640
rect 798 42096 429210 42360
rect 880 41816 429210 42096
rect 798 41552 429210 41816
rect 880 41272 429210 41552
rect 798 41008 429210 41272
rect 880 40728 429210 41008
rect 798 40464 429210 40728
rect 880 40184 429210 40464
rect 798 39920 429210 40184
rect 880 39640 429210 39920
rect 798 39376 429210 39640
rect 880 39096 429210 39376
rect 798 38832 429210 39096
rect 880 38552 429210 38832
rect 798 38288 429210 38552
rect 880 38008 429210 38288
rect 798 37744 429210 38008
rect 880 37464 429210 37744
rect 798 37200 429210 37464
rect 880 36920 429210 37200
rect 798 36656 429210 36920
rect 880 36376 429210 36656
rect 798 36112 429210 36376
rect 880 35832 429210 36112
rect 798 35568 429210 35832
rect 880 35288 429120 35568
rect 798 35024 429210 35288
rect 880 34744 429120 35024
rect 798 34480 429210 34744
rect 880 34200 429120 34480
rect 798 33936 429210 34200
rect 880 33656 429120 33936
rect 798 33392 429210 33656
rect 880 33112 429120 33392
rect 798 32848 429210 33112
rect 880 32568 429120 32848
rect 798 32304 429210 32568
rect 880 32024 429120 32304
rect 798 31760 429210 32024
rect 880 31480 429120 31760
rect 798 31216 429210 31480
rect 880 30936 429120 31216
rect 798 30672 429210 30936
rect 880 30392 429120 30672
rect 798 30128 429210 30392
rect 880 29848 429120 30128
rect 798 29584 429210 29848
rect 880 29304 429120 29584
rect 798 29040 429210 29304
rect 880 28760 429120 29040
rect 798 28496 429210 28760
rect 880 28216 429120 28496
rect 798 27952 429210 28216
rect 880 27672 429120 27952
rect 798 27408 429210 27672
rect 880 27128 429120 27408
rect 798 26864 429210 27128
rect 880 26584 429120 26864
rect 798 26320 429210 26584
rect 880 26040 429120 26320
rect 798 25776 429210 26040
rect 880 25496 429120 25776
rect 798 25232 429210 25496
rect 880 24952 429120 25232
rect 798 24688 429210 24952
rect 880 24408 429120 24688
rect 798 24144 429210 24408
rect 880 23864 429120 24144
rect 798 23600 429210 23864
rect 880 23320 429120 23600
rect 798 23056 429210 23320
rect 880 22776 429120 23056
rect 798 22512 429210 22776
rect 880 22232 429120 22512
rect 798 21968 429210 22232
rect 880 21688 429120 21968
rect 798 21424 429210 21688
rect 880 21144 429120 21424
rect 798 20880 429210 21144
rect 880 20600 429120 20880
rect 798 20336 429210 20600
rect 880 20056 429120 20336
rect 798 19792 429210 20056
rect 880 19512 429120 19792
rect 798 19248 429210 19512
rect 880 18968 429120 19248
rect 798 18704 429210 18968
rect 880 18424 429120 18704
rect 798 18160 429210 18424
rect 880 17880 429210 18160
rect 798 17616 429210 17880
rect 880 17336 429210 17616
rect 798 17072 429210 17336
rect 880 16792 429210 17072
rect 798 16528 429210 16792
rect 880 16248 429210 16528
rect 798 15984 429210 16248
rect 880 15704 429210 15984
rect 798 15440 429210 15704
rect 880 15160 429210 15440
rect 798 14896 429210 15160
rect 880 14616 429210 14896
rect 798 14352 429210 14616
rect 880 14072 429210 14352
rect 798 13808 429210 14072
rect 880 13528 429210 13808
rect 798 13264 429210 13528
rect 880 12984 429210 13264
rect 798 12720 429210 12984
rect 880 12440 429210 12720
rect 798 12176 429210 12440
rect 880 11896 429210 12176
rect 798 11632 429210 11896
rect 880 11352 429210 11632
rect 798 11088 429210 11352
rect 880 10808 429210 11088
rect 798 10544 429210 10808
rect 880 10264 429210 10544
rect 798 10000 429210 10264
rect 880 9720 429210 10000
rect 798 9456 429210 9720
rect 880 9176 429210 9456
rect 798 8912 429210 9176
rect 880 8632 429210 8912
rect 798 8368 429210 8632
rect 880 8088 429210 8368
rect 798 7824 429210 8088
rect 880 7544 429210 7824
rect 798 7280 429210 7544
rect 880 7000 429210 7280
rect 798 6736 429210 7000
rect 880 6456 429210 6736
rect 798 6192 429210 6456
rect 880 5912 429210 6192
rect 798 5648 429210 5912
rect 880 5368 429210 5648
rect 798 5104 429210 5368
rect 880 4824 429210 5104
rect 798 4560 429210 4824
rect 880 4280 429210 4560
rect 798 4016 429210 4280
rect 880 3736 429210 4016
rect 798 3472 429210 3736
rect 880 3192 429210 3472
rect 798 2928 429210 3192
rect 880 2648 429210 2928
rect 798 2384 429210 2648
rect 880 2104 429210 2384
rect 798 1840 429210 2104
rect 880 1560 429210 1840
rect 798 1296 429210 1560
rect 880 1016 429210 1296
rect 798 851 429210 1016
<< metal4 >>
rect 4208 2128 4528 177392
rect 9208 2128 9528 177392
rect 14208 2128 14528 177392
rect 19208 2128 19528 177392
rect 24208 2128 24528 177392
rect 29208 2128 29528 177392
rect 34208 2128 34528 177392
rect 39208 2128 39528 177392
rect 44208 2128 44528 177392
rect 49208 2128 49528 177392
rect 54208 2128 54528 177392
rect 59208 2128 59528 177392
rect 64208 137232 64528 177392
rect 69208 137232 69528 177392
rect 74208 137232 74528 177392
rect 79208 137232 79528 177392
rect 84208 137232 84528 177392
rect 89208 137232 89528 177392
rect 94208 137232 94528 177392
rect 99208 137232 99528 177392
rect 104208 137232 104528 177392
rect 109208 137232 109528 177392
rect 114208 137232 114528 177392
rect 119208 137232 119528 177392
rect 124208 137232 124528 177392
rect 129208 137232 129528 177392
rect 134208 137232 134528 177392
rect 139208 137232 139528 177392
rect 144208 137232 144528 177392
rect 149208 137232 149528 177392
rect 154208 137232 154528 177392
rect 159208 137232 159528 177392
rect 164208 137232 164528 177392
rect 169208 137232 169528 177392
rect 174208 137232 174528 177392
rect 179208 137232 179528 177392
rect 184208 137232 184528 177392
rect 189208 137232 189528 177392
rect 194208 137232 194528 177392
rect 199208 137232 199528 177392
rect 204208 137232 204528 177392
rect 209208 137232 209528 177392
rect 64208 2128 64528 30328
rect 69208 2128 69528 30328
rect 74208 2128 74528 30328
rect 79208 2128 79528 30328
rect 84208 2128 84528 30328
rect 89208 2128 89528 30328
rect 94208 2128 94528 30328
rect 99208 2128 99528 30328
rect 104208 2128 104528 30328
rect 109208 2128 109528 30328
rect 114208 2128 114528 30328
rect 119208 2128 119528 30328
rect 124208 2128 124528 30328
rect 129208 2128 129528 30328
rect 134208 2128 134528 30328
rect 139208 2128 139528 30328
rect 144208 2128 144528 30328
rect 149208 2128 149528 30328
rect 154208 2128 154528 30328
rect 159208 2128 159528 30328
rect 164208 2128 164528 30328
rect 169208 2128 169528 30328
rect 174208 2128 174528 30328
rect 179208 2128 179528 30328
rect 184208 2128 184528 30328
rect 189208 2128 189528 30328
rect 194208 2128 194528 30328
rect 199208 2128 199528 30328
rect 204208 2128 204528 30328
rect 209208 2128 209528 30328
rect 214208 2128 214528 177392
rect 219208 2128 219528 177392
rect 224208 2128 224528 177392
rect 229208 2128 229528 177392
rect 234208 2128 234528 177392
rect 239208 2128 239528 177392
rect 244208 2128 244528 177392
rect 249208 2128 249528 177392
rect 254208 2128 254528 177392
rect 259208 2128 259528 177392
rect 264208 2128 264528 177392
rect 269208 2128 269528 177392
rect 274208 2128 274528 177392
rect 279208 2128 279528 177392
rect 284208 2128 284528 177392
rect 289208 2128 289528 177392
rect 294208 2128 294528 177392
rect 299208 2128 299528 177392
rect 304208 2128 304528 177392
rect 309208 2128 309528 177392
rect 314208 2128 314528 177392
rect 319208 2128 319528 177392
rect 324208 2128 324528 177392
rect 329208 2128 329528 177392
rect 334208 2128 334528 177392
rect 339208 44168 339528 177392
rect 344208 44168 344528 177392
rect 349208 44168 349528 177392
rect 354208 44168 354528 177392
rect 359208 44168 359528 177392
rect 364208 44168 364528 177392
rect 369208 44168 369528 177392
rect 374208 44168 374528 177392
rect 379208 44168 379528 177392
rect 384208 2128 384528 177392
rect 389208 2128 389528 177392
rect 394208 2128 394528 177392
rect 399208 2128 399528 177392
rect 404208 2128 404528 177392
rect 409208 2128 409528 177392
rect 414208 2128 414528 177392
rect 419208 2128 419528 177392
rect 424208 2128 424528 177392
<< obsm4 >>
rect 3187 177472 425717 178669
rect 3187 2048 4128 177472
rect 4608 2048 9128 177472
rect 9608 2048 14128 177472
rect 14608 2048 19128 177472
rect 19608 2048 24128 177472
rect 24608 2048 29128 177472
rect 29608 2048 34128 177472
rect 34608 2048 39128 177472
rect 39608 2048 44128 177472
rect 44608 2048 49128 177472
rect 49608 2048 54128 177472
rect 54608 2048 59128 177472
rect 59608 137152 64128 177472
rect 64608 137152 69128 177472
rect 69608 137152 74128 177472
rect 74608 137152 79128 177472
rect 79608 137152 84128 177472
rect 84608 137152 89128 177472
rect 89608 137152 94128 177472
rect 94608 137152 99128 177472
rect 99608 137152 104128 177472
rect 104608 137152 109128 177472
rect 109608 137152 114128 177472
rect 114608 137152 119128 177472
rect 119608 137152 124128 177472
rect 124608 137152 129128 177472
rect 129608 137152 134128 177472
rect 134608 137152 139128 177472
rect 139608 137152 144128 177472
rect 144608 137152 149128 177472
rect 149608 137152 154128 177472
rect 154608 137152 159128 177472
rect 159608 137152 164128 177472
rect 164608 137152 169128 177472
rect 169608 137152 174128 177472
rect 174608 137152 179128 177472
rect 179608 137152 184128 177472
rect 184608 137152 189128 177472
rect 189608 137152 194128 177472
rect 194608 137152 199128 177472
rect 199608 137152 204128 177472
rect 204608 137152 209128 177472
rect 209608 137152 214128 177472
rect 59608 30408 214128 137152
rect 59608 2048 64128 30408
rect 64608 2048 69128 30408
rect 69608 2048 74128 30408
rect 74608 2048 79128 30408
rect 79608 2048 84128 30408
rect 84608 2048 89128 30408
rect 89608 2048 94128 30408
rect 94608 2048 99128 30408
rect 99608 2048 104128 30408
rect 104608 2048 109128 30408
rect 109608 2048 114128 30408
rect 114608 2048 119128 30408
rect 119608 2048 124128 30408
rect 124608 2048 129128 30408
rect 129608 2048 134128 30408
rect 134608 2048 139128 30408
rect 139608 2048 144128 30408
rect 144608 2048 149128 30408
rect 149608 2048 154128 30408
rect 154608 2048 159128 30408
rect 159608 2048 164128 30408
rect 164608 2048 169128 30408
rect 169608 2048 174128 30408
rect 174608 2048 179128 30408
rect 179608 2048 184128 30408
rect 184608 2048 189128 30408
rect 189608 2048 194128 30408
rect 194608 2048 199128 30408
rect 199608 2048 204128 30408
rect 204608 2048 209128 30408
rect 209608 2048 214128 30408
rect 214608 2048 219128 177472
rect 219608 2048 224128 177472
rect 224608 2048 229128 177472
rect 229608 2048 234128 177472
rect 234608 2048 239128 177472
rect 239608 2048 244128 177472
rect 244608 2048 249128 177472
rect 249608 2048 254128 177472
rect 254608 2048 259128 177472
rect 259608 2048 264128 177472
rect 264608 2048 269128 177472
rect 269608 2048 274128 177472
rect 274608 2048 279128 177472
rect 279608 2048 284128 177472
rect 284608 2048 289128 177472
rect 289608 2048 294128 177472
rect 294608 2048 299128 177472
rect 299608 2048 304128 177472
rect 304608 2048 309128 177472
rect 309608 2048 314128 177472
rect 314608 2048 319128 177472
rect 319608 2048 324128 177472
rect 324608 2048 329128 177472
rect 329608 2048 334128 177472
rect 334608 44088 339128 177472
rect 339608 44088 344128 177472
rect 344608 44088 349128 177472
rect 349608 44088 354128 177472
rect 354608 44088 359128 177472
rect 359608 44088 364128 177472
rect 364608 44088 369128 177472
rect 369608 44088 374128 177472
rect 374608 44088 379128 177472
rect 379608 44088 384128 177472
rect 334608 2048 384128 44088
rect 384608 2048 389128 177472
rect 389608 2048 394128 177472
rect 394608 2048 399128 177472
rect 399608 2048 404128 177472
rect 404608 2048 409128 177472
rect 409608 2048 414128 177472
rect 414608 2048 419128 177472
rect 419608 2048 424128 177472
rect 424608 2048 425717 177472
rect 3187 851 425717 2048
<< metal5 >>
rect 1104 173796 428812 174116
rect 1104 158478 428812 158798
rect 1104 143160 428812 143480
rect 1104 127842 428812 128162
rect 1104 112524 428812 112844
rect 1104 97206 428812 97526
rect 1104 81888 428812 82208
rect 1104 66570 428812 66890
rect 1104 51252 428812 51572
rect 1104 35934 428812 36254
rect 1104 20616 428812 20936
rect 1104 5298 428812 5618
<< obsm5 >>
rect 60652 174436 350036 175260
rect 60652 159118 350036 173476
rect 60652 143800 350036 158158
rect 60652 128482 350036 142840
rect 60652 113164 350036 127522
rect 60652 97846 350036 112204
rect 60652 82528 350036 96886
rect 60652 67210 350036 81568
rect 60652 51892 350036 66250
rect 60652 47100 350036 50932
<< labels >>
rlabel metal2 s 570 0 626 800 6 clock
port 1 nsew signal input
rlabel metal2 s 11794 179200 11850 180000 6 core_clk
port 2 nsew signal output
rlabel metal2 s 77298 179200 77354 180000 6 core_rstn
port 3 nsew signal output
rlabel metal2 s 938 0 994 800 6 flash_clk
port 4 nsew signal output
rlabel metal3 s 0 1096 800 1216 6 flash_clk_ieb
port 5 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 flash_clk_oeb
port 6 nsew signal output
rlabel metal3 s 0 1640 800 1760 6 flash_csb
port 7 nsew signal output
rlabel metal2 s 1674 0 1730 800 6 flash_csb_ieb
port 8 nsew signal output
rlabel metal2 s 2042 0 2098 800 6 flash_csb_oeb
port 9 nsew signal output
rlabel metal3 s 0 2184 800 2304 6 flash_io0_di
port 10 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 flash_io0_do
port 11 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 flash_io0_ieb
port 12 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 flash_io0_oeb
port 13 nsew signal output
rlabel metal2 s 3146 0 3202 800 6 flash_io1_di
port 14 nsew signal input
rlabel metal3 s 0 3272 800 3392 6 flash_io1_do
port 15 nsew signal output
rlabel metal2 s 3514 0 3570 800 6 flash_io1_ieb
port 16 nsew signal output
rlabel metal3 s 0 3816 800 3936 6 flash_io1_oeb
port 17 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 gpio_in_pad
port 18 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 gpio_inenb_pad
port 19 nsew signal output
rlabel metal3 s 0 4360 800 4480 6 gpio_mode0_pad
port 20 nsew signal output
rlabel metal2 s 4618 0 4674 800 6 gpio_mode1_pad
port 21 nsew signal output
rlabel metal3 s 0 4904 800 5024 6 gpio_out_pad
port 22 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 gpio_outenb_pad
port 23 nsew signal output
rlabel metal3 s 429200 67464 430000 67584 6 jtag_out
port 24 nsew signal output
rlabel metal3 s 429200 66920 430000 67040 6 jtag_outenb
port 25 nsew signal output
rlabel metal2 s 77666 179200 77722 180000 6 la_input[0]
port 26 nsew signal input
rlabel metal2 s 76930 179200 76986 180000 6 la_input[100]
port 27 nsew signal input
rlabel metal2 s 78034 179200 78090 180000 6 la_input[101]
port 28 nsew signal input
rlabel metal2 s 76562 179200 76618 180000 6 la_input[102]
port 29 nsew signal input
rlabel metal2 s 78402 179200 78458 180000 6 la_input[103]
port 30 nsew signal input
rlabel metal2 s 76194 179200 76250 180000 6 la_input[104]
port 31 nsew signal input
rlabel metal2 s 78770 179200 78826 180000 6 la_input[105]
port 32 nsew signal input
rlabel metal2 s 75826 179200 75882 180000 6 la_input[106]
port 33 nsew signal input
rlabel metal2 s 79138 179200 79194 180000 6 la_input[107]
port 34 nsew signal input
rlabel metal2 s 75458 179200 75514 180000 6 la_input[108]
port 35 nsew signal input
rlabel metal2 s 79506 179200 79562 180000 6 la_input[109]
port 36 nsew signal input
rlabel metal2 s 75090 179200 75146 180000 6 la_input[10]
port 37 nsew signal input
rlabel metal2 s 79874 179200 79930 180000 6 la_input[110]
port 38 nsew signal input
rlabel metal2 s 74722 179200 74778 180000 6 la_input[111]
port 39 nsew signal input
rlabel metal2 s 80242 179200 80298 180000 6 la_input[112]
port 40 nsew signal input
rlabel metal2 s 74354 179200 74410 180000 6 la_input[113]
port 41 nsew signal input
rlabel metal2 s 80610 179200 80666 180000 6 la_input[114]
port 42 nsew signal input
rlabel metal2 s 73986 179200 74042 180000 6 la_input[115]
port 43 nsew signal input
rlabel metal2 s 80978 179200 81034 180000 6 la_input[116]
port 44 nsew signal input
rlabel metal2 s 73618 179200 73674 180000 6 la_input[117]
port 45 nsew signal input
rlabel metal2 s 81346 179200 81402 180000 6 la_input[118]
port 46 nsew signal input
rlabel metal2 s 73250 179200 73306 180000 6 la_input[119]
port 47 nsew signal input
rlabel metal2 s 81714 179200 81770 180000 6 la_input[11]
port 48 nsew signal input
rlabel metal2 s 72882 179200 72938 180000 6 la_input[120]
port 49 nsew signal input
rlabel metal2 s 82082 179200 82138 180000 6 la_input[121]
port 50 nsew signal input
rlabel metal2 s 72514 179200 72570 180000 6 la_input[122]
port 51 nsew signal input
rlabel metal2 s 82450 179200 82506 180000 6 la_input[123]
port 52 nsew signal input
rlabel metal2 s 72146 179200 72202 180000 6 la_input[124]
port 53 nsew signal input
rlabel metal2 s 82818 179200 82874 180000 6 la_input[125]
port 54 nsew signal input
rlabel metal2 s 71778 179200 71834 180000 6 la_input[126]
port 55 nsew signal input
rlabel metal2 s 83186 179200 83242 180000 6 la_input[127]
port 56 nsew signal input
rlabel metal2 s 71410 179200 71466 180000 6 la_input[12]
port 57 nsew signal input
rlabel metal2 s 83554 179200 83610 180000 6 la_input[13]
port 58 nsew signal input
rlabel metal2 s 71042 179200 71098 180000 6 la_input[14]
port 59 nsew signal input
rlabel metal2 s 83922 179200 83978 180000 6 la_input[15]
port 60 nsew signal input
rlabel metal2 s 70674 179200 70730 180000 6 la_input[16]
port 61 nsew signal input
rlabel metal2 s 84290 179200 84346 180000 6 la_input[17]
port 62 nsew signal input
rlabel metal2 s 70306 179200 70362 180000 6 la_input[18]
port 63 nsew signal input
rlabel metal2 s 84658 179200 84714 180000 6 la_input[19]
port 64 nsew signal input
rlabel metal2 s 69938 179200 69994 180000 6 la_input[1]
port 65 nsew signal input
rlabel metal2 s 85026 179200 85082 180000 6 la_input[20]
port 66 nsew signal input
rlabel metal2 s 69570 179200 69626 180000 6 la_input[21]
port 67 nsew signal input
rlabel metal2 s 85394 179200 85450 180000 6 la_input[22]
port 68 nsew signal input
rlabel metal2 s 69202 179200 69258 180000 6 la_input[23]
port 69 nsew signal input
rlabel metal2 s 85762 179200 85818 180000 6 la_input[24]
port 70 nsew signal input
rlabel metal2 s 68834 179200 68890 180000 6 la_input[25]
port 71 nsew signal input
rlabel metal2 s 86130 179200 86186 180000 6 la_input[26]
port 72 nsew signal input
rlabel metal2 s 68466 179200 68522 180000 6 la_input[27]
port 73 nsew signal input
rlabel metal2 s 86498 179200 86554 180000 6 la_input[28]
port 74 nsew signal input
rlabel metal2 s 68098 179200 68154 180000 6 la_input[29]
port 75 nsew signal input
rlabel metal2 s 86866 179200 86922 180000 6 la_input[2]
port 76 nsew signal input
rlabel metal2 s 67730 179200 67786 180000 6 la_input[30]
port 77 nsew signal input
rlabel metal2 s 87234 179200 87290 180000 6 la_input[31]
port 78 nsew signal input
rlabel metal2 s 67362 179200 67418 180000 6 la_input[32]
port 79 nsew signal input
rlabel metal2 s 87602 179200 87658 180000 6 la_input[33]
port 80 nsew signal input
rlabel metal2 s 66994 179200 67050 180000 6 la_input[34]
port 81 nsew signal input
rlabel metal2 s 87970 179200 88026 180000 6 la_input[35]
port 82 nsew signal input
rlabel metal2 s 66626 179200 66682 180000 6 la_input[36]
port 83 nsew signal input
rlabel metal2 s 88338 179200 88394 180000 6 la_input[37]
port 84 nsew signal input
rlabel metal2 s 66258 179200 66314 180000 6 la_input[38]
port 85 nsew signal input
rlabel metal2 s 88706 179200 88762 180000 6 la_input[39]
port 86 nsew signal input
rlabel metal2 s 65890 179200 65946 180000 6 la_input[3]
port 87 nsew signal input
rlabel metal2 s 89074 179200 89130 180000 6 la_input[40]
port 88 nsew signal input
rlabel metal2 s 65522 179200 65578 180000 6 la_input[41]
port 89 nsew signal input
rlabel metal2 s 89442 179200 89498 180000 6 la_input[42]
port 90 nsew signal input
rlabel metal2 s 65154 179200 65210 180000 6 la_input[43]
port 91 nsew signal input
rlabel metal2 s 89810 179200 89866 180000 6 la_input[44]
port 92 nsew signal input
rlabel metal2 s 64786 179200 64842 180000 6 la_input[45]
port 93 nsew signal input
rlabel metal2 s 90178 179200 90234 180000 6 la_input[46]
port 94 nsew signal input
rlabel metal2 s 64418 179200 64474 180000 6 la_input[47]
port 95 nsew signal input
rlabel metal2 s 90546 179200 90602 180000 6 la_input[48]
port 96 nsew signal input
rlabel metal2 s 64050 179200 64106 180000 6 la_input[49]
port 97 nsew signal input
rlabel metal2 s 90914 179200 90970 180000 6 la_input[4]
port 98 nsew signal input
rlabel metal2 s 63682 179200 63738 180000 6 la_input[50]
port 99 nsew signal input
rlabel metal2 s 91282 179200 91338 180000 6 la_input[51]
port 100 nsew signal input
rlabel metal2 s 63314 179200 63370 180000 6 la_input[52]
port 101 nsew signal input
rlabel metal2 s 91650 179200 91706 180000 6 la_input[53]
port 102 nsew signal input
rlabel metal2 s 62946 179200 63002 180000 6 la_input[54]
port 103 nsew signal input
rlabel metal2 s 92018 179200 92074 180000 6 la_input[55]
port 104 nsew signal input
rlabel metal2 s 62578 179200 62634 180000 6 la_input[56]
port 105 nsew signal input
rlabel metal2 s 92386 179200 92442 180000 6 la_input[57]
port 106 nsew signal input
rlabel metal2 s 62210 179200 62266 180000 6 la_input[58]
port 107 nsew signal input
rlabel metal2 s 92754 179200 92810 180000 6 la_input[59]
port 108 nsew signal input
rlabel metal2 s 61842 179200 61898 180000 6 la_input[5]
port 109 nsew signal input
rlabel metal2 s 93122 179200 93178 180000 6 la_input[60]
port 110 nsew signal input
rlabel metal2 s 61474 179200 61530 180000 6 la_input[61]
port 111 nsew signal input
rlabel metal2 s 93490 179200 93546 180000 6 la_input[62]
port 112 nsew signal input
rlabel metal2 s 61106 179200 61162 180000 6 la_input[63]
port 113 nsew signal input
rlabel metal2 s 93858 179200 93914 180000 6 la_input[64]
port 114 nsew signal input
rlabel metal2 s 60738 179200 60794 180000 6 la_input[65]
port 115 nsew signal input
rlabel metal2 s 94226 179200 94282 180000 6 la_input[66]
port 116 nsew signal input
rlabel metal2 s 60370 179200 60426 180000 6 la_input[67]
port 117 nsew signal input
rlabel metal2 s 94594 179200 94650 180000 6 la_input[68]
port 118 nsew signal input
rlabel metal2 s 60002 179200 60058 180000 6 la_input[69]
port 119 nsew signal input
rlabel metal2 s 94962 179200 95018 180000 6 la_input[6]
port 120 nsew signal input
rlabel metal2 s 59634 179200 59690 180000 6 la_input[70]
port 121 nsew signal input
rlabel metal2 s 95330 179200 95386 180000 6 la_input[71]
port 122 nsew signal input
rlabel metal2 s 59266 179200 59322 180000 6 la_input[72]
port 123 nsew signal input
rlabel metal2 s 95698 179200 95754 180000 6 la_input[73]
port 124 nsew signal input
rlabel metal2 s 58898 179200 58954 180000 6 la_input[74]
port 125 nsew signal input
rlabel metal2 s 96066 179200 96122 180000 6 la_input[75]
port 126 nsew signal input
rlabel metal2 s 58530 179200 58586 180000 6 la_input[76]
port 127 nsew signal input
rlabel metal2 s 96434 179200 96490 180000 6 la_input[77]
port 128 nsew signal input
rlabel metal2 s 58162 179200 58218 180000 6 la_input[78]
port 129 nsew signal input
rlabel metal2 s 96802 179200 96858 180000 6 la_input[79]
port 130 nsew signal input
rlabel metal2 s 57794 179200 57850 180000 6 la_input[7]
port 131 nsew signal input
rlabel metal2 s 97170 179200 97226 180000 6 la_input[80]
port 132 nsew signal input
rlabel metal2 s 57426 179200 57482 180000 6 la_input[81]
port 133 nsew signal input
rlabel metal2 s 97538 179200 97594 180000 6 la_input[82]
port 134 nsew signal input
rlabel metal2 s 57058 179200 57114 180000 6 la_input[83]
port 135 nsew signal input
rlabel metal2 s 97906 179200 97962 180000 6 la_input[84]
port 136 nsew signal input
rlabel metal2 s 56690 179200 56746 180000 6 la_input[85]
port 137 nsew signal input
rlabel metal2 s 98274 179200 98330 180000 6 la_input[86]
port 138 nsew signal input
rlabel metal2 s 56322 179200 56378 180000 6 la_input[87]
port 139 nsew signal input
rlabel metal2 s 98642 179200 98698 180000 6 la_input[88]
port 140 nsew signal input
rlabel metal2 s 55954 179200 56010 180000 6 la_input[89]
port 141 nsew signal input
rlabel metal2 s 99010 179200 99066 180000 6 la_input[8]
port 142 nsew signal input
rlabel metal2 s 55586 179200 55642 180000 6 la_input[90]
port 143 nsew signal input
rlabel metal2 s 99378 179200 99434 180000 6 la_input[91]
port 144 nsew signal input
rlabel metal2 s 55218 179200 55274 180000 6 la_input[92]
port 145 nsew signal input
rlabel metal2 s 99746 179200 99802 180000 6 la_input[93]
port 146 nsew signal input
rlabel metal2 s 54850 179200 54906 180000 6 la_input[94]
port 147 nsew signal input
rlabel metal2 s 100114 179200 100170 180000 6 la_input[95]
port 148 nsew signal input
rlabel metal2 s 54482 179200 54538 180000 6 la_input[96]
port 149 nsew signal input
rlabel metal2 s 100482 179200 100538 180000 6 la_input[97]
port 150 nsew signal input
rlabel metal2 s 54114 179200 54170 180000 6 la_input[98]
port 151 nsew signal input
rlabel metal2 s 100850 179200 100906 180000 6 la_input[99]
port 152 nsew signal input
rlabel metal2 s 53746 179200 53802 180000 6 la_input[9]
port 153 nsew signal input
rlabel metal2 s 101218 179200 101274 180000 6 la_oen[0]
port 154 nsew signal output
rlabel metal2 s 53378 179200 53434 180000 6 la_oen[100]
port 155 nsew signal output
rlabel metal2 s 101586 179200 101642 180000 6 la_oen[101]
port 156 nsew signal output
rlabel metal2 s 53010 179200 53066 180000 6 la_oen[102]
port 157 nsew signal output
rlabel metal2 s 101954 179200 102010 180000 6 la_oen[103]
port 158 nsew signal output
rlabel metal2 s 52642 179200 52698 180000 6 la_oen[104]
port 159 nsew signal output
rlabel metal2 s 102322 179200 102378 180000 6 la_oen[105]
port 160 nsew signal output
rlabel metal2 s 52274 179200 52330 180000 6 la_oen[106]
port 161 nsew signal output
rlabel metal2 s 102690 179200 102746 180000 6 la_oen[107]
port 162 nsew signal output
rlabel metal2 s 51906 179200 51962 180000 6 la_oen[108]
port 163 nsew signal output
rlabel metal2 s 103058 179200 103114 180000 6 la_oen[109]
port 164 nsew signal output
rlabel metal2 s 51538 179200 51594 180000 6 la_oen[10]
port 165 nsew signal output
rlabel metal2 s 103426 179200 103482 180000 6 la_oen[110]
port 166 nsew signal output
rlabel metal2 s 51170 179200 51226 180000 6 la_oen[111]
port 167 nsew signal output
rlabel metal2 s 103794 179200 103850 180000 6 la_oen[112]
port 168 nsew signal output
rlabel metal2 s 50802 179200 50858 180000 6 la_oen[113]
port 169 nsew signal output
rlabel metal2 s 104162 179200 104218 180000 6 la_oen[114]
port 170 nsew signal output
rlabel metal2 s 50434 179200 50490 180000 6 la_oen[115]
port 171 nsew signal output
rlabel metal2 s 104530 179200 104586 180000 6 la_oen[116]
port 172 nsew signal output
rlabel metal2 s 50066 179200 50122 180000 6 la_oen[117]
port 173 nsew signal output
rlabel metal2 s 104898 179200 104954 180000 6 la_oen[118]
port 174 nsew signal output
rlabel metal2 s 49698 179200 49754 180000 6 la_oen[119]
port 175 nsew signal output
rlabel metal2 s 105266 179200 105322 180000 6 la_oen[11]
port 176 nsew signal output
rlabel metal2 s 49330 179200 49386 180000 6 la_oen[120]
port 177 nsew signal output
rlabel metal2 s 105634 179200 105690 180000 6 la_oen[121]
port 178 nsew signal output
rlabel metal2 s 48962 179200 49018 180000 6 la_oen[122]
port 179 nsew signal output
rlabel metal2 s 106002 179200 106058 180000 6 la_oen[123]
port 180 nsew signal output
rlabel metal2 s 48594 179200 48650 180000 6 la_oen[124]
port 181 nsew signal output
rlabel metal2 s 106370 179200 106426 180000 6 la_oen[125]
port 182 nsew signal output
rlabel metal2 s 48226 179200 48282 180000 6 la_oen[126]
port 183 nsew signal output
rlabel metal2 s 106738 179200 106794 180000 6 la_oen[127]
port 184 nsew signal output
rlabel metal2 s 47858 179200 47914 180000 6 la_oen[12]
port 185 nsew signal output
rlabel metal2 s 107106 179200 107162 180000 6 la_oen[13]
port 186 nsew signal output
rlabel metal2 s 47490 179200 47546 180000 6 la_oen[14]
port 187 nsew signal output
rlabel metal2 s 107474 179200 107530 180000 6 la_oen[15]
port 188 nsew signal output
rlabel metal2 s 47122 179200 47178 180000 6 la_oen[16]
port 189 nsew signal output
rlabel metal2 s 107842 179200 107898 180000 6 la_oen[17]
port 190 nsew signal output
rlabel metal2 s 46754 179200 46810 180000 6 la_oen[18]
port 191 nsew signal output
rlabel metal2 s 108210 179200 108266 180000 6 la_oen[19]
port 192 nsew signal output
rlabel metal2 s 46386 179200 46442 180000 6 la_oen[1]
port 193 nsew signal output
rlabel metal2 s 108578 179200 108634 180000 6 la_oen[20]
port 194 nsew signal output
rlabel metal2 s 46018 179200 46074 180000 6 la_oen[21]
port 195 nsew signal output
rlabel metal2 s 108946 179200 109002 180000 6 la_oen[22]
port 196 nsew signal output
rlabel metal2 s 45650 179200 45706 180000 6 la_oen[23]
port 197 nsew signal output
rlabel metal2 s 109314 179200 109370 180000 6 la_oen[24]
port 198 nsew signal output
rlabel metal2 s 45282 179200 45338 180000 6 la_oen[25]
port 199 nsew signal output
rlabel metal2 s 109682 179200 109738 180000 6 la_oen[26]
port 200 nsew signal output
rlabel metal2 s 44914 179200 44970 180000 6 la_oen[27]
port 201 nsew signal output
rlabel metal2 s 110050 179200 110106 180000 6 la_oen[28]
port 202 nsew signal output
rlabel metal2 s 44546 179200 44602 180000 6 la_oen[29]
port 203 nsew signal output
rlabel metal2 s 110418 179200 110474 180000 6 la_oen[2]
port 204 nsew signal output
rlabel metal2 s 44178 179200 44234 180000 6 la_oen[30]
port 205 nsew signal output
rlabel metal2 s 110786 179200 110842 180000 6 la_oen[31]
port 206 nsew signal output
rlabel metal2 s 43810 179200 43866 180000 6 la_oen[32]
port 207 nsew signal output
rlabel metal2 s 111154 179200 111210 180000 6 la_oen[33]
port 208 nsew signal output
rlabel metal2 s 43442 179200 43498 180000 6 la_oen[34]
port 209 nsew signal output
rlabel metal2 s 111522 179200 111578 180000 6 la_oen[35]
port 210 nsew signal output
rlabel metal2 s 43074 179200 43130 180000 6 la_oen[36]
port 211 nsew signal output
rlabel metal2 s 111890 179200 111946 180000 6 la_oen[37]
port 212 nsew signal output
rlabel metal2 s 42706 179200 42762 180000 6 la_oen[38]
port 213 nsew signal output
rlabel metal2 s 112258 179200 112314 180000 6 la_oen[39]
port 214 nsew signal output
rlabel metal2 s 42338 179200 42394 180000 6 la_oen[3]
port 215 nsew signal output
rlabel metal2 s 112626 179200 112682 180000 6 la_oen[40]
port 216 nsew signal output
rlabel metal2 s 41970 179200 42026 180000 6 la_oen[41]
port 217 nsew signal output
rlabel metal2 s 112994 179200 113050 180000 6 la_oen[42]
port 218 nsew signal output
rlabel metal2 s 41602 179200 41658 180000 6 la_oen[43]
port 219 nsew signal output
rlabel metal2 s 113362 179200 113418 180000 6 la_oen[44]
port 220 nsew signal output
rlabel metal2 s 41234 179200 41290 180000 6 la_oen[45]
port 221 nsew signal output
rlabel metal2 s 113730 179200 113786 180000 6 la_oen[46]
port 222 nsew signal output
rlabel metal2 s 40866 179200 40922 180000 6 la_oen[47]
port 223 nsew signal output
rlabel metal2 s 114098 179200 114154 180000 6 la_oen[48]
port 224 nsew signal output
rlabel metal2 s 40498 179200 40554 180000 6 la_oen[49]
port 225 nsew signal output
rlabel metal2 s 114466 179200 114522 180000 6 la_oen[4]
port 226 nsew signal output
rlabel metal2 s 40130 179200 40186 180000 6 la_oen[50]
port 227 nsew signal output
rlabel metal2 s 114834 179200 114890 180000 6 la_oen[51]
port 228 nsew signal output
rlabel metal2 s 39762 179200 39818 180000 6 la_oen[52]
port 229 nsew signal output
rlabel metal2 s 115202 179200 115258 180000 6 la_oen[53]
port 230 nsew signal output
rlabel metal2 s 39394 179200 39450 180000 6 la_oen[54]
port 231 nsew signal output
rlabel metal2 s 115570 179200 115626 180000 6 la_oen[55]
port 232 nsew signal output
rlabel metal2 s 39026 179200 39082 180000 6 la_oen[56]
port 233 nsew signal output
rlabel metal2 s 115938 179200 115994 180000 6 la_oen[57]
port 234 nsew signal output
rlabel metal2 s 38658 179200 38714 180000 6 la_oen[58]
port 235 nsew signal output
rlabel metal2 s 116306 179200 116362 180000 6 la_oen[59]
port 236 nsew signal output
rlabel metal2 s 38290 179200 38346 180000 6 la_oen[5]
port 237 nsew signal output
rlabel metal2 s 116674 179200 116730 180000 6 la_oen[60]
port 238 nsew signal output
rlabel metal2 s 37922 179200 37978 180000 6 la_oen[61]
port 239 nsew signal output
rlabel metal2 s 117042 179200 117098 180000 6 la_oen[62]
port 240 nsew signal output
rlabel metal2 s 37554 179200 37610 180000 6 la_oen[63]
port 241 nsew signal output
rlabel metal2 s 117410 179200 117466 180000 6 la_oen[64]
port 242 nsew signal output
rlabel metal2 s 37186 179200 37242 180000 6 la_oen[65]
port 243 nsew signal output
rlabel metal2 s 117778 179200 117834 180000 6 la_oen[66]
port 244 nsew signal output
rlabel metal2 s 36818 179200 36874 180000 6 la_oen[67]
port 245 nsew signal output
rlabel metal2 s 118146 179200 118202 180000 6 la_oen[68]
port 246 nsew signal output
rlabel metal2 s 36450 179200 36506 180000 6 la_oen[69]
port 247 nsew signal output
rlabel metal2 s 118514 179200 118570 180000 6 la_oen[6]
port 248 nsew signal output
rlabel metal2 s 36082 179200 36138 180000 6 la_oen[70]
port 249 nsew signal output
rlabel metal2 s 118882 179200 118938 180000 6 la_oen[71]
port 250 nsew signal output
rlabel metal2 s 35714 179200 35770 180000 6 la_oen[72]
port 251 nsew signal output
rlabel metal2 s 119250 179200 119306 180000 6 la_oen[73]
port 252 nsew signal output
rlabel metal2 s 35346 179200 35402 180000 6 la_oen[74]
port 253 nsew signal output
rlabel metal2 s 119618 179200 119674 180000 6 la_oen[75]
port 254 nsew signal output
rlabel metal2 s 34978 179200 35034 180000 6 la_oen[76]
port 255 nsew signal output
rlabel metal2 s 119986 179200 120042 180000 6 la_oen[77]
port 256 nsew signal output
rlabel metal2 s 34610 179200 34666 180000 6 la_oen[78]
port 257 nsew signal output
rlabel metal2 s 120354 179200 120410 180000 6 la_oen[79]
port 258 nsew signal output
rlabel metal2 s 34242 179200 34298 180000 6 la_oen[7]
port 259 nsew signal output
rlabel metal2 s 120722 179200 120778 180000 6 la_oen[80]
port 260 nsew signal output
rlabel metal2 s 33874 179200 33930 180000 6 la_oen[81]
port 261 nsew signal output
rlabel metal2 s 121090 179200 121146 180000 6 la_oen[82]
port 262 nsew signal output
rlabel metal2 s 33506 179200 33562 180000 6 la_oen[83]
port 263 nsew signal output
rlabel metal2 s 121458 179200 121514 180000 6 la_oen[84]
port 264 nsew signal output
rlabel metal2 s 33138 179200 33194 180000 6 la_oen[85]
port 265 nsew signal output
rlabel metal2 s 121826 179200 121882 180000 6 la_oen[86]
port 266 nsew signal output
rlabel metal2 s 32770 179200 32826 180000 6 la_oen[87]
port 267 nsew signal output
rlabel metal2 s 122194 179200 122250 180000 6 la_oen[88]
port 268 nsew signal output
rlabel metal2 s 32402 179200 32458 180000 6 la_oen[89]
port 269 nsew signal output
rlabel metal2 s 122562 179200 122618 180000 6 la_oen[8]
port 270 nsew signal output
rlabel metal2 s 32034 179200 32090 180000 6 la_oen[90]
port 271 nsew signal output
rlabel metal2 s 122930 179200 122986 180000 6 la_oen[91]
port 272 nsew signal output
rlabel metal2 s 31666 179200 31722 180000 6 la_oen[92]
port 273 nsew signal output
rlabel metal2 s 123298 179200 123354 180000 6 la_oen[93]
port 274 nsew signal output
rlabel metal2 s 31298 179200 31354 180000 6 la_oen[94]
port 275 nsew signal output
rlabel metal2 s 123666 179200 123722 180000 6 la_oen[95]
port 276 nsew signal output
rlabel metal2 s 30930 179200 30986 180000 6 la_oen[96]
port 277 nsew signal output
rlabel metal2 s 124034 179200 124090 180000 6 la_oen[97]
port 278 nsew signal output
rlabel metal2 s 30562 179200 30618 180000 6 la_oen[98]
port 279 nsew signal output
rlabel metal2 s 124402 179200 124458 180000 6 la_oen[99]
port 280 nsew signal output
rlabel metal2 s 30194 179200 30250 180000 6 la_oen[9]
port 281 nsew signal output
rlabel metal2 s 124770 179200 124826 180000 6 la_output[0]
port 282 nsew signal output
rlabel metal2 s 29826 179200 29882 180000 6 la_output[100]
port 283 nsew signal output
rlabel metal2 s 125138 179200 125194 180000 6 la_output[101]
port 284 nsew signal output
rlabel metal2 s 29458 179200 29514 180000 6 la_output[102]
port 285 nsew signal output
rlabel metal2 s 125506 179200 125562 180000 6 la_output[103]
port 286 nsew signal output
rlabel metal2 s 29090 179200 29146 180000 6 la_output[104]
port 287 nsew signal output
rlabel metal2 s 125874 179200 125930 180000 6 la_output[105]
port 288 nsew signal output
rlabel metal2 s 28722 179200 28778 180000 6 la_output[106]
port 289 nsew signal output
rlabel metal2 s 126242 179200 126298 180000 6 la_output[107]
port 290 nsew signal output
rlabel metal2 s 28354 179200 28410 180000 6 la_output[108]
port 291 nsew signal output
rlabel metal2 s 126610 179200 126666 180000 6 la_output[109]
port 292 nsew signal output
rlabel metal2 s 27986 179200 28042 180000 6 la_output[10]
port 293 nsew signal output
rlabel metal2 s 126978 179200 127034 180000 6 la_output[110]
port 294 nsew signal output
rlabel metal2 s 27618 179200 27674 180000 6 la_output[111]
port 295 nsew signal output
rlabel metal2 s 127346 179200 127402 180000 6 la_output[112]
port 296 nsew signal output
rlabel metal2 s 27250 179200 27306 180000 6 la_output[113]
port 297 nsew signal output
rlabel metal2 s 127714 179200 127770 180000 6 la_output[114]
port 298 nsew signal output
rlabel metal2 s 26882 179200 26938 180000 6 la_output[115]
port 299 nsew signal output
rlabel metal2 s 128082 179200 128138 180000 6 la_output[116]
port 300 nsew signal output
rlabel metal2 s 26514 179200 26570 180000 6 la_output[117]
port 301 nsew signal output
rlabel metal2 s 128450 179200 128506 180000 6 la_output[118]
port 302 nsew signal output
rlabel metal2 s 26146 179200 26202 180000 6 la_output[119]
port 303 nsew signal output
rlabel metal2 s 128818 179200 128874 180000 6 la_output[11]
port 304 nsew signal output
rlabel metal2 s 25778 179200 25834 180000 6 la_output[120]
port 305 nsew signal output
rlabel metal2 s 129186 179200 129242 180000 6 la_output[121]
port 306 nsew signal output
rlabel metal2 s 25410 179200 25466 180000 6 la_output[122]
port 307 nsew signal output
rlabel metal2 s 129554 179200 129610 180000 6 la_output[123]
port 308 nsew signal output
rlabel metal2 s 25042 179200 25098 180000 6 la_output[124]
port 309 nsew signal output
rlabel metal2 s 129922 179200 129978 180000 6 la_output[125]
port 310 nsew signal output
rlabel metal2 s 24674 179200 24730 180000 6 la_output[126]
port 311 nsew signal output
rlabel metal2 s 130290 179200 130346 180000 6 la_output[127]
port 312 nsew signal output
rlabel metal2 s 24306 179200 24362 180000 6 la_output[12]
port 313 nsew signal output
rlabel metal2 s 130658 179200 130714 180000 6 la_output[13]
port 314 nsew signal output
rlabel metal2 s 23938 179200 23994 180000 6 la_output[14]
port 315 nsew signal output
rlabel metal2 s 131026 179200 131082 180000 6 la_output[15]
port 316 nsew signal output
rlabel metal2 s 23570 179200 23626 180000 6 la_output[16]
port 317 nsew signal output
rlabel metal2 s 131394 179200 131450 180000 6 la_output[17]
port 318 nsew signal output
rlabel metal2 s 23202 179200 23258 180000 6 la_output[18]
port 319 nsew signal output
rlabel metal2 s 131762 179200 131818 180000 6 la_output[19]
port 320 nsew signal output
rlabel metal2 s 22834 179200 22890 180000 6 la_output[1]
port 321 nsew signal output
rlabel metal2 s 132130 179200 132186 180000 6 la_output[20]
port 322 nsew signal output
rlabel metal2 s 22466 179200 22522 180000 6 la_output[21]
port 323 nsew signal output
rlabel metal2 s 132498 179200 132554 180000 6 la_output[22]
port 324 nsew signal output
rlabel metal2 s 22098 179200 22154 180000 6 la_output[23]
port 325 nsew signal output
rlabel metal2 s 132866 179200 132922 180000 6 la_output[24]
port 326 nsew signal output
rlabel metal2 s 21730 179200 21786 180000 6 la_output[25]
port 327 nsew signal output
rlabel metal2 s 133234 179200 133290 180000 6 la_output[26]
port 328 nsew signal output
rlabel metal2 s 21362 179200 21418 180000 6 la_output[27]
port 329 nsew signal output
rlabel metal2 s 133602 179200 133658 180000 6 la_output[28]
port 330 nsew signal output
rlabel metal2 s 20994 179200 21050 180000 6 la_output[29]
port 331 nsew signal output
rlabel metal2 s 133970 179200 134026 180000 6 la_output[2]
port 332 nsew signal output
rlabel metal2 s 20626 179200 20682 180000 6 la_output[30]
port 333 nsew signal output
rlabel metal2 s 134338 179200 134394 180000 6 la_output[31]
port 334 nsew signal output
rlabel metal2 s 20258 179200 20314 180000 6 la_output[32]
port 335 nsew signal output
rlabel metal2 s 134706 179200 134762 180000 6 la_output[33]
port 336 nsew signal output
rlabel metal2 s 19890 179200 19946 180000 6 la_output[34]
port 337 nsew signal output
rlabel metal2 s 135074 179200 135130 180000 6 la_output[35]
port 338 nsew signal output
rlabel metal2 s 19522 179200 19578 180000 6 la_output[36]
port 339 nsew signal output
rlabel metal2 s 135442 179200 135498 180000 6 la_output[37]
port 340 nsew signal output
rlabel metal2 s 19154 179200 19210 180000 6 la_output[38]
port 341 nsew signal output
rlabel metal2 s 135810 179200 135866 180000 6 la_output[39]
port 342 nsew signal output
rlabel metal2 s 18786 179200 18842 180000 6 la_output[3]
port 343 nsew signal output
rlabel metal2 s 136178 179200 136234 180000 6 la_output[40]
port 344 nsew signal output
rlabel metal2 s 18418 179200 18474 180000 6 la_output[41]
port 345 nsew signal output
rlabel metal2 s 136546 179200 136602 180000 6 la_output[42]
port 346 nsew signal output
rlabel metal2 s 18050 179200 18106 180000 6 la_output[43]
port 347 nsew signal output
rlabel metal2 s 136914 179200 136970 180000 6 la_output[44]
port 348 nsew signal output
rlabel metal2 s 17682 179200 17738 180000 6 la_output[45]
port 349 nsew signal output
rlabel metal2 s 137282 179200 137338 180000 6 la_output[46]
port 350 nsew signal output
rlabel metal2 s 17314 179200 17370 180000 6 la_output[47]
port 351 nsew signal output
rlabel metal2 s 137650 179200 137706 180000 6 la_output[48]
port 352 nsew signal output
rlabel metal2 s 16946 179200 17002 180000 6 la_output[49]
port 353 nsew signal output
rlabel metal2 s 138018 179200 138074 180000 6 la_output[4]
port 354 nsew signal output
rlabel metal2 s 16578 179200 16634 180000 6 la_output[50]
port 355 nsew signal output
rlabel metal2 s 138386 179200 138442 180000 6 la_output[51]
port 356 nsew signal output
rlabel metal2 s 16210 179200 16266 180000 6 la_output[52]
port 357 nsew signal output
rlabel metal2 s 138754 179200 138810 180000 6 la_output[53]
port 358 nsew signal output
rlabel metal2 s 15842 179200 15898 180000 6 la_output[54]
port 359 nsew signal output
rlabel metal2 s 139122 179200 139178 180000 6 la_output[55]
port 360 nsew signal output
rlabel metal2 s 15474 179200 15530 180000 6 la_output[56]
port 361 nsew signal output
rlabel metal2 s 139490 179200 139546 180000 6 la_output[57]
port 362 nsew signal output
rlabel metal2 s 15106 179200 15162 180000 6 la_output[58]
port 363 nsew signal output
rlabel metal2 s 139858 179200 139914 180000 6 la_output[59]
port 364 nsew signal output
rlabel metal2 s 14738 179200 14794 180000 6 la_output[5]
port 365 nsew signal output
rlabel metal2 s 140226 179200 140282 180000 6 la_output[60]
port 366 nsew signal output
rlabel metal2 s 14370 179200 14426 180000 6 la_output[61]
port 367 nsew signal output
rlabel metal2 s 140594 179200 140650 180000 6 la_output[62]
port 368 nsew signal output
rlabel metal2 s 14002 179200 14058 180000 6 la_output[63]
port 369 nsew signal output
rlabel metal2 s 140962 179200 141018 180000 6 la_output[64]
port 370 nsew signal output
rlabel metal2 s 13634 179200 13690 180000 6 la_output[65]
port 371 nsew signal output
rlabel metal2 s 141330 179200 141386 180000 6 la_output[66]
port 372 nsew signal output
rlabel metal2 s 13266 179200 13322 180000 6 la_output[67]
port 373 nsew signal output
rlabel metal2 s 141698 179200 141754 180000 6 la_output[68]
port 374 nsew signal output
rlabel metal2 s 12898 179200 12954 180000 6 la_output[69]
port 375 nsew signal output
rlabel metal2 s 142066 179200 142122 180000 6 la_output[6]
port 376 nsew signal output
rlabel metal2 s 12530 179200 12586 180000 6 la_output[70]
port 377 nsew signal output
rlabel metal2 s 142434 179200 142490 180000 6 la_output[71]
port 378 nsew signal output
rlabel metal2 s 12162 179200 12218 180000 6 la_output[72]
port 379 nsew signal output
rlabel metal2 s 142802 179200 142858 180000 6 la_output[73]
port 380 nsew signal output
rlabel metal2 s 143170 179200 143226 180000 6 la_output[74]
port 381 nsew signal output
rlabel metal2 s 11426 179200 11482 180000 6 la_output[75]
port 382 nsew signal output
rlabel metal2 s 143538 179200 143594 180000 6 la_output[76]
port 383 nsew signal output
rlabel metal2 s 11058 179200 11114 180000 6 la_output[77]
port 384 nsew signal output
rlabel metal2 s 143906 179200 143962 180000 6 la_output[78]
port 385 nsew signal output
rlabel metal2 s 10690 179200 10746 180000 6 la_output[79]
port 386 nsew signal output
rlabel metal2 s 144274 179200 144330 180000 6 la_output[7]
port 387 nsew signal output
rlabel metal2 s 10322 179200 10378 180000 6 la_output[80]
port 388 nsew signal output
rlabel metal2 s 144642 179200 144698 180000 6 la_output[81]
port 389 nsew signal output
rlabel metal2 s 9954 179200 10010 180000 6 la_output[82]
port 390 nsew signal output
rlabel metal2 s 145010 179200 145066 180000 6 la_output[83]
port 391 nsew signal output
rlabel metal2 s 9586 179200 9642 180000 6 la_output[84]
port 392 nsew signal output
rlabel metal2 s 145378 179200 145434 180000 6 la_output[85]
port 393 nsew signal output
rlabel metal2 s 9218 179200 9274 180000 6 la_output[86]
port 394 nsew signal output
rlabel metal2 s 145746 179200 145802 180000 6 la_output[87]
port 395 nsew signal output
rlabel metal2 s 8850 179200 8906 180000 6 la_output[88]
port 396 nsew signal output
rlabel metal2 s 146114 179200 146170 180000 6 la_output[89]
port 397 nsew signal output
rlabel metal2 s 8482 179200 8538 180000 6 la_output[8]
port 398 nsew signal output
rlabel metal2 s 146482 179200 146538 180000 6 la_output[90]
port 399 nsew signal output
rlabel metal2 s 8114 179200 8170 180000 6 la_output[91]
port 400 nsew signal output
rlabel metal2 s 146850 179200 146906 180000 6 la_output[92]
port 401 nsew signal output
rlabel metal2 s 7746 179200 7802 180000 6 la_output[93]
port 402 nsew signal output
rlabel metal2 s 147218 179200 147274 180000 6 la_output[94]
port 403 nsew signal output
rlabel metal2 s 7378 179200 7434 180000 6 la_output[95]
port 404 nsew signal output
rlabel metal2 s 147586 179200 147642 180000 6 la_output[96]
port 405 nsew signal output
rlabel metal2 s 7010 179200 7066 180000 6 la_output[97]
port 406 nsew signal output
rlabel metal2 s 147954 179200 148010 180000 6 la_output[98]
port 407 nsew signal output
rlabel metal2 s 6642 179200 6698 180000 6 la_output[99]
port 408 nsew signal output
rlabel metal2 s 148322 179200 148378 180000 6 la_output[9]
port 409 nsew signal output
rlabel metal3 s 429200 27208 430000 27328 6 mask_rev[0]
port 410 nsew signal input
rlabel metal3 s 429200 26664 430000 26784 6 mask_rev[10]
port 411 nsew signal input
rlabel metal3 s 429200 27752 430000 27872 6 mask_rev[11]
port 412 nsew signal input
rlabel metal3 s 429200 26120 430000 26240 6 mask_rev[12]
port 413 nsew signal input
rlabel metal3 s 429200 28296 430000 28416 6 mask_rev[13]
port 414 nsew signal input
rlabel metal3 s 429200 25576 430000 25696 6 mask_rev[14]
port 415 nsew signal input
rlabel metal3 s 429200 28840 430000 28960 6 mask_rev[15]
port 416 nsew signal input
rlabel metal3 s 429200 25032 430000 25152 6 mask_rev[16]
port 417 nsew signal input
rlabel metal3 s 429200 29384 430000 29504 6 mask_rev[17]
port 418 nsew signal input
rlabel metal3 s 429200 24488 430000 24608 6 mask_rev[18]
port 419 nsew signal input
rlabel metal3 s 429200 29928 430000 30048 6 mask_rev[19]
port 420 nsew signal input
rlabel metal3 s 429200 23944 430000 24064 6 mask_rev[1]
port 421 nsew signal input
rlabel metal3 s 429200 30472 430000 30592 6 mask_rev[20]
port 422 nsew signal input
rlabel metal3 s 429200 23400 430000 23520 6 mask_rev[21]
port 423 nsew signal input
rlabel metal3 s 429200 31016 430000 31136 6 mask_rev[22]
port 424 nsew signal input
rlabel metal3 s 429200 22856 430000 22976 6 mask_rev[23]
port 425 nsew signal input
rlabel metal3 s 429200 31560 430000 31680 6 mask_rev[24]
port 426 nsew signal input
rlabel metal3 s 429200 22312 430000 22432 6 mask_rev[25]
port 427 nsew signal input
rlabel metal3 s 429200 32104 430000 32224 6 mask_rev[26]
port 428 nsew signal input
rlabel metal3 s 429200 21768 430000 21888 6 mask_rev[27]
port 429 nsew signal input
rlabel metal3 s 429200 32648 430000 32768 6 mask_rev[28]
port 430 nsew signal input
rlabel metal3 s 429200 21224 430000 21344 6 mask_rev[29]
port 431 nsew signal input
rlabel metal3 s 429200 33192 430000 33312 6 mask_rev[2]
port 432 nsew signal input
rlabel metal3 s 429200 20680 430000 20800 6 mask_rev[30]
port 433 nsew signal input
rlabel metal3 s 429200 33736 430000 33856 6 mask_rev[31]
port 434 nsew signal input
rlabel metal3 s 429200 20136 430000 20256 6 mask_rev[3]
port 435 nsew signal input
rlabel metal3 s 429200 34280 430000 34400 6 mask_rev[4]
port 436 nsew signal input
rlabel metal3 s 429200 19592 430000 19712 6 mask_rev[5]
port 437 nsew signal input
rlabel metal3 s 429200 34824 430000 34944 6 mask_rev[6]
port 438 nsew signal input
rlabel metal3 s 429200 19048 430000 19168 6 mask_rev[7]
port 439 nsew signal input
rlabel metal3 s 429200 35368 430000 35488 6 mask_rev[8]
port 440 nsew signal input
rlabel metal3 s 429200 18504 430000 18624 6 mask_rev[9]
port 441 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 mgmt_addr[0]
port 442 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 mgmt_addr[1]
port 443 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 mgmt_addr[2]
port 444 nsew signal output
rlabel metal3 s 0 8712 800 8832 6 mgmt_addr[3]
port 445 nsew signal output
rlabel metal3 s 0 6536 800 6656 6 mgmt_addr[4]
port 446 nsew signal output
rlabel metal3 s 0 9256 800 9376 6 mgmt_addr[5]
port 447 nsew signal output
rlabel metal3 s 0 5992 800 6112 6 mgmt_addr[6]
port 448 nsew signal output
rlabel metal3 s 0 9800 800 9920 6 mgmt_addr[7]
port 449 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 mgmt_addr_ro[0]
port 450 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 mgmt_addr_ro[1]
port 451 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 mgmt_addr_ro[2]
port 452 nsew signal output
rlabel metal3 s 0 11432 800 11552 6 mgmt_addr_ro[3]
port 453 nsew signal output
rlabel metal3 s 0 11976 800 12096 6 mgmt_addr_ro[4]
port 454 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 mgmt_addr_ro[5]
port 455 nsew signal output
rlabel metal3 s 0 13064 800 13184 6 mgmt_addr_ro[6]
port 456 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 mgmt_addr_ro[7]
port 457 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 mgmt_ena[0]
port 458 nsew signal output
rlabel metal3 s 0 14696 800 14816 6 mgmt_ena[1]
port 459 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 mgmt_ena_ro
port 460 nsew signal output
rlabel metal3 s 429200 68008 430000 68128 6 mgmt_in_data[0]
port 461 nsew signal input
rlabel metal2 s 754 0 810 800 6 mgmt_in_data[10]
port 462 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 mgmt_in_data[11]
port 463 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 mgmt_in_data[12]
port 464 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 mgmt_in_data[13]
port 465 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 mgmt_in_data[14]
port 466 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 mgmt_in_data[15]
port 467 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 mgmt_in_data[16]
port 468 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 mgmt_in_data[17]
port 469 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 mgmt_in_data[18]
port 470 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 mgmt_in_data[19]
port 471 nsew signal input
rlabel metal3 s 429200 112616 430000 112736 6 mgmt_in_data[1]
port 472 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 mgmt_in_data[20]
port 473 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 mgmt_in_data[21]
port 474 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 mgmt_in_data[22]
port 475 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 mgmt_in_data[23]
port 476 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 mgmt_in_data[24]
port 477 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 mgmt_in_data[25]
port 478 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 mgmt_in_data[26]
port 479 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 mgmt_in_data[27]
port 480 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 mgmt_in_data[28]
port 481 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 mgmt_in_data[29]
port 482 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 mgmt_in_data[2]
port 483 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 mgmt_in_data[30]
port 484 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 mgmt_in_data[31]
port 485 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 mgmt_in_data[32]
port 486 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 mgmt_in_data[33]
port 487 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 mgmt_in_data[34]
port 488 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 mgmt_in_data[35]
port 489 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 mgmt_in_data[36]
port 490 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 mgmt_in_data[37]
port 491 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 mgmt_in_data[3]
port 492 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 mgmt_in_data[4]
port 493 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 mgmt_in_data[5]
port 494 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 mgmt_in_data[6]
port 495 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 mgmt_in_data[7]
port 496 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 mgmt_in_data[8]
port 497 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 mgmt_in_data[9]
port 498 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 mgmt_out_data[0]
port 499 nsew signal output
rlabel metal2 s 429106 179200 429162 180000 6 mgmt_out_data[10]
port 500 nsew signal output
rlabel metal3 s 429200 178984 430000 179104 6 mgmt_out_data[11]
port 501 nsew signal output
rlabel metal2 s 428738 179200 428794 180000 6 mgmt_out_data[12]
port 502 nsew signal output
rlabel metal3 s 429200 178440 430000 178560 6 mgmt_out_data[13]
port 503 nsew signal output
rlabel metal2 s 428370 179200 428426 180000 6 mgmt_out_data[14]
port 504 nsew signal output
rlabel metal2 s 338578 179200 338634 180000 6 mgmt_out_data[15]
port 505 nsew signal output
rlabel metal2 s 287058 179200 287114 180000 6 mgmt_out_data[16]
port 506 nsew signal output
rlabel metal2 s 210146 179200 210202 180000 6 mgmt_out_data[17]
port 507 nsew signal output
rlabel metal2 s 148690 179200 148746 180000 6 mgmt_out_data[18]
port 508 nsew signal output
rlabel metal2 s 149058 179200 149114 180000 6 mgmt_out_data[19]
port 509 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 mgmt_out_data[1]
port 510 nsew signal output
rlabel metal2 s 6274 179200 6330 180000 6 mgmt_out_data[20]
port 511 nsew signal output
rlabel metal2 s 754 179200 810 180000 6 mgmt_out_data[21]
port 512 nsew signal output
rlabel metal3 s 0 178984 800 179104 6 mgmt_out_data[22]
port 513 nsew signal output
rlabel metal2 s 1122 179200 1178 180000 6 mgmt_out_data[23]
port 514 nsew signal output
rlabel metal3 s 0 178440 800 178560 6 mgmt_out_data[24]
port 515 nsew signal output
rlabel metal2 s 1490 179200 1546 180000 6 mgmt_out_data[25]
port 516 nsew signal output
rlabel metal2 s 1858 179200 1914 180000 6 mgmt_out_data[26]
port 517 nsew signal output
rlabel metal3 s 0 177896 800 178016 6 mgmt_out_data[27]
port 518 nsew signal output
rlabel metal2 s 2226 179200 2282 180000 6 mgmt_out_data[28]
port 519 nsew signal output
rlabel metal3 s 0 177352 800 177472 6 mgmt_out_data[29]
port 520 nsew signal output
rlabel metal3 s 429200 157224 430000 157344 6 mgmt_out_data[2]
port 521 nsew signal output
rlabel metal2 s 2594 179200 2650 180000 6 mgmt_out_data[30]
port 522 nsew signal output
rlabel metal2 s 2962 179200 3018 180000 6 mgmt_out_data[31]
port 523 nsew signal output
rlabel metal3 s 0 176808 800 176928 6 mgmt_out_data[32]
port 524 nsew signal output
rlabel metal2 s 3330 179200 3386 180000 6 mgmt_out_data[33]
port 525 nsew signal output
rlabel metal3 s 0 176264 800 176384 6 mgmt_out_data[34]
port 526 nsew signal output
rlabel metal2 s 3698 179200 3754 180000 6 mgmt_out_data[35]
port 527 nsew signal output
rlabel metal2 s 4066 179200 4122 180000 6 mgmt_out_data[36]
port 528 nsew signal output
rlabel metal3 s 0 149064 800 149184 6 mgmt_out_data[37]
port 529 nsew signal output
rlabel metal2 s 428002 179200 428058 180000 6 mgmt_out_data[3]
port 530 nsew signal output
rlabel metal3 s 429200 177896 430000 178016 6 mgmt_out_data[4]
port 531 nsew signal output
rlabel metal2 s 427634 179200 427690 180000 6 mgmt_out_data[5]
port 532 nsew signal output
rlabel metal3 s 429200 177352 430000 177472 6 mgmt_out_data[6]
port 533 nsew signal output
rlabel metal2 s 427266 179200 427322 180000 6 mgmt_out_data[7]
port 534 nsew signal output
rlabel metal2 s 426898 179200 426954 180000 6 mgmt_out_data[8]
port 535 nsew signal output
rlabel metal3 s 429200 176808 430000 176928 6 mgmt_out_data[9]
port 536 nsew signal output
rlabel metal3 s 0 15784 800 15904 6 mgmt_rdata[0]
port 537 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 mgmt_rdata[10]
port 538 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 mgmt_rdata[11]
port 539 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 mgmt_rdata[12]
port 540 nsew signal input
rlabel metal3 s 0 17960 800 18080 6 mgmt_rdata[13]
port 541 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 mgmt_rdata[14]
port 542 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 mgmt_rdata[15]
port 543 nsew signal input
rlabel metal3 s 0 19592 800 19712 6 mgmt_rdata[16]
port 544 nsew signal input
rlabel metal3 s 0 20136 800 20256 6 mgmt_rdata[17]
port 545 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 mgmt_rdata[18]
port 546 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 mgmt_rdata[19]
port 547 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 mgmt_rdata[1]
port 548 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 mgmt_rdata[20]
port 549 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 mgmt_rdata[21]
port 550 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 mgmt_rdata[22]
port 551 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 mgmt_rdata[23]
port 552 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 mgmt_rdata[24]
port 553 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 mgmt_rdata[25]
port 554 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 mgmt_rdata[26]
port 555 nsew signal input
rlabel metal3 s 0 22856 800 22976 6 mgmt_rdata[27]
port 556 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 mgmt_rdata[28]
port 557 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 mgmt_rdata[29]
port 558 nsew signal input
rlabel metal3 s 0 23400 800 23520 6 mgmt_rdata[2]
port 559 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 mgmt_rdata[30]
port 560 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 mgmt_rdata[31]
port 561 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 mgmt_rdata[32]
port 562 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 mgmt_rdata[33]
port 563 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 mgmt_rdata[34]
port 564 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 mgmt_rdata[35]
port 565 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 mgmt_rdata[36]
port 566 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 mgmt_rdata[37]
port 567 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 mgmt_rdata[38]
port 568 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 mgmt_rdata[39]
port 569 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 mgmt_rdata[3]
port 570 nsew signal input
rlabel metal3 s 0 26120 800 26240 6 mgmt_rdata[40]
port 571 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 mgmt_rdata[41]
port 572 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 mgmt_rdata[42]
port 573 nsew signal input
rlabel metal3 s 0 26664 800 26784 6 mgmt_rdata[43]
port 574 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 mgmt_rdata[44]
port 575 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 mgmt_rdata[45]
port 576 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 mgmt_rdata[46]
port 577 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 mgmt_rdata[47]
port 578 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 mgmt_rdata[48]
port 579 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 mgmt_rdata[49]
port 580 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 mgmt_rdata[4]
port 581 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 mgmt_rdata[50]
port 582 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 mgmt_rdata[51]
port 583 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 mgmt_rdata[52]
port 584 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 mgmt_rdata[53]
port 585 nsew signal input
rlabel metal3 s 0 29384 800 29504 6 mgmt_rdata[54]
port 586 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 mgmt_rdata[55]
port 587 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 mgmt_rdata[56]
port 588 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 mgmt_rdata[57]
port 589 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 mgmt_rdata[58]
port 590 nsew signal input
rlabel metal3 s 0 30472 800 30592 6 mgmt_rdata[59]
port 591 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 mgmt_rdata[5]
port 592 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 mgmt_rdata[60]
port 593 nsew signal input
rlabel metal3 s 0 31016 800 31136 6 mgmt_rdata[61]
port 594 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 mgmt_rdata[62]
port 595 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 mgmt_rdata[63]
port 596 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 mgmt_rdata[6]
port 597 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 mgmt_rdata[7]
port 598 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 mgmt_rdata[8]
port 599 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 mgmt_rdata[9]
port 600 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 mgmt_rdata_ro[0]
port 601 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 mgmt_rdata_ro[10]
port 602 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 mgmt_rdata_ro[11]
port 603 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 mgmt_rdata_ro[12]
port 604 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 mgmt_rdata_ro[13]
port 605 nsew signal input
rlabel metal3 s 0 33736 800 33856 6 mgmt_rdata_ro[14]
port 606 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 mgmt_rdata_ro[15]
port 607 nsew signal input
rlabel metal3 s 0 34280 800 34400 6 mgmt_rdata_ro[16]
port 608 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 mgmt_rdata_ro[17]
port 609 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 mgmt_rdata_ro[18]
port 610 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 mgmt_rdata_ro[19]
port 611 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 mgmt_rdata_ro[1]
port 612 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 mgmt_rdata_ro[20]
port 613 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 mgmt_rdata_ro[21]
port 614 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 mgmt_rdata_ro[22]
port 615 nsew signal input
rlabel metal3 s 0 35912 800 36032 6 mgmt_rdata_ro[23]
port 616 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 mgmt_rdata_ro[24]
port 617 nsew signal input
rlabel metal3 s 0 36456 800 36576 6 mgmt_rdata_ro[25]
port 618 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 mgmt_rdata_ro[26]
port 619 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 mgmt_rdata_ro[27]
port 620 nsew signal input
rlabel metal3 s 0 37000 800 37120 6 mgmt_rdata_ro[28]
port 621 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 mgmt_rdata_ro[29]
port 622 nsew signal input
rlabel metal3 s 0 37544 800 37664 6 mgmt_rdata_ro[2]
port 623 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 mgmt_rdata_ro[30]
port 624 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 mgmt_rdata_ro[31]
port 625 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 mgmt_rdata_ro[3]
port 626 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 mgmt_rdata_ro[4]
port 627 nsew signal input
rlabel metal3 s 0 38632 800 38752 6 mgmt_rdata_ro[5]
port 628 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 mgmt_rdata_ro[6]
port 629 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 mgmt_rdata_ro[7]
port 630 nsew signal input
rlabel metal3 s 0 39176 800 39296 6 mgmt_rdata_ro[8]
port 631 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 mgmt_rdata_ro[9]
port 632 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 mgmt_wdata[0]
port 633 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 mgmt_wdata[10]
port 634 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 mgmt_wdata[11]
port 635 nsew signal output
rlabel metal3 s 0 40264 800 40384 6 mgmt_wdata[12]
port 636 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 mgmt_wdata[13]
port 637 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 mgmt_wdata[14]
port 638 nsew signal output
rlabel metal2 s 25594 0 25650 800 6 mgmt_wdata[15]
port 639 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 mgmt_wdata[16]
port 640 nsew signal output
rlabel metal3 s 0 41352 800 41472 6 mgmt_wdata[17]
port 641 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 mgmt_wdata[18]
port 642 nsew signal output
rlabel metal3 s 0 41896 800 42016 6 mgmt_wdata[19]
port 643 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 mgmt_wdata[1]
port 644 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 mgmt_wdata[20]
port 645 nsew signal output
rlabel metal3 s 0 42440 800 42560 6 mgmt_wdata[21]
port 646 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 mgmt_wdata[22]
port 647 nsew signal output
rlabel metal3 s 0 42984 800 43104 6 mgmt_wdata[23]
port 648 nsew signal output
rlabel metal2 s 27802 0 27858 800 6 mgmt_wdata[24]
port 649 nsew signal output
rlabel metal2 s 28170 0 28226 800 6 mgmt_wdata[25]
port 650 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 mgmt_wdata[26]
port 651 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 mgmt_wdata[27]
port 652 nsew signal output
rlabel metal3 s 0 44072 800 44192 6 mgmt_wdata[28]
port 653 nsew signal output
rlabel metal2 s 28906 0 28962 800 6 mgmt_wdata[29]
port 654 nsew signal output
rlabel metal3 s 0 44616 800 44736 6 mgmt_wdata[2]
port 655 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 mgmt_wdata[30]
port 656 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 mgmt_wdata[31]
port 657 nsew signal output
rlabel metal3 s 0 45160 800 45280 6 mgmt_wdata[3]
port 658 nsew signal output
rlabel metal2 s 30010 0 30066 800 6 mgmt_wdata[4]
port 659 nsew signal output
rlabel metal3 s 0 45704 800 45824 6 mgmt_wdata[5]
port 660 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 mgmt_wdata[6]
port 661 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 mgmt_wdata[7]
port 662 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 mgmt_wdata[8]
port 663 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 mgmt_wdata[9]
port 664 nsew signal output
rlabel metal3 s 0 46792 800 46912 6 mgmt_wen[0]
port 665 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 mgmt_wen[1]
port 666 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 mgmt_wen_mask[0]
port 667 nsew signal output
rlabel metal3 s 0 47336 800 47456 6 mgmt_wen_mask[1]
port 668 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 mgmt_wen_mask[2]
port 669 nsew signal output
rlabel metal3 s 0 47880 800 48000 6 mgmt_wen_mask[3]
port 670 nsew signal output
rlabel metal2 s 32586 0 32642 800 6 mgmt_wen_mask[4]
port 671 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 mgmt_wen_mask[5]
port 672 nsew signal output
rlabel metal3 s 0 48424 800 48544 6 mgmt_wen_mask[6]
port 673 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 mgmt_wen_mask[7]
port 674 nsew signal output
rlabel metal2 s 5906 179200 5962 180000 6 mprj2_vcc_pwrgood
port 675 nsew signal input
rlabel metal2 s 5538 179200 5594 180000 6 mprj2_vdd_pwrgood
port 676 nsew signal input
rlabel metal3 s 0 175720 800 175840 6 mprj_ack_i
port 677 nsew signal input
rlabel metal2 s 149426 179200 149482 180000 6 mprj_adr_o[0]
port 678 nsew signal output
rlabel metal2 s 5170 179200 5226 180000 6 mprj_adr_o[10]
port 679 nsew signal output
rlabel metal2 s 149794 179200 149850 180000 6 mprj_adr_o[11]
port 680 nsew signal output
rlabel metal2 s 4802 179200 4858 180000 6 mprj_adr_o[12]
port 681 nsew signal output
rlabel metal2 s 150162 179200 150218 180000 6 mprj_adr_o[13]
port 682 nsew signal output
rlabel metal2 s 4434 179200 4490 180000 6 mprj_adr_o[14]
port 683 nsew signal output
rlabel metal2 s 150530 179200 150586 180000 6 mprj_adr_o[15]
port 684 nsew signal output
rlabel metal2 s 150898 179200 150954 180000 6 mprj_adr_o[16]
port 685 nsew signal output
rlabel metal2 s 151266 179200 151322 180000 6 mprj_adr_o[17]
port 686 nsew signal output
rlabel metal2 s 151634 179200 151690 180000 6 mprj_adr_o[18]
port 687 nsew signal output
rlabel metal2 s 152002 179200 152058 180000 6 mprj_adr_o[19]
port 688 nsew signal output
rlabel metal2 s 152370 179200 152426 180000 6 mprj_adr_o[1]
port 689 nsew signal output
rlabel metal2 s 152738 179200 152794 180000 6 mprj_adr_o[20]
port 690 nsew signal output
rlabel metal2 s 153106 179200 153162 180000 6 mprj_adr_o[21]
port 691 nsew signal output
rlabel metal2 s 153474 179200 153530 180000 6 mprj_adr_o[22]
port 692 nsew signal output
rlabel metal2 s 153842 179200 153898 180000 6 mprj_adr_o[23]
port 693 nsew signal output
rlabel metal2 s 154210 179200 154266 180000 6 mprj_adr_o[24]
port 694 nsew signal output
rlabel metal2 s 154578 179200 154634 180000 6 mprj_adr_o[25]
port 695 nsew signal output
rlabel metal2 s 154946 179200 155002 180000 6 mprj_adr_o[26]
port 696 nsew signal output
rlabel metal2 s 155314 179200 155370 180000 6 mprj_adr_o[27]
port 697 nsew signal output
rlabel metal2 s 155682 179200 155738 180000 6 mprj_adr_o[28]
port 698 nsew signal output
rlabel metal2 s 156050 179200 156106 180000 6 mprj_adr_o[29]
port 699 nsew signal output
rlabel metal2 s 156418 179200 156474 180000 6 mprj_adr_o[2]
port 700 nsew signal output
rlabel metal2 s 156786 179200 156842 180000 6 mprj_adr_o[30]
port 701 nsew signal output
rlabel metal2 s 157154 179200 157210 180000 6 mprj_adr_o[31]
port 702 nsew signal output
rlabel metal2 s 157522 179200 157578 180000 6 mprj_adr_o[3]
port 703 nsew signal output
rlabel metal2 s 157890 179200 157946 180000 6 mprj_adr_o[4]
port 704 nsew signal output
rlabel metal2 s 158258 179200 158314 180000 6 mprj_adr_o[5]
port 705 nsew signal output
rlabel metal2 s 158626 179200 158682 180000 6 mprj_adr_o[6]
port 706 nsew signal output
rlabel metal2 s 158994 179200 159050 180000 6 mprj_adr_o[7]
port 707 nsew signal output
rlabel metal2 s 159362 179200 159418 180000 6 mprj_adr_o[8]
port 708 nsew signal output
rlabel metal2 s 159730 179200 159786 180000 6 mprj_adr_o[9]
port 709 nsew signal output
rlabel metal3 s 0 175176 800 175296 6 mprj_cyc_o
port 710 nsew signal output
rlabel metal3 s 0 174632 800 174752 6 mprj_dat_i[0]
port 711 nsew signal input
rlabel metal3 s 0 174088 800 174208 6 mprj_dat_i[10]
port 712 nsew signal input
rlabel metal3 s 0 173544 800 173664 6 mprj_dat_i[11]
port 713 nsew signal input
rlabel metal3 s 0 173000 800 173120 6 mprj_dat_i[12]
port 714 nsew signal input
rlabel metal3 s 0 172456 800 172576 6 mprj_dat_i[13]
port 715 nsew signal input
rlabel metal3 s 0 171912 800 172032 6 mprj_dat_i[14]
port 716 nsew signal input
rlabel metal3 s 0 171368 800 171488 6 mprj_dat_i[15]
port 717 nsew signal input
rlabel metal3 s 0 170824 800 170944 6 mprj_dat_i[16]
port 718 nsew signal input
rlabel metal3 s 0 170280 800 170400 6 mprj_dat_i[17]
port 719 nsew signal input
rlabel metal3 s 0 169736 800 169856 6 mprj_dat_i[18]
port 720 nsew signal input
rlabel metal3 s 0 169192 800 169312 6 mprj_dat_i[19]
port 721 nsew signal input
rlabel metal3 s 0 168648 800 168768 6 mprj_dat_i[1]
port 722 nsew signal input
rlabel metal3 s 0 168104 800 168224 6 mprj_dat_i[20]
port 723 nsew signal input
rlabel metal3 s 0 167560 800 167680 6 mprj_dat_i[21]
port 724 nsew signal input
rlabel metal3 s 0 167016 800 167136 6 mprj_dat_i[22]
port 725 nsew signal input
rlabel metal3 s 0 166472 800 166592 6 mprj_dat_i[23]
port 726 nsew signal input
rlabel metal3 s 0 165928 800 166048 6 mprj_dat_i[24]
port 727 nsew signal input
rlabel metal3 s 0 165384 800 165504 6 mprj_dat_i[25]
port 728 nsew signal input
rlabel metal3 s 0 164840 800 164960 6 mprj_dat_i[26]
port 729 nsew signal input
rlabel metal3 s 0 164296 800 164416 6 mprj_dat_i[27]
port 730 nsew signal input
rlabel metal3 s 0 163752 800 163872 6 mprj_dat_i[28]
port 731 nsew signal input
rlabel metal3 s 0 163208 800 163328 6 mprj_dat_i[29]
port 732 nsew signal input
rlabel metal3 s 0 162664 800 162784 6 mprj_dat_i[2]
port 733 nsew signal input
rlabel metal3 s 0 162120 800 162240 6 mprj_dat_i[30]
port 734 nsew signal input
rlabel metal3 s 0 161576 800 161696 6 mprj_dat_i[31]
port 735 nsew signal input
rlabel metal3 s 0 161032 800 161152 6 mprj_dat_i[3]
port 736 nsew signal input
rlabel metal3 s 0 160488 800 160608 6 mprj_dat_i[4]
port 737 nsew signal input
rlabel metal3 s 0 159944 800 160064 6 mprj_dat_i[5]
port 738 nsew signal input
rlabel metal3 s 0 159400 800 159520 6 mprj_dat_i[6]
port 739 nsew signal input
rlabel metal3 s 0 158856 800 158976 6 mprj_dat_i[7]
port 740 nsew signal input
rlabel metal3 s 0 158312 800 158432 6 mprj_dat_i[8]
port 741 nsew signal input
rlabel metal3 s 0 157768 800 157888 6 mprj_dat_i[9]
port 742 nsew signal input
rlabel metal2 s 160098 179200 160154 180000 6 mprj_dat_o[0]
port 743 nsew signal output
rlabel metal2 s 160466 179200 160522 180000 6 mprj_dat_o[10]
port 744 nsew signal output
rlabel metal2 s 160834 179200 160890 180000 6 mprj_dat_o[11]
port 745 nsew signal output
rlabel metal2 s 161202 179200 161258 180000 6 mprj_dat_o[12]
port 746 nsew signal output
rlabel metal2 s 161570 179200 161626 180000 6 mprj_dat_o[13]
port 747 nsew signal output
rlabel metal2 s 161938 179200 161994 180000 6 mprj_dat_o[14]
port 748 nsew signal output
rlabel metal2 s 162306 179200 162362 180000 6 mprj_dat_o[15]
port 749 nsew signal output
rlabel metal2 s 162674 179200 162730 180000 6 mprj_dat_o[16]
port 750 nsew signal output
rlabel metal2 s 163042 179200 163098 180000 6 mprj_dat_o[17]
port 751 nsew signal output
rlabel metal2 s 163410 179200 163466 180000 6 mprj_dat_o[18]
port 752 nsew signal output
rlabel metal2 s 163778 179200 163834 180000 6 mprj_dat_o[19]
port 753 nsew signal output
rlabel metal2 s 164146 179200 164202 180000 6 mprj_dat_o[1]
port 754 nsew signal output
rlabel metal2 s 164514 179200 164570 180000 6 mprj_dat_o[20]
port 755 nsew signal output
rlabel metal2 s 164882 179200 164938 180000 6 mprj_dat_o[21]
port 756 nsew signal output
rlabel metal2 s 165250 179200 165306 180000 6 mprj_dat_o[22]
port 757 nsew signal output
rlabel metal2 s 165618 179200 165674 180000 6 mprj_dat_o[23]
port 758 nsew signal output
rlabel metal2 s 165986 179200 166042 180000 6 mprj_dat_o[24]
port 759 nsew signal output
rlabel metal2 s 166354 179200 166410 180000 6 mprj_dat_o[25]
port 760 nsew signal output
rlabel metal2 s 166722 179200 166778 180000 6 mprj_dat_o[26]
port 761 nsew signal output
rlabel metal2 s 167090 179200 167146 180000 6 mprj_dat_o[27]
port 762 nsew signal output
rlabel metal2 s 167458 179200 167514 180000 6 mprj_dat_o[28]
port 763 nsew signal output
rlabel metal2 s 167826 179200 167882 180000 6 mprj_dat_o[29]
port 764 nsew signal output
rlabel metal2 s 168194 179200 168250 180000 6 mprj_dat_o[2]
port 765 nsew signal output
rlabel metal2 s 168562 179200 168618 180000 6 mprj_dat_o[30]
port 766 nsew signal output
rlabel metal2 s 168930 179200 168986 180000 6 mprj_dat_o[31]
port 767 nsew signal output
rlabel metal2 s 169298 179200 169354 180000 6 mprj_dat_o[3]
port 768 nsew signal output
rlabel metal2 s 169666 179200 169722 180000 6 mprj_dat_o[4]
port 769 nsew signal output
rlabel metal2 s 170034 179200 170090 180000 6 mprj_dat_o[5]
port 770 nsew signal output
rlabel metal2 s 170402 179200 170458 180000 6 mprj_dat_o[6]
port 771 nsew signal output
rlabel metal2 s 170770 179200 170826 180000 6 mprj_dat_o[7]
port 772 nsew signal output
rlabel metal2 s 171138 179200 171194 180000 6 mprj_dat_o[8]
port 773 nsew signal output
rlabel metal2 s 171506 179200 171562 180000 6 mprj_dat_o[9]
port 774 nsew signal output
rlabel metal2 s 295154 179200 295210 180000 6 mprj_io_loader_clock
port 775 nsew signal output
rlabel metal3 s 429200 66376 430000 66496 6 mprj_io_loader_data
port 776 nsew signal output
rlabel metal2 s 299938 179200 299994 180000 6 mprj_io_loader_resetn
port 777 nsew signal output
rlabel metal2 s 171874 179200 171930 180000 6 mprj_sel_o[0]
port 778 nsew signal output
rlabel metal2 s 172242 179200 172298 180000 6 mprj_sel_o[1]
port 779 nsew signal output
rlabel metal2 s 172610 179200 172666 180000 6 mprj_sel_o[2]
port 780 nsew signal output
rlabel metal2 s 172978 179200 173034 180000 6 mprj_sel_o[3]
port 781 nsew signal output
rlabel metal2 s 173346 179200 173402 180000 6 mprj_stb_o
port 782 nsew signal output
rlabel metal2 s 173714 179200 173770 180000 6 mprj_vcc_pwrgood
port 783 nsew signal input
rlabel metal2 s 174082 179200 174138 180000 6 mprj_vdd_pwrgood
port 784 nsew signal input
rlabel metal2 s 174450 179200 174506 180000 6 mprj_we_o
port 785 nsew signal output
rlabel metal3 s 429200 50600 430000 50720 6 porb
port 786 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 pwr_ctrl_out[0]
port 787 nsew signal output
rlabel metal2 s 15106 0 15162 800 6 pwr_ctrl_out[1]
port 788 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 pwr_ctrl_out[2]
port 789 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 pwr_ctrl_out[3]
port 790 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 resetb
port 791 nsew signal input
rlabel metal3 s 429200 112072 430000 112192 6 sdo_out
port 792 nsew signal output
rlabel metal3 s 429200 113160 430000 113280 6 sdo_outenb
port 793 nsew signal output
rlabel metal2 s 174818 179200 174874 180000 6 user_clk
port 794 nsew signal output
rlabel metal4 s 424208 2128 424528 177392 6 VPWR
port 795 nsew power bidirectional
rlabel metal4 s 414208 2128 414528 177392 6 VPWR
port 796 nsew power bidirectional
rlabel metal4 s 404208 2128 404528 177392 6 VPWR
port 797 nsew power bidirectional
rlabel metal4 s 394208 2128 394528 177392 6 VPWR
port 798 nsew power bidirectional
rlabel metal4 s 384208 2128 384528 177392 6 VPWR
port 799 nsew power bidirectional
rlabel metal4 s 374208 44168 374528 177392 6 VPWR
port 800 nsew power bidirectional
rlabel metal4 s 364208 44168 364528 177392 6 VPWR
port 801 nsew power bidirectional
rlabel metal4 s 354208 44168 354528 177392 6 VPWR
port 802 nsew power bidirectional
rlabel metal4 s 344208 44168 344528 177392 6 VPWR
port 803 nsew power bidirectional
rlabel metal4 s 334208 2128 334528 177392 6 VPWR
port 804 nsew power bidirectional
rlabel metal4 s 324208 2128 324528 177392 6 VPWR
port 805 nsew power bidirectional
rlabel metal4 s 314208 2128 314528 177392 6 VPWR
port 806 nsew power bidirectional
rlabel metal4 s 304208 2128 304528 177392 6 VPWR
port 807 nsew power bidirectional
rlabel metal4 s 294208 2128 294528 177392 6 VPWR
port 808 nsew power bidirectional
rlabel metal4 s 284208 2128 284528 177392 6 VPWR
port 809 nsew power bidirectional
rlabel metal4 s 274208 2128 274528 177392 6 VPWR
port 810 nsew power bidirectional
rlabel metal4 s 264208 2128 264528 177392 6 VPWR
port 811 nsew power bidirectional
rlabel metal4 s 254208 2128 254528 177392 6 VPWR
port 812 nsew power bidirectional
rlabel metal4 s 244208 2128 244528 177392 6 VPWR
port 813 nsew power bidirectional
rlabel metal4 s 234208 2128 234528 177392 6 VPWR
port 814 nsew power bidirectional
rlabel metal4 s 224208 2128 224528 177392 6 VPWR
port 815 nsew power bidirectional
rlabel metal4 s 214208 2128 214528 177392 6 VPWR
port 816 nsew power bidirectional
rlabel metal4 s 204208 137232 204528 177392 6 VPWR
port 817 nsew power bidirectional
rlabel metal4 s 194208 137232 194528 177392 6 VPWR
port 818 nsew power bidirectional
rlabel metal4 s 184208 137232 184528 177392 6 VPWR
port 819 nsew power bidirectional
rlabel metal4 s 174208 137232 174528 177392 6 VPWR
port 820 nsew power bidirectional
rlabel metal4 s 164208 137232 164528 177392 6 VPWR
port 821 nsew power bidirectional
rlabel metal4 s 154208 137232 154528 177392 6 VPWR
port 822 nsew power bidirectional
rlabel metal4 s 144208 137232 144528 177392 6 VPWR
port 823 nsew power bidirectional
rlabel metal4 s 134208 137232 134528 177392 6 VPWR
port 824 nsew power bidirectional
rlabel metal4 s 124208 137232 124528 177392 6 VPWR
port 825 nsew power bidirectional
rlabel metal4 s 114208 137232 114528 177392 6 VPWR
port 826 nsew power bidirectional
rlabel metal4 s 104208 137232 104528 177392 6 VPWR
port 827 nsew power bidirectional
rlabel metal4 s 94208 137232 94528 177392 6 VPWR
port 828 nsew power bidirectional
rlabel metal4 s 84208 137232 84528 177392 6 VPWR
port 829 nsew power bidirectional
rlabel metal4 s 74208 137232 74528 177392 6 VPWR
port 830 nsew power bidirectional
rlabel metal4 s 64208 137232 64528 177392 6 VPWR
port 831 nsew power bidirectional
rlabel metal4 s 54208 2128 54528 177392 6 VPWR
port 832 nsew power bidirectional
rlabel metal4 s 44208 2128 44528 177392 6 VPWR
port 833 nsew power bidirectional
rlabel metal4 s 34208 2128 34528 177392 6 VPWR
port 834 nsew power bidirectional
rlabel metal4 s 24208 2128 24528 177392 6 VPWR
port 835 nsew power bidirectional
rlabel metal4 s 14208 2128 14528 177392 6 VPWR
port 836 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 177392 6 VPWR
port 837 nsew power bidirectional
rlabel metal4 s 204208 2128 204528 30328 6 VPWR
port 838 nsew power bidirectional
rlabel metal4 s 194208 2128 194528 30328 6 VPWR
port 839 nsew power bidirectional
rlabel metal4 s 184208 2128 184528 30328 6 VPWR
port 840 nsew power bidirectional
rlabel metal4 s 174208 2128 174528 30328 6 VPWR
port 841 nsew power bidirectional
rlabel metal4 s 164208 2128 164528 30328 6 VPWR
port 842 nsew power bidirectional
rlabel metal4 s 154208 2128 154528 30328 6 VPWR
port 843 nsew power bidirectional
rlabel metal4 s 144208 2128 144528 30328 6 VPWR
port 844 nsew power bidirectional
rlabel metal4 s 134208 2128 134528 30328 6 VPWR
port 845 nsew power bidirectional
rlabel metal4 s 124208 2128 124528 30328 6 VPWR
port 846 nsew power bidirectional
rlabel metal4 s 114208 2128 114528 30328 6 VPWR
port 847 nsew power bidirectional
rlabel metal4 s 104208 2128 104528 30328 6 VPWR
port 848 nsew power bidirectional
rlabel metal4 s 94208 2128 94528 30328 6 VPWR
port 849 nsew power bidirectional
rlabel metal4 s 84208 2128 84528 30328 6 VPWR
port 850 nsew power bidirectional
rlabel metal4 s 74208 2128 74528 30328 6 VPWR
port 851 nsew power bidirectional
rlabel metal4 s 64208 2128 64528 30328 6 VPWR
port 852 nsew power bidirectional
rlabel metal5 s 1104 158478 428812 158798 6 VPWR
port 853 nsew power bidirectional
rlabel metal5 s 1104 127842 428812 128162 6 VPWR
port 854 nsew power bidirectional
rlabel metal5 s 1104 97206 428812 97526 6 VPWR
port 855 nsew power bidirectional
rlabel metal5 s 1104 66570 428812 66890 6 VPWR
port 856 nsew power bidirectional
rlabel metal5 s 1104 35934 428812 36254 6 VPWR
port 857 nsew power bidirectional
rlabel metal5 s 1104 5298 428812 5618 6 VPWR
port 858 nsew power bidirectional
rlabel metal4 s 419208 2128 419528 177392 6 VGND
port 859 nsew ground bidirectional
rlabel metal4 s 409208 2128 409528 177392 6 VGND
port 860 nsew ground bidirectional
rlabel metal4 s 399208 2128 399528 177392 6 VGND
port 861 nsew ground bidirectional
rlabel metal4 s 389208 2128 389528 177392 6 VGND
port 862 nsew ground bidirectional
rlabel metal4 s 379208 44168 379528 177392 6 VGND
port 863 nsew ground bidirectional
rlabel metal4 s 369208 44168 369528 177392 6 VGND
port 864 nsew ground bidirectional
rlabel metal4 s 359208 44168 359528 177392 6 VGND
port 865 nsew ground bidirectional
rlabel metal4 s 349208 44168 349528 177392 6 VGND
port 866 nsew ground bidirectional
rlabel metal4 s 339208 44168 339528 177392 6 VGND
port 867 nsew ground bidirectional
rlabel metal4 s 329208 2128 329528 177392 6 VGND
port 868 nsew ground bidirectional
rlabel metal4 s 319208 2128 319528 177392 6 VGND
port 869 nsew ground bidirectional
rlabel metal4 s 309208 2128 309528 177392 6 VGND
port 870 nsew ground bidirectional
rlabel metal4 s 299208 2128 299528 177392 6 VGND
port 871 nsew ground bidirectional
rlabel metal4 s 289208 2128 289528 177392 6 VGND
port 872 nsew ground bidirectional
rlabel metal4 s 279208 2128 279528 177392 6 VGND
port 873 nsew ground bidirectional
rlabel metal4 s 269208 2128 269528 177392 6 VGND
port 874 nsew ground bidirectional
rlabel metal4 s 259208 2128 259528 177392 6 VGND
port 875 nsew ground bidirectional
rlabel metal4 s 249208 2128 249528 177392 6 VGND
port 876 nsew ground bidirectional
rlabel metal4 s 239208 2128 239528 177392 6 VGND
port 877 nsew ground bidirectional
rlabel metal4 s 229208 2128 229528 177392 6 VGND
port 878 nsew ground bidirectional
rlabel metal4 s 219208 2128 219528 177392 6 VGND
port 879 nsew ground bidirectional
rlabel metal4 s 209208 137232 209528 177392 6 VGND
port 880 nsew ground bidirectional
rlabel metal4 s 199208 137232 199528 177392 6 VGND
port 881 nsew ground bidirectional
rlabel metal4 s 189208 137232 189528 177392 6 VGND
port 882 nsew ground bidirectional
rlabel metal4 s 179208 137232 179528 177392 6 VGND
port 883 nsew ground bidirectional
rlabel metal4 s 169208 137232 169528 177392 6 VGND
port 884 nsew ground bidirectional
rlabel metal4 s 159208 137232 159528 177392 6 VGND
port 885 nsew ground bidirectional
rlabel metal4 s 149208 137232 149528 177392 6 VGND
port 886 nsew ground bidirectional
rlabel metal4 s 139208 137232 139528 177392 6 VGND
port 887 nsew ground bidirectional
rlabel metal4 s 129208 137232 129528 177392 6 VGND
port 888 nsew ground bidirectional
rlabel metal4 s 119208 137232 119528 177392 6 VGND
port 889 nsew ground bidirectional
rlabel metal4 s 109208 137232 109528 177392 6 VGND
port 890 nsew ground bidirectional
rlabel metal4 s 99208 137232 99528 177392 6 VGND
port 891 nsew ground bidirectional
rlabel metal4 s 89208 137232 89528 177392 6 VGND
port 892 nsew ground bidirectional
rlabel metal4 s 79208 137232 79528 177392 6 VGND
port 893 nsew ground bidirectional
rlabel metal4 s 69208 137232 69528 177392 6 VGND
port 894 nsew ground bidirectional
rlabel metal4 s 59208 2128 59528 177392 6 VGND
port 895 nsew ground bidirectional
rlabel metal4 s 49208 2128 49528 177392 6 VGND
port 896 nsew ground bidirectional
rlabel metal4 s 39208 2128 39528 177392 6 VGND
port 897 nsew ground bidirectional
rlabel metal4 s 29208 2128 29528 177392 6 VGND
port 898 nsew ground bidirectional
rlabel metal4 s 19208 2128 19528 177392 6 VGND
port 899 nsew ground bidirectional
rlabel metal4 s 9208 2128 9528 177392 6 VGND
port 900 nsew ground bidirectional
rlabel metal4 s 209208 2128 209528 30328 6 VGND
port 901 nsew ground bidirectional
rlabel metal4 s 199208 2128 199528 30328 6 VGND
port 902 nsew ground bidirectional
rlabel metal4 s 189208 2128 189528 30328 6 VGND
port 903 nsew ground bidirectional
rlabel metal4 s 179208 2128 179528 30328 6 VGND
port 904 nsew ground bidirectional
rlabel metal4 s 169208 2128 169528 30328 6 VGND
port 905 nsew ground bidirectional
rlabel metal4 s 159208 2128 159528 30328 6 VGND
port 906 nsew ground bidirectional
rlabel metal4 s 149208 2128 149528 30328 6 VGND
port 907 nsew ground bidirectional
rlabel metal4 s 139208 2128 139528 30328 6 VGND
port 908 nsew ground bidirectional
rlabel metal4 s 129208 2128 129528 30328 6 VGND
port 909 nsew ground bidirectional
rlabel metal4 s 119208 2128 119528 30328 6 VGND
port 910 nsew ground bidirectional
rlabel metal4 s 109208 2128 109528 30328 6 VGND
port 911 nsew ground bidirectional
rlabel metal4 s 99208 2128 99528 30328 6 VGND
port 912 nsew ground bidirectional
rlabel metal4 s 89208 2128 89528 30328 6 VGND
port 913 nsew ground bidirectional
rlabel metal4 s 79208 2128 79528 30328 6 VGND
port 914 nsew ground bidirectional
rlabel metal4 s 69208 2128 69528 30328 6 VGND
port 915 nsew ground bidirectional
rlabel metal5 s 1104 173796 428812 174116 6 VGND
port 916 nsew ground bidirectional
rlabel metal5 s 1104 143160 428812 143480 6 VGND
port 917 nsew ground bidirectional
rlabel metal5 s 1104 112524 428812 112844 6 VGND
port 918 nsew ground bidirectional
rlabel metal5 s 1104 81888 428812 82208 6 VGND
port 919 nsew ground bidirectional
rlabel metal5 s 1104 51252 428812 51572 6 VGND
port 920 nsew ground bidirectional
rlabel metal5 s 1104 20616 428812 20936 6 VGND
port 921 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 430000 180000
string LEFview TRUE
string GDS_FILE ../gds/mgmt_core.gds
string GDS_END 176095322
string GDS_START 49314066
<< end >>

