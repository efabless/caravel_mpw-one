VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mprj_logic_high
  CLASS BLOCK ;
  FOREIGN mprj_logic_high ;
  ORIGIN 0.000 0.000 ;
  SIZE 370.000 BY 25.000 ;
  PIN HI[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 5.000 ;
    END
  END HI[0]
  PIN HI[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 5.000 ;
    END
  END HI[100]
  PIN HI[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 5.000 ;
    END
  END HI[101]
  PIN HI[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 5.000 ;
    END
  END HI[102]
  PIN HI[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 5.000 ;
    END
  END HI[103]
  PIN HI[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 5.000 ;
    END
  END HI[104]
  PIN HI[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 5.000 ;
    END
  END HI[105]
  PIN HI[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 5.000 ;
    END
  END HI[106]
  PIN HI[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 5.000 ;
    END
  END HI[107]
  PIN HI[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 5.000 ;
    END
  END HI[108]
  PIN HI[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 5.000 ;
    END
  END HI[109]
  PIN HI[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 5.000 ;
    END
  END HI[10]
  PIN HI[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 5.000 ;
    END
  END HI[110]
  PIN HI[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 5.000 ;
    END
  END HI[111]
  PIN HI[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 5.000 ;
    END
  END HI[112]
  PIN HI[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 5.000 ;
    END
  END HI[113]
  PIN HI[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 5.000 ;
    END
  END HI[114]
  PIN HI[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 5.000 ;
    END
  END HI[115]
  PIN HI[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 5.000 ;
    END
  END HI[116]
  PIN HI[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 5.000 ;
    END
  END HI[117]
  PIN HI[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 5.000 ;
    END
  END HI[118]
  PIN HI[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 5.000 ;
    END
  END HI[119]
  PIN HI[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 5.000 ;
    END
  END HI[11]
  PIN HI[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 5.000 ;
    END
  END HI[120]
  PIN HI[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 5.000 ;
    END
  END HI[121]
  PIN HI[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 5.000 ;
    END
  END HI[122]
  PIN HI[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 5.000 ;
    END
  END HI[123]
  PIN HI[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 5.000 ;
    END
  END HI[124]
  PIN HI[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 5.000 ;
    END
  END HI[125]
  PIN HI[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 5.000 ;
    END
  END HI[126]
  PIN HI[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 5.000 ;
    END
  END HI[127]
  PIN HI[128]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 5.000 ;
    END
  END HI[128]
  PIN HI[129]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 5.000 ;
    END
  END HI[129]
  PIN HI[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 5.000 ;
    END
  END HI[12]
  PIN HI[130]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 5.000 ;
    END
  END HI[130]
  PIN HI[131]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 5.000 ;
    END
  END HI[131]
  PIN HI[132]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 5.000 ;
    END
  END HI[132]
  PIN HI[133]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 5.000 ;
    END
  END HI[133]
  PIN HI[134]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 5.000 ;
    END
  END HI[134]
  PIN HI[135]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 5.000 ;
    END
  END HI[135]
  PIN HI[136]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 5.000 ;
    END
  END HI[136]
  PIN HI[137]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 5.000 ;
    END
  END HI[137]
  PIN HI[138]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 5.000 ;
    END
  END HI[138]
  PIN HI[139]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 5.000 ;
    END
  END HI[139]
  PIN HI[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 5.000 ;
    END
  END HI[13]
  PIN HI[140]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 5.000 ;
    END
  END HI[140]
  PIN HI[141]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 5.000 ;
    END
  END HI[141]
  PIN HI[142]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 5.000 ;
    END
  END HI[142]
  PIN HI[143]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 5.000 ;
    END
  END HI[143]
  PIN HI[144]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 5.000 ;
    END
  END HI[144]
  PIN HI[145]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 5.000 ;
    END
  END HI[145]
  PIN HI[146]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 5.000 ;
    END
  END HI[146]
  PIN HI[147]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 5.000 ;
    END
  END HI[147]
  PIN HI[148]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 5.000 ;
    END
  END HI[148]
  PIN HI[149]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 5.000 ;
    END
  END HI[149]
  PIN HI[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 5.000 ;
    END
  END HI[14]
  PIN HI[150]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 5.000 ;
    END
  END HI[150]
  PIN HI[151]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 5.000 ;
    END
  END HI[151]
  PIN HI[152]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 5.000 ;
    END
  END HI[152]
  PIN HI[153]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 5.000 ;
    END
  END HI[153]
  PIN HI[154]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 5.000 ;
    END
  END HI[154]
  PIN HI[155]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 5.000 ;
    END
  END HI[155]
  PIN HI[156]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 5.000 ;
    END
  END HI[156]
  PIN HI[157]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 5.000 ;
    END
  END HI[157]
  PIN HI[158]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 5.000 ;
    END
  END HI[158]
  PIN HI[159]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 5.000 ;
    END
  END HI[159]
  PIN HI[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 5.000 ;
    END
  END HI[15]
  PIN HI[160]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 5.000 ;
    END
  END HI[160]
  PIN HI[161]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 5.000 ;
    END
  END HI[161]
  PIN HI[162]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 5.000 ;
    END
  END HI[162]
  PIN HI[163]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 5.000 ;
    END
  END HI[163]
  PIN HI[164]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 5.000 ;
    END
  END HI[164]
  PIN HI[165]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 5.000 ;
    END
  END HI[165]
  PIN HI[166]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 5.000 ;
    END
  END HI[166]
  PIN HI[167]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 5.000 ;
    END
  END HI[167]
  PIN HI[168]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 5.000 ;
    END
  END HI[168]
  PIN HI[169]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 5.000 ;
    END
  END HI[169]
  PIN HI[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 5.000 ;
    END
  END HI[16]
  PIN HI[170]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 5.000 ;
    END
  END HI[170]
  PIN HI[171]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 5.000 ;
    END
  END HI[171]
  PIN HI[172]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 5.000 ;
    END
  END HI[172]
  PIN HI[173]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 5.000 ;
    END
  END HI[173]
  PIN HI[174]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 5.000 ;
    END
  END HI[174]
  PIN HI[175]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 5.000 ;
    END
  END HI[175]
  PIN HI[176]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 5.000 ;
    END
  END HI[176]
  PIN HI[177]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 5.000 ;
    END
  END HI[177]
  PIN HI[178]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 5.000 ;
    END
  END HI[178]
  PIN HI[179]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 5.000 ;
    END
  END HI[179]
  PIN HI[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 5.000 ;
    END
  END HI[17]
  PIN HI[180]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 5.000 ;
    END
  END HI[180]
  PIN HI[181]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 5.000 ;
    END
  END HI[181]
  PIN HI[182]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 5.000 ;
    END
  END HI[182]
  PIN HI[183]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 5.000 ;
    END
  END HI[183]
  PIN HI[184]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 5.000 ;
    END
  END HI[184]
  PIN HI[185]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 5.000 ;
    END
  END HI[185]
  PIN HI[186]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 5.000 ;
    END
  END HI[186]
  PIN HI[187]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 5.000 ;
    END
  END HI[187]
  PIN HI[188]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 5.000 ;
    END
  END HI[188]
  PIN HI[189]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 5.000 ;
    END
  END HI[189]
  PIN HI[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 5.000 ;
    END
  END HI[18]
  PIN HI[190]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 5.000 ;
    END
  END HI[190]
  PIN HI[191]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 5.000 ;
    END
  END HI[191]
  PIN HI[192]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 5.000 ;
    END
  END HI[192]
  PIN HI[193]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 5.000 ;
    END
  END HI[193]
  PIN HI[194]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 5.000 ;
    END
  END HI[194]
  PIN HI[195]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 5.000 ;
    END
  END HI[195]
  PIN HI[196]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 5.000 ;
    END
  END HI[196]
  PIN HI[197]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 5.000 ;
    END
  END HI[197]
  PIN HI[198]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 5.000 ;
    END
  END HI[198]
  PIN HI[199]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 5.000 ;
    END
  END HI[199]
  PIN HI[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 5.000 ;
    END
  END HI[19]
  PIN HI[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 5.000 ;
    END
  END HI[1]
  PIN HI[200]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 5.000 ;
    END
  END HI[200]
  PIN HI[201]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 5.000 ;
    END
  END HI[201]
  PIN HI[202]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 5.000 ;
    END
  END HI[202]
  PIN HI[203]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 5.000 ;
    END
  END HI[203]
  PIN HI[204]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 20.000 152.170 25.000 ;
    END
  END HI[204]
  PIN HI[205]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 5.000 6.760 ;
    END
  END HI[205]
  PIN HI[206]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 5.000 8.800 ;
    END
  END HI[206]
  PIN HI[207]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 5.000 10.840 ;
    END
  END HI[207]
  PIN HI[208]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 5.000 12.880 ;
    END
  END HI[208]
  PIN HI[209]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 5.000 14.920 ;
    END
  END HI[209]
  PIN HI[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 5.000 16.960 ;
    END
  END HI[20]
  PIN HI[210]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 5.000 19.000 ;
    END
  END HI[210]
  PIN HI[211]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 20.000 3.130 25.000 ;
    END
  END HI[211]
  PIN HI[212]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 20.000 4.510 25.000 ;
    END
  END HI[212]
  PIN HI[213]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 20.000 5.890 25.000 ;
    END
  END HI[213]
  PIN HI[214]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 20.000 7.270 25.000 ;
    END
  END HI[214]
  PIN HI[215]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 20.000 8.650 25.000 ;
    END
  END HI[215]
  PIN HI[216]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 20.000 10.030 25.000 ;
    END
  END HI[216]
  PIN HI[217]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 20.000 11.410 25.000 ;
    END
  END HI[217]
  PIN HI[218]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 20.000 12.790 25.000 ;
    END
  END HI[218]
  PIN HI[219]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 20.000 14.170 25.000 ;
    END
  END HI[219]
  PIN HI[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 20.000 15.550 25.000 ;
    END
  END HI[21]
  PIN HI[220]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 20.000 16.930 25.000 ;
    END
  END HI[220]
  PIN HI[221]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 20.000 18.310 25.000 ;
    END
  END HI[221]
  PIN HI[222]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 20.000 19.690 25.000 ;
    END
  END HI[222]
  PIN HI[223]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 20.000 21.070 25.000 ;
    END
  END HI[223]
  PIN HI[224]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 20.000 22.450 25.000 ;
    END
  END HI[224]
  PIN HI[225]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 20.000 23.830 25.000 ;
    END
  END HI[225]
  PIN HI[226]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 20.000 25.210 25.000 ;
    END
  END HI[226]
  PIN HI[227]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 20.000 26.590 25.000 ;
    END
  END HI[227]
  PIN HI[228]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 20.000 27.970 25.000 ;
    END
  END HI[228]
  PIN HI[229]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 20.000 29.350 25.000 ;
    END
  END HI[229]
  PIN HI[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 20.000 30.730 25.000 ;
    END
  END HI[22]
  PIN HI[230]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 20.000 32.110 25.000 ;
    END
  END HI[230]
  PIN HI[231]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 20.000 33.490 25.000 ;
    END
  END HI[231]
  PIN HI[232]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 20.000 34.870 25.000 ;
    END
  END HI[232]
  PIN HI[233]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 20.000 36.250 25.000 ;
    END
  END HI[233]
  PIN HI[234]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 20.000 37.630 25.000 ;
    END
  END HI[234]
  PIN HI[235]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 20.000 39.010 25.000 ;
    END
  END HI[235]
  PIN HI[236]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 20.000 40.390 25.000 ;
    END
  END HI[236]
  PIN HI[237]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 20.000 41.770 25.000 ;
    END
  END HI[237]
  PIN HI[238]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 20.000 43.150 25.000 ;
    END
  END HI[238]
  PIN HI[239]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 20.000 44.530 25.000 ;
    END
  END HI[239]
  PIN HI[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 20.000 45.910 25.000 ;
    END
  END HI[23]
  PIN HI[240]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 20.000 47.290 25.000 ;
    END
  END HI[240]
  PIN HI[241]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 20.000 48.670 25.000 ;
    END
  END HI[241]
  PIN HI[242]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 20.000 50.050 25.000 ;
    END
  END HI[242]
  PIN HI[243]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 20.000 51.430 25.000 ;
    END
  END HI[243]
  PIN HI[244]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 20.000 52.810 25.000 ;
    END
  END HI[244]
  PIN HI[245]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 20.000 54.190 25.000 ;
    END
  END HI[245]
  PIN HI[246]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 20.000 55.570 25.000 ;
    END
  END HI[246]
  PIN HI[247]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 20.000 56.950 25.000 ;
    END
  END HI[247]
  PIN HI[248]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 20.000 58.330 25.000 ;
    END
  END HI[248]
  PIN HI[249]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 20.000 59.710 25.000 ;
    END
  END HI[249]
  PIN HI[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 20.000 61.090 25.000 ;
    END
  END HI[24]
  PIN HI[250]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 20.000 62.470 25.000 ;
    END
  END HI[250]
  PIN HI[251]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 20.000 63.850 25.000 ;
    END
  END HI[251]
  PIN HI[252]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 20.000 65.230 25.000 ;
    END
  END HI[252]
  PIN HI[253]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 20.000 66.610 25.000 ;
    END
  END HI[253]
  PIN HI[254]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 20.000 67.990 25.000 ;
    END
  END HI[254]
  PIN HI[255]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 20.000 69.370 25.000 ;
    END
  END HI[255]
  PIN HI[256]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 20.000 70.750 25.000 ;
    END
  END HI[256]
  PIN HI[257]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 20.000 72.130 25.000 ;
    END
  END HI[257]
  PIN HI[258]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 20.000 73.510 25.000 ;
    END
  END HI[258]
  PIN HI[259]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 20.000 74.890 25.000 ;
    END
  END HI[259]
  PIN HI[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 20.000 76.270 25.000 ;
    END
  END HI[25]
  PIN HI[260]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 20.000 77.650 25.000 ;
    END
  END HI[260]
  PIN HI[261]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 20.000 79.030 25.000 ;
    END
  END HI[261]
  PIN HI[262]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 20.000 80.410 25.000 ;
    END
  END HI[262]
  PIN HI[263]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 20.000 81.790 25.000 ;
    END
  END HI[263]
  PIN HI[264]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 20.000 83.170 25.000 ;
    END
  END HI[264]
  PIN HI[265]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 20.000 84.550 25.000 ;
    END
  END HI[265]
  PIN HI[266]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 20.000 85.930 25.000 ;
    END
  END HI[266]
  PIN HI[267]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 20.000 87.310 25.000 ;
    END
  END HI[267]
  PIN HI[268]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 20.000 88.690 25.000 ;
    END
  END HI[268]
  PIN HI[269]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 20.000 90.070 25.000 ;
    END
  END HI[269]
  PIN HI[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 20.000 91.450 25.000 ;
    END
  END HI[26]
  PIN HI[270]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 20.000 92.830 25.000 ;
    END
  END HI[270]
  PIN HI[271]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 20.000 94.210 25.000 ;
    END
  END HI[271]
  PIN HI[272]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 20.000 95.590 25.000 ;
    END
  END HI[272]
  PIN HI[273]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 20.000 96.970 25.000 ;
    END
  END HI[273]
  PIN HI[274]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 20.000 98.350 25.000 ;
    END
  END HI[274]
  PIN HI[275]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 20.000 99.730 25.000 ;
    END
  END HI[275]
  PIN HI[276]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 20.000 101.110 25.000 ;
    END
  END HI[276]
  PIN HI[277]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 20.000 102.490 25.000 ;
    END
  END HI[277]
  PIN HI[278]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 20.000 103.870 25.000 ;
    END
  END HI[278]
  PIN HI[279]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 20.000 105.250 25.000 ;
    END
  END HI[279]
  PIN HI[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 20.000 106.630 25.000 ;
    END
  END HI[27]
  PIN HI[280]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 20.000 108.010 25.000 ;
    END
  END HI[280]
  PIN HI[281]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 20.000 109.390 25.000 ;
    END
  END HI[281]
  PIN HI[282]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 20.000 110.770 25.000 ;
    END
  END HI[282]
  PIN HI[283]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 20.000 112.150 25.000 ;
    END
  END HI[283]
  PIN HI[284]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 20.000 113.530 25.000 ;
    END
  END HI[284]
  PIN HI[285]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 20.000 114.910 25.000 ;
    END
  END HI[285]
  PIN HI[286]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 20.000 116.290 25.000 ;
    END
  END HI[286]
  PIN HI[287]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 20.000 117.670 25.000 ;
    END
  END HI[287]
  PIN HI[288]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 20.000 119.050 25.000 ;
    END
  END HI[288]
  PIN HI[289]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 20.000 120.430 25.000 ;
    END
  END HI[289]
  PIN HI[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 20.000 121.810 25.000 ;
    END
  END HI[28]
  PIN HI[290]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 20.000 123.190 25.000 ;
    END
  END HI[290]
  PIN HI[291]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 20.000 124.570 25.000 ;
    END
  END HI[291]
  PIN HI[292]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 20.000 125.950 25.000 ;
    END
  END HI[292]
  PIN HI[293]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 20.000 127.330 25.000 ;
    END
  END HI[293]
  PIN HI[294]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 20.000 128.710 25.000 ;
    END
  END HI[294]
  PIN HI[295]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 20.000 130.090 25.000 ;
    END
  END HI[295]
  PIN HI[296]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 20.000 131.470 25.000 ;
    END
  END HI[296]
  PIN HI[297]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 20.000 132.850 25.000 ;
    END
  END HI[297]
  PIN HI[298]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 20.000 134.230 25.000 ;
    END
  END HI[298]
  PIN HI[299]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 20.000 135.610 25.000 ;
    END
  END HI[299]
  PIN HI[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 20.000 136.990 25.000 ;
    END
  END HI[29]
  PIN HI[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 20.000 138.370 25.000 ;
    END
  END HI[2]
  PIN HI[300]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 20.000 139.750 25.000 ;
    END
  END HI[300]
  PIN HI[301]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 20.000 141.130 25.000 ;
    END
  END HI[301]
  PIN HI[302]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 20.000 142.510 25.000 ;
    END
  END HI[302]
  PIN HI[303]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 20.000 143.890 25.000 ;
    END
  END HI[303]
  PIN HI[304]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 20.000 145.270 25.000 ;
    END
  END HI[304]
  PIN HI[305]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 20.000 146.650 25.000 ;
    END
  END HI[305]
  PIN HI[306]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 20.000 148.030 25.000 ;
    END
  END HI[306]
  PIN HI[307]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 20.000 149.410 25.000 ;
    END
  END HI[307]
  PIN HI[308]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 20.000 150.790 25.000 ;
    END
  END HI[308]
  PIN HI[309]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 0.000 349.510 5.000 ;
    END
  END HI[309]
  PIN HI[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 5.000 ;
    END
  END HI[30]
  PIN HI[310]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 5.000 ;
    END
  END HI[310]
  PIN HI[311]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 0.000 239.110 5.000 ;
    END
  END HI[311]
  PIN HI[312]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 5.000 ;
    END
  END HI[312]
  PIN HI[313]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 5.000 ;
    END
  END HI[313]
  PIN HI[314]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 5.000 ;
    END
  END HI[314]
  PIN HI[315]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 5.000 ;
    END
  END HI[315]
  PIN HI[316]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 0.000 346.750 5.000 ;
    END
  END HI[316]
  PIN HI[317]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 5.000 ;
    END
  END HI[317]
  PIN HI[318]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 5.000 ;
    END
  END HI[318]
  PIN HI[319]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 5.000 ;
    END
  END HI[319]
  PIN HI[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 5.000 ;
    END
  END HI[31]
  PIN HI[320]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 5.000 ;
    END
  END HI[320]
  PIN HI[321]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 5.000 ;
    END
  END HI[321]
  PIN HI[322]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 5.000 ;
    END
  END HI[322]
  PIN HI[323]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 5.000 ;
    END
  END HI[323]
  PIN HI[324]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 5.000 ;
    END
  END HI[324]
  PIN HI[325]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 5.000 ;
    END
  END HI[325]
  PIN HI[326]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 5.000 ;
    END
  END HI[326]
  PIN HI[327]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 5.000 ;
    END
  END HI[327]
  PIN HI[328]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 5.000 ;
    END
  END HI[328]
  PIN HI[329]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 0.000 324.670 5.000 ;
    END
  END HI[329]
  PIN HI[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 5.000 ;
    END
  END HI[32]
  PIN HI[330]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 5.000 ;
    END
  END HI[330]
  PIN HI[331]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 5.000 ;
    END
  END HI[331]
  PIN HI[332]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 5.000 ;
    END
  END HI[332]
  PIN HI[333]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 5.000 ;
    END
  END HI[333]
  PIN HI[334]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 5.000 ;
    END
  END HI[334]
  PIN HI[335]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 5.000 ;
    END
  END HI[335]
  PIN HI[336]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 5.000 ;
    END
  END HI[336]
  PIN HI[337]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 5.000 ;
    END
  END HI[337]
  PIN HI[338]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 5.000 ;
    END
  END HI[338]
  PIN HI[339]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 0.000 277.750 5.000 ;
    END
  END HI[339]
  PIN HI[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 5.000 ;
    END
  END HI[33]
  PIN HI[340]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 0.000 286.030 5.000 ;
    END
  END HI[340]
  PIN HI[341]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 5.000 ;
    END
  END HI[341]
  PIN HI[342]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 5.000 ;
    END
  END HI[342]
  PIN HI[343]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 5.000 ;
    END
  END HI[343]
  PIN HI[344]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 5.000 ;
    END
  END HI[344]
  PIN HI[345]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 5.000 ;
    END
  END HI[345]
  PIN HI[346]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 5.000 ;
    END
  END HI[346]
  PIN HI[347]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 5.000 ;
    END
  END HI[347]
  PIN HI[348]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 5.000 ;
    END
  END HI[348]
  PIN HI[349]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 0.000 294.310 5.000 ;
    END
  END HI[349]
  PIN HI[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 5.000 ;
    END
  END HI[34]
  PIN HI[350]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 5.000 ;
    END
  END HI[350]
  PIN HI[351]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 5.000 ;
    END
  END HI[351]
  PIN HI[352]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 5.000 ;
    END
  END HI[352]
  PIN HI[353]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 5.000 ;
    END
  END HI[353]
  PIN HI[354]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 5.000 ;
    END
  END HI[354]
  PIN HI[355]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 5.000 ;
    END
  END HI[355]
  PIN HI[356]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 5.000 ;
    END
  END HI[356]
  PIN HI[357]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 5.000 ;
    END
  END HI[357]
  PIN HI[358]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 5.000 ;
    END
  END HI[358]
  PIN HI[359]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 5.000 ;
    END
  END HI[359]
  PIN HI[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 5.000 ;
    END
  END HI[35]
  PIN HI[360]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 5.000 ;
    END
  END HI[360]
  PIN HI[361]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 5.000 ;
    END
  END HI[361]
  PIN HI[362]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 5.000 ;
    END
  END HI[362]
  PIN HI[363]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 5.000 ;
    END
  END HI[363]
  PIN HI[364]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 5.000 ;
    END
  END HI[364]
  PIN HI[365]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 5.000 ;
    END
  END HI[365]
  PIN HI[366]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 5.000 ;
    END
  END HI[366]
  PIN HI[367]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 5.000 ;
    END
  END HI[367]
  PIN HI[368]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 5.000 ;
    END
  END HI[368]
  PIN HI[369]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 5.000 ;
    END
  END HI[369]
  PIN HI[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 5.000 ;
    END
  END HI[36]
  PIN HI[370]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 5.000 ;
    END
  END HI[370]
  PIN HI[371]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 5.000 ;
    END
  END HI[371]
  PIN HI[372]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 5.000 ;
    END
  END HI[372]
  PIN HI[373]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 5.000 ;
    END
  END HI[373]
  PIN HI[374]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 5.000 ;
    END
  END HI[374]
  PIN HI[375]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 5.000 ;
    END
  END HI[375]
  PIN HI[376]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 5.000 ;
    END
  END HI[376]
  PIN HI[377]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 5.000 ;
    END
  END HI[377]
  PIN HI[378]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 5.000 ;
    END
  END HI[378]
  PIN HI[379]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 5.000 ;
    END
  END HI[379]
  PIN HI[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 5.000 ;
    END
  END HI[37]
  PIN HI[380]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 0.000 305.350 5.000 ;
    END
  END HI[380]
  PIN HI[381]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 5.000 ;
    END
  END HI[381]
  PIN HI[382]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 5.000 ;
    END
  END HI[382]
  PIN HI[383]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 5.000 ;
    END
  END HI[383]
  PIN HI[384]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 5.000 ;
    END
  END HI[384]
  PIN HI[385]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 5.000 ;
    END
  END HI[385]
  PIN HI[386]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 5.000 ;
    END
  END HI[386]
  PIN HI[387]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 5.000 ;
    END
  END HI[387]
  PIN HI[388]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 0.000 308.110 5.000 ;
    END
  END HI[388]
  PIN HI[389]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 5.000 ;
    END
  END HI[389]
  PIN HI[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 0.000 335.710 5.000 ;
    END
  END HI[38]
  PIN HI[390]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 5.000 ;
    END
  END HI[390]
  PIN HI[391]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 5.000 ;
    END
  END HI[391]
  PIN HI[392]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 5.000 ;
    END
  END HI[392]
  PIN HI[393]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 5.000 ;
    END
  END HI[393]
  PIN HI[394]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 5.000 ;
    END
  END HI[394]
  PIN HI[395]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 0.000 310.870 5.000 ;
    END
  END HI[395]
  PIN HI[396]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 5.000 ;
    END
  END HI[396]
  PIN HI[397]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 5.000 ;
    END
  END HI[397]
  PIN HI[398]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 5.000 ;
    END
  END HI[398]
  PIN HI[399]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 5.000 ;
    END
  END HI[399]
  PIN HI[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 5.000 ;
    END
  END HI[39]
  PIN HI[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 5.000 ;
    END
  END HI[3]
  PIN HI[400]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 5.000 ;
    END
  END HI[400]
  PIN HI[401]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 5.000 ;
    END
  END HI[401]
  PIN HI[402]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 5.000 ;
    END
  END HI[402]
  PIN HI[403]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 5.000 ;
    END
  END HI[403]
  PIN HI[404]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 5.000 ;
    END
  END HI[404]
  PIN HI[405]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 5.000 ;
    END
  END HI[405]
  PIN HI[406]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 5.000 ;
    END
  END HI[406]
  PIN HI[407]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 5.000 ;
    END
  END HI[407]
  PIN HI[408]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 5.000 ;
    END
  END HI[408]
  PIN HI[409]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 5.000 ;
    END
  END HI[409]
  PIN HI[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 5.000 ;
    END
  END HI[40]
  PIN HI[410]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 5.000 ;
    END
  END HI[410]
  PIN HI[411]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 0.000 252.910 5.000 ;
    END
  END HI[411]
  PIN HI[412]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 5.000 ;
    END
  END HI[412]
  PIN HI[413]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 20.000 337.090 25.000 ;
    END
  END HI[413]
  PIN HI[414]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 20.000 181.150 25.000 ;
    END
  END HI[414]
  PIN HI[415]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 20.000 182.530 25.000 ;
    END
  END HI[415]
  PIN HI[416]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 20.000 183.910 25.000 ;
    END
  END HI[416]
  PIN HI[417]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 20.000 185.290 25.000 ;
    END
  END HI[417]
  PIN HI[418]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 20.000 186.670 25.000 ;
    END
  END HI[418]
  PIN HI[419]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 20.000 188.050 25.000 ;
    END
  END HI[419]
  PIN HI[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 20.000 189.430 25.000 ;
    END
  END HI[41]
  PIN HI[420]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 20.000 190.810 25.000 ;
    END
  END HI[420]
  PIN HI[421]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 20.000 192.190 25.000 ;
    END
  END HI[421]
  PIN HI[422]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 20.000 193.570 25.000 ;
    END
  END HI[422]
  PIN HI[423]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 20.000 194.950 25.000 ;
    END
  END HI[423]
  PIN HI[424]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 20.000 196.330 25.000 ;
    END
  END HI[424]
  PIN HI[425]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 20.000 197.710 25.000 ;
    END
  END HI[425]
  PIN HI[426]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 20.000 199.090 25.000 ;
    END
  END HI[426]
  PIN HI[427]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 20.000 200.470 25.000 ;
    END
  END HI[427]
  PIN HI[428]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 20.000 201.850 25.000 ;
    END
  END HI[428]
  PIN HI[429]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 20.000 203.230 25.000 ;
    END
  END HI[429]
  PIN HI[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 20.000 204.610 25.000 ;
    END
  END HI[42]
  PIN HI[430]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 20.000 205.990 25.000 ;
    END
  END HI[430]
  PIN HI[431]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 20.000 207.370 25.000 ;
    END
  END HI[431]
  PIN HI[432]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 20.000 208.750 25.000 ;
    END
  END HI[432]
  PIN HI[433]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 20.000 210.130 25.000 ;
    END
  END HI[433]
  PIN HI[434]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 20.000 211.510 25.000 ;
    END
  END HI[434]
  PIN HI[435]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 20.000 212.890 25.000 ;
    END
  END HI[435]
  PIN HI[436]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 20.000 214.270 25.000 ;
    END
  END HI[436]
  PIN HI[437]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 20.000 215.650 25.000 ;
    END
  END HI[437]
  PIN HI[438]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 20.000 217.030 25.000 ;
    END
  END HI[438]
  PIN HI[439]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 20.000 218.410 25.000 ;
    END
  END HI[439]
  PIN HI[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 20.000 219.790 25.000 ;
    END
  END HI[43]
  PIN HI[440]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 20.000 221.170 25.000 ;
    END
  END HI[440]
  PIN HI[441]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 20.000 222.550 25.000 ;
    END
  END HI[441]
  PIN HI[442]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 20.000 223.930 25.000 ;
    END
  END HI[442]
  PIN HI[443]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 20.000 225.310 25.000 ;
    END
  END HI[443]
  PIN HI[444]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 20.000 226.690 25.000 ;
    END
  END HI[444]
  PIN HI[445]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 20.000 228.070 25.000 ;
    END
  END HI[445]
  PIN HI[446]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 20.000 229.450 25.000 ;
    END
  END HI[446]
  PIN HI[447]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 20.000 230.830 25.000 ;
    END
  END HI[447]
  PIN HI[448]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 20.000 232.210 25.000 ;
    END
  END HI[448]
  PIN HI[449]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 20.000 233.590 25.000 ;
    END
  END HI[449]
  PIN HI[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 20.000 234.970 25.000 ;
    END
  END HI[44]
  PIN HI[450]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 20.000 236.350 25.000 ;
    END
  END HI[450]
  PIN HI[451]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 20.000 237.730 25.000 ;
    END
  END HI[451]
  PIN HI[452]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 20.000 239.110 25.000 ;
    END
  END HI[452]
  PIN HI[453]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 20.000 240.490 25.000 ;
    END
  END HI[453]
  PIN HI[454]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 20.000 241.870 25.000 ;
    END
  END HI[454]
  PIN HI[455]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 20.000 243.250 25.000 ;
    END
  END HI[455]
  PIN HI[456]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 20.000 244.630 25.000 ;
    END
  END HI[456]
  PIN HI[457]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 20.000 246.010 25.000 ;
    END
  END HI[457]
  PIN HI[458]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 20.000 247.390 25.000 ;
    END
  END HI[458]
  PIN HI[459]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 20.000 248.770 25.000 ;
    END
  END HI[459]
  PIN HI[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 20.000 250.150 25.000 ;
    END
  END HI[45]
  PIN HI[460]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 20.000 251.530 25.000 ;
    END
  END HI[460]
  PIN HI[461]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 20.000 252.910 25.000 ;
    END
  END HI[461]
  PIN HI[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 20.000 254.290 25.000 ;
    END
  END HI[46]
  PIN HI[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 20.000 255.670 25.000 ;
    END
  END HI[47]
  PIN HI[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 20.000 257.050 25.000 ;
    END
  END HI[48]
  PIN HI[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 20.000 258.430 25.000 ;
    END
  END HI[49]
  PIN HI[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 20.000 259.810 25.000 ;
    END
  END HI[4]
  PIN HI[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 20.000 261.190 25.000 ;
    END
  END HI[50]
  PIN HI[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 20.000 262.570 25.000 ;
    END
  END HI[51]
  PIN HI[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 20.000 263.950 25.000 ;
    END
  END HI[52]
  PIN HI[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 20.000 265.330 25.000 ;
    END
  END HI[53]
  PIN HI[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 20.000 266.710 25.000 ;
    END
  END HI[54]
  PIN HI[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 20.000 268.090 25.000 ;
    END
  END HI[55]
  PIN HI[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 20.000 269.470 25.000 ;
    END
  END HI[56]
  PIN HI[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 20.000 270.850 25.000 ;
    END
  END HI[57]
  PIN HI[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 20.000 272.230 25.000 ;
    END
  END HI[58]
  PIN HI[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 20.000 273.610 25.000 ;
    END
  END HI[59]
  PIN HI[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 20.000 274.990 25.000 ;
    END
  END HI[5]
  PIN HI[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 20.000 276.370 25.000 ;
    END
  END HI[60]
  PIN HI[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 20.000 277.750 25.000 ;
    END
  END HI[61]
  PIN HI[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 20.000 279.130 25.000 ;
    END
  END HI[62]
  PIN HI[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 20.000 280.510 25.000 ;
    END
  END HI[63]
  PIN HI[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 20.000 281.890 25.000 ;
    END
  END HI[64]
  PIN HI[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 20.000 283.270 25.000 ;
    END
  END HI[65]
  PIN HI[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 20.000 284.650 25.000 ;
    END
  END HI[66]
  PIN HI[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 20.000 286.030 25.000 ;
    END
  END HI[67]
  PIN HI[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 20.000 287.410 25.000 ;
    END
  END HI[68]
  PIN HI[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 20.000 288.790 25.000 ;
    END
  END HI[69]
  PIN HI[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 20.000 290.170 25.000 ;
    END
  END HI[6]
  PIN HI[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 20.000 291.550 25.000 ;
    END
  END HI[70]
  PIN HI[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 20.000 292.930 25.000 ;
    END
  END HI[71]
  PIN HI[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 20.000 294.310 25.000 ;
    END
  END HI[72]
  PIN HI[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 20.000 295.690 25.000 ;
    END
  END HI[73]
  PIN HI[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 20.000 297.070 25.000 ;
    END
  END HI[74]
  PIN HI[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 20.000 298.450 25.000 ;
    END
  END HI[75]
  PIN HI[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 20.000 299.830 25.000 ;
    END
  END HI[76]
  PIN HI[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 20.000 301.210 25.000 ;
    END
  END HI[77]
  PIN HI[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 20.000 302.590 25.000 ;
    END
  END HI[78]
  PIN HI[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 20.000 303.970 25.000 ;
    END
  END HI[79]
  PIN HI[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 20.000 305.350 25.000 ;
    END
  END HI[7]
  PIN HI[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 20.000 306.730 25.000 ;
    END
  END HI[80]
  PIN HI[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 20.000 308.110 25.000 ;
    END
  END HI[81]
  PIN HI[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 20.000 309.490 25.000 ;
    END
  END HI[82]
  PIN HI[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 20.000 310.870 25.000 ;
    END
  END HI[83]
  PIN HI[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 20.000 312.250 25.000 ;
    END
  END HI[84]
  PIN HI[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 20.000 313.630 25.000 ;
    END
  END HI[85]
  PIN HI[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 20.000 315.010 25.000 ;
    END
  END HI[86]
  PIN HI[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 20.000 316.390 25.000 ;
    END
  END HI[87]
  PIN HI[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 20.000 317.770 25.000 ;
    END
  END HI[88]
  PIN HI[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 20.000 319.150 25.000 ;
    END
  END HI[89]
  PIN HI[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 20.000 320.530 25.000 ;
    END
  END HI[8]
  PIN HI[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 20.000 321.910 25.000 ;
    END
  END HI[90]
  PIN HI[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 20.000 323.290 25.000 ;
    END
  END HI[91]
  PIN HI[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 20.000 324.670 25.000 ;
    END
  END HI[92]
  PIN HI[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 20.000 326.050 25.000 ;
    END
  END HI[93]
  PIN HI[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 20.000 327.430 25.000 ;
    END
  END HI[94]
  PIN HI[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 20.000 328.810 25.000 ;
    END
  END HI[95]
  PIN HI[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 20.000 330.190 25.000 ;
    END
  END HI[96]
  PIN HI[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 20.000 331.570 25.000 ;
    END
  END HI[97]
  PIN HI[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 20.000 332.950 25.000 ;
    END
  END HI[98]
  PIN HI[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 20.000 334.330 25.000 ;
    END
  END HI[99]
  PIN HI[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 20.000 335.710 25.000 ;
    END
  END HI[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 315.270 5.200 315.770 19.280 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 255.270 5.200 255.770 19.280 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 195.270 5.200 195.770 19.280 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 135.270 5.200 135.770 19.280 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 75.270 5.200 75.770 19.280 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 15.270 5.200 15.770 19.280 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 5.520 16.750 364.320 17.250 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 5.520 5.950 364.320 6.450 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 345.270 5.200 345.770 19.280 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 285.270 5.200 285.770 19.280 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 225.270 5.200 225.770 19.280 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 165.270 5.200 165.770 19.280 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 105.270 5.200 105.770 19.280 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 45.270 5.200 45.770 19.280 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 5.520 11.350 364.320 11.850 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 364.320 19.125 ;
      LAYER met1 ;
        RECT 2.830 5.200 364.320 20.020 ;
      LAYER met2 ;
        RECT 3.410 19.720 3.950 20.050 ;
        RECT 4.790 19.720 5.330 20.050 ;
        RECT 6.170 19.720 6.710 20.050 ;
        RECT 7.550 19.720 8.090 20.050 ;
        RECT 8.930 19.720 9.470 20.050 ;
        RECT 10.310 19.720 10.850 20.050 ;
        RECT 11.690 19.720 12.230 20.050 ;
        RECT 13.070 19.720 13.610 20.050 ;
        RECT 14.450 19.720 14.990 20.050 ;
        RECT 15.830 19.720 16.370 20.050 ;
        RECT 17.210 19.720 17.750 20.050 ;
        RECT 18.590 19.720 19.130 20.050 ;
        RECT 19.970 19.720 20.510 20.050 ;
        RECT 21.350 19.720 21.890 20.050 ;
        RECT 22.730 19.720 23.270 20.050 ;
        RECT 24.110 19.720 24.650 20.050 ;
        RECT 25.490 19.720 26.030 20.050 ;
        RECT 26.870 19.720 27.410 20.050 ;
        RECT 28.250 19.720 28.790 20.050 ;
        RECT 29.630 19.720 30.170 20.050 ;
        RECT 31.010 19.720 31.550 20.050 ;
        RECT 32.390 19.720 32.930 20.050 ;
        RECT 33.770 19.720 34.310 20.050 ;
        RECT 35.150 19.720 35.690 20.050 ;
        RECT 36.530 19.720 37.070 20.050 ;
        RECT 37.910 19.720 38.450 20.050 ;
        RECT 39.290 19.720 39.830 20.050 ;
        RECT 40.670 19.720 41.210 20.050 ;
        RECT 42.050 19.720 42.590 20.050 ;
        RECT 43.430 19.720 43.970 20.050 ;
        RECT 44.810 19.720 45.350 20.050 ;
        RECT 46.190 19.720 46.730 20.050 ;
        RECT 47.570 19.720 48.110 20.050 ;
        RECT 48.950 19.720 49.490 20.050 ;
        RECT 50.330 19.720 50.870 20.050 ;
        RECT 51.710 19.720 52.250 20.050 ;
        RECT 53.090 19.720 53.630 20.050 ;
        RECT 54.470 19.720 55.010 20.050 ;
        RECT 55.850 19.720 56.390 20.050 ;
        RECT 57.230 19.720 57.770 20.050 ;
        RECT 58.610 19.720 59.150 20.050 ;
        RECT 59.990 19.720 60.530 20.050 ;
        RECT 61.370 19.720 61.910 20.050 ;
        RECT 62.750 19.720 63.290 20.050 ;
        RECT 64.130 19.720 64.670 20.050 ;
        RECT 65.510 19.720 66.050 20.050 ;
        RECT 66.890 19.720 67.430 20.050 ;
        RECT 68.270 19.720 68.810 20.050 ;
        RECT 69.650 19.720 70.190 20.050 ;
        RECT 71.030 19.720 71.570 20.050 ;
        RECT 72.410 19.720 72.950 20.050 ;
        RECT 73.790 19.720 74.330 20.050 ;
        RECT 75.170 19.720 75.710 20.050 ;
        RECT 76.550 19.720 77.090 20.050 ;
        RECT 77.930 19.720 78.470 20.050 ;
        RECT 79.310 19.720 79.850 20.050 ;
        RECT 80.690 19.720 81.230 20.050 ;
        RECT 82.070 19.720 82.610 20.050 ;
        RECT 83.450 19.720 83.990 20.050 ;
        RECT 84.830 19.720 85.370 20.050 ;
        RECT 86.210 19.720 86.750 20.050 ;
        RECT 87.590 19.720 88.130 20.050 ;
        RECT 88.970 19.720 89.510 20.050 ;
        RECT 90.350 19.720 90.890 20.050 ;
        RECT 91.730 19.720 92.270 20.050 ;
        RECT 93.110 19.720 93.650 20.050 ;
        RECT 94.490 19.720 95.030 20.050 ;
        RECT 95.870 19.720 96.410 20.050 ;
        RECT 97.250 19.720 97.790 20.050 ;
        RECT 98.630 19.720 99.170 20.050 ;
        RECT 100.010 19.720 100.550 20.050 ;
        RECT 101.390 19.720 101.930 20.050 ;
        RECT 102.770 19.720 103.310 20.050 ;
        RECT 104.150 19.720 104.690 20.050 ;
        RECT 105.530 19.720 106.070 20.050 ;
        RECT 106.910 19.720 107.450 20.050 ;
        RECT 108.290 19.720 108.830 20.050 ;
        RECT 109.670 19.720 110.210 20.050 ;
        RECT 111.050 19.720 111.590 20.050 ;
        RECT 112.430 19.720 112.970 20.050 ;
        RECT 113.810 19.720 114.350 20.050 ;
        RECT 115.190 19.720 115.730 20.050 ;
        RECT 116.570 19.720 117.110 20.050 ;
        RECT 117.950 19.720 118.490 20.050 ;
        RECT 119.330 19.720 119.870 20.050 ;
        RECT 120.710 19.720 121.250 20.050 ;
        RECT 122.090 19.720 122.630 20.050 ;
        RECT 123.470 19.720 124.010 20.050 ;
        RECT 124.850 19.720 125.390 20.050 ;
        RECT 126.230 19.720 126.770 20.050 ;
        RECT 127.610 19.720 128.150 20.050 ;
        RECT 128.990 19.720 129.530 20.050 ;
        RECT 130.370 19.720 130.910 20.050 ;
        RECT 131.750 19.720 132.290 20.050 ;
        RECT 133.130 19.720 133.670 20.050 ;
        RECT 134.510 19.720 135.050 20.050 ;
        RECT 135.890 19.720 136.430 20.050 ;
        RECT 137.270 19.720 137.810 20.050 ;
        RECT 138.650 19.720 139.190 20.050 ;
        RECT 140.030 19.720 140.570 20.050 ;
        RECT 141.410 19.720 141.950 20.050 ;
        RECT 142.790 19.720 143.330 20.050 ;
        RECT 144.170 19.720 144.710 20.050 ;
        RECT 145.550 19.720 146.090 20.050 ;
        RECT 146.930 19.720 147.470 20.050 ;
        RECT 148.310 19.720 148.850 20.050 ;
        RECT 149.690 19.720 150.230 20.050 ;
        RECT 151.070 19.720 151.610 20.050 ;
        RECT 152.450 19.720 180.590 20.050 ;
        RECT 181.430 19.720 181.970 20.050 ;
        RECT 182.810 19.720 183.350 20.050 ;
        RECT 184.190 19.720 184.730 20.050 ;
        RECT 185.570 19.720 186.110 20.050 ;
        RECT 186.950 19.720 187.490 20.050 ;
        RECT 188.330 19.720 188.870 20.050 ;
        RECT 189.710 19.720 190.250 20.050 ;
        RECT 191.090 19.720 191.630 20.050 ;
        RECT 192.470 19.720 193.010 20.050 ;
        RECT 193.850 19.720 194.390 20.050 ;
        RECT 195.230 19.720 195.770 20.050 ;
        RECT 196.610 19.720 197.150 20.050 ;
        RECT 197.990 19.720 198.530 20.050 ;
        RECT 199.370 19.720 199.910 20.050 ;
        RECT 200.750 19.720 201.290 20.050 ;
        RECT 202.130 19.720 202.670 20.050 ;
        RECT 203.510 19.720 204.050 20.050 ;
        RECT 204.890 19.720 205.430 20.050 ;
        RECT 206.270 19.720 206.810 20.050 ;
        RECT 207.650 19.720 208.190 20.050 ;
        RECT 209.030 19.720 209.570 20.050 ;
        RECT 210.410 19.720 210.950 20.050 ;
        RECT 211.790 19.720 212.330 20.050 ;
        RECT 213.170 19.720 213.710 20.050 ;
        RECT 214.550 19.720 215.090 20.050 ;
        RECT 215.930 19.720 216.470 20.050 ;
        RECT 217.310 19.720 217.850 20.050 ;
        RECT 218.690 19.720 219.230 20.050 ;
        RECT 220.070 19.720 220.610 20.050 ;
        RECT 221.450 19.720 221.990 20.050 ;
        RECT 222.830 19.720 223.370 20.050 ;
        RECT 224.210 19.720 224.750 20.050 ;
        RECT 225.590 19.720 226.130 20.050 ;
        RECT 226.970 19.720 227.510 20.050 ;
        RECT 228.350 19.720 228.890 20.050 ;
        RECT 229.730 19.720 230.270 20.050 ;
        RECT 231.110 19.720 231.650 20.050 ;
        RECT 232.490 19.720 233.030 20.050 ;
        RECT 233.870 19.720 234.410 20.050 ;
        RECT 235.250 19.720 235.790 20.050 ;
        RECT 236.630 19.720 237.170 20.050 ;
        RECT 238.010 19.720 238.550 20.050 ;
        RECT 239.390 19.720 239.930 20.050 ;
        RECT 240.770 19.720 241.310 20.050 ;
        RECT 242.150 19.720 242.690 20.050 ;
        RECT 243.530 19.720 244.070 20.050 ;
        RECT 244.910 19.720 245.450 20.050 ;
        RECT 246.290 19.720 246.830 20.050 ;
        RECT 247.670 19.720 248.210 20.050 ;
        RECT 249.050 19.720 249.590 20.050 ;
        RECT 250.430 19.720 250.970 20.050 ;
        RECT 251.810 19.720 252.350 20.050 ;
        RECT 253.190 19.720 253.730 20.050 ;
        RECT 254.570 19.720 255.110 20.050 ;
        RECT 255.950 19.720 256.490 20.050 ;
        RECT 257.330 19.720 257.870 20.050 ;
        RECT 258.710 19.720 259.250 20.050 ;
        RECT 260.090 19.720 260.630 20.050 ;
        RECT 261.470 19.720 262.010 20.050 ;
        RECT 262.850 19.720 263.390 20.050 ;
        RECT 264.230 19.720 264.770 20.050 ;
        RECT 265.610 19.720 266.150 20.050 ;
        RECT 266.990 19.720 267.530 20.050 ;
        RECT 268.370 19.720 268.910 20.050 ;
        RECT 269.750 19.720 270.290 20.050 ;
        RECT 271.130 19.720 271.670 20.050 ;
        RECT 272.510 19.720 273.050 20.050 ;
        RECT 273.890 19.720 274.430 20.050 ;
        RECT 275.270 19.720 275.810 20.050 ;
        RECT 276.650 19.720 277.190 20.050 ;
        RECT 278.030 19.720 278.570 20.050 ;
        RECT 279.410 19.720 279.950 20.050 ;
        RECT 280.790 19.720 281.330 20.050 ;
        RECT 282.170 19.720 282.710 20.050 ;
        RECT 283.550 19.720 284.090 20.050 ;
        RECT 284.930 19.720 285.470 20.050 ;
        RECT 286.310 19.720 286.850 20.050 ;
        RECT 287.690 19.720 288.230 20.050 ;
        RECT 289.070 19.720 289.610 20.050 ;
        RECT 290.450 19.720 290.990 20.050 ;
        RECT 291.830 19.720 292.370 20.050 ;
        RECT 293.210 19.720 293.750 20.050 ;
        RECT 294.590 19.720 295.130 20.050 ;
        RECT 295.970 19.720 296.510 20.050 ;
        RECT 297.350 19.720 297.890 20.050 ;
        RECT 298.730 19.720 299.270 20.050 ;
        RECT 300.110 19.720 300.650 20.050 ;
        RECT 301.490 19.720 302.030 20.050 ;
        RECT 302.870 19.720 303.410 20.050 ;
        RECT 304.250 19.720 304.790 20.050 ;
        RECT 305.630 19.720 306.170 20.050 ;
        RECT 307.010 19.720 307.550 20.050 ;
        RECT 308.390 19.720 308.930 20.050 ;
        RECT 309.770 19.720 310.310 20.050 ;
        RECT 311.150 19.720 311.690 20.050 ;
        RECT 312.530 19.720 313.070 20.050 ;
        RECT 313.910 19.720 314.450 20.050 ;
        RECT 315.290 19.720 315.830 20.050 ;
        RECT 316.670 19.720 317.210 20.050 ;
        RECT 318.050 19.720 318.590 20.050 ;
        RECT 319.430 19.720 319.970 20.050 ;
        RECT 320.810 19.720 321.350 20.050 ;
        RECT 322.190 19.720 322.730 20.050 ;
        RECT 323.570 19.720 324.110 20.050 ;
        RECT 324.950 19.720 325.490 20.050 ;
        RECT 326.330 19.720 326.870 20.050 ;
        RECT 327.710 19.720 328.250 20.050 ;
        RECT 329.090 19.720 329.630 20.050 ;
        RECT 330.470 19.720 331.010 20.050 ;
        RECT 331.850 19.720 332.390 20.050 ;
        RECT 333.230 19.720 333.770 20.050 ;
        RECT 334.610 19.720 335.150 20.050 ;
        RECT 335.990 19.720 336.530 20.050 ;
        RECT 337.370 19.720 349.500 20.050 ;
        RECT 2.860 19.560 349.500 19.720 ;
        RECT 2.860 5.280 14.990 19.560 ;
        RECT 3.410 4.350 3.950 5.280 ;
        RECT 4.790 4.350 5.330 5.280 ;
        RECT 6.170 4.350 6.710 5.280 ;
        RECT 7.550 4.350 8.090 5.280 ;
        RECT 8.930 4.350 9.470 5.280 ;
        RECT 10.310 4.350 10.850 5.280 ;
        RECT 11.690 4.350 12.230 5.280 ;
        RECT 13.070 4.350 13.610 5.280 ;
        RECT 14.450 4.350 14.990 5.280 ;
        RECT 16.050 5.280 44.990 19.560 ;
        RECT 46.050 5.280 74.990 19.560 ;
        RECT 76.050 5.280 104.990 19.560 ;
        RECT 106.050 5.280 134.990 19.560 ;
        RECT 16.050 4.920 16.370 5.280 ;
        RECT 15.830 4.350 16.370 4.920 ;
        RECT 17.210 4.350 17.750 5.280 ;
        RECT 18.590 4.350 19.130 5.280 ;
        RECT 19.970 4.350 20.510 5.280 ;
        RECT 21.350 4.350 21.890 5.280 ;
        RECT 22.730 4.350 23.270 5.280 ;
        RECT 24.110 4.350 24.650 5.280 ;
        RECT 25.490 4.350 26.030 5.280 ;
        RECT 26.870 4.350 27.410 5.280 ;
        RECT 28.250 4.350 28.790 5.280 ;
        RECT 29.630 4.350 30.170 5.280 ;
        RECT 31.010 4.350 31.550 5.280 ;
        RECT 32.390 4.350 32.930 5.280 ;
        RECT 33.770 4.350 34.310 5.280 ;
        RECT 35.150 4.350 35.690 5.280 ;
        RECT 36.530 4.350 37.070 5.280 ;
        RECT 37.910 4.350 38.450 5.280 ;
        RECT 39.290 4.350 39.830 5.280 ;
        RECT 40.670 4.350 41.210 5.280 ;
        RECT 42.050 4.350 42.590 5.280 ;
        RECT 43.430 4.350 43.970 5.280 ;
        RECT 44.810 4.920 44.990 5.280 ;
        RECT 44.810 4.350 45.350 4.920 ;
        RECT 46.190 4.350 46.730 5.280 ;
        RECT 47.570 4.350 48.110 5.280 ;
        RECT 48.950 4.350 49.490 5.280 ;
        RECT 50.330 4.350 50.870 5.280 ;
        RECT 51.710 4.350 52.250 5.280 ;
        RECT 53.090 4.350 53.630 5.280 ;
        RECT 54.470 4.350 55.010 5.280 ;
        RECT 55.850 4.350 56.390 5.280 ;
        RECT 57.230 4.350 57.770 5.280 ;
        RECT 58.610 4.350 59.150 5.280 ;
        RECT 59.990 4.350 60.530 5.280 ;
        RECT 61.370 4.350 61.910 5.280 ;
        RECT 62.750 4.350 63.290 5.280 ;
        RECT 64.130 4.350 64.670 5.280 ;
        RECT 65.510 4.350 66.050 5.280 ;
        RECT 66.890 4.350 67.430 5.280 ;
        RECT 68.270 4.350 68.810 5.280 ;
        RECT 69.650 4.350 70.190 5.280 ;
        RECT 71.030 4.350 71.570 5.280 ;
        RECT 72.410 4.350 72.950 5.280 ;
        RECT 73.790 4.350 74.330 5.280 ;
        RECT 75.170 4.350 75.710 4.920 ;
        RECT 76.550 4.350 77.090 5.280 ;
        RECT 77.930 4.350 78.470 5.280 ;
        RECT 79.310 4.350 79.850 5.280 ;
        RECT 80.690 4.350 81.230 5.280 ;
        RECT 82.070 4.350 82.610 5.280 ;
        RECT 83.450 4.350 83.990 5.280 ;
        RECT 84.830 4.350 85.370 5.280 ;
        RECT 86.210 4.350 86.750 5.280 ;
        RECT 87.590 4.350 88.130 5.280 ;
        RECT 88.970 4.350 89.510 5.280 ;
        RECT 90.350 4.350 90.890 5.280 ;
        RECT 91.730 4.350 92.270 5.280 ;
        RECT 93.110 4.350 93.650 5.280 ;
        RECT 94.490 4.350 95.030 5.280 ;
        RECT 95.870 4.350 96.410 5.280 ;
        RECT 97.250 4.350 97.790 5.280 ;
        RECT 98.630 4.350 99.170 5.280 ;
        RECT 100.010 4.350 100.550 5.280 ;
        RECT 101.390 4.350 101.930 5.280 ;
        RECT 102.770 4.350 103.310 5.280 ;
        RECT 104.150 4.350 104.690 5.280 ;
        RECT 106.050 4.920 106.070 5.280 ;
        RECT 105.530 4.350 106.070 4.920 ;
        RECT 106.910 4.350 107.450 5.280 ;
        RECT 108.290 4.350 108.830 5.280 ;
        RECT 109.670 4.350 110.210 5.280 ;
        RECT 111.050 4.350 111.590 5.280 ;
        RECT 112.430 4.350 112.970 5.280 ;
        RECT 113.810 4.350 114.350 5.280 ;
        RECT 115.190 4.350 115.730 5.280 ;
        RECT 116.570 4.350 117.110 5.280 ;
        RECT 117.950 4.350 118.490 5.280 ;
        RECT 119.330 4.350 119.870 5.280 ;
        RECT 120.710 4.350 121.250 5.280 ;
        RECT 122.090 4.350 122.630 5.280 ;
        RECT 123.470 4.350 124.010 5.280 ;
        RECT 124.850 4.350 125.390 5.280 ;
        RECT 126.230 4.350 126.770 5.280 ;
        RECT 127.610 4.350 128.150 5.280 ;
        RECT 128.990 4.350 129.530 5.280 ;
        RECT 130.370 4.350 130.910 5.280 ;
        RECT 131.750 4.350 132.290 5.280 ;
        RECT 133.130 4.350 133.670 5.280 ;
        RECT 134.510 4.920 134.990 5.280 ;
        RECT 136.050 5.280 164.990 19.560 ;
        RECT 136.050 4.920 136.430 5.280 ;
        RECT 134.510 4.350 135.050 4.920 ;
        RECT 135.890 4.350 136.430 4.920 ;
        RECT 137.270 4.350 137.810 5.280 ;
        RECT 138.650 4.350 139.190 5.280 ;
        RECT 140.030 4.350 140.570 5.280 ;
        RECT 141.410 4.350 141.950 5.280 ;
        RECT 142.790 4.350 143.330 5.280 ;
        RECT 144.170 4.350 144.710 5.280 ;
        RECT 145.550 4.350 146.090 5.280 ;
        RECT 146.930 4.350 147.470 5.280 ;
        RECT 148.310 4.350 148.850 5.280 ;
        RECT 149.690 4.350 150.230 5.280 ;
        RECT 151.070 4.350 151.610 5.280 ;
        RECT 152.450 4.350 152.990 5.280 ;
        RECT 153.830 4.350 154.370 5.280 ;
        RECT 155.210 4.350 155.750 5.280 ;
        RECT 156.590 4.350 157.130 5.280 ;
        RECT 157.970 4.350 158.510 5.280 ;
        RECT 159.350 4.350 159.890 5.280 ;
        RECT 160.730 4.350 161.270 5.280 ;
        RECT 162.110 4.920 164.990 5.280 ;
        RECT 166.050 5.280 194.990 19.560 ;
        RECT 196.050 5.280 224.990 19.560 ;
        RECT 226.050 5.280 254.990 19.560 ;
        RECT 166.050 4.920 190.250 5.280 ;
        RECT 162.110 4.350 190.250 4.920 ;
        RECT 191.090 4.350 191.630 5.280 ;
        RECT 192.470 4.350 193.010 5.280 ;
        RECT 193.850 4.350 194.390 5.280 ;
        RECT 195.230 4.350 195.770 4.920 ;
        RECT 196.610 4.350 197.150 5.280 ;
        RECT 197.990 4.350 198.530 5.280 ;
        RECT 199.370 4.350 199.910 5.280 ;
        RECT 200.750 4.350 201.290 5.280 ;
        RECT 202.130 4.350 202.670 5.280 ;
        RECT 203.510 4.350 204.050 5.280 ;
        RECT 204.890 4.350 205.430 5.280 ;
        RECT 206.270 4.350 206.810 5.280 ;
        RECT 207.650 4.350 208.190 5.280 ;
        RECT 209.030 4.350 209.570 5.280 ;
        RECT 210.410 4.350 210.950 5.280 ;
        RECT 211.790 4.350 212.330 5.280 ;
        RECT 213.170 4.350 213.710 5.280 ;
        RECT 214.550 4.350 215.090 5.280 ;
        RECT 215.930 4.350 216.470 5.280 ;
        RECT 217.310 4.350 217.850 5.280 ;
        RECT 218.690 4.350 219.230 5.280 ;
        RECT 220.070 4.350 220.610 5.280 ;
        RECT 221.450 4.350 221.990 5.280 ;
        RECT 222.830 4.350 223.370 5.280 ;
        RECT 224.210 4.350 224.750 5.280 ;
        RECT 226.050 4.920 226.130 5.280 ;
        RECT 225.590 4.350 226.130 4.920 ;
        RECT 226.970 4.350 227.510 5.280 ;
        RECT 228.350 4.350 228.890 5.280 ;
        RECT 229.730 4.350 230.270 5.280 ;
        RECT 231.110 4.350 231.650 5.280 ;
        RECT 232.490 4.350 233.030 5.280 ;
        RECT 233.870 4.350 234.410 5.280 ;
        RECT 235.250 4.350 235.790 5.280 ;
        RECT 236.630 4.350 237.170 5.280 ;
        RECT 238.010 4.350 238.550 5.280 ;
        RECT 239.390 4.350 239.930 5.280 ;
        RECT 240.770 4.350 241.310 5.280 ;
        RECT 242.150 4.350 242.690 5.280 ;
        RECT 243.530 4.350 244.070 5.280 ;
        RECT 244.910 4.350 245.450 5.280 ;
        RECT 246.290 4.350 246.830 5.280 ;
        RECT 247.670 4.350 248.210 5.280 ;
        RECT 249.050 4.350 249.590 5.280 ;
        RECT 250.430 4.350 250.970 5.280 ;
        RECT 251.810 4.350 252.350 5.280 ;
        RECT 253.190 4.350 253.730 5.280 ;
        RECT 254.570 4.920 254.990 5.280 ;
        RECT 256.050 5.280 284.990 19.560 ;
        RECT 286.050 5.280 314.990 19.560 ;
        RECT 316.050 5.280 344.990 19.560 ;
        RECT 346.050 5.280 349.500 19.560 ;
        RECT 256.050 4.920 256.490 5.280 ;
        RECT 254.570 4.350 255.110 4.920 ;
        RECT 255.950 4.350 256.490 4.920 ;
        RECT 257.330 4.350 257.870 5.280 ;
        RECT 258.710 4.350 259.250 5.280 ;
        RECT 260.090 4.350 260.630 5.280 ;
        RECT 261.470 4.350 262.010 5.280 ;
        RECT 262.850 4.350 263.390 5.280 ;
        RECT 264.230 4.350 264.770 5.280 ;
        RECT 265.610 4.350 266.150 5.280 ;
        RECT 266.990 4.350 267.530 5.280 ;
        RECT 268.370 4.350 268.910 5.280 ;
        RECT 269.750 4.350 270.290 5.280 ;
        RECT 271.130 4.350 271.670 5.280 ;
        RECT 272.510 4.350 273.050 5.280 ;
        RECT 273.890 4.350 274.430 5.280 ;
        RECT 275.270 4.350 275.810 5.280 ;
        RECT 276.650 4.350 277.190 5.280 ;
        RECT 278.030 4.350 278.570 5.280 ;
        RECT 279.410 4.350 279.950 5.280 ;
        RECT 280.790 4.350 281.330 5.280 ;
        RECT 282.170 4.350 282.710 5.280 ;
        RECT 283.550 4.350 284.090 5.280 ;
        RECT 284.930 4.920 284.990 5.280 ;
        RECT 284.930 4.350 285.470 4.920 ;
        RECT 286.310 4.350 286.850 5.280 ;
        RECT 287.690 4.350 288.230 5.280 ;
        RECT 289.070 4.350 289.610 5.280 ;
        RECT 290.450 4.350 290.990 5.280 ;
        RECT 291.830 4.350 292.370 5.280 ;
        RECT 293.210 4.350 293.750 5.280 ;
        RECT 294.590 4.350 295.130 5.280 ;
        RECT 295.970 4.350 296.510 5.280 ;
        RECT 297.350 4.350 297.890 5.280 ;
        RECT 298.730 4.350 299.270 5.280 ;
        RECT 300.110 4.350 300.650 5.280 ;
        RECT 301.490 4.350 302.030 5.280 ;
        RECT 302.870 4.350 303.410 5.280 ;
        RECT 304.250 4.350 304.790 5.280 ;
        RECT 305.630 4.350 306.170 5.280 ;
        RECT 307.010 4.350 307.550 5.280 ;
        RECT 308.390 4.350 308.930 5.280 ;
        RECT 309.770 4.350 310.310 5.280 ;
        RECT 311.150 4.350 311.690 5.280 ;
        RECT 312.530 4.350 313.070 5.280 ;
        RECT 313.910 4.350 314.450 5.280 ;
        RECT 315.290 4.350 315.830 4.920 ;
        RECT 316.670 4.350 317.210 5.280 ;
        RECT 318.050 4.350 318.590 5.280 ;
        RECT 319.430 4.350 319.970 5.280 ;
        RECT 320.810 4.350 321.350 5.280 ;
        RECT 322.190 4.350 322.730 5.280 ;
        RECT 323.570 4.350 324.110 5.280 ;
        RECT 324.950 4.350 325.490 5.280 ;
        RECT 326.330 4.350 326.870 5.280 ;
        RECT 327.710 4.350 328.250 5.280 ;
        RECT 329.090 4.350 329.630 5.280 ;
        RECT 330.470 4.350 331.010 5.280 ;
        RECT 331.850 4.350 332.390 5.280 ;
        RECT 333.230 4.350 333.770 5.280 ;
        RECT 334.610 4.350 335.150 5.280 ;
        RECT 335.990 4.350 336.530 5.280 ;
        RECT 337.370 4.350 337.910 5.280 ;
        RECT 338.750 4.350 339.290 5.280 ;
        RECT 340.130 4.350 340.670 5.280 ;
        RECT 341.510 4.350 342.050 5.280 ;
        RECT 342.890 4.350 343.430 5.280 ;
        RECT 344.270 4.350 344.810 5.280 ;
        RECT 346.050 4.920 346.190 5.280 ;
        RECT 345.650 4.350 346.190 4.920 ;
        RECT 347.030 4.350 347.570 5.280 ;
        RECT 348.410 4.350 348.950 5.280 ;
      LAYER met3 ;
        RECT 5.400 18.000 142.995 18.865 ;
        RECT 4.910 17.650 142.995 18.000 ;
        RECT 4.910 17.360 5.120 17.650 ;
        RECT 5.400 15.960 142.995 16.350 ;
        RECT 4.910 15.320 142.995 15.960 ;
        RECT 5.400 13.920 142.995 15.320 ;
        RECT 4.910 13.280 142.995 13.920 ;
        RECT 5.400 12.250 142.995 13.280 ;
        RECT 4.910 11.240 5.120 11.880 ;
        RECT 5.400 9.840 142.995 10.950 ;
        RECT 4.910 9.200 142.995 9.840 ;
        RECT 5.400 7.800 142.995 9.200 ;
        RECT 4.910 7.160 142.995 7.800 ;
        RECT 5.400 6.850 142.995 7.160 ;
  END
END mprj_logic_high
END LIBRARY

