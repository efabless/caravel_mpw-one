magic
tech sky130A
magscale 1 2
timestamp 1622561373
<< obsli1 >>
rect 1104 1071 5888 5457
<< obsm1 >>
rect 474 1040 6518 5488
<< metal2 >>
rect 938 6200 994 7000
rect 1398 6200 1454 7000
rect 1858 6200 1914 7000
rect 2778 6200 2834 7000
rect 3238 6200 3294 7000
rect 4158 6200 4214 7000
rect 4618 6200 4674 7000
rect 5538 6200 5594 7000
rect 5998 6200 6054 7000
rect 6458 6200 6514 7000
rect 478 0 534 800
rect 938 0 994 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 3698 0 3754 800
rect 4158 0 4214 800
rect 5078 0 5134 800
rect 5538 0 5594 800
rect 5998 0 6054 800
<< obsm2 >>
rect 480 6144 882 6225
rect 1050 6144 1342 6225
rect 1510 6144 1802 6225
rect 1970 6144 2722 6225
rect 2890 6144 3182 6225
rect 3350 6144 4102 6225
rect 4270 6144 4562 6225
rect 4730 6144 5482 6225
rect 5650 6144 5942 6225
rect 6110 6144 6402 6225
rect 480 856 6512 6144
rect 590 711 882 856
rect 1050 711 1342 856
rect 1510 711 2262 856
rect 2430 711 2722 856
rect 2890 711 3642 856
rect 3810 711 4102 856
rect 4270 711 5022 856
rect 5190 711 5482 856
rect 5650 711 5942 856
rect 6110 711 6512 856
<< metal3 >>
rect 0 6128 800 6248
rect 0 5448 800 5568
rect 6200 5448 7000 5568
rect 6200 4768 7000 4888
rect 0 4088 800 4208
rect 0 3408 800 3528
rect 6200 3408 7000 3528
rect 6200 2728 7000 2848
rect 0 2048 800 2168
rect 0 1368 800 1488
rect 6200 1368 7000 1488
rect 6200 688 7000 808
<< obsm3 >>
rect 880 6048 6200 6221
rect 800 5648 6200 6048
rect 880 5368 6120 5648
rect 800 4968 6200 5368
rect 800 4688 6120 4968
rect 800 4288 6200 4688
rect 880 4008 6200 4288
rect 800 3608 6200 4008
rect 880 3328 6120 3608
rect 800 2928 6200 3328
rect 800 2648 6120 2928
rect 800 2248 6200 2648
rect 880 1968 6200 2248
rect 800 1568 6200 1968
rect 880 1288 6120 1568
rect 800 888 6200 1288
rect 800 715 6120 888
<< metal4 >>
rect 1743 1040 2063 5488
rect 2541 1040 2861 5488
rect 3340 1040 3660 5488
rect 4139 1040 4459 5488
rect 4937 1040 5257 5488
<< obsm4 >>
rect 2143 1040 2461 5488
rect 2941 1040 3260 5488
rect 3740 1040 4059 5488
<< metal5 >>
rect 1104 4900 5888 5220
rect 1104 4096 5888 4416
rect 1104 3292 5888 3612
rect 1104 2488 5888 2808
rect 1104 1684 5888 2004
<< labels >>
rlabel metal2 s 938 0 994 800 6 mask_rev[0]
port 1 nsew signal output
rlabel metal2 s 1398 6200 1454 7000 6 mask_rev[10]
port 2 nsew signal output
rlabel metal2 s 2778 6200 2834 7000 6 mask_rev[11]
port 3 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 mask_rev[12]
port 4 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 mask_rev[13]
port 5 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 mask_rev[14]
port 6 nsew signal output
rlabel metal2 s 3238 6200 3294 7000 6 mask_rev[15]
port 7 nsew signal output
rlabel metal2 s 1858 6200 1914 7000 6 mask_rev[16]
port 8 nsew signal output
rlabel metal2 s 5538 6200 5594 7000 6 mask_rev[17]
port 9 nsew signal output
rlabel metal2 s 4618 6200 4674 7000 6 mask_rev[18]
port 10 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 mask_rev[19]
port 11 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 mask_rev[1]
port 12 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 mask_rev[20]
port 13 nsew signal output
rlabel metal2 s 2318 0 2374 800 6 mask_rev[21]
port 14 nsew signal output
rlabel metal3 s 6200 688 7000 808 6 mask_rev[22]
port 15 nsew signal output
rlabel metal3 s 6200 5448 7000 5568 6 mask_rev[23]
port 16 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 mask_rev[24]
port 17 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 mask_rev[25]
port 18 nsew signal output
rlabel metal3 s 6200 4768 7000 4888 6 mask_rev[26]
port 19 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 mask_rev[27]
port 20 nsew signal output
rlabel metal2 s 478 0 534 800 6 mask_rev[28]
port 21 nsew signal output
rlabel metal3 s 6200 1368 7000 1488 6 mask_rev[29]
port 22 nsew signal output
rlabel metal2 s 6458 6200 6514 7000 6 mask_rev[2]
port 23 nsew signal output
rlabel metal3 s 6200 2728 7000 2848 6 mask_rev[30]
port 24 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 mask_rev[31]
port 25 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 mask_rev[3]
port 26 nsew signal output
rlabel metal2 s 1398 0 1454 800 6 mask_rev[4]
port 27 nsew signal output
rlabel metal2 s 938 6200 994 7000 6 mask_rev[5]
port 28 nsew signal output
rlabel metal2 s 5998 6200 6054 7000 6 mask_rev[6]
port 29 nsew signal output
rlabel metal2 s 4158 6200 4214 7000 6 mask_rev[7]
port 30 nsew signal output
rlabel metal3 s 6200 3408 7000 3528 6 mask_rev[8]
port 31 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 mask_rev[9]
port 32 nsew signal output
rlabel metal4 s 4937 1040 5257 5488 6 VPWR
port 33 nsew power bidirectional
rlabel metal4 s 3340 1040 3660 5488 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 1743 1040 2063 5488 6 VPWR
port 35 nsew power bidirectional
rlabel metal5 s 1104 4900 5888 5220 6 VPWR
port 36 nsew power bidirectional
rlabel metal5 s 1104 3292 5888 3612 6 VPWR
port 37 nsew power bidirectional
rlabel metal5 s 1104 1684 5888 2004 6 VPWR
port 38 nsew power bidirectional
rlabel metal4 s 4139 1040 4459 5488 6 VGND
port 39 nsew ground bidirectional
rlabel metal4 s 2541 1040 2861 5488 6 VGND
port 40 nsew ground bidirectional
rlabel metal5 s 1104 4096 5888 4416 6 VGND
port 41 nsew ground bidirectional
rlabel metal5 s 1104 2488 5888 2808 6 VGND
port 42 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 7000 7000
string LEFview TRUE
string GDS_FILE /project/openlane/user_id_programming/runs/user_id_programming/results/magic/user_id_programming.gds
string GDS_END 90386
string GDS_START 24124
<< end >>

