VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gpio_control_block
  CLASS BLOCK ;
  FOREIGN gpio_control_block ;
  ORIGIN 0.000 0.000 ;
  SIZE 169.670 BY 91.720 ;
  PIN mgmt_gpio_in
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.670 0.000 169.670 0.600 ;
    END
  END mgmt_gpio_in
  PIN mgmt_gpio_oeb
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.670 3.400 169.670 4.000 ;
    END
  END mgmt_gpio_oeb
  PIN mgmt_gpio_out
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.670 7.480 169.670 8.080 ;
    END
  END mgmt_gpio_out
  PIN pad_gpio_ana_en
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.670 11.560 169.670 12.160 ;
    END
  END pad_gpio_ana_en
  PIN pad_gpio_ana_pol
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.670 15.640 169.670 16.240 ;
    END
  END pad_gpio_ana_pol
  PIN pad_gpio_ana_sel
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.670 19.720 169.670 20.320 ;
    END
  END pad_gpio_ana_sel
  PIN pad_gpio_dm[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.670 23.800 169.670 24.400 ;
    END
  END pad_gpio_dm[0]
  PIN pad_gpio_dm[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.670 27.200 169.670 27.800 ;
    END
  END pad_gpio_dm[1]
  PIN pad_gpio_dm[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.670 31.280 169.670 31.880 ;
    END
  END pad_gpio_dm[2]
  PIN pad_gpio_holdover
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.670 35.360 169.670 35.960 ;
    END
  END pad_gpio_holdover
  PIN pad_gpio_ib_mode_sel
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.670 39.440 169.670 40.040 ;
    END
  END pad_gpio_ib_mode_sel
  PIN pad_gpio_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.670 43.520 169.670 44.120 ;
    END
  END pad_gpio_in
  PIN pad_gpio_inenb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.670 47.600 169.670 48.200 ;
    END
  END pad_gpio_inenb
  PIN pad_gpio_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.670 51.000 169.670 51.600 ;
    END
  END pad_gpio_out
  PIN pad_gpio_outenb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.670 55.080 169.670 55.680 ;
    END
  END pad_gpio_outenb
  PIN pad_gpio_slow_sel
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.670 59.160 169.670 59.760 ;
    END
  END pad_gpio_slow_sel
  PIN pad_gpio_vtrip_sel
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.670 63.240 169.670 63.840 ;
    END
  END pad_gpio_vtrip_sel
  PIN resetn
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.670 67.320 169.670 67.920 ;
    END
  END resetn
  PIN serial_clock
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.670 71.400 169.670 72.000 ;
    END
  END serial_clock
  PIN serial_data_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.670 74.800 169.670 75.400 ;
    END
  END serial_data_in
  PIN serial_data_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.670 78.880 169.670 79.480 ;
    END
  END serial_data_out
  PIN user_gpio_in
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.670 82.960 169.670 83.560 ;
    END
  END user_gpio_in
  PIN user_gpio_oeb
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.670 87.040 169.670 87.640 ;
    END
  END user_gpio_oeb
  PIN user_gpio_out
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.670 91.120 169.670 91.720 ;
    END
  END user_gpio_out
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.190 20.645 44.350 22.245 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.190 32.855 44.350 34.455 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.190 9.395 57.085 80.285 ;
      LAYER met1 ;
        RECT 0.190 9.240 120.640 81.860 ;
      LAYER met2 ;
        RECT 2.590 0.115 120.620 91.605 ;
      LAYER met3 ;
        RECT 6.780 79.880 49.670 80.365 ;
        RECT 6.780 78.480 49.270 79.880 ;
        RECT 6.780 75.800 49.670 78.480 ;
        RECT 6.780 74.400 49.270 75.800 ;
        RECT 6.780 72.400 49.670 74.400 ;
        RECT 6.780 71.000 49.270 72.400 ;
        RECT 6.780 68.320 49.670 71.000 ;
        RECT 6.780 66.920 49.270 68.320 ;
        RECT 6.780 64.240 49.670 66.920 ;
        RECT 6.780 62.840 49.270 64.240 ;
        RECT 6.780 60.160 49.670 62.840 ;
        RECT 6.780 58.760 49.270 60.160 ;
        RECT 6.780 56.080 49.670 58.760 ;
        RECT 6.780 54.680 49.270 56.080 ;
        RECT 6.780 52.000 49.670 54.680 ;
        RECT 6.780 50.600 49.270 52.000 ;
        RECT 6.780 48.600 49.670 50.600 ;
        RECT 6.780 47.200 49.270 48.600 ;
        RECT 6.780 44.520 49.670 47.200 ;
        RECT 6.780 43.120 49.270 44.520 ;
        RECT 6.780 40.440 49.670 43.120 ;
        RECT 6.780 39.040 49.270 40.440 ;
        RECT 6.780 36.360 49.670 39.040 ;
        RECT 6.780 34.960 49.270 36.360 ;
        RECT 6.780 32.280 49.670 34.960 ;
        RECT 6.780 30.880 49.270 32.280 ;
        RECT 6.780 28.200 49.670 30.880 ;
        RECT 6.780 26.800 49.270 28.200 ;
        RECT 6.780 24.800 49.670 26.800 ;
        RECT 6.780 23.400 49.270 24.800 ;
        RECT 6.780 20.720 49.670 23.400 ;
        RECT 6.780 19.320 49.270 20.720 ;
        RECT 6.780 16.640 49.670 19.320 ;
        RECT 6.780 15.240 49.270 16.640 ;
        RECT 6.780 12.560 49.670 15.240 ;
        RECT 6.780 11.160 49.270 12.560 ;
        RECT 6.780 9.315 49.670 11.160 ;
      LAYER met4 ;
        RECT 6.780 9.240 37.955 80.440 ;
      LAYER met5 ;
        RECT 0.190 36.055 44.350 71.070 ;
  END
END gpio_control_block
END LIBRARY

