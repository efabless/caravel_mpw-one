VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_core
  CLASS BLOCK ;
  FOREIGN mgmt_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 2150.000 BY 850.000 ;
  PIN clock
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END clock
  PIN core_clk
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 571.410 846.000 571.690 850.000 ;
    END
  END core_clk
  PIN core_rstn
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1127.090 846.000 1127.370 850.000 ;
    END
  END core_rstn
  PIN flash_clk
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END flash_clk
  PIN flash_clk_ieb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END flash_clk_ieb
  PIN flash_clk_oeb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END flash_clk_oeb
  PIN flash_csb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END flash_csb
  PIN flash_csb_ieb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END flash_csb_ieb
  PIN flash_csb_oeb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END flash_csb_oeb
  PIN flash_io0_di
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END flash_io0_di
  PIN flash_io0_do
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END flash_io0_do
  PIN flash_io0_ieb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END flash_io0_ieb
  PIN flash_io0_oeb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END flash_io0_oeb
  PIN flash_io1_di
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END flash_io1_di
  PIN flash_io1_do
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END flash_io1_do
  PIN flash_io1_ieb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END flash_io1_ieb
  PIN flash_io1_oeb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END flash_io1_oeb
  PIN gpio_in_pad
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END gpio_in_pad
  PIN gpio_inenb_pad
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END gpio_inenb_pad
  PIN gpio_mode0_pad
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END gpio_mode0_pad
  PIN gpio_mode1_pad
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END gpio_mode1_pad
  PIN gpio_out_pad
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END gpio_out_pad
  PIN gpio_outenb_pad
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END gpio_outenb_pad
  PIN jtag_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2146.000 337.320 2150.000 337.920 ;
    END
  END jtag_out
  PIN jtag_outenb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2146.000 334.600 2150.000 335.200 ;
    END
  END jtag_outenb
  PIN la_input[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1125.250 846.000 1125.530 850.000 ;
    END
  END la_input[0]
  PIN la_input[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1128.930 846.000 1129.210 850.000 ;
    END
  END la_input[100]
  PIN la_input[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1123.410 846.000 1123.690 850.000 ;
    END
  END la_input[101]
  PIN la_input[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1130.770 846.000 1131.050 850.000 ;
    END
  END la_input[102]
  PIN la_input[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1121.570 846.000 1121.850 850.000 ;
    END
  END la_input[103]
  PIN la_input[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.610 846.000 1132.890 850.000 ;
    END
  END la_input[104]
  PIN la_input[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1119.730 846.000 1120.010 850.000 ;
    END
  END la_input[105]
  PIN la_input[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1134.450 846.000 1134.730 850.000 ;
    END
  END la_input[106]
  PIN la_input[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1117.890 846.000 1118.170 850.000 ;
    END
  END la_input[107]
  PIN la_input[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1136.290 846.000 1136.570 850.000 ;
    END
  END la_input[108]
  PIN la_input[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1116.050 846.000 1116.330 850.000 ;
    END
  END la_input[109]
  PIN la_input[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1138.130 846.000 1138.410 850.000 ;
    END
  END la_input[10]
  PIN la_input[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1114.210 846.000 1114.490 850.000 ;
    END
  END la_input[110]
  PIN la_input[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1139.970 846.000 1140.250 850.000 ;
    END
  END la_input[111]
  PIN la_input[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1112.370 846.000 1112.650 850.000 ;
    END
  END la_input[112]
  PIN la_input[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1141.810 846.000 1142.090 850.000 ;
    END
  END la_input[113]
  PIN la_input[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1110.530 846.000 1110.810 850.000 ;
    END
  END la_input[114]
  PIN la_input[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1143.650 846.000 1143.930 850.000 ;
    END
  END la_input[115]
  PIN la_input[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1108.690 846.000 1108.970 850.000 ;
    END
  END la_input[116]
  PIN la_input[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1145.490 846.000 1145.770 850.000 ;
    END
  END la_input[117]
  PIN la_input[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1106.850 846.000 1107.130 850.000 ;
    END
  END la_input[118]
  PIN la_input[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1147.330 846.000 1147.610 850.000 ;
    END
  END la_input[119]
  PIN la_input[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1105.010 846.000 1105.290 850.000 ;
    END
  END la_input[11]
  PIN la_input[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1149.170 846.000 1149.450 850.000 ;
    END
  END la_input[120]
  PIN la_input[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1103.170 846.000 1103.450 850.000 ;
    END
  END la_input[121]
  PIN la_input[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1151.010 846.000 1151.290 850.000 ;
    END
  END la_input[122]
  PIN la_input[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1101.330 846.000 1101.610 850.000 ;
    END
  END la_input[123]
  PIN la_input[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1152.850 846.000 1153.130 850.000 ;
    END
  END la_input[124]
  PIN la_input[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1099.490 846.000 1099.770 850.000 ;
    END
  END la_input[125]
  PIN la_input[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1154.690 846.000 1154.970 850.000 ;
    END
  END la_input[126]
  PIN la_input[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1097.650 846.000 1097.930 850.000 ;
    END
  END la_input[127]
  PIN la_input[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1156.530 846.000 1156.810 850.000 ;
    END
  END la_input[12]
  PIN la_input[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1095.810 846.000 1096.090 850.000 ;
    END
  END la_input[13]
  PIN la_input[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1158.370 846.000 1158.650 850.000 ;
    END
  END la_input[14]
  PIN la_input[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1093.970 846.000 1094.250 850.000 ;
    END
  END la_input[15]
  PIN la_input[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1160.210 846.000 1160.490 850.000 ;
    END
  END la_input[16]
  PIN la_input[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1092.130 846.000 1092.410 850.000 ;
    END
  END la_input[17]
  PIN la_input[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.050 846.000 1162.330 850.000 ;
    END
  END la_input[18]
  PIN la_input[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.290 846.000 1090.570 850.000 ;
    END
  END la_input[19]
  PIN la_input[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1163.890 846.000 1164.170 850.000 ;
    END
  END la_input[1]
  PIN la_input[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1088.450 846.000 1088.730 850.000 ;
    END
  END la_input[20]
  PIN la_input[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1165.730 846.000 1166.010 850.000 ;
    END
  END la_input[21]
  PIN la_input[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1086.610 846.000 1086.890 850.000 ;
    END
  END la_input[22]
  PIN la_input[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1167.570 846.000 1167.850 850.000 ;
    END
  END la_input[23]
  PIN la_input[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1084.770 846.000 1085.050 850.000 ;
    END
  END la_input[24]
  PIN la_input[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1169.410 846.000 1169.690 850.000 ;
    END
  END la_input[25]
  PIN la_input[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1082.930 846.000 1083.210 850.000 ;
    END
  END la_input[26]
  PIN la_input[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1171.250 846.000 1171.530 850.000 ;
    END
  END la_input[27]
  PIN la_input[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1081.090 846.000 1081.370 850.000 ;
    END
  END la_input[28]
  PIN la_input[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1173.090 846.000 1173.370 850.000 ;
    END
  END la_input[29]
  PIN la_input[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1079.250 846.000 1079.530 850.000 ;
    END
  END la_input[2]
  PIN la_input[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1174.930 846.000 1175.210 850.000 ;
    END
  END la_input[30]
  PIN la_input[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1077.410 846.000 1077.690 850.000 ;
    END
  END la_input[31]
  PIN la_input[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1176.770 846.000 1177.050 850.000 ;
    END
  END la_input[32]
  PIN la_input[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1075.570 846.000 1075.850 850.000 ;
    END
  END la_input[33]
  PIN la_input[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1178.610 846.000 1178.890 850.000 ;
    END
  END la_input[34]
  PIN la_input[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.730 846.000 1074.010 850.000 ;
    END
  END la_input[35]
  PIN la_input[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1180.450 846.000 1180.730 850.000 ;
    END
  END la_input[36]
  PIN la_input[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1071.890 846.000 1072.170 850.000 ;
    END
  END la_input[37]
  PIN la_input[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1182.290 846.000 1182.570 850.000 ;
    END
  END la_input[38]
  PIN la_input[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1070.050 846.000 1070.330 850.000 ;
    END
  END la_input[39]
  PIN la_input[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1184.130 846.000 1184.410 850.000 ;
    END
  END la_input[3]
  PIN la_input[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1068.210 846.000 1068.490 850.000 ;
    END
  END la_input[40]
  PIN la_input[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.970 846.000 1186.250 850.000 ;
    END
  END la_input[41]
  PIN la_input[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1066.370 846.000 1066.650 850.000 ;
    END
  END la_input[42]
  PIN la_input[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1187.810 846.000 1188.090 850.000 ;
    END
  END la_input[43]
  PIN la_input[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1064.530 846.000 1064.810 850.000 ;
    END
  END la_input[44]
  PIN la_input[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1189.650 846.000 1189.930 850.000 ;
    END
  END la_input[45]
  PIN la_input[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1062.690 846.000 1062.970 850.000 ;
    END
  END la_input[46]
  PIN la_input[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1191.490 846.000 1191.770 850.000 ;
    END
  END la_input[47]
  PIN la_input[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1060.850 846.000 1061.130 850.000 ;
    END
  END la_input[48]
  PIN la_input[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1193.330 846.000 1193.610 850.000 ;
    END
  END la_input[49]
  PIN la_input[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1059.010 846.000 1059.290 850.000 ;
    END
  END la_input[4]
  PIN la_input[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1195.170 846.000 1195.450 850.000 ;
    END
  END la_input[50]
  PIN la_input[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1057.170 846.000 1057.450 850.000 ;
    END
  END la_input[51]
  PIN la_input[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.010 846.000 1197.290 850.000 ;
    END
  END la_input[52]
  PIN la_input[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.330 846.000 1055.610 850.000 ;
    END
  END la_input[53]
  PIN la_input[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1198.850 846.000 1199.130 850.000 ;
    END
  END la_input[54]
  PIN la_input[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1053.490 846.000 1053.770 850.000 ;
    END
  END la_input[55]
  PIN la_input[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1200.690 846.000 1200.970 850.000 ;
    END
  END la_input[56]
  PIN la_input[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1051.650 846.000 1051.930 850.000 ;
    END
  END la_input[57]
  PIN la_input[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1202.530 846.000 1202.810 850.000 ;
    END
  END la_input[58]
  PIN la_input[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1049.810 846.000 1050.090 850.000 ;
    END
  END la_input[59]
  PIN la_input[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1204.370 846.000 1204.650 850.000 ;
    END
  END la_input[5]
  PIN la_input[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1047.970 846.000 1048.250 850.000 ;
    END
  END la_input[60]
  PIN la_input[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1206.210 846.000 1206.490 850.000 ;
    END
  END la_input[61]
  PIN la_input[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1046.130 846.000 1046.410 850.000 ;
    END
  END la_input[62]
  PIN la_input[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1208.050 846.000 1208.330 850.000 ;
    END
  END la_input[63]
  PIN la_input[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1044.290 846.000 1044.570 850.000 ;
    END
  END la_input[64]
  PIN la_input[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1209.890 846.000 1210.170 850.000 ;
    END
  END la_input[65]
  PIN la_input[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1042.450 846.000 1042.730 850.000 ;
    END
  END la_input[66]
  PIN la_input[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1211.730 846.000 1212.010 850.000 ;
    END
  END la_input[67]
  PIN la_input[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1040.610 846.000 1040.890 850.000 ;
    END
  END la_input[68]
  PIN la_input[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1213.570 846.000 1213.850 850.000 ;
    END
  END la_input[69]
  PIN la_input[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1038.770 846.000 1039.050 850.000 ;
    END
  END la_input[6]
  PIN la_input[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.410 846.000 1215.690 850.000 ;
    END
  END la_input[70]
  PIN la_input[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1036.930 846.000 1037.210 850.000 ;
    END
  END la_input[71]
  PIN la_input[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1217.250 846.000 1217.530 850.000 ;
    END
  END la_input[72]
  PIN la_input[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1035.090 846.000 1035.370 850.000 ;
    END
  END la_input[73]
  PIN la_input[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1219.090 846.000 1219.370 850.000 ;
    END
  END la_input[74]
  PIN la_input[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1033.250 846.000 1033.530 850.000 ;
    END
  END la_input[75]
  PIN la_input[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1220.930 846.000 1221.210 850.000 ;
    END
  END la_input[76]
  PIN la_input[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1031.410 846.000 1031.690 850.000 ;
    END
  END la_input[77]
  PIN la_input[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1222.770 846.000 1223.050 850.000 ;
    END
  END la_input[78]
  PIN la_input[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1029.570 846.000 1029.850 850.000 ;
    END
  END la_input[79]
  PIN la_input[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1224.610 846.000 1224.890 850.000 ;
    END
  END la_input[7]
  PIN la_input[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1027.730 846.000 1028.010 850.000 ;
    END
  END la_input[80]
  PIN la_input[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1226.450 846.000 1226.730 850.000 ;
    END
  END la_input[81]
  PIN la_input[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.890 846.000 1026.170 850.000 ;
    END
  END la_input[82]
  PIN la_input[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1228.290 846.000 1228.570 850.000 ;
    END
  END la_input[83]
  PIN la_input[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1024.050 846.000 1024.330 850.000 ;
    END
  END la_input[84]
  PIN la_input[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1230.130 846.000 1230.410 850.000 ;
    END
  END la_input[85]
  PIN la_input[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1022.210 846.000 1022.490 850.000 ;
    END
  END la_input[86]
  PIN la_input[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1231.970 846.000 1232.250 850.000 ;
    END
  END la_input[87]
  PIN la_input[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1020.370 846.000 1020.650 850.000 ;
    END
  END la_input[88]
  PIN la_input[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1233.810 846.000 1234.090 850.000 ;
    END
  END la_input[89]
  PIN la_input[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1018.530 846.000 1018.810 850.000 ;
    END
  END la_input[8]
  PIN la_input[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1235.650 846.000 1235.930 850.000 ;
    END
  END la_input[90]
  PIN la_input[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1016.690 846.000 1016.970 850.000 ;
    END
  END la_input[91]
  PIN la_input[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1237.490 846.000 1237.770 850.000 ;
    END
  END la_input[92]
  PIN la_input[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1014.850 846.000 1015.130 850.000 ;
    END
  END la_input[93]
  PIN la_input[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1239.330 846.000 1239.610 850.000 ;
    END
  END la_input[94]
  PIN la_input[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1013.010 846.000 1013.290 850.000 ;
    END
  END la_input[95]
  PIN la_input[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1241.170 846.000 1241.450 850.000 ;
    END
  END la_input[96]
  PIN la_input[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1011.170 846.000 1011.450 850.000 ;
    END
  END la_input[97]
  PIN la_input[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1243.010 846.000 1243.290 850.000 ;
    END
  END la_input[98]
  PIN la_input[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1009.330 846.000 1009.610 850.000 ;
    END
  END la_input[99]
  PIN la_input[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1244.850 846.000 1245.130 850.000 ;
    END
  END la_input[9]
  PIN la_oen[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1007.490 846.000 1007.770 850.000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1246.690 846.000 1246.970 850.000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1005.650 846.000 1005.930 850.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1248.530 846.000 1248.810 850.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1003.810 846.000 1004.090 850.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1250.370 846.000 1250.650 850.000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1001.970 846.000 1002.250 850.000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1252.210 846.000 1252.490 850.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1000.130 846.000 1000.410 850.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1254.050 846.000 1254.330 850.000 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 998.290 846.000 998.570 850.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1255.890 846.000 1256.170 850.000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 996.450 846.000 996.730 850.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1257.730 846.000 1258.010 850.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 994.610 846.000 994.890 850.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1259.570 846.000 1259.850 850.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 992.770 846.000 993.050 850.000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1261.410 846.000 1261.690 850.000 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 990.930 846.000 991.210 850.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1263.250 846.000 1263.530 850.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 989.090 846.000 989.370 850.000 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1265.090 846.000 1265.370 850.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 987.250 846.000 987.530 850.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1266.930 846.000 1267.210 850.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 985.410 846.000 985.690 850.000 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1268.770 846.000 1269.050 850.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 983.570 846.000 983.850 850.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1270.610 846.000 1270.890 850.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 981.730 846.000 982.010 850.000 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1272.450 846.000 1272.730 850.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 979.890 846.000 980.170 850.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1274.290 846.000 1274.570 850.000 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 978.050 846.000 978.330 850.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1276.130 846.000 1276.410 850.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 976.210 846.000 976.490 850.000 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1277.970 846.000 1278.250 850.000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 974.370 846.000 974.650 850.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1279.810 846.000 1280.090 850.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 972.530 846.000 972.810 850.000 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1281.650 846.000 1281.930 850.000 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 970.690 846.000 970.970 850.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1283.490 846.000 1283.770 850.000 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 968.850 846.000 969.130 850.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1285.330 846.000 1285.610 850.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 967.010 846.000 967.290 850.000 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1287.170 846.000 1287.450 850.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 965.170 846.000 965.450 850.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1289.010 846.000 1289.290 850.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 963.330 846.000 963.610 850.000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1290.850 846.000 1291.130 850.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 961.490 846.000 961.770 850.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1292.690 846.000 1292.970 850.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 959.650 846.000 959.930 850.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1294.530 846.000 1294.810 850.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 957.810 846.000 958.090 850.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1296.370 846.000 1296.650 850.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 955.970 846.000 956.250 850.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1298.210 846.000 1298.490 850.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 954.130 846.000 954.410 850.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1300.050 846.000 1300.330 850.000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 952.290 846.000 952.570 850.000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1301.890 846.000 1302.170 850.000 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 950.450 846.000 950.730 850.000 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1303.730 846.000 1304.010 850.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 948.610 846.000 948.890 850.000 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1305.570 846.000 1305.850 850.000 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 946.770 846.000 947.050 850.000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1307.410 846.000 1307.690 850.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 944.930 846.000 945.210 850.000 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1309.250 846.000 1309.530 850.000 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 943.090 846.000 943.370 850.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1311.090 846.000 1311.370 850.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 941.250 846.000 941.530 850.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1312.930 846.000 1313.210 850.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 939.410 846.000 939.690 850.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1314.770 846.000 1315.050 850.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 937.570 846.000 937.850 850.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1316.610 846.000 1316.890 850.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 935.730 846.000 936.010 850.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1318.450 846.000 1318.730 850.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 933.890 846.000 934.170 850.000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1320.290 846.000 1320.570 850.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 932.050 846.000 932.330 850.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1322.130 846.000 1322.410 850.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 930.210 846.000 930.490 850.000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1323.970 846.000 1324.250 850.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 928.370 846.000 928.650 850.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1325.810 846.000 1326.090 850.000 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 926.530 846.000 926.810 850.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1327.650 846.000 1327.930 850.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.690 846.000 924.970 850.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1329.490 846.000 1329.770 850.000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 922.850 846.000 923.130 850.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1331.330 846.000 1331.610 850.000 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 921.010 846.000 921.290 850.000 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1333.170 846.000 1333.450 850.000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 919.170 846.000 919.450 850.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1335.010 846.000 1335.290 850.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 917.330 846.000 917.610 850.000 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1336.850 846.000 1337.130 850.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 915.490 846.000 915.770 850.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1338.690 846.000 1338.970 850.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 913.650 846.000 913.930 850.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1340.530 846.000 1340.810 850.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 911.810 846.000 912.090 850.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1342.370 846.000 1342.650 850.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 909.970 846.000 910.250 850.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1344.210 846.000 1344.490 850.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 908.130 846.000 908.410 850.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1346.050 846.000 1346.330 850.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 906.290 846.000 906.570 850.000 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1347.890 846.000 1348.170 850.000 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 904.450 846.000 904.730 850.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1349.730 846.000 1350.010 850.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 902.610 846.000 902.890 850.000 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1351.570 846.000 1351.850 850.000 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 900.770 846.000 901.050 850.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1353.410 846.000 1353.690 850.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 898.930 846.000 899.210 850.000 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1355.250 846.000 1355.530 850.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 897.090 846.000 897.370 850.000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1357.090 846.000 1357.370 850.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 895.250 846.000 895.530 850.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1358.930 846.000 1359.210 850.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 893.410 846.000 893.690 850.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1360.770 846.000 1361.050 850.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 891.570 846.000 891.850 850.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1362.610 846.000 1362.890 850.000 ;
    END
  END la_oen[9]
  PIN la_output[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 889.730 846.000 890.010 850.000 ;
    END
  END la_output[0]
  PIN la_output[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1364.450 846.000 1364.730 850.000 ;
    END
  END la_output[100]
  PIN la_output[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 887.890 846.000 888.170 850.000 ;
    END
  END la_output[101]
  PIN la_output[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1366.290 846.000 1366.570 850.000 ;
    END
  END la_output[102]
  PIN la_output[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 886.050 846.000 886.330 850.000 ;
    END
  END la_output[103]
  PIN la_output[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1368.130 846.000 1368.410 850.000 ;
    END
  END la_output[104]
  PIN la_output[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 884.210 846.000 884.490 850.000 ;
    END
  END la_output[105]
  PIN la_output[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1369.970 846.000 1370.250 850.000 ;
    END
  END la_output[106]
  PIN la_output[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 882.370 846.000 882.650 850.000 ;
    END
  END la_output[107]
  PIN la_output[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1371.810 846.000 1372.090 850.000 ;
    END
  END la_output[108]
  PIN la_output[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 880.530 846.000 880.810 850.000 ;
    END
  END la_output[109]
  PIN la_output[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1373.650 846.000 1373.930 850.000 ;
    END
  END la_output[10]
  PIN la_output[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 878.690 846.000 878.970 850.000 ;
    END
  END la_output[110]
  PIN la_output[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1375.490 846.000 1375.770 850.000 ;
    END
  END la_output[111]
  PIN la_output[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 876.850 846.000 877.130 850.000 ;
    END
  END la_output[112]
  PIN la_output[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1377.330 846.000 1377.610 850.000 ;
    END
  END la_output[113]
  PIN la_output[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 875.010 846.000 875.290 850.000 ;
    END
  END la_output[114]
  PIN la_output[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1379.170 846.000 1379.450 850.000 ;
    END
  END la_output[115]
  PIN la_output[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 873.170 846.000 873.450 850.000 ;
    END
  END la_output[116]
  PIN la_output[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1381.010 846.000 1381.290 850.000 ;
    END
  END la_output[117]
  PIN la_output[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 871.330 846.000 871.610 850.000 ;
    END
  END la_output[118]
  PIN la_output[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1382.850 846.000 1383.130 850.000 ;
    END
  END la_output[119]
  PIN la_output[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 869.490 846.000 869.770 850.000 ;
    END
  END la_output[11]
  PIN la_output[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1384.690 846.000 1384.970 850.000 ;
    END
  END la_output[120]
  PIN la_output[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 867.650 846.000 867.930 850.000 ;
    END
  END la_output[121]
  PIN la_output[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1386.530 846.000 1386.810 850.000 ;
    END
  END la_output[122]
  PIN la_output[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 865.810 846.000 866.090 850.000 ;
    END
  END la_output[123]
  PIN la_output[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1388.370 846.000 1388.650 850.000 ;
    END
  END la_output[124]
  PIN la_output[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 863.970 846.000 864.250 850.000 ;
    END
  END la_output[125]
  PIN la_output[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1390.210 846.000 1390.490 850.000 ;
    END
  END la_output[126]
  PIN la_output[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 862.130 846.000 862.410 850.000 ;
    END
  END la_output[127]
  PIN la_output[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1392.050 846.000 1392.330 850.000 ;
    END
  END la_output[12]
  PIN la_output[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 860.290 846.000 860.570 850.000 ;
    END
  END la_output[13]
  PIN la_output[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1393.890 846.000 1394.170 850.000 ;
    END
  END la_output[14]
  PIN la_output[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 858.450 846.000 858.730 850.000 ;
    END
  END la_output[15]
  PIN la_output[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1395.730 846.000 1396.010 850.000 ;
    END
  END la_output[16]
  PIN la_output[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 856.610 846.000 856.890 850.000 ;
    END
  END la_output[17]
  PIN la_output[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1397.570 846.000 1397.850 850.000 ;
    END
  END la_output[18]
  PIN la_output[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 854.770 846.000 855.050 850.000 ;
    END
  END la_output[19]
  PIN la_output[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1399.410 846.000 1399.690 850.000 ;
    END
  END la_output[1]
  PIN la_output[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.930 846.000 853.210 850.000 ;
    END
  END la_output[20]
  PIN la_output[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1401.250 846.000 1401.530 850.000 ;
    END
  END la_output[21]
  PIN la_output[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 851.090 846.000 851.370 850.000 ;
    END
  END la_output[22]
  PIN la_output[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1403.090 846.000 1403.370 850.000 ;
    END
  END la_output[23]
  PIN la_output[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 849.250 846.000 849.530 850.000 ;
    END
  END la_output[24]
  PIN la_output[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1404.930 846.000 1405.210 850.000 ;
    END
  END la_output[25]
  PIN la_output[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 847.410 846.000 847.690 850.000 ;
    END
  END la_output[26]
  PIN la_output[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1406.770 846.000 1407.050 850.000 ;
    END
  END la_output[27]
  PIN la_output[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 845.570 846.000 845.850 850.000 ;
    END
  END la_output[28]
  PIN la_output[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1408.610 846.000 1408.890 850.000 ;
    END
  END la_output[29]
  PIN la_output[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 843.730 846.000 844.010 850.000 ;
    END
  END la_output[2]
  PIN la_output[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1410.450 846.000 1410.730 850.000 ;
    END
  END la_output[30]
  PIN la_output[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 841.890 846.000 842.170 850.000 ;
    END
  END la_output[31]
  PIN la_output[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1412.290 846.000 1412.570 850.000 ;
    END
  END la_output[32]
  PIN la_output[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 840.050 846.000 840.330 850.000 ;
    END
  END la_output[33]
  PIN la_output[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1414.130 846.000 1414.410 850.000 ;
    END
  END la_output[34]
  PIN la_output[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 838.210 846.000 838.490 850.000 ;
    END
  END la_output[35]
  PIN la_output[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1415.970 846.000 1416.250 850.000 ;
    END
  END la_output[36]
  PIN la_output[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 836.370 846.000 836.650 850.000 ;
    END
  END la_output[37]
  PIN la_output[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1417.810 846.000 1418.090 850.000 ;
    END
  END la_output[38]
  PIN la_output[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 834.530 846.000 834.810 850.000 ;
    END
  END la_output[39]
  PIN la_output[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1419.650 846.000 1419.930 850.000 ;
    END
  END la_output[3]
  PIN la_output[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 832.690 846.000 832.970 850.000 ;
    END
  END la_output[40]
  PIN la_output[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1421.490 846.000 1421.770 850.000 ;
    END
  END la_output[41]
  PIN la_output[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 830.850 846.000 831.130 850.000 ;
    END
  END la_output[42]
  PIN la_output[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1423.330 846.000 1423.610 850.000 ;
    END
  END la_output[43]
  PIN la_output[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 829.010 846.000 829.290 850.000 ;
    END
  END la_output[44]
  PIN la_output[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1425.170 846.000 1425.450 850.000 ;
    END
  END la_output[45]
  PIN la_output[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 827.170 846.000 827.450 850.000 ;
    END
  END la_output[46]
  PIN la_output[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1427.010 846.000 1427.290 850.000 ;
    END
  END la_output[47]
  PIN la_output[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 825.330 846.000 825.610 850.000 ;
    END
  END la_output[48]
  PIN la_output[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1428.850 846.000 1429.130 850.000 ;
    END
  END la_output[49]
  PIN la_output[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 823.490 846.000 823.770 850.000 ;
    END
  END la_output[4]
  PIN la_output[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1430.690 846.000 1430.970 850.000 ;
    END
  END la_output[50]
  PIN la_output[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 821.650 846.000 821.930 850.000 ;
    END
  END la_output[51]
  PIN la_output[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1432.530 846.000 1432.810 850.000 ;
    END
  END la_output[52]
  PIN la_output[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 819.810 846.000 820.090 850.000 ;
    END
  END la_output[53]
  PIN la_output[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1434.370 846.000 1434.650 850.000 ;
    END
  END la_output[54]
  PIN la_output[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.970 846.000 818.250 850.000 ;
    END
  END la_output[55]
  PIN la_output[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1436.210 846.000 1436.490 850.000 ;
    END
  END la_output[56]
  PIN la_output[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 816.130 846.000 816.410 850.000 ;
    END
  END la_output[57]
  PIN la_output[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1438.050 846.000 1438.330 850.000 ;
    END
  END la_output[58]
  PIN la_output[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 814.290 846.000 814.570 850.000 ;
    END
  END la_output[59]
  PIN la_output[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1439.890 846.000 1440.170 850.000 ;
    END
  END la_output[5]
  PIN la_output[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 812.450 846.000 812.730 850.000 ;
    END
  END la_output[60]
  PIN la_output[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1441.730 846.000 1442.010 850.000 ;
    END
  END la_output[61]
  PIN la_output[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 810.610 846.000 810.890 850.000 ;
    END
  END la_output[62]
  PIN la_output[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1443.570 846.000 1443.850 850.000 ;
    END
  END la_output[63]
  PIN la_output[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 808.770 846.000 809.050 850.000 ;
    END
  END la_output[64]
  PIN la_output[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1445.410 846.000 1445.690 850.000 ;
    END
  END la_output[65]
  PIN la_output[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 806.930 846.000 807.210 850.000 ;
    END
  END la_output[66]
  PIN la_output[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1447.250 846.000 1447.530 850.000 ;
    END
  END la_output[67]
  PIN la_output[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 805.090 846.000 805.370 850.000 ;
    END
  END la_output[68]
  PIN la_output[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1449.090 846.000 1449.370 850.000 ;
    END
  END la_output[69]
  PIN la_output[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 803.250 846.000 803.530 850.000 ;
    END
  END la_output[6]
  PIN la_output[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1450.930 846.000 1451.210 850.000 ;
    END
  END la_output[70]
  PIN la_output[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 801.410 846.000 801.690 850.000 ;
    END
  END la_output[71]
  PIN la_output[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1452.770 846.000 1453.050 850.000 ;
    END
  END la_output[72]
  PIN la_output[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 799.570 846.000 799.850 850.000 ;
    END
  END la_output[73]
  PIN la_output[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1454.610 846.000 1454.890 850.000 ;
    END
  END la_output[74]
  PIN la_output[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 797.730 846.000 798.010 850.000 ;
    END
  END la_output[75]
  PIN la_output[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1456.450 846.000 1456.730 850.000 ;
    END
  END la_output[76]
  PIN la_output[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 795.890 846.000 796.170 850.000 ;
    END
  END la_output[77]
  PIN la_output[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1458.290 846.000 1458.570 850.000 ;
    END
  END la_output[78]
  PIN la_output[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 794.050 846.000 794.330 850.000 ;
    END
  END la_output[79]
  PIN la_output[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1460.130 846.000 1460.410 850.000 ;
    END
  END la_output[7]
  PIN la_output[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 792.210 846.000 792.490 850.000 ;
    END
  END la_output[80]
  PIN la_output[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1461.970 846.000 1462.250 850.000 ;
    END
  END la_output[81]
  PIN la_output[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 790.370 846.000 790.650 850.000 ;
    END
  END la_output[82]
  PIN la_output[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1463.810 846.000 1464.090 850.000 ;
    END
  END la_output[83]
  PIN la_output[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 788.530 846.000 788.810 850.000 ;
    END
  END la_output[84]
  PIN la_output[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1465.650 846.000 1465.930 850.000 ;
    END
  END la_output[85]
  PIN la_output[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 786.690 846.000 786.970 850.000 ;
    END
  END la_output[86]
  PIN la_output[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1467.490 846.000 1467.770 850.000 ;
    END
  END la_output[87]
  PIN la_output[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 784.850 846.000 785.130 850.000 ;
    END
  END la_output[88]
  PIN la_output[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1469.330 846.000 1469.610 850.000 ;
    END
  END la_output[89]
  PIN la_output[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 783.010 846.000 783.290 850.000 ;
    END
  END la_output[8]
  PIN la_output[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1471.170 846.000 1471.450 850.000 ;
    END
  END la_output[90]
  PIN la_output[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 781.170 846.000 781.450 850.000 ;
    END
  END la_output[91]
  PIN la_output[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1473.010 846.000 1473.290 850.000 ;
    END
  END la_output[92]
  PIN la_output[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 779.330 846.000 779.610 850.000 ;
    END
  END la_output[93]
  PIN la_output[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1474.850 846.000 1475.130 850.000 ;
    END
  END la_output[94]
  PIN la_output[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 777.490 846.000 777.770 850.000 ;
    END
  END la_output[95]
  PIN la_output[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1476.690 846.000 1476.970 850.000 ;
    END
  END la_output[96]
  PIN la_output[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 775.650 846.000 775.930 850.000 ;
    END
  END la_output[97]
  PIN la_output[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1478.530 846.000 1478.810 850.000 ;
    END
  END la_output[98]
  PIN la_output[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 773.810 846.000 774.090 850.000 ;
    END
  END la_output[99]
  PIN la_output[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1480.370 846.000 1480.650 850.000 ;
    END
  END la_output[9]
  PIN mask_rev[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2146.450 0.000 2146.730 4.000 ;
    END
  END mask_rev[0]
  PIN mask_rev[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2144.610 0.000 2144.890 4.000 ;
    END
  END mask_rev[10]
  PIN mask_rev[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2146.000 5.480 2150.000 6.080 ;
    END
  END mask_rev[11]
  PIN mask_rev[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2142.770 0.000 2143.050 4.000 ;
    END
  END mask_rev[12]
  PIN mask_rev[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2146.000 8.200 2150.000 8.800 ;
    END
  END mask_rev[13]
  PIN mask_rev[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2140.930 0.000 2141.210 4.000 ;
    END
  END mask_rev[14]
  PIN mask_rev[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2139.090 0.000 2139.370 4.000 ;
    END
  END mask_rev[15]
  PIN mask_rev[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2146.000 10.920 2150.000 11.520 ;
    END
  END mask_rev[16]
  PIN mask_rev[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2137.250 0.000 2137.530 4.000 ;
    END
  END mask_rev[17]
  PIN mask_rev[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2146.000 13.640 2150.000 14.240 ;
    END
  END mask_rev[18]
  PIN mask_rev[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2135.410 0.000 2135.690 4.000 ;
    END
  END mask_rev[19]
  PIN mask_rev[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2133.570 0.000 2133.850 4.000 ;
    END
  END mask_rev[1]
  PIN mask_rev[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2146.000 16.360 2150.000 16.960 ;
    END
  END mask_rev[20]
  PIN mask_rev[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2131.730 0.000 2132.010 4.000 ;
    END
  END mask_rev[21]
  PIN mask_rev[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2146.000 19.080 2150.000 19.680 ;
    END
  END mask_rev[22]
  PIN mask_rev[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2129.890 0.000 2130.170 4.000 ;
    END
  END mask_rev[23]
  PIN mask_rev[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2128.050 0.000 2128.330 4.000 ;
    END
  END mask_rev[24]
  PIN mask_rev[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2146.000 21.800 2150.000 22.400 ;
    END
  END mask_rev[25]
  PIN mask_rev[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2126.210 0.000 2126.490 4.000 ;
    END
  END mask_rev[26]
  PIN mask_rev[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2146.000 24.520 2150.000 25.120 ;
    END
  END mask_rev[27]
  PIN mask_rev[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2124.370 0.000 2124.650 4.000 ;
    END
  END mask_rev[28]
  PIN mask_rev[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2122.530 0.000 2122.810 4.000 ;
    END
  END mask_rev[29]
  PIN mask_rev[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2146.000 27.240 2150.000 27.840 ;
    END
  END mask_rev[2]
  PIN mask_rev[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2120.690 0.000 2120.970 4.000 ;
    END
  END mask_rev[30]
  PIN mask_rev[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2146.000 29.960 2150.000 30.560 ;
    END
  END mask_rev[31]
  PIN mask_rev[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2118.850 0.000 2119.130 4.000 ;
    END
  END mask_rev[3]
  PIN mask_rev[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2117.010 0.000 2117.290 4.000 ;
    END
  END mask_rev[4]
  PIN mask_rev[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2146.000 32.680 2150.000 33.280 ;
    END
  END mask_rev[5]
  PIN mask_rev[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2115.170 0.000 2115.450 4.000 ;
    END
  END mask_rev[6]
  PIN mask_rev[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2146.000 35.400 2150.000 36.000 ;
    END
  END mask_rev[7]
  PIN mask_rev[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2113.330 0.000 2113.610 4.000 ;
    END
  END mask_rev[8]
  PIN mask_rev[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2111.490 0.000 2111.770 4.000 ;
    END
  END mask_rev[9]
  PIN mgmt_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END mgmt_addr[0]
  PIN mgmt_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END mgmt_addr[1]
  PIN mgmt_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END mgmt_addr[2]
  PIN mgmt_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END mgmt_addr[3]
  PIN mgmt_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END mgmt_addr[4]
  PIN mgmt_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END mgmt_addr[5]
  PIN mgmt_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END mgmt_addr[6]
  PIN mgmt_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END mgmt_addr[7]
  PIN mgmt_addr_ro[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END mgmt_addr_ro[0]
  PIN mgmt_addr_ro[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END mgmt_addr_ro[1]
  PIN mgmt_addr_ro[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END mgmt_addr_ro[2]
  PIN mgmt_addr_ro[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END mgmt_addr_ro[3]
  PIN mgmt_addr_ro[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END mgmt_addr_ro[4]
  PIN mgmt_addr_ro[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END mgmt_addr_ro[5]
  PIN mgmt_addr_ro[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END mgmt_addr_ro[6]
  PIN mgmt_addr_ro[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END mgmt_addr_ro[7]
  PIN mgmt_ena[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END mgmt_ena[0]
  PIN mgmt_ena[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END mgmt_ena[1]
  PIN mgmt_ena_ro
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END mgmt_ena_ro
  PIN mgmt_in_data[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2146.000 340.040 2150.000 340.640 ;
    END
  END mgmt_in_data[0]
  PIN mgmt_in_data[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END mgmt_in_data[10]
  PIN mgmt_in_data[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END mgmt_in_data[11]
  PIN mgmt_in_data[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END mgmt_in_data[12]
  PIN mgmt_in_data[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END mgmt_in_data[13]
  PIN mgmt_in_data[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END mgmt_in_data[14]
  PIN mgmt_in_data[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END mgmt_in_data[15]
  PIN mgmt_in_data[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END mgmt_in_data[16]
  PIN mgmt_in_data[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END mgmt_in_data[17]
  PIN mgmt_in_data[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END mgmt_in_data[18]
  PIN mgmt_in_data[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END mgmt_in_data[19]
  PIN mgmt_in_data[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2146.000 563.080 2150.000 563.680 ;
    END
  END mgmt_in_data[1]
  PIN mgmt_in_data[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END mgmt_in_data[20]
  PIN mgmt_in_data[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END mgmt_in_data[21]
  PIN mgmt_in_data[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END mgmt_in_data[22]
  PIN mgmt_in_data[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END mgmt_in_data[23]
  PIN mgmt_in_data[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END mgmt_in_data[24]
  PIN mgmt_in_data[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END mgmt_in_data[25]
  PIN mgmt_in_data[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END mgmt_in_data[26]
  PIN mgmt_in_data[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END mgmt_in_data[27]
  PIN mgmt_in_data[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END mgmt_in_data[28]
  PIN mgmt_in_data[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END mgmt_in_data[29]
  PIN mgmt_in_data[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END mgmt_in_data[2]
  PIN mgmt_in_data[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END mgmt_in_data[30]
  PIN mgmt_in_data[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END mgmt_in_data[31]
  PIN mgmt_in_data[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END mgmt_in_data[32]
  PIN mgmt_in_data[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END mgmt_in_data[33]
  PIN mgmt_in_data[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END mgmt_in_data[34]
  PIN mgmt_in_data[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END mgmt_in_data[35]
  PIN mgmt_in_data[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END mgmt_in_data[36]
  PIN mgmt_in_data[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END mgmt_in_data[37]
  PIN mgmt_in_data[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END mgmt_in_data[3]
  PIN mgmt_in_data[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END mgmt_in_data[4]
  PIN mgmt_in_data[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END mgmt_in_data[5]
  PIN mgmt_in_data[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END mgmt_in_data[6]
  PIN mgmt_in_data[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END mgmt_in_data[7]
  PIN mgmt_in_data[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END mgmt_in_data[8]
  PIN mgmt_in_data[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END mgmt_in_data[9]
  PIN mgmt_out_data[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END mgmt_out_data[0]
  PIN mgmt_out_data[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2146.450 846.000 2146.730 850.000 ;
    END
  END mgmt_out_data[10]
  PIN mgmt_out_data[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2144.610 846.000 2144.890 850.000 ;
    END
  END mgmt_out_data[11]
  PIN mgmt_out_data[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2146.000 843.240 2150.000 843.840 ;
    END
  END mgmt_out_data[12]
  PIN mgmt_out_data[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2142.770 846.000 2143.050 850.000 ;
    END
  END mgmt_out_data[13]
  PIN mgmt_out_data[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2140.930 846.000 2141.210 850.000 ;
    END
  END mgmt_out_data[14]
  PIN mgmt_out_data[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1675.410 846.000 1675.690 850.000 ;
    END
  END mgmt_out_data[15]
  PIN mgmt_out_data[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1482.210 846.000 1482.490 850.000 ;
    END
  END mgmt_out_data[16]
  PIN mgmt_out_data[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 771.970 846.000 772.250 850.000 ;
    END
  END mgmt_out_data[17]
  PIN mgmt_out_data[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 696.530 846.000 696.810 850.000 ;
    END
  END mgmt_out_data[18]
  PIN mgmt_out_data[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 444.450 846.000 444.730 850.000 ;
    END
  END mgmt_out_data[19]
  PIN mgmt_out_data[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END mgmt_out_data[1]
  PIN mgmt_out_data[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 186.850 846.000 187.130 850.000 ;
    END
  END mgmt_out_data[20]
  PIN mgmt_out_data[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 846.000 3.130 850.000 ;
    END
  END mgmt_out_data[21]
  PIN mgmt_out_data[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4.690 846.000 4.970 850.000 ;
    END
  END mgmt_out_data[22]
  PIN mgmt_out_data[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END mgmt_out_data[23]
  PIN mgmt_out_data[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.530 846.000 6.810 850.000 ;
    END
  END mgmt_out_data[24]
  PIN mgmt_out_data[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 8.370 846.000 8.650 850.000 ;
    END
  END mgmt_out_data[25]
  PIN mgmt_out_data[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 840.520 4.000 841.120 ;
    END
  END mgmt_out_data[26]
  PIN mgmt_out_data[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 10.210 846.000 10.490 850.000 ;
    END
  END mgmt_out_data[27]
  PIN mgmt_out_data[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 837.800 4.000 838.400 ;
    END
  END mgmt_out_data[28]
  PIN mgmt_out_data[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.050 846.000 12.330 850.000 ;
    END
  END mgmt_out_data[29]
  PIN mgmt_out_data[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2146.000 786.120 2150.000 786.720 ;
    END
  END mgmt_out_data[2]
  PIN mgmt_out_data[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.890 846.000 14.170 850.000 ;
    END
  END mgmt_out_data[30]
  PIN mgmt_out_data[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 835.080 4.000 835.680 ;
    END
  END mgmt_out_data[31]
  PIN mgmt_out_data[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.730 846.000 16.010 850.000 ;
    END
  END mgmt_out_data[32]
  PIN mgmt_out_data[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 832.360 4.000 832.960 ;
    END
  END mgmt_out_data[33]
  PIN mgmt_out_data[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.570 846.000 17.850 850.000 ;
    END
  END mgmt_out_data[34]
  PIN mgmt_out_data[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.410 846.000 19.690 850.000 ;
    END
  END mgmt_out_data[35]
  PIN mgmt_out_data[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END mgmt_out_data[36]
  PIN mgmt_out_data[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 745.320 4.000 745.920 ;
    END
  END mgmt_out_data[37]
  PIN mgmt_out_data[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2146.000 840.520 2150.000 841.120 ;
    END
  END mgmt_out_data[3]
  PIN mgmt_out_data[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2139.090 846.000 2139.370 850.000 ;
    END
  END mgmt_out_data[4]
  PIN mgmt_out_data[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2146.000 837.800 2150.000 838.400 ;
    END
  END mgmt_out_data[5]
  PIN mgmt_out_data[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2137.250 846.000 2137.530 850.000 ;
    END
  END mgmt_out_data[6]
  PIN mgmt_out_data[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2135.410 846.000 2135.690 850.000 ;
    END
  END mgmt_out_data[7]
  PIN mgmt_out_data[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2146.000 835.080 2150.000 835.680 ;
    END
  END mgmt_out_data[8]
  PIN mgmt_out_data[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2133.570 846.000 2133.850 850.000 ;
    END
  END mgmt_out_data[9]
  PIN mgmt_rdata[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END mgmt_rdata[0]
  PIN mgmt_rdata[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END mgmt_rdata[10]
  PIN mgmt_rdata[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END mgmt_rdata[11]
  PIN mgmt_rdata[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END mgmt_rdata[12]
  PIN mgmt_rdata[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END mgmt_rdata[13]
  PIN mgmt_rdata[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END mgmt_rdata[14]
  PIN mgmt_rdata[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END mgmt_rdata[15]
  PIN mgmt_rdata[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END mgmt_rdata[16]
  PIN mgmt_rdata[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END mgmt_rdata[17]
  PIN mgmt_rdata[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END mgmt_rdata[18]
  PIN mgmt_rdata[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END mgmt_rdata[19]
  PIN mgmt_rdata[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END mgmt_rdata[1]
  PIN mgmt_rdata[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END mgmt_rdata[20]
  PIN mgmt_rdata[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END mgmt_rdata[21]
  PIN mgmt_rdata[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END mgmt_rdata[22]
  PIN mgmt_rdata[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END mgmt_rdata[23]
  PIN mgmt_rdata[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END mgmt_rdata[24]
  PIN mgmt_rdata[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END mgmt_rdata[25]
  PIN mgmt_rdata[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END mgmt_rdata[26]
  PIN mgmt_rdata[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END mgmt_rdata[27]
  PIN mgmt_rdata[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END mgmt_rdata[28]
  PIN mgmt_rdata[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END mgmt_rdata[29]
  PIN mgmt_rdata[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END mgmt_rdata[2]
  PIN mgmt_rdata[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END mgmt_rdata[30]
  PIN mgmt_rdata[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END mgmt_rdata[31]
  PIN mgmt_rdata[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END mgmt_rdata[32]
  PIN mgmt_rdata[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END mgmt_rdata[33]
  PIN mgmt_rdata[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END mgmt_rdata[34]
  PIN mgmt_rdata[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END mgmt_rdata[35]
  PIN mgmt_rdata[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END mgmt_rdata[36]
  PIN mgmt_rdata[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END mgmt_rdata[37]
  PIN mgmt_rdata[38]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END mgmt_rdata[38]
  PIN mgmt_rdata[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END mgmt_rdata[39]
  PIN mgmt_rdata[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END mgmt_rdata[3]
  PIN mgmt_rdata[40]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END mgmt_rdata[40]
  PIN mgmt_rdata[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END mgmt_rdata[41]
  PIN mgmt_rdata[42]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END mgmt_rdata[42]
  PIN mgmt_rdata[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END mgmt_rdata[43]
  PIN mgmt_rdata[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END mgmt_rdata[44]
  PIN mgmt_rdata[45]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END mgmt_rdata[45]
  PIN mgmt_rdata[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END mgmt_rdata[46]
  PIN mgmt_rdata[47]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END mgmt_rdata[47]
  PIN mgmt_rdata[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END mgmt_rdata[48]
  PIN mgmt_rdata[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END mgmt_rdata[49]
  PIN mgmt_rdata[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END mgmt_rdata[4]
  PIN mgmt_rdata[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END mgmt_rdata[50]
  PIN mgmt_rdata[51]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END mgmt_rdata[51]
  PIN mgmt_rdata[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END mgmt_rdata[52]
  PIN mgmt_rdata[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END mgmt_rdata[53]
  PIN mgmt_rdata[54]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END mgmt_rdata[54]
  PIN mgmt_rdata[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END mgmt_rdata[55]
  PIN mgmt_rdata[56]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END mgmt_rdata[56]
  PIN mgmt_rdata[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END mgmt_rdata[57]
  PIN mgmt_rdata[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END mgmt_rdata[58]
  PIN mgmt_rdata[59]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END mgmt_rdata[59]
  PIN mgmt_rdata[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END mgmt_rdata[5]
  PIN mgmt_rdata[60]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END mgmt_rdata[60]
  PIN mgmt_rdata[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END mgmt_rdata[61]
  PIN mgmt_rdata[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END mgmt_rdata[62]
  PIN mgmt_rdata[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END mgmt_rdata[63]
  PIN mgmt_rdata[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END mgmt_rdata[6]
  PIN mgmt_rdata[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END mgmt_rdata[7]
  PIN mgmt_rdata[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END mgmt_rdata[8]
  PIN mgmt_rdata[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END mgmt_rdata[9]
  PIN mgmt_rdata_ro[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END mgmt_rdata_ro[0]
  PIN mgmt_rdata_ro[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END mgmt_rdata_ro[10]
  PIN mgmt_rdata_ro[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END mgmt_rdata_ro[11]
  PIN mgmt_rdata_ro[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END mgmt_rdata_ro[12]
  PIN mgmt_rdata_ro[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END mgmt_rdata_ro[13]
  PIN mgmt_rdata_ro[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END mgmt_rdata_ro[14]
  PIN mgmt_rdata_ro[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END mgmt_rdata_ro[15]
  PIN mgmt_rdata_ro[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END mgmt_rdata_ro[16]
  PIN mgmt_rdata_ro[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END mgmt_rdata_ro[17]
  PIN mgmt_rdata_ro[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END mgmt_rdata_ro[18]
  PIN mgmt_rdata_ro[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END mgmt_rdata_ro[19]
  PIN mgmt_rdata_ro[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END mgmt_rdata_ro[1]
  PIN mgmt_rdata_ro[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END mgmt_rdata_ro[20]
  PIN mgmt_rdata_ro[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END mgmt_rdata_ro[21]
  PIN mgmt_rdata_ro[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END mgmt_rdata_ro[22]
  PIN mgmt_rdata_ro[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END mgmt_rdata_ro[23]
  PIN mgmt_rdata_ro[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END mgmt_rdata_ro[24]
  PIN mgmt_rdata_ro[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END mgmt_rdata_ro[25]
  PIN mgmt_rdata_ro[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END mgmt_rdata_ro[26]
  PIN mgmt_rdata_ro[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END mgmt_rdata_ro[27]
  PIN mgmt_rdata_ro[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END mgmt_rdata_ro[28]
  PIN mgmt_rdata_ro[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END mgmt_rdata_ro[29]
  PIN mgmt_rdata_ro[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END mgmt_rdata_ro[2]
  PIN mgmt_rdata_ro[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END mgmt_rdata_ro[30]
  PIN mgmt_rdata_ro[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END mgmt_rdata_ro[31]
  PIN mgmt_rdata_ro[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END mgmt_rdata_ro[3]
  PIN mgmt_rdata_ro[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END mgmt_rdata_ro[4]
  PIN mgmt_rdata_ro[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END mgmt_rdata_ro[5]
  PIN mgmt_rdata_ro[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END mgmt_rdata_ro[6]
  PIN mgmt_rdata_ro[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END mgmt_rdata_ro[7]
  PIN mgmt_rdata_ro[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END mgmt_rdata_ro[8]
  PIN mgmt_rdata_ro[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END mgmt_rdata_ro[9]
  PIN mgmt_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END mgmt_wdata[0]
  PIN mgmt_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END mgmt_wdata[10]
  PIN mgmt_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END mgmt_wdata[11]
  PIN mgmt_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END mgmt_wdata[12]
  PIN mgmt_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END mgmt_wdata[13]
  PIN mgmt_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END mgmt_wdata[14]
  PIN mgmt_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END mgmt_wdata[15]
  PIN mgmt_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END mgmt_wdata[16]
  PIN mgmt_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END mgmt_wdata[17]
  PIN mgmt_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END mgmt_wdata[18]
  PIN mgmt_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END mgmt_wdata[19]
  PIN mgmt_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END mgmt_wdata[1]
  PIN mgmt_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END mgmt_wdata[20]
  PIN mgmt_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END mgmt_wdata[21]
  PIN mgmt_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END mgmt_wdata[22]
  PIN mgmt_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END mgmt_wdata[23]
  PIN mgmt_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END mgmt_wdata[24]
  PIN mgmt_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END mgmt_wdata[25]
  PIN mgmt_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END mgmt_wdata[26]
  PIN mgmt_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END mgmt_wdata[27]
  PIN mgmt_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END mgmt_wdata[28]
  PIN mgmt_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END mgmt_wdata[29]
  PIN mgmt_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END mgmt_wdata[2]
  PIN mgmt_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END mgmt_wdata[30]
  PIN mgmt_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END mgmt_wdata[31]
  PIN mgmt_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END mgmt_wdata[3]
  PIN mgmt_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END mgmt_wdata[4]
  PIN mgmt_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END mgmt_wdata[5]
  PIN mgmt_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END mgmt_wdata[6]
  PIN mgmt_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END mgmt_wdata[7]
  PIN mgmt_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END mgmt_wdata[8]
  PIN mgmt_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END mgmt_wdata[9]
  PIN mgmt_wen[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END mgmt_wen[0]
  PIN mgmt_wen[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END mgmt_wen[1]
  PIN mgmt_wen_mask[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END mgmt_wen_mask[0]
  PIN mgmt_wen_mask[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END mgmt_wen_mask[1]
  PIN mgmt_wen_mask[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END mgmt_wen_mask[2]
  PIN mgmt_wen_mask[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END mgmt_wen_mask[3]
  PIN mgmt_wen_mask[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END mgmt_wen_mask[4]
  PIN mgmt_wen_mask[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END mgmt_wen_mask[5]
  PIN mgmt_wen_mask[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 4.000 ;
    END
  END mgmt_wen_mask[6]
  PIN mgmt_wen_mask[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END mgmt_wen_mask[7]
  PIN mprj2_vcc_pwrgood
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 770.130 846.000 770.410 850.000 ;
    END
  END mprj2_vcc_pwrgood
  PIN mprj2_vdd_pwrgood
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1484.050 846.000 1484.330 850.000 ;
    END
  END mprj2_vdd_pwrgood
  PIN mprj_ack_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.250 846.000 21.530 850.000 ;
    END
  END mprj_ack_i
  PIN mprj_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 768.290 846.000 768.570 850.000 ;
    END
  END mprj_adr_o[0]
  PIN mprj_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1485.890 846.000 1486.170 850.000 ;
    END
  END mprj_adr_o[10]
  PIN mprj_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 766.450 846.000 766.730 850.000 ;
    END
  END mprj_adr_o[11]
  PIN mprj_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1487.730 846.000 1488.010 850.000 ;
    END
  END mprj_adr_o[12]
  PIN mprj_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 764.610 846.000 764.890 850.000 ;
    END
  END mprj_adr_o[13]
  PIN mprj_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1489.570 846.000 1489.850 850.000 ;
    END
  END mprj_adr_o[14]
  PIN mprj_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 762.770 846.000 763.050 850.000 ;
    END
  END mprj_adr_o[15]
  PIN mprj_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1491.410 846.000 1491.690 850.000 ;
    END
  END mprj_adr_o[16]
  PIN mprj_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 760.930 846.000 761.210 850.000 ;
    END
  END mprj_adr_o[17]
  PIN mprj_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1493.250 846.000 1493.530 850.000 ;
    END
  END mprj_adr_o[18]
  PIN mprj_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 759.090 846.000 759.370 850.000 ;
    END
  END mprj_adr_o[19]
  PIN mprj_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1495.090 846.000 1495.370 850.000 ;
    END
  END mprj_adr_o[1]
  PIN mprj_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 757.250 846.000 757.530 850.000 ;
    END
  END mprj_adr_o[20]
  PIN mprj_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1496.930 846.000 1497.210 850.000 ;
    END
  END mprj_adr_o[21]
  PIN mprj_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 755.410 846.000 755.690 850.000 ;
    END
  END mprj_adr_o[22]
  PIN mprj_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1498.770 846.000 1499.050 850.000 ;
    END
  END mprj_adr_o[23]
  PIN mprj_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 753.570 846.000 753.850 850.000 ;
    END
  END mprj_adr_o[24]
  PIN mprj_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1500.610 846.000 1500.890 850.000 ;
    END
  END mprj_adr_o[25]
  PIN mprj_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 751.730 846.000 752.010 850.000 ;
    END
  END mprj_adr_o[26]
  PIN mprj_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1502.450 846.000 1502.730 850.000 ;
    END
  END mprj_adr_o[27]
  PIN mprj_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 749.890 846.000 750.170 850.000 ;
    END
  END mprj_adr_o[28]
  PIN mprj_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1504.290 846.000 1504.570 850.000 ;
    END
  END mprj_adr_o[29]
  PIN mprj_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 748.050 846.000 748.330 850.000 ;
    END
  END mprj_adr_o[2]
  PIN mprj_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1506.130 846.000 1506.410 850.000 ;
    END
  END mprj_adr_o[30]
  PIN mprj_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 746.210 846.000 746.490 850.000 ;
    END
  END mprj_adr_o[31]
  PIN mprj_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1507.970 846.000 1508.250 850.000 ;
    END
  END mprj_adr_o[3]
  PIN mprj_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 744.370 846.000 744.650 850.000 ;
    END
  END mprj_adr_o[4]
  PIN mprj_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1509.810 846.000 1510.090 850.000 ;
    END
  END mprj_adr_o[5]
  PIN mprj_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 742.530 846.000 742.810 850.000 ;
    END
  END mprj_adr_o[6]
  PIN mprj_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1511.650 846.000 1511.930 850.000 ;
    END
  END mprj_adr_o[7]
  PIN mprj_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 740.690 846.000 740.970 850.000 ;
    END
  END mprj_adr_o[8]
  PIN mprj_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1513.490 846.000 1513.770 850.000 ;
    END
  END mprj_adr_o[9]
  PIN mprj_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 738.850 846.000 739.130 850.000 ;
    END
  END mprj_cyc_o
  PIN mprj_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.920 4.000 827.520 ;
    END
  END mprj_dat_i[0]
  PIN mprj_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 846.000 23.370 850.000 ;
    END
  END mprj_dat_i[10]
  PIN mprj_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.930 846.000 25.210 850.000 ;
    END
  END mprj_dat_i[11]
  PIN mprj_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 824.200 4.000 824.800 ;
    END
  END mprj_dat_i[12]
  PIN mprj_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 846.000 27.050 850.000 ;
    END
  END mprj_dat_i[13]
  PIN mprj_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 821.480 4.000 822.080 ;
    END
  END mprj_dat_i[14]
  PIN mprj_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 846.000 28.890 850.000 ;
    END
  END mprj_dat_i[15]
  PIN mprj_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.450 846.000 30.730 850.000 ;
    END
  END mprj_dat_i[16]
  PIN mprj_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 818.760 4.000 819.360 ;
    END
  END mprj_dat_i[17]
  PIN mprj_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.290 846.000 32.570 850.000 ;
    END
  END mprj_dat_i[18]
  PIN mprj_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 816.040 4.000 816.640 ;
    END
  END mprj_dat_i[19]
  PIN mprj_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.130 846.000 34.410 850.000 ;
    END
  END mprj_dat_i[1]
  PIN mprj_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.970 846.000 36.250 850.000 ;
    END
  END mprj_dat_i[20]
  PIN mprj_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 813.320 4.000 813.920 ;
    END
  END mprj_dat_i[21]
  PIN mprj_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.810 846.000 38.090 850.000 ;
    END
  END mprj_dat_i[22]
  PIN mprj_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 810.600 4.000 811.200 ;
    END
  END mprj_dat_i[23]
  PIN mprj_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.650 846.000 39.930 850.000 ;
    END
  END mprj_dat_i[24]
  PIN mprj_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.490 846.000 41.770 850.000 ;
    END
  END mprj_dat_i[25]
  PIN mprj_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.880 4.000 808.480 ;
    END
  END mprj_dat_i[26]
  PIN mprj_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.330 846.000 43.610 850.000 ;
    END
  END mprj_dat_i[27]
  PIN mprj_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.160 4.000 805.760 ;
    END
  END mprj_dat_i[28]
  PIN mprj_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.170 846.000 45.450 850.000 ;
    END
  END mprj_dat_i[29]
  PIN mprj_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 846.000 47.290 850.000 ;
    END
  END mprj_dat_i[2]
  PIN mprj_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.440 4.000 803.040 ;
    END
  END mprj_dat_i[30]
  PIN mprj_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 846.000 49.130 850.000 ;
    END
  END mprj_dat_i[31]
  PIN mprj_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.720 4.000 800.320 ;
    END
  END mprj_dat_i[3]
  PIN mprj_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 846.000 50.970 850.000 ;
    END
  END mprj_dat_i[4]
  PIN mprj_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 846.000 52.810 850.000 ;
    END
  END mprj_dat_i[5]
  PIN mprj_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.000 4.000 797.600 ;
    END
  END mprj_dat_i[6]
  PIN mprj_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.370 846.000 54.650 850.000 ;
    END
  END mprj_dat_i[7]
  PIN mprj_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 794.280 4.000 794.880 ;
    END
  END mprj_dat_i[8]
  PIN mprj_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.210 846.000 56.490 850.000 ;
    END
  END mprj_dat_i[9]
  PIN mprj_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1515.330 846.000 1515.610 850.000 ;
    END
  END mprj_dat_o[0]
  PIN mprj_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 737.010 846.000 737.290 850.000 ;
    END
  END mprj_dat_o[10]
  PIN mprj_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1517.170 846.000 1517.450 850.000 ;
    END
  END mprj_dat_o[11]
  PIN mprj_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 735.170 846.000 735.450 850.000 ;
    END
  END mprj_dat_o[12]
  PIN mprj_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1519.010 846.000 1519.290 850.000 ;
    END
  END mprj_dat_o[13]
  PIN mprj_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 733.330 846.000 733.610 850.000 ;
    END
  END mprj_dat_o[14]
  PIN mprj_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1520.850 846.000 1521.130 850.000 ;
    END
  END mprj_dat_o[15]
  PIN mprj_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 731.490 846.000 731.770 850.000 ;
    END
  END mprj_dat_o[16]
  PIN mprj_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1522.690 846.000 1522.970 850.000 ;
    END
  END mprj_dat_o[17]
  PIN mprj_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 729.650 846.000 729.930 850.000 ;
    END
  END mprj_dat_o[18]
  PIN mprj_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1524.530 846.000 1524.810 850.000 ;
    END
  END mprj_dat_o[19]
  PIN mprj_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 727.810 846.000 728.090 850.000 ;
    END
  END mprj_dat_o[1]
  PIN mprj_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1526.370 846.000 1526.650 850.000 ;
    END
  END mprj_dat_o[20]
  PIN mprj_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 725.970 846.000 726.250 850.000 ;
    END
  END mprj_dat_o[21]
  PIN mprj_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1528.210 846.000 1528.490 850.000 ;
    END
  END mprj_dat_o[22]
  PIN mprj_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 724.130 846.000 724.410 850.000 ;
    END
  END mprj_dat_o[23]
  PIN mprj_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1530.050 846.000 1530.330 850.000 ;
    END
  END mprj_dat_o[24]
  PIN mprj_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 722.290 846.000 722.570 850.000 ;
    END
  END mprj_dat_o[25]
  PIN mprj_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1531.890 846.000 1532.170 850.000 ;
    END
  END mprj_dat_o[26]
  PIN mprj_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 720.450 846.000 720.730 850.000 ;
    END
  END mprj_dat_o[27]
  PIN mprj_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1533.730 846.000 1534.010 850.000 ;
    END
  END mprj_dat_o[28]
  PIN mprj_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 718.610 846.000 718.890 850.000 ;
    END
  END mprj_dat_o[29]
  PIN mprj_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1535.570 846.000 1535.850 850.000 ;
    END
  END mprj_dat_o[2]
  PIN mprj_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 716.770 846.000 717.050 850.000 ;
    END
  END mprj_dat_o[30]
  PIN mprj_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1537.410 846.000 1537.690 850.000 ;
    END
  END mprj_dat_o[31]
  PIN mprj_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 714.930 846.000 715.210 850.000 ;
    END
  END mprj_dat_o[3]
  PIN mprj_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1539.250 846.000 1539.530 850.000 ;
    END
  END mprj_dat_o[4]
  PIN mprj_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 713.090 846.000 713.370 850.000 ;
    END
  END mprj_dat_o[5]
  PIN mprj_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1541.090 846.000 1541.370 850.000 ;
    END
  END mprj_dat_o[6]
  PIN mprj_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 711.250 846.000 711.530 850.000 ;
    END
  END mprj_dat_o[7]
  PIN mprj_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1542.930 846.000 1543.210 850.000 ;
    END
  END mprj_dat_o[8]
  PIN mprj_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 709.410 846.000 709.690 850.000 ;
    END
  END mprj_dat_o[9]
  PIN mprj_io_loader_clock
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2146.000 448.840 2150.000 449.440 ;
    END
  END mprj_io_loader_clock
  PIN mprj_io_loader_data
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2146.000 331.880 2150.000 332.480 ;
    END
  END mprj_io_loader_data
  PIN mprj_io_loader_resetn
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2146.000 481.480 2150.000 482.080 ;
    END
  END mprj_io_loader_resetn
  PIN mprj_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1544.770 846.000 1545.050 850.000 ;
    END
  END mprj_sel_o[0]
  PIN mprj_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 707.570 846.000 707.850 850.000 ;
    END
  END mprj_sel_o[1]
  PIN mprj_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1546.610 846.000 1546.890 850.000 ;
    END
  END mprj_sel_o[2]
  PIN mprj_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 705.730 846.000 706.010 850.000 ;
    END
  END mprj_sel_o[3]
  PIN mprj_stb_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1548.450 846.000 1548.730 850.000 ;
    END
  END mprj_stb_o
  PIN mprj_vcc_pwrgood
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 703.890 846.000 704.170 850.000 ;
    END
  END mprj_vcc_pwrgood
  PIN mprj_vdd_pwrgood
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1550.290 846.000 1550.570 850.000 ;
    END
  END mprj_vdd_pwrgood
  PIN mprj_we_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 702.050 846.000 702.330 850.000 ;
    END
  END mprj_we_o
  PIN porb
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2146.000 108.840 2150.000 109.440 ;
    END
  END porb
  PIN pwr_ctrl_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END pwr_ctrl_out[0]
  PIN pwr_ctrl_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END pwr_ctrl_out[1]
  PIN pwr_ctrl_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END pwr_ctrl_out[2]
  PIN pwr_ctrl_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END pwr_ctrl_out[3]
  PIN resetb
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END resetb
  PIN sdo_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2146.000 560.360 2150.000 560.960 ;
    END
  END sdo_out
  PIN sdo_outenb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2146.000 565.800 2150.000 566.400 ;
    END
  END sdo_outenb
  PIN user_clk
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1552.130 846.000 1552.410 850.000 ;
    END
  END user_clk
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 5.520 837.520 2144.060 838.000 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 5.520 834.800 2144.060 835.280 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2144.060 849.915 ;
      LAYER met1 ;
        RECT 2.830 838.280 2146.750 849.960 ;
        RECT 2.830 837.240 5.240 838.280 ;
        RECT 2144.340 837.240 2146.750 838.280 ;
        RECT 2.830 835.560 2146.750 837.240 ;
        RECT 2.830 834.520 5.240 835.560 ;
        RECT 2144.340 834.520 2146.750 835.560 ;
        RECT 2.830 3.100 2146.750 834.520 ;
      LAYER met2 ;
        RECT 3.410 845.720 4.410 849.990 ;
        RECT 5.250 845.720 6.250 849.990 ;
        RECT 7.090 845.720 8.090 849.990 ;
        RECT 8.930 845.720 9.930 849.990 ;
        RECT 10.770 845.720 11.770 849.990 ;
        RECT 12.610 845.720 13.610 849.990 ;
        RECT 14.450 845.720 15.450 849.990 ;
        RECT 16.290 845.720 17.290 849.990 ;
        RECT 18.130 845.720 19.130 849.990 ;
        RECT 19.970 845.720 20.970 849.990 ;
        RECT 21.810 845.720 22.810 849.990 ;
        RECT 23.650 845.720 24.650 849.990 ;
        RECT 25.490 845.720 26.490 849.990 ;
        RECT 27.330 845.720 28.330 849.990 ;
        RECT 29.170 845.720 30.170 849.990 ;
        RECT 31.010 845.720 32.010 849.990 ;
        RECT 32.850 845.720 33.850 849.990 ;
        RECT 34.690 845.720 35.690 849.990 ;
        RECT 36.530 845.720 37.530 849.990 ;
        RECT 38.370 845.720 39.370 849.990 ;
        RECT 40.210 845.720 41.210 849.990 ;
        RECT 42.050 845.720 43.050 849.990 ;
        RECT 43.890 845.720 44.890 849.990 ;
        RECT 45.730 845.720 46.730 849.990 ;
        RECT 47.570 845.720 48.570 849.990 ;
        RECT 49.410 845.720 50.410 849.990 ;
        RECT 51.250 845.720 52.250 849.990 ;
        RECT 53.090 845.720 54.090 849.990 ;
        RECT 54.930 845.720 55.930 849.990 ;
        RECT 56.770 845.720 186.570 849.990 ;
        RECT 187.410 845.720 444.170 849.990 ;
        RECT 445.010 845.720 571.130 849.990 ;
        RECT 571.970 845.720 696.250 849.990 ;
        RECT 697.090 845.720 701.770 849.990 ;
        RECT 702.610 845.720 703.610 849.990 ;
        RECT 704.450 845.720 705.450 849.990 ;
        RECT 706.290 845.720 707.290 849.990 ;
        RECT 708.130 845.720 709.130 849.990 ;
        RECT 709.970 845.720 710.970 849.990 ;
        RECT 711.810 845.720 712.810 849.990 ;
        RECT 713.650 845.720 714.650 849.990 ;
        RECT 715.490 845.720 716.490 849.990 ;
        RECT 717.330 845.720 718.330 849.990 ;
        RECT 719.170 845.720 720.170 849.990 ;
        RECT 721.010 845.720 722.010 849.990 ;
        RECT 722.850 845.720 723.850 849.990 ;
        RECT 724.690 845.720 725.690 849.990 ;
        RECT 726.530 845.720 727.530 849.990 ;
        RECT 728.370 845.720 729.370 849.990 ;
        RECT 730.210 845.720 731.210 849.990 ;
        RECT 732.050 845.720 733.050 849.990 ;
        RECT 733.890 845.720 734.890 849.990 ;
        RECT 735.730 845.720 736.730 849.990 ;
        RECT 737.570 845.720 738.570 849.990 ;
        RECT 739.410 845.720 740.410 849.990 ;
        RECT 741.250 845.720 742.250 849.990 ;
        RECT 743.090 845.720 744.090 849.990 ;
        RECT 744.930 845.720 745.930 849.990 ;
        RECT 746.770 845.720 747.770 849.990 ;
        RECT 748.610 845.720 749.610 849.990 ;
        RECT 750.450 845.720 751.450 849.990 ;
        RECT 752.290 845.720 753.290 849.990 ;
        RECT 754.130 845.720 755.130 849.990 ;
        RECT 755.970 845.720 756.970 849.990 ;
        RECT 757.810 845.720 758.810 849.990 ;
        RECT 759.650 845.720 760.650 849.990 ;
        RECT 761.490 845.720 762.490 849.990 ;
        RECT 763.330 845.720 764.330 849.990 ;
        RECT 765.170 845.720 766.170 849.990 ;
        RECT 767.010 845.720 768.010 849.990 ;
        RECT 768.850 845.720 769.850 849.990 ;
        RECT 770.690 845.720 771.690 849.990 ;
        RECT 772.530 845.720 773.530 849.990 ;
        RECT 774.370 845.720 775.370 849.990 ;
        RECT 776.210 845.720 777.210 849.990 ;
        RECT 778.050 845.720 779.050 849.990 ;
        RECT 779.890 845.720 780.890 849.990 ;
        RECT 781.730 845.720 782.730 849.990 ;
        RECT 783.570 845.720 784.570 849.990 ;
        RECT 785.410 845.720 786.410 849.990 ;
        RECT 787.250 845.720 788.250 849.990 ;
        RECT 789.090 845.720 790.090 849.990 ;
        RECT 790.930 845.720 791.930 849.990 ;
        RECT 792.770 845.720 793.770 849.990 ;
        RECT 794.610 845.720 795.610 849.990 ;
        RECT 796.450 845.720 797.450 849.990 ;
        RECT 798.290 845.720 799.290 849.990 ;
        RECT 800.130 845.720 801.130 849.990 ;
        RECT 801.970 845.720 802.970 849.990 ;
        RECT 803.810 845.720 804.810 849.990 ;
        RECT 805.650 845.720 806.650 849.990 ;
        RECT 807.490 845.720 808.490 849.990 ;
        RECT 809.330 845.720 810.330 849.990 ;
        RECT 811.170 845.720 812.170 849.990 ;
        RECT 813.010 845.720 814.010 849.990 ;
        RECT 814.850 845.720 815.850 849.990 ;
        RECT 816.690 845.720 817.690 849.990 ;
        RECT 818.530 845.720 819.530 849.990 ;
        RECT 820.370 845.720 821.370 849.990 ;
        RECT 822.210 845.720 823.210 849.990 ;
        RECT 824.050 845.720 825.050 849.990 ;
        RECT 825.890 845.720 826.890 849.990 ;
        RECT 827.730 845.720 828.730 849.990 ;
        RECT 829.570 845.720 830.570 849.990 ;
        RECT 831.410 845.720 832.410 849.990 ;
        RECT 833.250 845.720 834.250 849.990 ;
        RECT 835.090 845.720 836.090 849.990 ;
        RECT 836.930 845.720 837.930 849.990 ;
        RECT 838.770 845.720 839.770 849.990 ;
        RECT 840.610 845.720 841.610 849.990 ;
        RECT 842.450 845.720 843.450 849.990 ;
        RECT 844.290 845.720 845.290 849.990 ;
        RECT 846.130 845.720 847.130 849.990 ;
        RECT 847.970 845.720 848.970 849.990 ;
        RECT 849.810 845.720 850.810 849.990 ;
        RECT 851.650 845.720 852.650 849.990 ;
        RECT 853.490 845.720 854.490 849.990 ;
        RECT 855.330 845.720 856.330 849.990 ;
        RECT 857.170 845.720 858.170 849.990 ;
        RECT 859.010 845.720 860.010 849.990 ;
        RECT 860.850 845.720 861.850 849.990 ;
        RECT 862.690 845.720 863.690 849.990 ;
        RECT 864.530 845.720 865.530 849.990 ;
        RECT 866.370 845.720 867.370 849.990 ;
        RECT 868.210 845.720 869.210 849.990 ;
        RECT 870.050 845.720 871.050 849.990 ;
        RECT 871.890 845.720 872.890 849.990 ;
        RECT 873.730 845.720 874.730 849.990 ;
        RECT 875.570 845.720 876.570 849.990 ;
        RECT 877.410 845.720 878.410 849.990 ;
        RECT 879.250 845.720 880.250 849.990 ;
        RECT 881.090 845.720 882.090 849.990 ;
        RECT 882.930 845.720 883.930 849.990 ;
        RECT 884.770 845.720 885.770 849.990 ;
        RECT 886.610 845.720 887.610 849.990 ;
        RECT 888.450 845.720 889.450 849.990 ;
        RECT 890.290 845.720 891.290 849.990 ;
        RECT 892.130 845.720 893.130 849.990 ;
        RECT 893.970 845.720 894.970 849.990 ;
        RECT 895.810 845.720 896.810 849.990 ;
        RECT 897.650 845.720 898.650 849.990 ;
        RECT 899.490 845.720 900.490 849.990 ;
        RECT 901.330 845.720 902.330 849.990 ;
        RECT 903.170 845.720 904.170 849.990 ;
        RECT 905.010 845.720 906.010 849.990 ;
        RECT 906.850 845.720 907.850 849.990 ;
        RECT 908.690 845.720 909.690 849.990 ;
        RECT 910.530 845.720 911.530 849.990 ;
        RECT 912.370 845.720 913.370 849.990 ;
        RECT 914.210 845.720 915.210 849.990 ;
        RECT 916.050 845.720 917.050 849.990 ;
        RECT 917.890 845.720 918.890 849.990 ;
        RECT 919.730 845.720 920.730 849.990 ;
        RECT 921.570 845.720 922.570 849.990 ;
        RECT 923.410 845.720 924.410 849.990 ;
        RECT 925.250 845.720 926.250 849.990 ;
        RECT 927.090 845.720 928.090 849.990 ;
        RECT 928.930 845.720 929.930 849.990 ;
        RECT 930.770 845.720 931.770 849.990 ;
        RECT 932.610 845.720 933.610 849.990 ;
        RECT 934.450 845.720 935.450 849.990 ;
        RECT 936.290 845.720 937.290 849.990 ;
        RECT 938.130 845.720 939.130 849.990 ;
        RECT 939.970 845.720 940.970 849.990 ;
        RECT 941.810 845.720 942.810 849.990 ;
        RECT 943.650 845.720 944.650 849.990 ;
        RECT 945.490 845.720 946.490 849.990 ;
        RECT 947.330 845.720 948.330 849.990 ;
        RECT 949.170 845.720 950.170 849.990 ;
        RECT 951.010 845.720 952.010 849.990 ;
        RECT 952.850 845.720 953.850 849.990 ;
        RECT 954.690 845.720 955.690 849.990 ;
        RECT 956.530 845.720 957.530 849.990 ;
        RECT 958.370 845.720 959.370 849.990 ;
        RECT 960.210 845.720 961.210 849.990 ;
        RECT 962.050 845.720 963.050 849.990 ;
        RECT 963.890 845.720 964.890 849.990 ;
        RECT 965.730 845.720 966.730 849.990 ;
        RECT 967.570 845.720 968.570 849.990 ;
        RECT 969.410 845.720 970.410 849.990 ;
        RECT 971.250 845.720 972.250 849.990 ;
        RECT 973.090 845.720 974.090 849.990 ;
        RECT 974.930 845.720 975.930 849.990 ;
        RECT 976.770 845.720 977.770 849.990 ;
        RECT 978.610 845.720 979.610 849.990 ;
        RECT 980.450 845.720 981.450 849.990 ;
        RECT 982.290 845.720 983.290 849.990 ;
        RECT 984.130 845.720 985.130 849.990 ;
        RECT 985.970 845.720 986.970 849.990 ;
        RECT 987.810 845.720 988.810 849.990 ;
        RECT 989.650 845.720 990.650 849.990 ;
        RECT 991.490 845.720 992.490 849.990 ;
        RECT 993.330 845.720 994.330 849.990 ;
        RECT 995.170 845.720 996.170 849.990 ;
        RECT 997.010 845.720 998.010 849.990 ;
        RECT 998.850 845.720 999.850 849.990 ;
        RECT 1000.690 845.720 1001.690 849.990 ;
        RECT 1002.530 845.720 1003.530 849.990 ;
        RECT 1004.370 845.720 1005.370 849.990 ;
        RECT 1006.210 845.720 1007.210 849.990 ;
        RECT 1008.050 845.720 1009.050 849.990 ;
        RECT 1009.890 845.720 1010.890 849.990 ;
        RECT 1011.730 845.720 1012.730 849.990 ;
        RECT 1013.570 845.720 1014.570 849.990 ;
        RECT 1015.410 845.720 1016.410 849.990 ;
        RECT 1017.250 845.720 1018.250 849.990 ;
        RECT 1019.090 845.720 1020.090 849.990 ;
        RECT 1020.930 845.720 1021.930 849.990 ;
        RECT 1022.770 845.720 1023.770 849.990 ;
        RECT 1024.610 845.720 1025.610 849.990 ;
        RECT 1026.450 845.720 1027.450 849.990 ;
        RECT 1028.290 845.720 1029.290 849.990 ;
        RECT 1030.130 845.720 1031.130 849.990 ;
        RECT 1031.970 845.720 1032.970 849.990 ;
        RECT 1033.810 845.720 1034.810 849.990 ;
        RECT 1035.650 845.720 1036.650 849.990 ;
        RECT 1037.490 845.720 1038.490 849.990 ;
        RECT 1039.330 845.720 1040.330 849.990 ;
        RECT 1041.170 845.720 1042.170 849.990 ;
        RECT 1043.010 845.720 1044.010 849.990 ;
        RECT 1044.850 845.720 1045.850 849.990 ;
        RECT 1046.690 845.720 1047.690 849.990 ;
        RECT 1048.530 845.720 1049.530 849.990 ;
        RECT 1050.370 845.720 1051.370 849.990 ;
        RECT 1052.210 845.720 1053.210 849.990 ;
        RECT 1054.050 845.720 1055.050 849.990 ;
        RECT 1055.890 845.720 1056.890 849.990 ;
        RECT 1057.730 845.720 1058.730 849.990 ;
        RECT 1059.570 845.720 1060.570 849.990 ;
        RECT 1061.410 845.720 1062.410 849.990 ;
        RECT 1063.250 845.720 1064.250 849.990 ;
        RECT 1065.090 845.720 1066.090 849.990 ;
        RECT 1066.930 845.720 1067.930 849.990 ;
        RECT 1068.770 845.720 1069.770 849.990 ;
        RECT 1070.610 845.720 1071.610 849.990 ;
        RECT 1072.450 845.720 1073.450 849.990 ;
        RECT 1074.290 845.720 1075.290 849.990 ;
        RECT 1076.130 845.720 1077.130 849.990 ;
        RECT 1077.970 845.720 1078.970 849.990 ;
        RECT 1079.810 845.720 1080.810 849.990 ;
        RECT 1081.650 845.720 1082.650 849.990 ;
        RECT 1083.490 845.720 1084.490 849.990 ;
        RECT 1085.330 845.720 1086.330 849.990 ;
        RECT 1087.170 845.720 1088.170 849.990 ;
        RECT 1089.010 845.720 1090.010 849.990 ;
        RECT 1090.850 845.720 1091.850 849.990 ;
        RECT 1092.690 845.720 1093.690 849.990 ;
        RECT 1094.530 845.720 1095.530 849.990 ;
        RECT 1096.370 845.720 1097.370 849.990 ;
        RECT 1098.210 845.720 1099.210 849.990 ;
        RECT 1100.050 845.720 1101.050 849.990 ;
        RECT 1101.890 845.720 1102.890 849.990 ;
        RECT 1103.730 845.720 1104.730 849.990 ;
        RECT 1105.570 845.720 1106.570 849.990 ;
        RECT 1107.410 845.720 1108.410 849.990 ;
        RECT 1109.250 845.720 1110.250 849.990 ;
        RECT 1111.090 845.720 1112.090 849.990 ;
        RECT 1112.930 845.720 1113.930 849.990 ;
        RECT 1114.770 845.720 1115.770 849.990 ;
        RECT 1116.610 845.720 1117.610 849.990 ;
        RECT 1118.450 845.720 1119.450 849.990 ;
        RECT 1120.290 845.720 1121.290 849.990 ;
        RECT 1122.130 845.720 1123.130 849.990 ;
        RECT 1123.970 845.720 1124.970 849.990 ;
        RECT 1125.810 845.720 1126.810 849.990 ;
        RECT 1127.650 845.720 1128.650 849.990 ;
        RECT 1129.490 845.720 1130.490 849.990 ;
        RECT 1131.330 845.720 1132.330 849.990 ;
        RECT 1133.170 845.720 1134.170 849.990 ;
        RECT 1135.010 845.720 1136.010 849.990 ;
        RECT 1136.850 845.720 1137.850 849.990 ;
        RECT 1138.690 845.720 1139.690 849.990 ;
        RECT 1140.530 845.720 1141.530 849.990 ;
        RECT 1142.370 845.720 1143.370 849.990 ;
        RECT 1144.210 845.720 1145.210 849.990 ;
        RECT 1146.050 845.720 1147.050 849.990 ;
        RECT 1147.890 845.720 1148.890 849.990 ;
        RECT 1149.730 845.720 1150.730 849.990 ;
        RECT 1151.570 845.720 1152.570 849.990 ;
        RECT 1153.410 845.720 1154.410 849.990 ;
        RECT 1155.250 845.720 1156.250 849.990 ;
        RECT 1157.090 845.720 1158.090 849.990 ;
        RECT 1158.930 845.720 1159.930 849.990 ;
        RECT 1160.770 845.720 1161.770 849.990 ;
        RECT 1162.610 845.720 1163.610 849.990 ;
        RECT 1164.450 845.720 1165.450 849.990 ;
        RECT 1166.290 845.720 1167.290 849.990 ;
        RECT 1168.130 845.720 1169.130 849.990 ;
        RECT 1169.970 845.720 1170.970 849.990 ;
        RECT 1171.810 845.720 1172.810 849.990 ;
        RECT 1173.650 845.720 1174.650 849.990 ;
        RECT 1175.490 845.720 1176.490 849.990 ;
        RECT 1177.330 845.720 1178.330 849.990 ;
        RECT 1179.170 845.720 1180.170 849.990 ;
        RECT 1181.010 845.720 1182.010 849.990 ;
        RECT 1182.850 845.720 1183.850 849.990 ;
        RECT 1184.690 845.720 1185.690 849.990 ;
        RECT 1186.530 845.720 1187.530 849.990 ;
        RECT 1188.370 845.720 1189.370 849.990 ;
        RECT 1190.210 845.720 1191.210 849.990 ;
        RECT 1192.050 845.720 1193.050 849.990 ;
        RECT 1193.890 845.720 1194.890 849.990 ;
        RECT 1195.730 845.720 1196.730 849.990 ;
        RECT 1197.570 845.720 1198.570 849.990 ;
        RECT 1199.410 845.720 1200.410 849.990 ;
        RECT 1201.250 845.720 1202.250 849.990 ;
        RECT 1203.090 845.720 1204.090 849.990 ;
        RECT 1204.930 845.720 1205.930 849.990 ;
        RECT 1206.770 845.720 1207.770 849.990 ;
        RECT 1208.610 845.720 1209.610 849.990 ;
        RECT 1210.450 845.720 1211.450 849.990 ;
        RECT 1212.290 845.720 1213.290 849.990 ;
        RECT 1214.130 845.720 1215.130 849.990 ;
        RECT 1215.970 845.720 1216.970 849.990 ;
        RECT 1217.810 845.720 1218.810 849.990 ;
        RECT 1219.650 845.720 1220.650 849.990 ;
        RECT 1221.490 845.720 1222.490 849.990 ;
        RECT 1223.330 845.720 1224.330 849.990 ;
        RECT 1225.170 845.720 1226.170 849.990 ;
        RECT 1227.010 845.720 1228.010 849.990 ;
        RECT 1228.850 845.720 1229.850 849.990 ;
        RECT 1230.690 845.720 1231.690 849.990 ;
        RECT 1232.530 845.720 1233.530 849.990 ;
        RECT 1234.370 845.720 1235.370 849.990 ;
        RECT 1236.210 845.720 1237.210 849.990 ;
        RECT 1238.050 845.720 1239.050 849.990 ;
        RECT 1239.890 845.720 1240.890 849.990 ;
        RECT 1241.730 845.720 1242.730 849.990 ;
        RECT 1243.570 845.720 1244.570 849.990 ;
        RECT 1245.410 845.720 1246.410 849.990 ;
        RECT 1247.250 845.720 1248.250 849.990 ;
        RECT 1249.090 845.720 1250.090 849.990 ;
        RECT 1250.930 845.720 1251.930 849.990 ;
        RECT 1252.770 845.720 1253.770 849.990 ;
        RECT 1254.610 845.720 1255.610 849.990 ;
        RECT 1256.450 845.720 1257.450 849.990 ;
        RECT 1258.290 845.720 1259.290 849.990 ;
        RECT 1260.130 845.720 1261.130 849.990 ;
        RECT 1261.970 845.720 1262.970 849.990 ;
        RECT 1263.810 845.720 1264.810 849.990 ;
        RECT 1265.650 845.720 1266.650 849.990 ;
        RECT 1267.490 845.720 1268.490 849.990 ;
        RECT 1269.330 845.720 1270.330 849.990 ;
        RECT 1271.170 845.720 1272.170 849.990 ;
        RECT 1273.010 845.720 1274.010 849.990 ;
        RECT 1274.850 845.720 1275.850 849.990 ;
        RECT 1276.690 845.720 1277.690 849.990 ;
        RECT 1278.530 845.720 1279.530 849.990 ;
        RECT 1280.370 845.720 1281.370 849.990 ;
        RECT 1282.210 845.720 1283.210 849.990 ;
        RECT 1284.050 845.720 1285.050 849.990 ;
        RECT 1285.890 845.720 1286.890 849.990 ;
        RECT 1287.730 845.720 1288.730 849.990 ;
        RECT 1289.570 845.720 1290.570 849.990 ;
        RECT 1291.410 845.720 1292.410 849.990 ;
        RECT 1293.250 845.720 1294.250 849.990 ;
        RECT 1295.090 845.720 1296.090 849.990 ;
        RECT 1296.930 845.720 1297.930 849.990 ;
        RECT 1298.770 845.720 1299.770 849.990 ;
        RECT 1300.610 845.720 1301.610 849.990 ;
        RECT 1302.450 845.720 1303.450 849.990 ;
        RECT 1304.290 845.720 1305.290 849.990 ;
        RECT 1306.130 845.720 1307.130 849.990 ;
        RECT 1307.970 845.720 1308.970 849.990 ;
        RECT 1309.810 845.720 1310.810 849.990 ;
        RECT 1311.650 845.720 1312.650 849.990 ;
        RECT 1313.490 845.720 1314.490 849.990 ;
        RECT 1315.330 845.720 1316.330 849.990 ;
        RECT 1317.170 845.720 1318.170 849.990 ;
        RECT 1319.010 845.720 1320.010 849.990 ;
        RECT 1320.850 845.720 1321.850 849.990 ;
        RECT 1322.690 845.720 1323.690 849.990 ;
        RECT 1324.530 845.720 1325.530 849.990 ;
        RECT 1326.370 845.720 1327.370 849.990 ;
        RECT 1328.210 845.720 1329.210 849.990 ;
        RECT 1330.050 845.720 1331.050 849.990 ;
        RECT 1331.890 845.720 1332.890 849.990 ;
        RECT 1333.730 845.720 1334.730 849.990 ;
        RECT 1335.570 845.720 1336.570 849.990 ;
        RECT 1337.410 845.720 1338.410 849.990 ;
        RECT 1339.250 845.720 1340.250 849.990 ;
        RECT 1341.090 845.720 1342.090 849.990 ;
        RECT 1342.930 845.720 1343.930 849.990 ;
        RECT 1344.770 845.720 1345.770 849.990 ;
        RECT 1346.610 845.720 1347.610 849.990 ;
        RECT 1348.450 845.720 1349.450 849.990 ;
        RECT 1350.290 845.720 1351.290 849.990 ;
        RECT 1352.130 845.720 1353.130 849.990 ;
        RECT 1353.970 845.720 1354.970 849.990 ;
        RECT 1355.810 845.720 1356.810 849.990 ;
        RECT 1357.650 845.720 1358.650 849.990 ;
        RECT 1359.490 845.720 1360.490 849.990 ;
        RECT 1361.330 845.720 1362.330 849.990 ;
        RECT 1363.170 845.720 1364.170 849.990 ;
        RECT 1365.010 845.720 1366.010 849.990 ;
        RECT 1366.850 845.720 1367.850 849.990 ;
        RECT 1368.690 845.720 1369.690 849.990 ;
        RECT 1370.530 845.720 1371.530 849.990 ;
        RECT 1372.370 845.720 1373.370 849.990 ;
        RECT 1374.210 845.720 1375.210 849.990 ;
        RECT 1376.050 845.720 1377.050 849.990 ;
        RECT 1377.890 845.720 1378.890 849.990 ;
        RECT 1379.730 845.720 1380.730 849.990 ;
        RECT 1381.570 845.720 1382.570 849.990 ;
        RECT 1383.410 845.720 1384.410 849.990 ;
        RECT 1385.250 845.720 1386.250 849.990 ;
        RECT 1387.090 845.720 1388.090 849.990 ;
        RECT 1388.930 845.720 1389.930 849.990 ;
        RECT 1390.770 845.720 1391.770 849.990 ;
        RECT 1392.610 845.720 1393.610 849.990 ;
        RECT 1394.450 845.720 1395.450 849.990 ;
        RECT 1396.290 845.720 1397.290 849.990 ;
        RECT 1398.130 845.720 1399.130 849.990 ;
        RECT 1399.970 845.720 1400.970 849.990 ;
        RECT 1401.810 845.720 1402.810 849.990 ;
        RECT 1403.650 845.720 1404.650 849.990 ;
        RECT 1405.490 845.720 1406.490 849.990 ;
        RECT 1407.330 845.720 1408.330 849.990 ;
        RECT 1409.170 845.720 1410.170 849.990 ;
        RECT 1411.010 845.720 1412.010 849.990 ;
        RECT 1412.850 845.720 1413.850 849.990 ;
        RECT 1414.690 845.720 1415.690 849.990 ;
        RECT 1416.530 845.720 1417.530 849.990 ;
        RECT 1418.370 845.720 1419.370 849.990 ;
        RECT 1420.210 845.720 1421.210 849.990 ;
        RECT 1422.050 845.720 1423.050 849.990 ;
        RECT 1423.890 845.720 1424.890 849.990 ;
        RECT 1425.730 845.720 1426.730 849.990 ;
        RECT 1427.570 845.720 1428.570 849.990 ;
        RECT 1429.410 845.720 1430.410 849.990 ;
        RECT 1431.250 845.720 1432.250 849.990 ;
        RECT 1433.090 845.720 1434.090 849.990 ;
        RECT 1434.930 845.720 1435.930 849.990 ;
        RECT 1436.770 845.720 1437.770 849.990 ;
        RECT 1438.610 845.720 1439.610 849.990 ;
        RECT 1440.450 845.720 1441.450 849.990 ;
        RECT 1442.290 845.720 1443.290 849.990 ;
        RECT 1444.130 845.720 1445.130 849.990 ;
        RECT 1445.970 845.720 1446.970 849.990 ;
        RECT 1447.810 845.720 1448.810 849.990 ;
        RECT 1449.650 845.720 1450.650 849.990 ;
        RECT 1451.490 845.720 1452.490 849.990 ;
        RECT 1453.330 845.720 1454.330 849.990 ;
        RECT 1455.170 845.720 1456.170 849.990 ;
        RECT 1457.010 845.720 1458.010 849.990 ;
        RECT 1458.850 845.720 1459.850 849.990 ;
        RECT 1460.690 845.720 1461.690 849.990 ;
        RECT 1462.530 845.720 1463.530 849.990 ;
        RECT 1464.370 845.720 1465.370 849.990 ;
        RECT 1466.210 845.720 1467.210 849.990 ;
        RECT 1468.050 845.720 1469.050 849.990 ;
        RECT 1469.890 845.720 1470.890 849.990 ;
        RECT 1471.730 845.720 1472.730 849.990 ;
        RECT 1473.570 845.720 1474.570 849.990 ;
        RECT 1475.410 845.720 1476.410 849.990 ;
        RECT 1477.250 845.720 1478.250 849.990 ;
        RECT 1479.090 845.720 1480.090 849.990 ;
        RECT 1480.930 845.720 1481.930 849.990 ;
        RECT 1482.770 845.720 1483.770 849.990 ;
        RECT 1484.610 845.720 1485.610 849.990 ;
        RECT 1486.450 845.720 1487.450 849.990 ;
        RECT 1488.290 845.720 1489.290 849.990 ;
        RECT 1490.130 845.720 1491.130 849.990 ;
        RECT 1491.970 845.720 1492.970 849.990 ;
        RECT 1493.810 845.720 1494.810 849.990 ;
        RECT 1495.650 845.720 1496.650 849.990 ;
        RECT 1497.490 845.720 1498.490 849.990 ;
        RECT 1499.330 845.720 1500.330 849.990 ;
        RECT 1501.170 845.720 1502.170 849.990 ;
        RECT 1503.010 845.720 1504.010 849.990 ;
        RECT 1504.850 845.720 1505.850 849.990 ;
        RECT 1506.690 845.720 1507.690 849.990 ;
        RECT 1508.530 845.720 1509.530 849.990 ;
        RECT 1510.370 845.720 1511.370 849.990 ;
        RECT 1512.210 845.720 1513.210 849.990 ;
        RECT 1514.050 845.720 1515.050 849.990 ;
        RECT 1515.890 845.720 1516.890 849.990 ;
        RECT 1517.730 845.720 1518.730 849.990 ;
        RECT 1519.570 845.720 1520.570 849.990 ;
        RECT 1521.410 845.720 1522.410 849.990 ;
        RECT 1523.250 845.720 1524.250 849.990 ;
        RECT 1525.090 845.720 1526.090 849.990 ;
        RECT 1526.930 845.720 1527.930 849.990 ;
        RECT 1528.770 845.720 1529.770 849.990 ;
        RECT 1530.610 845.720 1531.610 849.990 ;
        RECT 1532.450 845.720 1533.450 849.990 ;
        RECT 1534.290 845.720 1535.290 849.990 ;
        RECT 1536.130 845.720 1537.130 849.990 ;
        RECT 1537.970 845.720 1538.970 849.990 ;
        RECT 1539.810 845.720 1540.810 849.990 ;
        RECT 1541.650 845.720 1542.650 849.990 ;
        RECT 1543.490 845.720 1544.490 849.990 ;
        RECT 1545.330 845.720 1546.330 849.990 ;
        RECT 1547.170 845.720 1548.170 849.990 ;
        RECT 1549.010 845.720 1550.010 849.990 ;
        RECT 1550.850 845.720 1551.850 849.990 ;
        RECT 1552.690 845.720 1675.130 849.990 ;
        RECT 1675.970 845.720 2133.290 849.990 ;
        RECT 2134.130 845.720 2135.130 849.990 ;
        RECT 2135.970 845.720 2136.970 849.990 ;
        RECT 2137.810 845.720 2138.810 849.990 ;
        RECT 2139.650 845.720 2140.650 849.990 ;
        RECT 2141.490 845.720 2142.490 849.990 ;
        RECT 2143.330 845.720 2144.330 849.990 ;
        RECT 2145.170 845.720 2146.170 849.990 ;
        RECT 2.850 4.280 2146.720 845.720 ;
        RECT 3.410 3.070 3.490 4.280 ;
        RECT 4.330 3.070 4.410 4.280 ;
        RECT 5.250 3.070 5.330 4.280 ;
        RECT 6.170 3.070 6.250 4.280 ;
        RECT 7.090 3.070 7.170 4.280 ;
        RECT 8.010 3.070 8.090 4.280 ;
        RECT 8.930 3.070 9.010 4.280 ;
        RECT 9.850 3.070 9.930 4.280 ;
        RECT 10.770 3.070 10.850 4.280 ;
        RECT 11.690 3.070 11.770 4.280 ;
        RECT 12.610 3.070 12.690 4.280 ;
        RECT 13.530 3.070 13.610 4.280 ;
        RECT 14.450 3.070 14.530 4.280 ;
        RECT 15.370 3.070 15.450 4.280 ;
        RECT 16.290 3.070 16.370 4.280 ;
        RECT 17.210 3.070 17.290 4.280 ;
        RECT 18.130 3.070 18.210 4.280 ;
        RECT 19.050 3.070 19.130 4.280 ;
        RECT 19.970 3.070 20.050 4.280 ;
        RECT 20.890 3.070 20.970 4.280 ;
        RECT 21.810 3.070 21.890 4.280 ;
        RECT 22.730 3.070 22.810 4.280 ;
        RECT 23.650 3.070 23.730 4.280 ;
        RECT 24.570 3.070 24.650 4.280 ;
        RECT 25.490 3.070 25.570 4.280 ;
        RECT 26.410 3.070 26.490 4.280 ;
        RECT 27.330 3.070 27.410 4.280 ;
        RECT 28.250 3.070 28.330 4.280 ;
        RECT 29.170 3.070 29.250 4.280 ;
        RECT 30.090 3.070 30.170 4.280 ;
        RECT 31.010 3.070 31.090 4.280 ;
        RECT 31.930 3.070 32.010 4.280 ;
        RECT 32.850 3.070 32.930 4.280 ;
        RECT 33.770 3.070 33.850 4.280 ;
        RECT 34.690 3.070 34.770 4.280 ;
        RECT 35.610 3.070 35.690 4.280 ;
        RECT 36.530 3.070 36.610 4.280 ;
        RECT 37.450 3.070 37.530 4.280 ;
        RECT 38.370 3.070 38.450 4.280 ;
        RECT 39.290 3.070 39.370 4.280 ;
        RECT 40.210 3.070 40.290 4.280 ;
        RECT 41.130 3.070 41.210 4.280 ;
        RECT 42.050 3.070 42.130 4.280 ;
        RECT 42.970 3.070 43.050 4.280 ;
        RECT 43.890 3.070 43.970 4.280 ;
        RECT 44.810 3.070 44.890 4.280 ;
        RECT 45.730 3.070 45.810 4.280 ;
        RECT 46.650 3.070 46.730 4.280 ;
        RECT 47.570 3.070 47.650 4.280 ;
        RECT 48.490 3.070 48.570 4.280 ;
        RECT 49.410 3.070 49.490 4.280 ;
        RECT 50.330 3.070 50.410 4.280 ;
        RECT 51.250 3.070 51.330 4.280 ;
        RECT 52.170 3.070 52.250 4.280 ;
        RECT 53.090 3.070 53.170 4.280 ;
        RECT 54.010 3.070 54.090 4.280 ;
        RECT 54.930 3.070 55.010 4.280 ;
        RECT 55.850 3.070 55.930 4.280 ;
        RECT 56.770 3.070 56.850 4.280 ;
        RECT 57.690 3.070 57.770 4.280 ;
        RECT 58.610 3.070 58.690 4.280 ;
        RECT 59.530 3.070 59.610 4.280 ;
        RECT 60.450 3.070 60.530 4.280 ;
        RECT 61.370 3.070 61.450 4.280 ;
        RECT 62.290 3.070 62.370 4.280 ;
        RECT 63.210 3.070 63.290 4.280 ;
        RECT 64.130 3.070 64.210 4.280 ;
        RECT 65.050 3.070 65.130 4.280 ;
        RECT 65.970 3.070 66.050 4.280 ;
        RECT 66.890 3.070 66.970 4.280 ;
        RECT 67.810 3.070 67.890 4.280 ;
        RECT 68.730 3.070 68.810 4.280 ;
        RECT 69.650 3.070 69.730 4.280 ;
        RECT 70.570 3.070 70.650 4.280 ;
        RECT 71.490 3.070 71.570 4.280 ;
        RECT 72.410 3.070 72.490 4.280 ;
        RECT 73.330 3.070 73.410 4.280 ;
        RECT 74.250 3.070 74.330 4.280 ;
        RECT 75.170 3.070 75.250 4.280 ;
        RECT 76.090 3.070 76.170 4.280 ;
        RECT 77.010 3.070 77.090 4.280 ;
        RECT 77.930 3.070 78.010 4.280 ;
        RECT 78.850 3.070 78.930 4.280 ;
        RECT 79.770 3.070 79.850 4.280 ;
        RECT 80.690 3.070 81.690 4.280 ;
        RECT 82.530 3.070 83.530 4.280 ;
        RECT 84.370 3.070 85.370 4.280 ;
        RECT 86.210 3.070 87.210 4.280 ;
        RECT 88.050 3.070 89.050 4.280 ;
        RECT 89.890 3.070 90.890 4.280 ;
        RECT 91.730 3.070 92.730 4.280 ;
        RECT 93.570 3.070 94.570 4.280 ;
        RECT 95.410 3.070 96.410 4.280 ;
        RECT 97.250 3.070 98.250 4.280 ;
        RECT 99.090 3.070 100.090 4.280 ;
        RECT 100.930 3.070 101.930 4.280 ;
        RECT 102.770 3.070 103.770 4.280 ;
        RECT 104.610 3.070 105.610 4.280 ;
        RECT 106.450 3.070 107.450 4.280 ;
        RECT 108.290 3.070 109.290 4.280 ;
        RECT 110.130 3.070 111.130 4.280 ;
        RECT 111.970 3.070 112.970 4.280 ;
        RECT 113.810 3.070 114.810 4.280 ;
        RECT 115.650 3.070 116.650 4.280 ;
        RECT 117.490 3.070 118.490 4.280 ;
        RECT 119.330 3.070 120.330 4.280 ;
        RECT 121.170 3.070 122.170 4.280 ;
        RECT 123.010 3.070 124.010 4.280 ;
        RECT 124.850 3.070 125.850 4.280 ;
        RECT 126.690 3.070 127.690 4.280 ;
        RECT 128.530 3.070 129.530 4.280 ;
        RECT 130.370 3.070 131.370 4.280 ;
        RECT 132.210 3.070 133.210 4.280 ;
        RECT 134.050 3.070 135.050 4.280 ;
        RECT 135.890 3.070 136.890 4.280 ;
        RECT 137.730 3.070 138.730 4.280 ;
        RECT 139.570 3.070 140.570 4.280 ;
        RECT 141.410 3.070 142.410 4.280 ;
        RECT 143.250 3.070 144.250 4.280 ;
        RECT 145.090 3.070 146.090 4.280 ;
        RECT 146.930 3.070 147.930 4.280 ;
        RECT 148.770 3.070 149.770 4.280 ;
        RECT 150.610 3.070 151.610 4.280 ;
        RECT 152.450 3.070 153.450 4.280 ;
        RECT 154.290 3.070 155.290 4.280 ;
        RECT 156.130 3.070 157.130 4.280 ;
        RECT 157.970 3.070 158.970 4.280 ;
        RECT 159.810 3.070 160.810 4.280 ;
        RECT 161.650 3.070 162.650 4.280 ;
        RECT 163.490 3.070 164.490 4.280 ;
        RECT 165.330 3.070 166.330 4.280 ;
        RECT 167.170 3.070 168.170 4.280 ;
        RECT 169.010 3.070 170.010 4.280 ;
        RECT 170.850 3.070 171.850 4.280 ;
        RECT 172.690 3.070 173.690 4.280 ;
        RECT 174.530 3.070 175.530 4.280 ;
        RECT 176.370 3.070 177.370 4.280 ;
        RECT 178.210 3.070 179.210 4.280 ;
        RECT 180.050 3.070 181.050 4.280 ;
        RECT 181.890 3.070 182.890 4.280 ;
        RECT 183.730 3.070 184.730 4.280 ;
        RECT 185.570 3.070 186.570 4.280 ;
        RECT 187.410 3.070 188.410 4.280 ;
        RECT 189.250 3.070 190.250 4.280 ;
        RECT 191.090 3.070 192.090 4.280 ;
        RECT 192.930 3.070 193.930 4.280 ;
        RECT 194.770 3.070 195.770 4.280 ;
        RECT 196.610 3.070 197.610 4.280 ;
        RECT 198.450 3.070 2111.210 4.280 ;
        RECT 2112.050 3.070 2113.050 4.280 ;
        RECT 2113.890 3.070 2114.890 4.280 ;
        RECT 2115.730 3.070 2116.730 4.280 ;
        RECT 2117.570 3.070 2118.570 4.280 ;
        RECT 2119.410 3.070 2120.410 4.280 ;
        RECT 2121.250 3.070 2122.250 4.280 ;
        RECT 2123.090 3.070 2124.090 4.280 ;
        RECT 2124.930 3.070 2125.930 4.280 ;
        RECT 2126.770 3.070 2127.770 4.280 ;
        RECT 2128.610 3.070 2129.610 4.280 ;
        RECT 2130.450 3.070 2131.450 4.280 ;
        RECT 2132.290 3.070 2133.290 4.280 ;
        RECT 2134.130 3.070 2135.130 4.280 ;
        RECT 2135.970 3.070 2136.970 4.280 ;
        RECT 2137.810 3.070 2138.810 4.280 ;
        RECT 2139.650 3.070 2140.650 4.280 ;
        RECT 2141.490 3.070 2142.490 4.280 ;
        RECT 2143.330 3.070 2144.330 4.280 ;
        RECT 2145.170 3.070 2146.170 4.280 ;
      LAYER met3 ;
        RECT 4.400 842.840 2145.600 843.705 ;
        RECT 2.825 841.520 2146.050 842.840 ;
        RECT 4.400 840.120 2145.600 841.520 ;
        RECT 2.825 838.800 2146.050 840.120 ;
        RECT 4.400 837.400 2145.600 838.800 ;
        RECT 2.825 836.080 2146.050 837.400 ;
        RECT 4.400 834.680 2145.600 836.080 ;
        RECT 2.825 833.360 2146.050 834.680 ;
        RECT 4.400 831.960 2146.050 833.360 ;
        RECT 2.825 830.640 2146.050 831.960 ;
        RECT 4.400 829.240 2146.050 830.640 ;
        RECT 2.825 827.920 2146.050 829.240 ;
        RECT 4.400 826.520 2146.050 827.920 ;
        RECT 2.825 825.200 2146.050 826.520 ;
        RECT 4.400 823.800 2146.050 825.200 ;
        RECT 2.825 822.480 2146.050 823.800 ;
        RECT 4.400 821.080 2146.050 822.480 ;
        RECT 2.825 819.760 2146.050 821.080 ;
        RECT 4.400 818.360 2146.050 819.760 ;
        RECT 2.825 817.040 2146.050 818.360 ;
        RECT 4.400 815.640 2146.050 817.040 ;
        RECT 2.825 814.320 2146.050 815.640 ;
        RECT 4.400 812.920 2146.050 814.320 ;
        RECT 2.825 811.600 2146.050 812.920 ;
        RECT 4.400 810.200 2146.050 811.600 ;
        RECT 2.825 808.880 2146.050 810.200 ;
        RECT 4.400 807.480 2146.050 808.880 ;
        RECT 2.825 806.160 2146.050 807.480 ;
        RECT 4.400 804.760 2146.050 806.160 ;
        RECT 2.825 803.440 2146.050 804.760 ;
        RECT 4.400 802.040 2146.050 803.440 ;
        RECT 2.825 800.720 2146.050 802.040 ;
        RECT 4.400 799.320 2146.050 800.720 ;
        RECT 2.825 798.000 2146.050 799.320 ;
        RECT 4.400 796.600 2146.050 798.000 ;
        RECT 2.825 795.280 2146.050 796.600 ;
        RECT 4.400 793.880 2146.050 795.280 ;
        RECT 2.825 787.120 2146.050 793.880 ;
        RECT 2.825 785.720 2145.600 787.120 ;
        RECT 2.825 746.320 2146.050 785.720 ;
        RECT 4.400 744.920 2146.050 746.320 ;
        RECT 2.825 566.800 2146.050 744.920 ;
        RECT 2.825 565.400 2145.600 566.800 ;
        RECT 2.825 564.080 2146.050 565.400 ;
        RECT 2.825 562.680 2145.600 564.080 ;
        RECT 2.825 561.360 2146.050 562.680 ;
        RECT 2.825 559.960 2145.600 561.360 ;
        RECT 2.825 482.480 2146.050 559.960 ;
        RECT 2.825 481.080 2145.600 482.480 ;
        RECT 2.825 449.840 2146.050 481.080 ;
        RECT 2.825 448.440 2145.600 449.840 ;
        RECT 2.825 341.040 2146.050 448.440 ;
        RECT 2.825 339.640 2145.600 341.040 ;
        RECT 2.825 338.320 2146.050 339.640 ;
        RECT 2.825 336.920 2145.600 338.320 ;
        RECT 2.825 335.600 2146.050 336.920 ;
        RECT 2.825 334.200 2145.600 335.600 ;
        RECT 2.825 332.880 2146.050 334.200 ;
        RECT 2.825 331.480 2145.600 332.880 ;
        RECT 2.825 199.600 2146.050 331.480 ;
        RECT 4.400 198.200 2146.050 199.600 ;
        RECT 2.825 196.880 2146.050 198.200 ;
        RECT 4.400 195.480 2146.050 196.880 ;
        RECT 2.825 194.160 2146.050 195.480 ;
        RECT 4.400 192.760 2146.050 194.160 ;
        RECT 2.825 191.440 2146.050 192.760 ;
        RECT 4.400 190.040 2146.050 191.440 ;
        RECT 2.825 188.720 2146.050 190.040 ;
        RECT 4.400 187.320 2146.050 188.720 ;
        RECT 2.825 186.000 2146.050 187.320 ;
        RECT 4.400 184.600 2146.050 186.000 ;
        RECT 2.825 183.280 2146.050 184.600 ;
        RECT 4.400 181.880 2146.050 183.280 ;
        RECT 2.825 180.560 2146.050 181.880 ;
        RECT 4.400 179.160 2146.050 180.560 ;
        RECT 2.825 177.840 2146.050 179.160 ;
        RECT 4.400 176.440 2146.050 177.840 ;
        RECT 2.825 175.120 2146.050 176.440 ;
        RECT 4.400 173.720 2146.050 175.120 ;
        RECT 2.825 172.400 2146.050 173.720 ;
        RECT 4.400 171.000 2146.050 172.400 ;
        RECT 2.825 169.680 2146.050 171.000 ;
        RECT 4.400 168.280 2146.050 169.680 ;
        RECT 2.825 166.960 2146.050 168.280 ;
        RECT 4.400 165.560 2146.050 166.960 ;
        RECT 2.825 164.240 2146.050 165.560 ;
        RECT 4.400 162.840 2146.050 164.240 ;
        RECT 2.825 161.520 2146.050 162.840 ;
        RECT 4.400 160.120 2146.050 161.520 ;
        RECT 2.825 158.800 2146.050 160.120 ;
        RECT 4.400 157.400 2146.050 158.800 ;
        RECT 2.825 156.080 2146.050 157.400 ;
        RECT 4.400 154.680 2146.050 156.080 ;
        RECT 2.825 153.360 2146.050 154.680 ;
        RECT 4.400 151.960 2146.050 153.360 ;
        RECT 2.825 150.640 2146.050 151.960 ;
        RECT 4.400 149.240 2146.050 150.640 ;
        RECT 2.825 147.920 2146.050 149.240 ;
        RECT 4.400 146.520 2146.050 147.920 ;
        RECT 2.825 145.200 2146.050 146.520 ;
        RECT 4.400 143.800 2146.050 145.200 ;
        RECT 2.825 142.480 2146.050 143.800 ;
        RECT 4.400 141.080 2146.050 142.480 ;
        RECT 2.825 139.760 2146.050 141.080 ;
        RECT 4.400 138.360 2146.050 139.760 ;
        RECT 2.825 137.040 2146.050 138.360 ;
        RECT 4.400 135.640 2146.050 137.040 ;
        RECT 2.825 134.320 2146.050 135.640 ;
        RECT 4.400 132.920 2146.050 134.320 ;
        RECT 2.825 131.600 2146.050 132.920 ;
        RECT 4.400 130.200 2146.050 131.600 ;
        RECT 2.825 128.880 2146.050 130.200 ;
        RECT 4.400 127.480 2146.050 128.880 ;
        RECT 2.825 126.160 2146.050 127.480 ;
        RECT 4.400 124.760 2146.050 126.160 ;
        RECT 2.825 123.440 2146.050 124.760 ;
        RECT 4.400 122.040 2146.050 123.440 ;
        RECT 2.825 120.720 2146.050 122.040 ;
        RECT 4.400 119.320 2146.050 120.720 ;
        RECT 2.825 118.000 2146.050 119.320 ;
        RECT 4.400 116.600 2146.050 118.000 ;
        RECT 2.825 115.280 2146.050 116.600 ;
        RECT 4.400 113.880 2146.050 115.280 ;
        RECT 2.825 112.560 2146.050 113.880 ;
        RECT 4.400 111.160 2146.050 112.560 ;
        RECT 2.825 109.840 2146.050 111.160 ;
        RECT 4.400 108.440 2145.600 109.840 ;
        RECT 2.825 107.120 2146.050 108.440 ;
        RECT 4.400 105.720 2146.050 107.120 ;
        RECT 2.825 104.400 2146.050 105.720 ;
        RECT 4.400 103.000 2146.050 104.400 ;
        RECT 2.825 101.680 2146.050 103.000 ;
        RECT 4.400 100.280 2146.050 101.680 ;
        RECT 2.825 98.960 2146.050 100.280 ;
        RECT 4.400 97.560 2146.050 98.960 ;
        RECT 2.825 96.240 2146.050 97.560 ;
        RECT 4.400 94.840 2146.050 96.240 ;
        RECT 2.825 93.520 2146.050 94.840 ;
        RECT 4.400 92.120 2146.050 93.520 ;
        RECT 2.825 90.800 2146.050 92.120 ;
        RECT 4.400 89.400 2146.050 90.800 ;
        RECT 2.825 88.080 2146.050 89.400 ;
        RECT 4.400 86.680 2146.050 88.080 ;
        RECT 2.825 85.360 2146.050 86.680 ;
        RECT 4.400 83.960 2146.050 85.360 ;
        RECT 2.825 82.640 2146.050 83.960 ;
        RECT 4.400 81.240 2146.050 82.640 ;
        RECT 2.825 79.920 2146.050 81.240 ;
        RECT 4.400 78.520 2146.050 79.920 ;
        RECT 2.825 77.200 2146.050 78.520 ;
        RECT 4.400 75.800 2146.050 77.200 ;
        RECT 2.825 74.480 2146.050 75.800 ;
        RECT 4.400 73.080 2146.050 74.480 ;
        RECT 2.825 71.760 2146.050 73.080 ;
        RECT 4.400 70.360 2146.050 71.760 ;
        RECT 2.825 69.040 2146.050 70.360 ;
        RECT 4.400 67.640 2146.050 69.040 ;
        RECT 2.825 66.320 2146.050 67.640 ;
        RECT 4.400 64.920 2146.050 66.320 ;
        RECT 2.825 63.600 2146.050 64.920 ;
        RECT 4.400 62.200 2146.050 63.600 ;
        RECT 2.825 60.880 2146.050 62.200 ;
        RECT 4.400 59.480 2146.050 60.880 ;
        RECT 2.825 58.160 2146.050 59.480 ;
        RECT 4.400 56.760 2146.050 58.160 ;
        RECT 2.825 55.440 2146.050 56.760 ;
        RECT 4.400 54.040 2146.050 55.440 ;
        RECT 2.825 52.720 2146.050 54.040 ;
        RECT 4.400 51.320 2146.050 52.720 ;
        RECT 2.825 50.000 2146.050 51.320 ;
        RECT 4.400 48.600 2146.050 50.000 ;
        RECT 2.825 47.280 2146.050 48.600 ;
        RECT 4.400 45.880 2146.050 47.280 ;
        RECT 2.825 44.560 2146.050 45.880 ;
        RECT 4.400 43.160 2146.050 44.560 ;
        RECT 2.825 41.840 2146.050 43.160 ;
        RECT 4.400 40.440 2146.050 41.840 ;
        RECT 2.825 39.120 2146.050 40.440 ;
        RECT 4.400 37.720 2146.050 39.120 ;
        RECT 2.825 36.400 2146.050 37.720 ;
        RECT 4.400 35.000 2145.600 36.400 ;
        RECT 2.825 33.680 2146.050 35.000 ;
        RECT 4.400 32.280 2145.600 33.680 ;
        RECT 2.825 30.960 2146.050 32.280 ;
        RECT 4.400 29.560 2145.600 30.960 ;
        RECT 2.825 28.240 2146.050 29.560 ;
        RECT 4.400 26.840 2145.600 28.240 ;
        RECT 2.825 25.520 2146.050 26.840 ;
        RECT 4.400 24.120 2145.600 25.520 ;
        RECT 2.825 22.800 2146.050 24.120 ;
        RECT 4.400 21.400 2145.600 22.800 ;
        RECT 2.825 20.080 2146.050 21.400 ;
        RECT 4.400 18.680 2145.600 20.080 ;
        RECT 2.825 17.360 2146.050 18.680 ;
        RECT 4.400 15.960 2145.600 17.360 ;
        RECT 2.825 14.640 2146.050 15.960 ;
        RECT 4.400 13.240 2145.600 14.640 ;
        RECT 2.825 11.920 2146.050 13.240 ;
        RECT 4.400 10.520 2145.600 11.920 ;
        RECT 2.825 9.200 2146.050 10.520 ;
        RECT 4.400 7.800 2145.600 9.200 ;
        RECT 2.825 6.480 2146.050 7.800 ;
        RECT 4.400 5.615 2145.600 6.480 ;
      LAYER met4 ;
        RECT 19.615 6.295 2137.290 841.665 ;
      LAYER met5 ;
        RECT 5.520 26.490 2144.060 835.500 ;
  END
END mgmt_core
END LIBRARY

