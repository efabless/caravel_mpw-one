magic
tech sky130A
magscale 1 2
timestamp 1623348513
<< pwell >>
rect 467 350 491 401
<< obsm1 >>
rect 0 852 876 918
rect 0 66 66 852
rect 113 491 141 824
rect 169 519 197 852
rect 225 491 253 824
rect 281 519 309 852
rect 337 491 365 824
rect 411 491 465 824
rect 511 491 539 824
rect 567 519 595 852
rect 623 491 651 824
rect 679 519 707 852
rect 735 491 763 824
rect 113 427 763 491
rect 113 94 141 427
rect 169 66 197 399
rect 225 94 253 427
rect 281 66 309 399
rect 337 94 365 427
rect 411 94 465 427
rect 511 94 539 427
rect 567 66 595 399
rect 623 94 651 427
rect 679 66 707 399
rect 735 94 763 427
rect 810 66 876 852
rect 0 0 876 66
<< metal2 >>
rect 0 852 383 918
rect 0 768 66 852
rect 411 824 465 918
rect 493 852 876 918
rect 94 796 782 824
rect 0 740 383 768
rect 0 656 66 740
rect 411 712 465 796
rect 810 768 876 852
rect 493 740 876 768
rect 94 684 782 712
rect 0 628 383 656
rect 0 544 66 628
rect 411 600 465 684
rect 810 656 876 740
rect 493 628 876 656
rect 94 572 782 600
rect 0 516 383 544
rect 411 488 465 572
rect 810 544 876 628
rect 493 516 876 544
rect 0 430 876 488
rect 0 374 383 402
rect 0 290 66 374
rect 411 346 465 430
rect 493 374 876 402
rect 94 318 782 346
rect 0 262 383 290
rect 0 178 66 262
rect 411 234 465 318
rect 810 290 876 374
rect 493 262 876 290
rect 94 206 782 234
rect 0 150 383 178
rect 0 66 66 150
rect 411 122 465 206
rect 810 178 876 262
rect 493 150 876 178
rect 94 94 782 122
rect 0 0 383 66
rect 411 0 465 94
rect 810 66 876 150
rect 493 0 876 66
<< labels >>
rlabel metal2 s 810 768 876 852 6 C0
port 1 nsew
rlabel metal2 s 810 656 876 740 6 C0
port 1 nsew
rlabel metal2 s 810 544 876 628 6 C0
port 1 nsew
rlabel metal2 s 810 290 876 374 6 C0
port 1 nsew
rlabel metal2 s 810 178 876 262 6 C0
port 1 nsew
rlabel metal2 s 810 66 876 150 6 C0
port 1 nsew
rlabel metal2 s 493 852 876 918 6 C0
port 1 nsew
rlabel metal2 s 493 740 876 768 6 C0
port 1 nsew
rlabel metal2 s 493 628 876 656 6 C0
port 1 nsew
rlabel metal2 s 493 516 876 544 6 C0
port 1 nsew
rlabel metal2 s 493 374 876 402 6 C0
port 1 nsew
rlabel metal2 s 493 262 876 290 6 C0
port 1 nsew
rlabel metal2 s 493 150 876 178 6 C0
port 1 nsew
rlabel metal2 s 493 0 876 66 6 C0
port 1 nsew
rlabel metal2 s 0 852 383 918 6 C0
port 1 nsew
rlabel metal2 s 0 768 66 852 6 C0
port 1 nsew
rlabel metal2 s 0 740 383 768 6 C0
port 1 nsew
rlabel metal2 s 0 656 66 740 6 C0
port 1 nsew
rlabel metal2 s 0 628 383 656 6 C0
port 1 nsew
rlabel metal2 s 0 544 66 628 6 C0
port 1 nsew
rlabel metal2 s 0 516 383 544 6 C0
port 1 nsew
rlabel metal2 s 0 374 383 402 6 C0
port 1 nsew
rlabel metal2 s 0 290 66 374 6 C0
port 1 nsew
rlabel metal2 s 0 262 383 290 6 C0
port 1 nsew
rlabel metal2 s 0 178 66 262 6 C0
port 1 nsew
rlabel metal2 s 0 150 383 178 6 C0
port 1 nsew
rlabel metal2 s 0 66 66 150 6 C0
port 1 nsew
rlabel metal2 s 0 0 383 66 6 C0
port 1 nsew
rlabel metal2 s 411 824 465 918 6 C1
port 2 nsew
rlabel metal2 s 411 712 465 796 6 C1
port 2 nsew
rlabel metal2 s 411 600 465 684 6 C1
port 2 nsew
rlabel metal2 s 411 488 465 572 6 C1
port 2 nsew
rlabel metal2 s 411 346 465 430 6 C1
port 2 nsew
rlabel metal2 s 411 234 465 318 6 C1
port 2 nsew
rlabel metal2 s 411 122 465 206 6 C1
port 2 nsew
rlabel metal2 s 411 0 465 94 6 C1
port 2 nsew
rlabel metal2 s 94 796 782 824 6 C1
port 2 nsew
rlabel metal2 s 94 684 782 712 6 C1
port 2 nsew
rlabel metal2 s 94 572 782 600 6 C1
port 2 nsew
rlabel metal2 s 94 318 782 346 6 C1
port 2 nsew
rlabel metal2 s 94 206 782 234 6 C1
port 2 nsew
rlabel metal2 s 94 94 782 122 6 C1
port 2 nsew
rlabel metal2 s 0 430 876 488 6 C1
port 2 nsew
rlabel pwell s 467 350 491 401 6 SUB
port 3 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 876 918
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 100224
string GDS_START 90816
<< end >>
