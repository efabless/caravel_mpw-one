magic
tech sky130A
magscale 1 2
timestamp 1623348512
<< checkpaint >>
rect -1260 -1260 1956 2066
<< nwell >>
rect 0 0 696 806
<< pmos >>
rect 204 102 234 704
rect 290 102 320 704
rect 376 102 406 704
rect 462 102 492 704
<< pdiff >>
rect 148 692 204 704
rect 148 658 159 692
rect 193 658 204 692
rect 148 624 204 658
rect 148 590 159 624
rect 193 590 204 624
rect 148 556 204 590
rect 148 522 159 556
rect 193 522 204 556
rect 148 488 204 522
rect 148 454 159 488
rect 193 454 204 488
rect 148 420 204 454
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 234 692 290 704
rect 234 658 245 692
rect 279 658 290 692
rect 234 624 290 658
rect 234 590 245 624
rect 279 590 290 624
rect 234 556 290 590
rect 234 522 245 556
rect 279 522 290 556
rect 234 488 290 522
rect 234 454 245 488
rect 279 454 290 488
rect 234 420 290 454
rect 234 386 245 420
rect 279 386 290 420
rect 234 352 290 386
rect 234 318 245 352
rect 279 318 290 352
rect 234 284 290 318
rect 234 250 245 284
rect 279 250 290 284
rect 234 216 290 250
rect 234 182 245 216
rect 279 182 290 216
rect 234 148 290 182
rect 234 114 245 148
rect 279 114 290 148
rect 234 102 290 114
rect 320 692 376 704
rect 320 658 331 692
rect 365 658 376 692
rect 320 624 376 658
rect 320 590 331 624
rect 365 590 376 624
rect 320 556 376 590
rect 320 522 331 556
rect 365 522 376 556
rect 320 488 376 522
rect 320 454 331 488
rect 365 454 376 488
rect 320 420 376 454
rect 320 386 331 420
rect 365 386 376 420
rect 320 352 376 386
rect 320 318 331 352
rect 365 318 376 352
rect 320 284 376 318
rect 320 250 331 284
rect 365 250 376 284
rect 320 216 376 250
rect 320 182 331 216
rect 365 182 376 216
rect 320 148 376 182
rect 320 114 331 148
rect 365 114 376 148
rect 320 102 376 114
rect 406 692 462 704
rect 406 658 417 692
rect 451 658 462 692
rect 406 624 462 658
rect 406 590 417 624
rect 451 590 462 624
rect 406 556 462 590
rect 406 522 417 556
rect 451 522 462 556
rect 406 488 462 522
rect 406 454 417 488
rect 451 454 462 488
rect 406 420 462 454
rect 406 386 417 420
rect 451 386 462 420
rect 406 352 462 386
rect 406 318 417 352
rect 451 318 462 352
rect 406 284 462 318
rect 406 250 417 284
rect 451 250 462 284
rect 406 216 462 250
rect 406 182 417 216
rect 451 182 462 216
rect 406 148 462 182
rect 406 114 417 148
rect 451 114 462 148
rect 406 102 462 114
rect 492 692 548 704
rect 492 658 503 692
rect 537 658 548 692
rect 492 624 548 658
rect 492 590 503 624
rect 537 590 548 624
rect 492 556 548 590
rect 492 522 503 556
rect 537 522 548 556
rect 492 488 548 522
rect 492 454 503 488
rect 537 454 548 488
rect 492 420 548 454
rect 492 386 503 420
rect 537 386 548 420
rect 492 352 548 386
rect 492 318 503 352
rect 537 318 548 352
rect 492 284 548 318
rect 492 250 503 284
rect 537 250 548 284
rect 492 216 548 250
rect 492 182 503 216
rect 537 182 548 216
rect 492 148 548 182
rect 492 114 503 148
rect 537 114 548 148
rect 492 102 548 114
<< pdiffc >>
rect 159 658 193 692
rect 159 590 193 624
rect 159 522 193 556
rect 159 454 193 488
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 245 658 279 692
rect 245 590 279 624
rect 245 522 279 556
rect 245 454 279 488
rect 245 386 279 420
rect 245 318 279 352
rect 245 250 279 284
rect 245 182 279 216
rect 245 114 279 148
rect 331 658 365 692
rect 331 590 365 624
rect 331 522 365 556
rect 331 454 365 488
rect 331 386 365 420
rect 331 318 365 352
rect 331 250 365 284
rect 331 182 365 216
rect 331 114 365 148
rect 417 658 451 692
rect 417 590 451 624
rect 417 522 451 556
rect 417 454 451 488
rect 417 386 451 420
rect 417 318 451 352
rect 417 250 451 284
rect 417 182 451 216
rect 417 114 451 148
rect 503 658 537 692
rect 503 590 537 624
rect 503 522 537 556
rect 503 454 537 488
rect 503 386 537 420
rect 503 318 537 352
rect 503 250 537 284
rect 503 182 537 216
rect 503 114 537 148
<< nsubdiff >>
rect 36 658 94 704
rect 36 624 48 658
rect 82 624 94 658
rect 36 590 94 624
rect 36 556 48 590
rect 82 556 94 590
rect 36 522 94 556
rect 36 488 48 522
rect 82 488 94 522
rect 36 454 94 488
rect 36 420 48 454
rect 82 420 94 454
rect 36 386 94 420
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 602 658 660 704
rect 602 624 614 658
rect 648 624 660 658
rect 602 590 660 624
rect 602 556 614 590
rect 648 556 660 590
rect 602 522 660 556
rect 602 488 614 522
rect 648 488 660 522
rect 602 454 660 488
rect 602 420 614 454
rect 648 420 660 454
rect 602 386 660 420
rect 602 352 614 386
rect 648 352 660 386
rect 602 318 660 352
rect 602 284 614 318
rect 648 284 660 318
rect 602 250 660 284
rect 602 216 614 250
rect 648 216 660 250
rect 602 182 660 216
rect 602 148 614 182
rect 648 148 660 182
rect 602 102 660 148
<< nsubdiffcont >>
rect 48 624 82 658
rect 48 556 82 590
rect 48 488 82 522
rect 48 420 82 454
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 614 624 648 658
rect 614 556 648 590
rect 614 488 648 522
rect 614 420 648 454
rect 614 352 648 386
rect 614 284 648 318
rect 614 216 648 250
rect 614 148 648 182
<< poly >>
rect 179 786 517 806
rect 179 752 195 786
rect 229 752 263 786
rect 297 752 331 786
rect 365 752 399 786
rect 433 752 467 786
rect 501 752 517 786
rect 179 736 517 752
rect 204 704 234 736
rect 290 704 320 736
rect 376 704 406 736
rect 462 704 492 736
rect 204 70 234 102
rect 290 70 320 102
rect 376 70 406 102
rect 462 70 492 102
rect 179 54 517 70
rect 179 20 195 54
rect 229 20 263 54
rect 297 20 331 54
rect 365 20 399 54
rect 433 20 467 54
rect 501 20 517 54
rect 179 0 517 20
<< polycont >>
rect 195 752 229 786
rect 263 752 297 786
rect 331 752 365 786
rect 399 752 433 786
rect 467 752 501 786
rect 195 20 229 54
rect 263 20 297 54
rect 331 20 365 54
rect 399 20 433 54
rect 467 20 501 54
<< locali >>
rect 179 752 187 786
rect 229 752 259 786
rect 297 752 331 786
rect 365 752 399 786
rect 437 752 467 786
rect 509 752 517 786
rect 159 692 193 708
rect 48 672 82 674
rect 48 600 82 624
rect 48 528 82 556
rect 48 456 82 488
rect 48 386 82 420
rect 48 318 82 350
rect 48 250 82 278
rect 48 182 82 206
rect 48 132 82 134
rect 159 624 193 638
rect 159 556 193 566
rect 159 488 193 494
rect 159 420 193 422
rect 159 384 193 386
rect 159 312 193 318
rect 159 240 193 250
rect 159 168 193 182
rect 159 98 193 114
rect 245 692 279 708
rect 245 624 279 638
rect 245 556 279 566
rect 245 488 279 494
rect 245 420 279 422
rect 245 384 279 386
rect 245 312 279 318
rect 245 240 279 250
rect 245 168 279 182
rect 245 98 279 114
rect 331 692 365 708
rect 331 624 365 638
rect 331 556 365 566
rect 331 488 365 494
rect 331 420 365 422
rect 331 384 365 386
rect 331 312 365 318
rect 331 240 365 250
rect 331 168 365 182
rect 331 98 365 114
rect 417 692 451 708
rect 417 624 451 638
rect 417 556 451 566
rect 417 488 451 494
rect 417 420 451 422
rect 417 384 451 386
rect 417 312 451 318
rect 417 240 451 250
rect 417 168 451 182
rect 417 98 451 114
rect 503 692 537 708
rect 503 624 537 638
rect 503 556 537 566
rect 503 488 537 494
rect 503 420 537 422
rect 503 384 537 386
rect 503 312 537 318
rect 503 240 537 250
rect 503 168 537 182
rect 614 672 648 674
rect 614 600 648 624
rect 614 528 648 556
rect 614 456 648 488
rect 614 386 648 420
rect 614 318 648 350
rect 614 250 648 278
rect 614 182 648 206
rect 614 132 648 134
rect 503 98 537 114
rect 179 20 187 54
rect 229 20 259 54
rect 297 20 331 54
rect 365 20 399 54
rect 437 20 467 54
rect 509 20 517 54
<< viali >>
rect 187 752 195 786
rect 195 752 221 786
rect 259 752 263 786
rect 263 752 293 786
rect 331 752 365 786
rect 403 752 433 786
rect 433 752 437 786
rect 475 752 501 786
rect 501 752 509 786
rect 48 658 82 672
rect 48 638 82 658
rect 48 590 82 600
rect 48 566 82 590
rect 48 522 82 528
rect 48 494 82 522
rect 48 454 82 456
rect 48 422 82 454
rect 48 352 82 384
rect 48 350 82 352
rect 48 284 82 312
rect 48 278 82 284
rect 48 216 82 240
rect 48 206 82 216
rect 48 148 82 168
rect 48 134 82 148
rect 159 658 193 672
rect 159 638 193 658
rect 159 590 193 600
rect 159 566 193 590
rect 159 522 193 528
rect 159 494 193 522
rect 159 454 193 456
rect 159 422 193 454
rect 159 352 193 384
rect 159 350 193 352
rect 159 284 193 312
rect 159 278 193 284
rect 159 216 193 240
rect 159 206 193 216
rect 159 148 193 168
rect 159 134 193 148
rect 245 658 279 672
rect 245 638 279 658
rect 245 590 279 600
rect 245 566 279 590
rect 245 522 279 528
rect 245 494 279 522
rect 245 454 279 456
rect 245 422 279 454
rect 245 352 279 384
rect 245 350 279 352
rect 245 284 279 312
rect 245 278 279 284
rect 245 216 279 240
rect 245 206 279 216
rect 245 148 279 168
rect 245 134 279 148
rect 331 658 365 672
rect 331 638 365 658
rect 331 590 365 600
rect 331 566 365 590
rect 331 522 365 528
rect 331 494 365 522
rect 331 454 365 456
rect 331 422 365 454
rect 331 352 365 384
rect 331 350 365 352
rect 331 284 365 312
rect 331 278 365 284
rect 331 216 365 240
rect 331 206 365 216
rect 331 148 365 168
rect 331 134 365 148
rect 417 658 451 672
rect 417 638 451 658
rect 417 590 451 600
rect 417 566 451 590
rect 417 522 451 528
rect 417 494 451 522
rect 417 454 451 456
rect 417 422 451 454
rect 417 352 451 384
rect 417 350 451 352
rect 417 284 451 312
rect 417 278 451 284
rect 417 216 451 240
rect 417 206 451 216
rect 417 148 451 168
rect 417 134 451 148
rect 503 658 537 672
rect 503 638 537 658
rect 503 590 537 600
rect 503 566 537 590
rect 503 522 537 528
rect 503 494 537 522
rect 503 454 537 456
rect 503 422 537 454
rect 503 352 537 384
rect 503 350 537 352
rect 503 284 537 312
rect 503 278 537 284
rect 503 216 537 240
rect 503 206 537 216
rect 503 148 537 168
rect 503 134 537 148
rect 614 658 648 672
rect 614 638 648 658
rect 614 590 648 600
rect 614 566 648 590
rect 614 522 648 528
rect 614 494 648 522
rect 614 454 648 456
rect 614 422 648 454
rect 614 352 648 384
rect 614 350 648 352
rect 614 284 648 312
rect 614 278 648 284
rect 614 216 648 240
rect 614 206 648 216
rect 614 148 648 168
rect 614 134 648 148
rect 187 20 195 54
rect 195 20 221 54
rect 259 20 263 54
rect 263 20 293 54
rect 331 20 365 54
rect 403 20 433 54
rect 433 20 437 54
rect 475 20 501 54
rect 501 20 509 54
<< metal1 >>
rect 175 786 521 806
rect 175 752 187 786
rect 221 752 259 786
rect 293 752 331 786
rect 365 752 403 786
rect 437 752 475 786
rect 509 752 521 786
rect 175 740 521 752
rect 36 672 94 684
rect 36 638 48 672
rect 82 638 94 672
rect 36 600 94 638
rect 36 566 48 600
rect 82 566 94 600
rect 36 528 94 566
rect 36 494 48 528
rect 82 494 94 528
rect 36 456 94 494
rect 36 422 48 456
rect 82 422 94 456
rect 36 384 94 422
rect 36 350 48 384
rect 82 350 94 384
rect 36 312 94 350
rect 36 278 48 312
rect 82 278 94 312
rect 36 240 94 278
rect 36 206 48 240
rect 82 206 94 240
rect 36 168 94 206
rect 36 134 48 168
rect 82 134 94 168
rect 36 122 94 134
rect 150 672 202 684
rect 150 638 159 672
rect 193 638 202 672
rect 150 600 202 638
rect 150 566 159 600
rect 193 566 202 600
rect 150 528 202 566
rect 150 494 159 528
rect 193 494 202 528
rect 150 456 202 494
rect 150 422 159 456
rect 193 422 202 456
rect 150 384 202 422
rect 150 372 159 384
rect 193 372 202 384
rect 150 312 202 320
rect 150 308 159 312
rect 193 308 202 312
rect 150 244 202 256
rect 150 180 202 192
rect 150 122 202 128
rect 236 678 288 684
rect 236 614 288 626
rect 236 550 288 562
rect 236 494 245 498
rect 279 494 288 498
rect 236 486 288 494
rect 236 422 245 434
rect 279 422 288 434
rect 236 384 288 422
rect 236 350 245 384
rect 279 350 288 384
rect 236 312 288 350
rect 236 278 245 312
rect 279 278 288 312
rect 236 240 288 278
rect 236 206 245 240
rect 279 206 288 240
rect 236 168 288 206
rect 236 134 245 168
rect 279 134 288 168
rect 236 122 288 134
rect 322 672 374 684
rect 322 638 331 672
rect 365 638 374 672
rect 322 600 374 638
rect 322 566 331 600
rect 365 566 374 600
rect 322 528 374 566
rect 322 494 331 528
rect 365 494 374 528
rect 322 456 374 494
rect 322 422 331 456
rect 365 422 374 456
rect 322 384 374 422
rect 322 372 331 384
rect 365 372 374 384
rect 322 312 374 320
rect 322 308 331 312
rect 365 308 374 312
rect 322 244 374 256
rect 322 180 374 192
rect 322 122 374 128
rect 408 678 460 684
rect 408 614 460 626
rect 408 550 460 562
rect 408 494 417 498
rect 451 494 460 498
rect 408 486 460 494
rect 408 422 417 434
rect 451 422 460 434
rect 408 384 460 422
rect 408 350 417 384
rect 451 350 460 384
rect 408 312 460 350
rect 408 278 417 312
rect 451 278 460 312
rect 408 240 460 278
rect 408 206 417 240
rect 451 206 460 240
rect 408 168 460 206
rect 408 134 417 168
rect 451 134 460 168
rect 408 122 460 134
rect 494 672 546 684
rect 494 638 503 672
rect 537 638 546 672
rect 494 600 546 638
rect 494 566 503 600
rect 537 566 546 600
rect 494 528 546 566
rect 494 494 503 528
rect 537 494 546 528
rect 494 456 546 494
rect 494 422 503 456
rect 537 422 546 456
rect 494 384 546 422
rect 494 372 503 384
rect 537 372 546 384
rect 494 312 546 320
rect 494 308 503 312
rect 537 308 546 312
rect 494 244 546 256
rect 494 180 546 192
rect 494 122 546 128
rect 602 672 660 684
rect 602 638 614 672
rect 648 638 660 672
rect 602 600 660 638
rect 602 566 614 600
rect 648 566 660 600
rect 602 528 660 566
rect 602 494 614 528
rect 648 494 660 528
rect 602 456 660 494
rect 602 422 614 456
rect 648 422 660 456
rect 602 384 660 422
rect 602 350 614 384
rect 648 350 660 384
rect 602 312 660 350
rect 602 278 614 312
rect 648 278 660 312
rect 602 240 660 278
rect 602 206 614 240
rect 648 206 660 240
rect 602 168 660 206
rect 602 134 614 168
rect 648 134 660 168
rect 602 122 660 134
rect 175 54 521 66
rect 175 20 187 54
rect 221 20 259 54
rect 293 20 331 54
rect 365 20 403 54
rect 437 20 475 54
rect 509 20 521 54
rect 175 0 521 20
<< via1 >>
rect 150 350 159 372
rect 159 350 193 372
rect 193 350 202 372
rect 150 320 202 350
rect 150 278 159 308
rect 159 278 193 308
rect 193 278 202 308
rect 150 256 202 278
rect 150 240 202 244
rect 150 206 159 240
rect 159 206 193 240
rect 193 206 202 240
rect 150 192 202 206
rect 150 168 202 180
rect 150 134 159 168
rect 159 134 193 168
rect 193 134 202 168
rect 150 128 202 134
rect 236 672 288 678
rect 236 638 245 672
rect 245 638 279 672
rect 279 638 288 672
rect 236 626 288 638
rect 236 600 288 614
rect 236 566 245 600
rect 245 566 279 600
rect 279 566 288 600
rect 236 562 288 566
rect 236 528 288 550
rect 236 498 245 528
rect 245 498 279 528
rect 279 498 288 528
rect 236 456 288 486
rect 236 434 245 456
rect 245 434 279 456
rect 279 434 288 456
rect 322 350 331 372
rect 331 350 365 372
rect 365 350 374 372
rect 322 320 374 350
rect 322 278 331 308
rect 331 278 365 308
rect 365 278 374 308
rect 322 256 374 278
rect 322 240 374 244
rect 322 206 331 240
rect 331 206 365 240
rect 365 206 374 240
rect 322 192 374 206
rect 322 168 374 180
rect 322 134 331 168
rect 331 134 365 168
rect 365 134 374 168
rect 322 128 374 134
rect 408 672 460 678
rect 408 638 417 672
rect 417 638 451 672
rect 451 638 460 672
rect 408 626 460 638
rect 408 600 460 614
rect 408 566 417 600
rect 417 566 451 600
rect 451 566 460 600
rect 408 562 460 566
rect 408 528 460 550
rect 408 498 417 528
rect 417 498 451 528
rect 451 498 460 528
rect 408 456 460 486
rect 408 434 417 456
rect 417 434 451 456
rect 451 434 460 456
rect 494 350 503 372
rect 503 350 537 372
rect 537 350 546 372
rect 494 320 546 350
rect 494 278 503 308
rect 503 278 537 308
rect 537 278 546 308
rect 494 256 546 278
rect 494 240 546 244
rect 494 206 503 240
rect 503 206 537 240
rect 537 206 546 240
rect 494 192 546 206
rect 494 168 546 180
rect 494 134 503 168
rect 503 134 537 168
rect 537 134 546 168
rect 494 128 546 134
<< metal2 >>
rect 10 678 686 684
rect 10 626 236 678
rect 288 626 408 678
rect 460 626 686 678
rect 10 614 686 626
rect 10 562 236 614
rect 288 562 408 614
rect 460 562 686 614
rect 10 550 686 562
rect 10 498 236 550
rect 288 498 408 550
rect 460 498 686 550
rect 10 486 686 498
rect 10 434 236 486
rect 288 434 408 486
rect 460 434 686 486
rect 10 428 686 434
rect 10 372 686 378
rect 10 320 150 372
rect 202 320 322 372
rect 374 320 494 372
rect 546 320 686 372
rect 10 308 686 320
rect 10 256 150 308
rect 202 256 322 308
rect 374 256 494 308
rect 546 256 686 308
rect 10 244 686 256
rect 10 192 150 244
rect 202 192 322 244
rect 374 192 494 244
rect 546 192 686 244
rect 10 180 686 192
rect 10 128 150 180
rect 202 128 322 180
rect 374 128 494 180
rect 546 128 686 180
rect 10 122 686 128
<< labels >>
flabel comment s 176 403 176 403 0 FreeSans 300 0 0 0 S
flabel comment s 262 403 262 403 0 FreeSans 300 0 0 0 S
flabel comment s 348 403 348 403 0 FreeSans 300 0 0 0 S
flabel comment s 434 403 434 403 0 FreeSans 300 0 0 0 S
flabel comment s 176 403 176 403 0 FreeSans 300 0 0 0 S
flabel comment s 262 403 262 403 0 FreeSans 300 0 0 0 D
flabel comment s 348 403 348 403 0 FreeSans 300 0 0 0 S
flabel comment s 434 403 434 403 0 FreeSans 300 0 0 0 D
flabel comment s 520 403 520 403 0 FreeSans 300 0 0 0 S
flabel metal1 s 319 761 377 786 0 FreeSans 100 0 0 0 GATE
port 3 nsew
flabel metal1 s 319 25 377 50 0 FreeSans 100 0 0 0 GATE
port 3 nsew
flabel metal1 s 614 397 648 408 0 FreeSans 100 0 0 0 BULK
port 1 nsew
flabel metal1 s 48 397 82 408 0 FreeSans 100 0 0 0 BULK
port 1 nsew
flabel metal2 s 16 213 30 276 0 FreeSans 100 0 0 0 SOURCE
port 4 nsew
flabel metal2 s 16 548 31 614 0 FreeSans 100 0 0 0 DRAIN
port 2 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 9494580
string GDS_START 9479142
<< end >>
