* SPICE NETLIST
***************************************

.SUBCKT drainOnly g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_g5v0d16v0 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_g5v0d16v0 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_var_lvt pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_var_hvt pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_var pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield_o1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield_o1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield_o1nhv pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield_o1phv pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_02p9x06p1_m1m2m3m4_shieldl1_fingercap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_05p9x05p9_m1m2m3m4_shieldl1_wafflecap pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_11p3x11p3_m1m2m3m4_shieldl1_wafflecap pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_02p7x41p1_m1m2m3m4_shieldl1_fingercap pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_02p7x21p1_m1m2m3m4_shieldl1_fingercap pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_02p7x11p1_m1m2m3m4_shieldl1_fingercap pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_02p7x06p1_m1m2m3m4_shieldl1_fingercap pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_55p8x23p1_pol1m1m2m3m4m5_noshield_m5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_55p8x23p1_pol1m1m2m3m4m5_noshield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_55p8x11p7_pol1m1m2m3m4m5_noshield_m5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_55p8x11p7_pol1m1m2m3m4m5_noshield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_44p7x23p1_pol1m1m2m3m4m5_noshield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_44p7x11p7_pol1m1m2m3m4m5_noshield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_33p6x23p1_pol1m1m2m3m4m5_noshield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_33p6x11p7_pol1m1m2m3m4m5_noshield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_22p5x23p1_pol1m1m2m3m4m5_noshield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_22p5x11p7_pol1m1m2m3m4m5_noshield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_11p5x23p1_pol1m1m2m3m4m5_noshield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_pol1m1m2m3m4m5_noshield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_11p3x11p8_l1m1m2m3m4_shieldm5_nhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5_x pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_04p4x04p6_m1m2m3_shieldl1m5_floatm4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1m5_floatm4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1m5_floatm4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldm5 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_06p8x06p1_m1m2m3_shieldl1m4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2m3_shieldpom4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldpom4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldm4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_01p8x01p8_m1m2_noshield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_04p4x04p6_m1m2m3_shieldl1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_shieldpom3 c0 c1 b term4
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3 c0 c1 b term4
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_shieldpo_floatm3 c0 c1 b term4
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_03p9x03p9_m1m2_shieldl1_floatm3 c0 c1 b term4
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldm5 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_m1m4_noshield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_noshield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_02p4x04p6_m1m2_noshield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield_o2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_noshield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT sky130_fd_pr__ind_04 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_55959141808669 2 3
**
R0 2 3 sky130_fd_pr__res_generic_po W=0.33 m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1__example_55959141808662
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1__example_55959141808663
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd__example_5595914180851
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__model__nfet_highvoltage__example_55959141808664 1 2
**
XM0 1 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__sio_clamp_pcap_4x5 1 2
**
X0 1 2 sky130_fd_pr__model__nfet_highvoltage__example_55959141808664
.ENDS
***************************************
.SUBCKT sky130_fd_io__esd_rcclamp_nfetcap 1 2
**
XM0 1 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=8 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd__example_55959141808678
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd2__example_55959141808679
**
.ENDS
***************************************
.SUBCKT ICV_1
**
.ENDS
***************************************
.SUBCKT ICV_2
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808677 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM1 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM2 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM3 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM4 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM5 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM6 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM7 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM8 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM9 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM10 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM11 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM12 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM13 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM14 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
.ENDS
***************************************
.SUBCKT ICV_3 1 2
**
X0 1 2 sky130_fd_io__esd_rcclamp_nfetcap
X1 1 2 sky130_fd_io__esd_rcclamp_nfetcap
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s__example_55959141808671
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s2__example_55959141808672
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808670 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM1 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM2 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM3 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM4 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM5 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM6 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM7 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM8 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM9 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM10 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM11 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM12 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM13 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM14 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM15 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM16 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM17 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s__example_55959141808675
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s2__example_55959141808676
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808674 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
XM1 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
XM2 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
XM3 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
XM4 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
XM5 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
XM6 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
XM7 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
XM8 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
XM9 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
XM10 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
XM11 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
XM12 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
XM13 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
XM14 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
XM15 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
XM16 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
XM17 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
XM18 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
XM19 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
XM20 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
XM21 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808673 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM1 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM2 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM3 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM4 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM5 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM6 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM7 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM8 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM9 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM10 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM11 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM12 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM13 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM14 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM15 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM16 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM17 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM18 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM19 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM20 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
XM21 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_55959141808668 2 3
**
R0 2 3 sky130_fd_pr__res_generic_po W=0.33 m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd__example_55959141808336
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd2__example_55959141808666
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_4
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_5
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_6
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_7
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808665 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM1 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM2 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM3 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM4 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM5 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM6 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM7 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM8 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM9 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM10 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM11 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM12 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM13 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM14 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM15 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM16 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM17 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM18 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM19 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM20 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM21 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM22 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM23 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM24 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM25 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM26 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM27 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM28 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM29 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM30 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM31 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM32 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM33 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM34 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM35 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM36 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM37 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM38 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM39 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM40 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM41 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM42 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM43 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM44 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM45 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM46 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM47 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM48 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM49 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_55959141808667 2 3
**
R0 2 3 sky130_fd_pr__res_generic_po W=0.33 m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_io__top_power_hvc_wpadv2 VSSD SRC_BDY_HVC DRN_HVC VDDIO P_CORE P_PAD
**
*.CALIBRE ISOLATED NETS: OGC_HVC VCCHIB VCCD VDDA VSSIO VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
R0 P_CORE P_PAD sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
X1 SRC_BDY_HVC VDDIO condiode m=1
X2 SRC_BDY_HVC VDDIO condiode m=1
X3 SRC_BDY_HVC VDDIO condiode m=1
X4 SRC_BDY_HVC VDDIO condiode m=1
X5 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X6 SRC_BDY_HVC VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X7 SRC_BDY_HVC VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X8 SRC_BDY_HVC VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X9 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2dn m=1
X10 VSSD DRN_HVC sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X11 19 20 sky130_fd_pr__res_bent_po__example_55959141808669
X83 SRC_BDY_HVC 19 sky130_fd_pr__model__nfet_highvoltage__example_55959141808664
X84 SRC_BDY_HVC 19 sky130_fd_io__sio_clamp_pcap_4x5
X85 SRC_BDY_HVC 19 sky130_fd_io__sio_clamp_pcap_4x5
X86 SRC_BDY_HVC 19 sky130_fd_io__sio_clamp_pcap_4x5
X87 SRC_BDY_HVC 19 sky130_fd_io__sio_clamp_pcap_4x5
X88 SRC_BDY_HVC 19 sky130_fd_io__esd_rcclamp_nfetcap
X89 SRC_BDY_HVC 19 sky130_fd_io__esd_rcclamp_nfetcap
X90 SRC_BDY_HVC 19 sky130_fd_io__esd_rcclamp_nfetcap
X91 SRC_BDY_HVC 19 21 sky130_fd_pr__nfet_01v8__example_55959141808677
X92 SRC_BDY_HVC 19 ICV_3
X93 SRC_BDY_HVC 19 ICV_3
X94 SRC_BDY_HVC 19 ICV_3
X95 SRC_BDY_HVC 19 ICV_3
X96 SRC_BDY_HVC 19 ICV_3
X97 SRC_BDY_HVC 19 ICV_3
X98 SRC_BDY_HVC 21 DRN_HVC sky130_fd_pr__nfet_01v8__example_55959141808670
X99 SRC_BDY_HVC 21 DRN_HVC sky130_fd_pr__nfet_01v8__example_55959141808670
X100 SRC_BDY_HVC 21 DRN_HVC sky130_fd_pr__nfet_01v8__example_55959141808670
X101 SRC_BDY_HVC 21 DRN_HVC sky130_fd_pr__nfet_01v8__example_55959141808674
X102 SRC_BDY_HVC 21 DRN_HVC sky130_fd_pr__nfet_01v8__example_55959141808673
X103 SRC_BDY_HVC 21 DRN_HVC sky130_fd_pr__nfet_01v8__example_55959141808673
X104 SRC_BDY_HVC 21 DRN_HVC sky130_fd_pr__nfet_01v8__example_55959141808673
X105 DRN_HVC 18 sky130_fd_pr__res_bent_po__example_55959141808668
X106 DRN_HVC 19 21 sky130_fd_pr__pfet_01v8__example_55959141808665
X107 18 20 sky130_fd_pr__res_bent_po__example_55959141808667
.ENDS
***************************************
.SUBCKT sky130_ef_io__vdda_hvc_clamped_pad VSSD VSSA VDDIO VDDA 13
**
*.CALIBRE ISOLATED NETS: VCCHIB VCCD VSSIO VSWITCH AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
X0 VSSD VSSA VDDA VDDIO VDDA 13 sky130_fd_io__top_power_hvc_wpadv2
*.CALIBRE WARNING OPEN Open circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT sky130_fd_io__top_ground_hvc_wpad VSSD SRC_BDY_HVC DRN_HVC VDDIO G_CORE G_PAD
**
*.CALIBRE ISOLATED NETS: OGC_HVC VCCHIB VCCD VDDA VSSIO VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
R0 G_CORE G_PAD sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
X1 SRC_BDY_HVC VDDIO condiode m=1
X2 SRC_BDY_HVC VDDIO condiode m=1
X3 SRC_BDY_HVC VDDIO condiode m=1
X4 SRC_BDY_HVC VDDIO condiode m=1
X5 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X6 SRC_BDY_HVC VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X7 SRC_BDY_HVC VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X8 SRC_BDY_HVC VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X9 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2dn m=1
X10 VSSD DRN_HVC sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X11 18 20 sky130_fd_pr__res_bent_po__example_55959141808669
X83 SRC_BDY_HVC 18 sky130_fd_pr__model__nfet_highvoltage__example_55959141808664
X84 SRC_BDY_HVC 18 sky130_fd_io__sio_clamp_pcap_4x5
X85 SRC_BDY_HVC 18 sky130_fd_io__sio_clamp_pcap_4x5
X86 SRC_BDY_HVC 18 sky130_fd_io__sio_clamp_pcap_4x5
X87 SRC_BDY_HVC 18 sky130_fd_io__sio_clamp_pcap_4x5
X88 SRC_BDY_HVC 18 sky130_fd_io__esd_rcclamp_nfetcap
X89 SRC_BDY_HVC 18 sky130_fd_io__esd_rcclamp_nfetcap
X90 SRC_BDY_HVC 18 sky130_fd_io__esd_rcclamp_nfetcap
X91 SRC_BDY_HVC 18 19 sky130_fd_pr__nfet_01v8__example_55959141808677
X92 SRC_BDY_HVC 18 ICV_3
X93 SRC_BDY_HVC 18 ICV_3
X94 SRC_BDY_HVC 18 ICV_3
X95 SRC_BDY_HVC 18 ICV_3
X96 SRC_BDY_HVC 18 ICV_3
X97 SRC_BDY_HVC 18 ICV_3
X98 SRC_BDY_HVC 19 DRN_HVC sky130_fd_pr__nfet_01v8__example_55959141808670
X99 SRC_BDY_HVC 19 DRN_HVC sky130_fd_pr__nfet_01v8__example_55959141808670
X100 SRC_BDY_HVC 19 DRN_HVC sky130_fd_pr__nfet_01v8__example_55959141808670
X101 SRC_BDY_HVC 19 DRN_HVC sky130_fd_pr__nfet_01v8__example_55959141808674
X102 SRC_BDY_HVC 19 DRN_HVC sky130_fd_pr__nfet_01v8__example_55959141808673
X103 SRC_BDY_HVC 19 DRN_HVC sky130_fd_pr__nfet_01v8__example_55959141808673
X104 SRC_BDY_HVC 19 DRN_HVC sky130_fd_pr__nfet_01v8__example_55959141808673
X105 DRN_HVC 21 sky130_fd_pr__res_bent_po__example_55959141808668
X106 DRN_HVC 18 19 sky130_fd_pr__pfet_01v8__example_55959141808665
X107 21 20 sky130_fd_pr__res_bent_po__example_55959141808667
.ENDS
***************************************
.SUBCKT sky130_ef_io__vssa_hvc_clamped_pad VSSD VDDIO VSSA VDDA 13
**
*.CALIBRE ISOLATED NETS: VCCHIB VCCD VSSIO VSWITCH AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
X0 VSSD VSSA VDDA VDDIO VSSA 13 sky130_fd_io__top_ground_hvc_wpad
*.CALIBRE WARNING OPEN Open circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_55959141808692 2 3
**
R0 3 2 sky130_fd_pr__res_generic_po W=0.33 m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808687 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 m=1
XM1 2 3 4 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 m=1
XM2 4 3 2 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 m=1
XM3 2 3 4 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 m=1
XM4 4 3 2 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 m=1
XM5 2 3 4 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 m=1
XM6 4 3 2 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 m=1
XM7 2 3 4 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 m=1
XM8 4 3 2 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 m=1
XM9 2 3 4 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1__example_55959141808682
**
.ENDS
***************************************
.SUBCKT ICV_8
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1__example_55959141808681
**
.ENDS
***************************************
.SUBCKT ICV_9
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_55959141808691 2 3
**
R0 3 2 sky130_fd_pr__res_generic_po W=0.33 m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd__example_55959141808700
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd2__example_55959141808559
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808699 1 2
**
XM0 1 2 1 1 sky130_fd_pr__nfet_01v8 L=8 W=7 m=1
XM1 1 2 1 1 sky130_fd_pr__nfet_01v8 L=8 W=7 m=1
XM2 1 2 1 1 sky130_fd_pr__nfet_01v8 L=8 W=7 m=1
XM3 1 2 1 1 sky130_fd_pr__nfet_01v8 L=8 W=7 m=1
XM4 1 2 1 1 sky130_fd_pr__nfet_01v8 L=8 W=7 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dftpl1s2__example_55959141808702
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808704 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM1 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM2 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM3 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM4 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM5 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM6 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM7 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM8 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM9 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM10 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM11 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM12 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM13 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM14 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM15 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM16 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM17 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM18 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM19 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
X20 1 1 sky130_fd_pr__diode_pw2nd_05v5 m=1
X21 1 1 sky130_fd_pr__diode_pw2nd_05v5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dftpl1s2__example_55959141808694
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808695 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM1 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM2 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM3 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM4 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM5 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM6 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM7 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM8 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM9 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM10 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM11 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM12 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM13 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM14 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM15 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM16 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM17 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM18 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM19 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
X20 1 1 sky130_fd_pr__diode_pw2nd_05v5 m=1
X21 1 1 sky130_fd_pr__diode_pw2nd_05v5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808696 1 2 3
**
XM0 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd2__example_55959141808378
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808698 1 2
**
XM0 1 2 1 1 sky130_fd_pr__nfet_01v8 L=8 W=5 m=1
XM1 1 2 1 1 sky130_fd_pr__nfet_01v8 L=8 W=5 m=1
XM2 1 2 1 1 sky130_fd_pr__nfet_01v8 L=8 W=5 m=1
XM3 1 2 1 1 sky130_fd_pr__nfet_01v8 L=8 W=5 m=1
XM4 1 2 1 1 sky130_fd_pr__nfet_01v8 L=8 W=5 m=1
XM5 1 2 1 1 sky130_fd_pr__nfet_01v8 L=8 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__tpl1__example_55959141808685
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__tpl1__example_55959141808686
**
.ENDS
***************************************
.SUBCKT sky130_fd_io__gnd2gnd_tap
**
.ENDS
***************************************
.SUBCKT sky130_fd_io__gnd2gnd_diff
**
.ENDS
***************************************
.SUBCKT sky130_fd_io__gnd2gnd_sub_dnwl 1 2
**
X0 1 2 sky130_fd_pr__model__parasitic__diode_ps2nw m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gnd2gnd_120x2_lv_isosub VSUB VSSI VSS_N
**
XD0 VSS_N VSSI sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
XD1 VSS_N VSSI sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
XD2 VSS_N VSSI sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
XD3 VSS_N VSSI sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
XD4 VSSI VSS_N sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
XD5 VSSI VSS_N sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
XD6 VSSI VSS_N sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
XD7 VSSI VSS_N sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
X8 VSUB VSSI sky130_fd_io__gnd2gnd_sub_dnwl
X9 VSUB VSS_N sky130_fd_io__gnd2gnd_sub_dnwl
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808701 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM1 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM2 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM3 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM4 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM5 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM6 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM7 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM8 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM9 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM10 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM11 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM12 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM13 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM14 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM15 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM16 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM17 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM18 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM19 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM20 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM21 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM22 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM23 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM24 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM25 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM26 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM27 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM28 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM29 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM30 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM31 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM32 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM33 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM34 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM35 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
X36 1 1 sky130_fd_pr__diode_pw2nd_05v5 m=1
X37 1 1 sky130_fd_pr__diode_pw2nd_05v5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808703 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM1 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM2 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM3 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM4 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM5 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM6 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM7 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM8 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM9 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM10 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM11 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM12 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM13 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM14 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM15 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM16 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM17 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM18 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM19 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM20 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM21 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM22 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM23 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
X24 1 1 sky130_fd_pr__diode_pw2nd_05v5 m=1
X25 1 1 sky130_fd_pr__diode_pw2nd_05v5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808705 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM1 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM2 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM3 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM4 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM5 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM6 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM7 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM8 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM9 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM10 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM11 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM12 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM13 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM14 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM15 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM16 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM17 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM18 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM19 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM20 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM21 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM22 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM23 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM24 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM25 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM26 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM27 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM28 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM29 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM30 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM31 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM32 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM33 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM34 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM35 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM36 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
XM37 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 m=1
X38 1 1 sky130_fd_pr__diode_pw2nd_05v5 m=1
X39 1 1 sky130_fd_pr__diode_pw2nd_05v5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808693 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM1 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM2 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM3 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM4 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM5 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM6 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM7 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM8 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM9 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM10 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM11 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM12 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM13 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM14 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM15 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM16 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM17 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM18 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM19 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM20 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM21 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM22 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM23 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM24 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM25 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM26 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM27 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM28 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM29 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM30 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM31 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM32 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM33 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM34 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM35 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM36 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
XM37 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 m=1
X38 1 1 sky130_fd_pr__diode_pw2nd_05v5 m=1
X39 1 1 sky130_fd_pr__diode_pw2nd_05v5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808697 1 2
**
XM0 1 2 1 1 sky130_fd_pr__nfet_01v8 L=4 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_55959141808688 2 3
**
R0 2 3 sky130_fd_pr__res_generic_po W=0.33 m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_55959141808690 2 3
**
R0 3 2 sky130_fd_pr__res_generic_po W=0.33 m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_io__top_power_lvc_wpad VSSD SRC_BDY_LVC2 SRC_BDY_LVC1 DRN_LVC1 VDDIO DRN_LVC2 BDY2_B2B P_CORE P_PAD
**
*.CALIBRE ISOLATED NETS: OGC_LVC VCCHIB VCCD VDDA VSSIO VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
R0 P_CORE P_PAD sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
X1 SRC_BDY_LVC1 VDDIO condiode m=1
X2 SRC_BDY_LVC2 VDDIO condiode m=1
X3 SRC_BDY_LVC1 VDDIO condiode m=1
R4 DRN_LVC1 21 sky130_fd_pr__res_generic_po W=0.33 m=1 w=480000u l=45000u
X5 SRC_BDY_LVC1 VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X6 SRC_BDY_LVC2 VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X7 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2dn m=1
X8 VSSD DRN_LVC1 sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X9 VSSD DRN_LVC2 sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X10 27 DRN_LVC2 sky130_fd_pr__res_bent_po__example_55959141808692
X11 DRN_LVC1 21 24 sky130_fd_pr__pfet_01v8__example_55959141808687
X12 DRN_LVC1 21 24 sky130_fd_pr__pfet_01v8__example_55959141808687
X13 DRN_LVC2 23 25 sky130_fd_pr__pfet_01v8__example_55959141808687
X14 DRN_LVC2 23 25 sky130_fd_pr__pfet_01v8__example_55959141808687
X203 23 26 sky130_fd_pr__res_bent_po__example_55959141808691
X204 SRC_BDY_LVC2 23 sky130_fd_pr__nfet_01v8__example_55959141808699
X205 SRC_BDY_LVC2 23 sky130_fd_pr__nfet_01v8__example_55959141808699
X206 SRC_BDY_LVC1 21 sky130_fd_pr__nfet_01v8__example_55959141808699
X207 SRC_BDY_LVC1 21 sky130_fd_pr__nfet_01v8__example_55959141808699
X208 SRC_BDY_LVC1 21 sky130_fd_pr__nfet_01v8__example_55959141808699
X209 SRC_BDY_LVC1 24 DRN_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808704
X210 SRC_BDY_LVC1 24 DRN_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808695
X211 SRC_BDY_LVC2 23 25 sky130_fd_pr__nfet_01v8__example_55959141808696
X212 SRC_BDY_LVC2 23 25 sky130_fd_pr__nfet_01v8__example_55959141808696
X213 SRC_BDY_LVC1 21 24 sky130_fd_pr__nfet_01v8__example_55959141808696
X214 SRC_BDY_LVC1 21 24 sky130_fd_pr__nfet_01v8__example_55959141808696
X215 SRC_BDY_LVC1 21 24 sky130_fd_pr__nfet_01v8__example_55959141808696
X216 SRC_BDY_LVC2 23 sky130_fd_pr__nfet_01v8__example_55959141808698
X217 VSSD BDY2_B2B SRC_BDY_LVC1 sky130_fd_io__gnd2gnd_120x2_lv_isosub
X218 SRC_BDY_LVC1 24 DRN_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808701
X219 SRC_BDY_LVC1 24 DRN_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808703
X220 SRC_BDY_LVC1 24 DRN_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808703
X221 SRC_BDY_LVC1 24 DRN_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808703
X222 SRC_BDY_LVC2 25 DRN_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705
X223 SRC_BDY_LVC2 25 DRN_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705
X224 SRC_BDY_LVC2 25 DRN_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705
X225 SRC_BDY_LVC2 25 DRN_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705
X226 SRC_BDY_LVC1 24 DRN_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808705
X227 SRC_BDY_LVC2 25 DRN_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808693
X228 SRC_BDY_LVC2 23 sky130_fd_pr__nfet_01v8__example_55959141808697
X229 22 26 sky130_fd_pr__res_bent_po__example_55959141808688
X230 27 22 sky130_fd_pr__res_bent_po__example_55959141808690
.ENDS
***************************************
.SUBCKT sky130_ef_io__vccd_lvc_clamped2_pad VSSD VSSA VSSIO VCCD VDDIO 13
**
*.CALIBRE ISOLATED NETS: VCCHIB VDDA VSWITCH AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
X0 VSSD VSSD VSSIO VCCD VDDIO VCCD VSSA VCCD 13 sky130_fd_io__top_power_lvc_wpad
*.CALIBRE WARNING OPEN Open circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT sky130_fd_io__top_ground_lvc_wpad VSSD SRC_BDY_LVC2 SRC_BDY_LVC1 DRN_LVC1 VDDIO DRN_LVC2 BDY2_B2B G_CORE G_PAD
**
*.CALIBRE ISOLATED NETS: OGC_LVC VCCHIB VCCD VDDA VSSIO VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
R0 G_CORE G_PAD sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
X1 SRC_BDY_LVC1 VDDIO condiode m=1
X2 SRC_BDY_LVC2 VDDIO condiode m=1
X3 SRC_BDY_LVC1 VDDIO condiode m=1
R4 DRN_LVC1 21 sky130_fd_pr__res_generic_po W=0.33 m=1 w=480000u l=45000u
X5 SRC_BDY_LVC1 VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X6 SRC_BDY_LVC2 VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X7 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2dn m=1
X8 VSSD DRN_LVC1 sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X9 VSSD DRN_LVC2 sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X10 27 DRN_LVC2 sky130_fd_pr__res_bent_po__example_55959141808692
X11 DRN_LVC1 21 24 sky130_fd_pr__pfet_01v8__example_55959141808687
X12 DRN_LVC1 21 24 sky130_fd_pr__pfet_01v8__example_55959141808687
X13 DRN_LVC2 23 25 sky130_fd_pr__pfet_01v8__example_55959141808687
X14 DRN_LVC2 23 25 sky130_fd_pr__pfet_01v8__example_55959141808687
X203 23 26 sky130_fd_pr__res_bent_po__example_55959141808691
X204 SRC_BDY_LVC2 23 sky130_fd_pr__nfet_01v8__example_55959141808699
X205 SRC_BDY_LVC2 23 sky130_fd_pr__nfet_01v8__example_55959141808699
X206 SRC_BDY_LVC1 21 sky130_fd_pr__nfet_01v8__example_55959141808699
X207 SRC_BDY_LVC1 21 sky130_fd_pr__nfet_01v8__example_55959141808699
X208 SRC_BDY_LVC1 21 sky130_fd_pr__nfet_01v8__example_55959141808699
X209 SRC_BDY_LVC1 24 DRN_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808704
X210 SRC_BDY_LVC1 24 DRN_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808695
X211 SRC_BDY_LVC2 23 25 sky130_fd_pr__nfet_01v8__example_55959141808696
X212 SRC_BDY_LVC2 23 25 sky130_fd_pr__nfet_01v8__example_55959141808696
X213 SRC_BDY_LVC1 21 24 sky130_fd_pr__nfet_01v8__example_55959141808696
X214 SRC_BDY_LVC1 21 24 sky130_fd_pr__nfet_01v8__example_55959141808696
X215 SRC_BDY_LVC1 21 24 sky130_fd_pr__nfet_01v8__example_55959141808696
X216 SRC_BDY_LVC2 23 sky130_fd_pr__nfet_01v8__example_55959141808698
X217 VSSD BDY2_B2B SRC_BDY_LVC1 sky130_fd_io__gnd2gnd_120x2_lv_isosub
X218 SRC_BDY_LVC1 24 DRN_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808701
X219 SRC_BDY_LVC1 24 DRN_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808703
X220 SRC_BDY_LVC1 24 DRN_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808703
X221 SRC_BDY_LVC1 24 DRN_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808703
X222 SRC_BDY_LVC2 25 DRN_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705
X223 SRC_BDY_LVC2 25 DRN_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705
X224 SRC_BDY_LVC2 25 DRN_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705
X225 SRC_BDY_LVC2 25 DRN_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705
X226 SRC_BDY_LVC1 24 DRN_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808705
X227 SRC_BDY_LVC2 25 DRN_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808693
X228 SRC_BDY_LVC2 23 sky130_fd_pr__nfet_01v8__example_55959141808697
X229 22 26 sky130_fd_pr__res_bent_po__example_55959141808688
X230 27 22 sky130_fd_pr__res_bent_po__example_55959141808690
.ENDS
***************************************
.SUBCKT sky130_ef_io__vssd_lvc_clamped2_pad VSSD VSSA VSSIO VCCD VDDIO 13
**
*.CALIBRE ISOLATED NETS: VCCHIB VDDA VSWITCH AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
X0 VSSD VSSD VSSIO VCCD VDDIO VCCD VSSA VSSD 13 sky130_fd_io__top_ground_lvc_wpad
*.CALIBRE WARNING OPEN Open circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808592 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd2__example_55959141808306
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808593 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 m=1
.ENDS
***************************************
.SUBCKT ICV_10
**
.ENDS
***************************************
.SUBCKT sky130_fd_io__res75only_small PAD ROUT
**
R0 PAD ROUT sky130_fd_pr__res_generic_po W=2 m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT ICV_11
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_55959141808251
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfm1sd2__example_55959141808561
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808560 1 2 3 4 5
**
XM0 5 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM1 3 2 5 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM2 5 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM3 4 2 5 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM4 5 2 4 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM5 4 2 5 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM6 5 2 4 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_55959141808563
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_12
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_io__amux_switch_1v2b VSSD 3 6 VDDIO VDDA PG_PAD_VDDIOQ_H_N PG_AMX_VDDA_H_N NG_AMX_VPMP_H NG_PAD_VPMP_H PAD_HV_P0 PAD_HV_P1 AMUXBUS_HV PAD_HV_N2 PAD_HV_N3 PAD_HV_N0 PAD_HV_N1
**
*.SEEDPROM
XM0 PAD_HV_N2 NG_PAD_VPMP_H 6 6 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM1 6 NG_PAD_VPMP_H PAD_HV_N2 6 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM2 PAD_HV_N2 NG_PAD_VPMP_H 6 6 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM3 6 NG_PAD_VPMP_H PAD_HV_N2 6 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM4 PAD_HV_N3 NG_PAD_VPMP_H 6 6 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM5 6 NG_PAD_VPMP_H PAD_HV_N3 6 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM6 PAD_HV_N3 NG_PAD_VPMP_H 6 6 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM7 6 NG_PAD_VPMP_H PAD_HV_N3 6 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 m=1
XM8 3 PG_PAD_VDDIOQ_H_N PAD_HV_P0 VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM9 PAD_HV_P0 PG_PAD_VDDIOQ_H_N 3 VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM10 3 PG_PAD_VDDIOQ_H_N PAD_HV_P0 VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM11 PAD_HV_P1 PG_PAD_VDDIOQ_H_N 3 VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM12 3 PG_PAD_VDDIOQ_H_N PAD_HV_P1 VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM13 PAD_HV_P1 PG_PAD_VDDIOQ_H_N 3 VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM14 3 PG_AMX_VDDA_H_N AMUXBUS_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM15 AMUXBUS_HV PG_AMX_VDDA_H_N 3 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM16 3 PG_AMX_VDDA_H_N AMUXBUS_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM17 AMUXBUS_HV PG_AMX_VDDA_H_N 3 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM18 3 PG_AMX_VDDA_H_N AMUXBUS_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
X19 3 VDDA condiode m=1
X20 6 VDDA condiode m=1
X21 VSSD VDDA sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X22 3 VDDA sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X23 6 VDDA sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X24 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X25 VSSD VDDA sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X31 3 NG_AMX_VPMP_H AMUXBUS_HV AMUXBUS_HV 3 sky130_fd_pr__nfet_01v8__example_55959141808560
X32 3 NG_PAD_VPMP_H PAD_HV_N0 PAD_HV_N1 3 sky130_fd_pr__nfet_01v8__example_55959141808560
X33 6 NG_AMX_VPMP_H 6 6 AMUXBUS_HV sky130_fd_pr__nfet_01v8__example_55959141808560
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd2__example_55959141808178
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd__example_55959141808278
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd2__example_55959141808462
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808583 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 m=1
XM1 3 2 4 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808498 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 m=1
XM1 1 2 3 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808580 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=0.7 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_amux_drvr_ls VGND VPWR_HV IN_B RST_H IN HLD_H_N OUT_H VPWR_LV OUT_H_N 10 11
**
XM0 OUT_H_N HLD_H_N 12 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 m=1
XM1 12 HLD_H_N OUT_H_N VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 m=1
XM2 13 VPWR_LV 10 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
XM3 10 VPWR_LV 13 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
XM4 11 VPWR_LV 12 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
XM5 12 VPWR_LV 11 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
X9 VGND RST_H OUT_H VGND sky130_fd_pr__nfet_01v8__example_55959141808583
X10 VGND HLD_H_N OUT_H 13 sky130_fd_pr__nfet_01v8__example_55959141808583
X11 VGND IN_B 10 sky130_fd_pr__nfet_01v8__example_55959141808498
X12 VGND IN 11 sky130_fd_pr__nfet_01v8__example_55959141808498
X13 VPWR_HV OUT_H OUT_H_N sky130_fd_pr__pfet_01v8__example_55959141808580
X14 VPWR_HV OUT_H_N OUT_H sky130_fd_pr__pfet_01v8__example_55959141808580
.ENDS
***************************************
.SUBCKT sky130_fd_pr__model__pfet_highvoltage__example_55959141808371 2 3 4
**
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__model__nfet_highvoltage__example_55959141808369 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__hvsbt_inv_x1 VGND VPWR 3 OUT
**
X0 VPWR 3 OUT sky130_fd_pr__model__pfet_highvoltage__example_55959141808371
X1 VPWR 3 OUT sky130_fd_pr__model__pfet_highvoltage__example_55959141808371
X2 VGND 3 OUT sky130_fd_pr__model__nfet_highvoltage__example_55959141808369
.ENDS
***************************************
.SUBCKT sky130_fd_pr__model__pfet_highvoltage__example_55959141808421 2 3 4 5 6
**
XM0 5 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
XM1 6 4 5 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__hvsbt_inv_x2 VGND VPWR IN OUT
**
XM0 OUT IN VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
XM1 VGND IN OUT VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
X2 VPWR IN IN OUT VPWR sky130_fd_pr__model__pfet_highvoltage__example_55959141808421
X3 VPWR IN IN OUT VPWR sky130_fd_pr__model__pfet_highvoltage__example_55959141808421
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_amx_inv4 VSSA VDA A Y
**
XM0 Y A VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 m=1
XM1 VSSA A Y VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 m=1
XM2 Y A VDA VDA sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
XM3 VDA A Y VDA sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808570 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd__example_55959141808106
**
.ENDS
***************************************
.SUBCKT sky130_fd_io__amx_inv1 1 2 3 4
**
XM0 4 3 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.75 m=1
XM1 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd__example_5595914180819
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd2__example_5595914180884
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808569 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 m=1
XM1 3 2 4 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 m=1
XM2 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd__example_55959141808242
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808579 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808568 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd__example_55959141808504
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808477 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__pfet_g5v0d10v5 L=1 W=0.42 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808567 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 m=1
XM1 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_amux_drvr VSSD VSSA VDDA VSWITCH VCCD VDDIO_Q 9 10 11 12 13 14 AMUX_EN_VDDA_H_N 16 AMUX_EN_VDDA_H 18 AMUX_EN_VDDIO_H_N 20 21 PD_CSD_VSWITCH_H
+ PU_CSD_VDDIOQ_H_N PGA_AMX_VDDA_H_N PGB_AMX_VDDA_H_N PD_CSD_VSWITCH_H_N NGA_PAD_VSWITCH_H NGA_PAD_VSWITCH_H_N AMUX_EN_VSWITCH_H NGA_AMX_VSWITCH_H NGB_AMX_VSWITCH_H NGB_PAD_VSWITCH_H NGB_PAD_VSWITCH_H_N D_B 35 36 NMIDA_ON_N NMIDA_VCCD NMIDA_VCCD_N AMUX_EN_VDDIO_H 41 42
+ 43 44 45 46 47 PGA_PAD_VDDIOQ_H_N PGB_PAD_VDDIOQ_H_N AMUXBUSA_ON_N AMUX_EN_VSWITCH_H_N AMUXBUSB_ON_N AMUXBUSA_ON AMUXBUSB_ON PU_ON_N PU_ON PD_ON_N PD_ON
**
*.SEEDPROM
XM0 PD_CSD_VSWITCH_H 13 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 m=1
XM1 VSSA VSSA PD_CSD_VSWITCH_H VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 m=1
XM2 PD_CSD_VSWITCH_H AMUX_EN_VDDIO_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 m=1
XM3 PU_CSD_VDDIOQ_H_N 21 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 m=1
XM4 VSSD 21 PU_CSD_VDDIOQ_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 m=1
XM5 PU_CSD_VDDIOQ_H_N 21 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 m=1
XM6 VSSD 21 PU_CSD_VDDIOQ_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 m=1
XM7 PU_CSD_VDDIOQ_H_N 21 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 m=1
XM8 VSSD 21 PU_CSD_VDDIOQ_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 m=1
XM9 PU_CSD_VDDIOQ_H_N 21 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 m=1
XM10 PD_CSD_VSWITCH_H 13 VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 L=2 W=0.75 m=1
XM11 VSWITCH 13 PD_CSD_VSWITCH_H VSWITCH sky130_fd_pr__pfet_g5v0d10v5 L=2 W=0.75 m=1
XM12 PU_CSD_VDDIOQ_H_N 21 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
XM13 VDDIO_Q 21 PU_CSD_VDDIOQ_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
XM14 PU_CSD_VDDIOQ_H_N 21 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
XM15 VDDIO_Q 21 PU_CSD_VDDIOQ_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
XM16 PU_CSD_VDDIOQ_H_N 21 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
XM17 VDDIO_Q 21 PU_CSD_VDDIOQ_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
XM18 PU_CSD_VDDIOQ_H_N 21 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
X19 VSSA VSWITCH sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X20 VSSA VSWITCH sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X21 VSSA VSWITCH sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X22 VSSD VSWITCH sky130_fd_pr__model__parasitic__diode_ps2dn m=1
X23 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X24 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X25 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X26 VSSD VDDIO_Q AMUXBUSA_ON_N AMUX_EN_VDDIO_H_N AMUXBUSA_ON AMUX_EN_VDDIO_H 16 VCCD 14 67 68 sky130_fd_io__gpiov2_amux_drvr_ls
X27 VSSA VSWITCH AMUXBUSA_ON_N AMUX_EN_VSWITCH_H_N AMUXBUSA_ON AMUX_EN_VSWITCH_H 70 VCCD 41 42 69 sky130_fd_io__gpiov2_amux_drvr_ls
X28 VSSA VSWITCH AMUXBUSB_ON_N AMUX_EN_VSWITCH_H_N AMUXBUSB_ON AMUX_EN_VSWITCH_H 72 VCCD 43 44 71 sky130_fd_io__gpiov2_amux_drvr_ls
X29 VSSA VSWITCH PD_ON_N AMUX_EN_VSWITCH_H_N PD_ON AMUX_EN_VSWITCH_H 74 VCCD 13 45 73 sky130_fd_io__gpiov2_amux_drvr_ls
X30 VSSD VDDIO_Q AMUXBUSB_ON_N AMUX_EN_VDDIO_H_N AMUXBUSB_ON AMUX_EN_VDDIO_H 18 VCCD 20 46 75 sky130_fd_io__gpiov2_amux_drvr_ls
X31 VSSD VDDIO_Q PU_ON_N AMUX_EN_VDDIO_H_N PU_ON AMUX_EN_VDDIO_H 21 VCCD 76 47 77 sky130_fd_io__gpiov2_amux_drvr_ls
X32 VSSD VCCD 35 D_B sky130_fd_io__hvsbt_inv_x1
X33 VSSD VCCD NMIDA_VCCD NMIDA_VCCD_N sky130_fd_io__hvsbt_inv_x1
X34 VSSD VCCD 36 35 sky130_fd_io__hvsbt_inv_x2
X35 VSSD VCCD NMIDA_ON_N NMIDA_VCCD sky130_fd_io__hvsbt_inv_x2
X36 VSSA VSWITCH 41 NGA_AMX_VSWITCH_H sky130_fd_io__gpiov2_amx_inv4
X37 VSSA VSWITCH 43 NGB_AMX_VSWITCH_H sky130_fd_io__gpiov2_amx_inv4
X38 VSSA VSWITCH 43 NGB_PAD_VSWITCH_H sky130_fd_io__gpiov2_amx_inv4
X39 VSSA VSWITCH 41 NGA_PAD_VSWITCH_H sky130_fd_io__gpiov2_amx_inv4
X40 VSSD VDDIO_Q 16 PGA_PAD_VDDIOQ_H_N sky130_fd_io__gpiov2_amx_inv4
X41 VSSD VDDIO_Q 18 PGB_PAD_VDDIOQ_H_N sky130_fd_io__gpiov2_amx_inv4
X42 VSSA 9 PGA_AMX_VDDA_H_N sky130_fd_pr__nfet_01v8__example_55959141808570
X43 VSSA AMUX_EN_VDDA_H_N 9 sky130_fd_pr__nfet_01v8__example_55959141808570
X44 VSSA AMUX_EN_VDDA_H_N 10 sky130_fd_pr__nfet_01v8__example_55959141808570
X45 VSSA 10 PGB_AMX_VDDA_H_N sky130_fd_pr__nfet_01v8__example_55959141808570
X46 VSSA VSWITCH PD_CSD_VSWITCH_H PD_CSD_VSWITCH_H_N sky130_fd_io__amx_inv1
X47 VSSA VSWITCH NGA_PAD_VSWITCH_H NGA_PAD_VSWITCH_H_N sky130_fd_io__amx_inv1
X48 VSSA VSWITCH NGB_PAD_VSWITCH_H NGB_PAD_VSWITCH_H_N sky130_fd_io__amx_inv1
X49 VSSA 14 65 9 sky130_fd_pr__nfet_01v8__example_55959141808569
X50 VSSA 16 65 11 sky130_fd_pr__nfet_01v8__example_55959141808569
X51 VSSA 18 66 12 sky130_fd_pr__nfet_01v8__example_55959141808569
X52 VSSA 20 66 10 sky130_fd_pr__nfet_01v8__example_55959141808569
X53 VSSA AMUX_EN_VDDA_H_N NGA_AMX_VSWITCH_H sky130_fd_pr__nfet_01v8__example_55959141808579
X54 VSSA AMUX_EN_VDDA_H_N NGB_AMX_VSWITCH_H sky130_fd_pr__nfet_01v8__example_55959141808579
X55 VSSA AMUX_EN_VDDIO_H_N NGB_PAD_VSWITCH_H sky130_fd_pr__nfet_01v8__example_55959141808579
X56 VSSA AMUX_EN_VDDIO_H_N NGA_PAD_VSWITCH_H sky130_fd_pr__nfet_01v8__example_55959141808579
X57 VSSA AMUX_EN_VDDA_H 65 sky130_fd_pr__nfet_01v8__example_55959141808568
X58 VSSA AMUX_EN_VDDA_H 66 sky130_fd_pr__nfet_01v8__example_55959141808568
X63 VDDA 11 9 sky130_fd_pr__pfet_01v8__example_55959141808477
X64 VDDA 12 10 sky130_fd_pr__pfet_01v8__example_55959141808477
X65 VDDA 9 11 sky130_fd_pr__pfet_01v8__example_55959141808477
X66 VDDA 10 12 sky130_fd_pr__pfet_01v8__example_55959141808477
X67 VDDA 9 PGA_AMX_VDDA_H_N sky130_fd_pr__pfet_01v8__example_55959141808567
X68 VDDA 10 PGB_AMX_VDDA_H_N sky130_fd_pr__pfet_01v8__example_55959141808567
*.CALIBRE WARNING OPEN Open circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808465 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808460 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.75 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_amux_ctl_inv_1 VNB VPB IN VPWR OUT VGND
**
*.SEEDPROM
XM0 OUT IN VGND VNB sky130_fd_pr__nfet_01v8 L=0.15 W=0.74 m=1
XM1 OUT IN VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=0.25 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd__example_55959141808476
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808590 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__tap_1
**
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VNB VPB VGND VPWR
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd__example_55959141808115
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808589 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808475 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__model__pfet_highvoltage__example_55959141808588 2 3 4 5
**
*.SEEDPROM
XM0 5 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_amux_ls VSSA VSSD VSWITCH VDDA VDDIO_Q VCCD ENABLE_VDDA_H AMUX_EN_VDDIO_H 15 ENABLE_VSWITCH_H AMUX_EN_VDDIO_H_N 18 19 20 21 HLD_I_H_N HLD_I_H AMUX_EN_VDDA_H_N AMUX_EN_VDDA_H AMUX_EN_VSWITCH_H_N
+ AMUX_EN_VSWITCH_H ANALOG_EN
**
*.SEEDPROM
XM0 35 32 34 VSSD sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 m=1
XM1 34 32 35 VSSD sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 m=1
XM2 35 32 34 VSSD sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 m=1
XM3 34 32 35 VSSD sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 m=1
XM4 36 33 34 VSSD sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 m=1
XM5 34 33 36 VSSD sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 m=1
XM6 36 33 34 VSSD sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 m=1
XM7 34 33 36 VSSD sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 m=1
XM8 18 ENABLE_VDDA_H VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 m=1
XM9 VSSA ENABLE_VSWITCH_H 21 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
XM10 34 HLD_I_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 m=1
XM11 VSSD HLD_I_H_N 34 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 m=1
XM12 34 HLD_I_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 m=1
XM13 VSSD HLD_I_H_N 34 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 m=1
XM14 30 VCCD 36 VSSD sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
XM15 31 VCCD 35 VSSD sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
XM16 36 VCCD 30 VSSD sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
XM17 35 VCCD 31 VSSD sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
XM18 30 VCCD 36 VSSD sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
XM19 31 VCCD 35 VSSD sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
XM20 36 VCCD 30 VSSD sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
XM21 35 VCCD 31 VSSD sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
X22 VSSD VSWITCH sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X23 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X24 VSSD VCCD sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X25 VSWITCH ENABLE_VSWITCH_H ENABLE_VSWITCH_H 21 VSWITCH sky130_fd_pr__model__pfet_highvoltage__example_55959141808421
X26 VSSA 15 AMUX_EN_VDDA_H_N sky130_fd_pr__nfet_01v8__example_55959141808570
X27 VSSA 29 AMUX_EN_VDDA_H sky130_fd_pr__nfet_01v8__example_55959141808570
X28 VSSA 18 15 sky130_fd_pr__nfet_01v8__example_55959141808570
X29 VSSA 20 AMUX_EN_VSWITCH_H sky130_fd_pr__nfet_01v8__example_55959141808570
X30 VSSA 19 AMUX_EN_VSWITCH_H_N sky130_fd_pr__nfet_01v8__example_55959141808570
X31 VSSA 21 19 sky130_fd_pr__nfet_01v8__example_55959141808570
X32 VSSA AMUX_EN_VDDIO_H 37 29 sky130_fd_pr__nfet_01v8__example_55959141808569
X33 VSSA AMUX_EN_VDDIO_H_N 37 15 sky130_fd_pr__nfet_01v8__example_55959141808569
X34 VSSA AMUX_EN_VDDIO_H 38 20 sky130_fd_pr__nfet_01v8__example_55959141808569
X35 VSSA AMUX_EN_VDDIO_H_N 38 19 sky130_fd_pr__nfet_01v8__example_55959141808569
X36 VSWITCH 19 20 sky130_fd_pr__pfet_01v8__example_55959141808477
X37 VDDA 15 29 sky130_fd_pr__pfet_01v8__example_55959141808477
X38 VSWITCH 20 19 sky130_fd_pr__pfet_01v8__example_55959141808477
X39 VDDA 29 15 sky130_fd_pr__pfet_01v8__example_55959141808477
X40 VSSD 31 AMUX_EN_VDDIO_H sky130_fd_pr__nfet_01v8__example_55959141808465
X41 VSSD HLD_I_H 30 sky130_fd_pr__nfet_01v8__example_55959141808465
X42 VSSD 30 AMUX_EN_VDDIO_H_N sky130_fd_pr__nfet_01v8__example_55959141808465
X43 VDDIO_Q 31 30 sky130_fd_pr__pfet_01v8__example_55959141808460
X44 VDDIO_Q 30 31 sky130_fd_pr__pfet_01v8__example_55959141808460
X45 VSSD VCCD 33 VCCD 32 VSSD sky130_fd_io__gpiov2_amux_ctl_inv_1
X46 VSSD VCCD ANALOG_EN VCCD 33 VSSD sky130_fd_io__gpiov2_amux_ctl_inv_1
X47 VDDIO_Q 30 AMUX_EN_VDDIO_H_N sky130_fd_pr__pfet_01v8__example_55959141808590
X48 VDDIO_Q 31 AMUX_EN_VDDIO_H sky130_fd_pr__pfet_01v8__example_55959141808590
X50 VSSA ENABLE_VDDA_H 37 sky130_fd_pr__nfet_01v8__example_55959141808589
X51 VSSA ENABLE_VSWITCH_H 38 sky130_fd_pr__nfet_01v8__example_55959141808589
X52 VDDA 15 AMUX_EN_VDDA_H_N sky130_fd_pr__pfet_01v8__example_55959141808475
X53 VDDA 29 AMUX_EN_VDDA_H sky130_fd_pr__pfet_01v8__example_55959141808475
X54 VSWITCH 19 AMUX_EN_VSWITCH_H_N sky130_fd_pr__pfet_01v8__example_55959141808475
X55 VSWITCH 20 AMUX_EN_VSWITCH_H sky130_fd_pr__pfet_01v8__example_55959141808475
X56 VDDA ENABLE_VDDA_H VDDA 18 sky130_fd_pr__model__pfet_highvoltage__example_55959141808588
X57 VDDA ENABLE_VDDA_H 18 VDDA sky130_fd_pr__model__pfet_highvoltage__example_55959141808588
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd__example_55959141808200
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_55959141808449
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808457 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
XM1 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd__example_55959141808233
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808445 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808450 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
XM1 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808447 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808451 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808248 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_amux_nand5 VGND VPWR OUT IN0 IN4 IN3 IN2 IN1
**
*.SEEDPROM
XM0 VGND 9 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 m=1
XM1 VGND OUT 9 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 m=1
X2 VPWR IN0 OUT sky130_fd_pr__pfet_01v8__example_55959141808457
X3 VGND IN0 10 sky130_fd_pr__nfet_01v8__example_55959141808445
X4 VPWR OUT 9 sky130_fd_pr__pfet_01v8__example_55959141808450
X5 VGND IN4 10 11 sky130_fd_pr__nfet_01v8__example_55959141808447
X6 VGND IN3 11 12 sky130_fd_pr__nfet_01v8__example_55959141808447
X7 VGND IN2 12 13 sky130_fd_pr__nfet_01v8__example_55959141808447
X8 VPWR 9 OUT sky130_fd_pr__pfet_01v8__example_55959141808451
X9 VGND IN1 13 OUT sky130_fd_pr__nfet_01v8__example_55959141808248
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_amux_nand4 VGND VPWR IN0 OUT IN3 IN2 IN1
**
*.SEEDPROM
XM0 VGND 8 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 m=1
XM1 VGND OUT 8 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 m=1
X2 VPWR IN0 OUT sky130_fd_pr__pfet_01v8__example_55959141808457
X3 VGND IN0 9 sky130_fd_pr__nfet_01v8__example_55959141808445
X4 VPWR OUT 8 sky130_fd_pr__pfet_01v8__example_55959141808450
X5 VGND IN3 9 10 sky130_fd_pr__nfet_01v8__example_55959141808447
X6 VGND IN2 10 11 sky130_fd_pr__nfet_01v8__example_55959141808447
X7 VPWR 8 OUT sky130_fd_pr__pfet_01v8__example_55959141808451
X8 VGND IN1 11 OUT sky130_fd_pr__nfet_01v8__example_55959141808248
.ENDS
***************************************
.SUBCKT sky130_fd_io__inv_1 VNB VPB A VPWR Y VGND
**
*.SEEDPROM
XM0 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=0.15 W=0.74 m=1
XM1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1.12 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__nand2_1 VNB VPB B A VPWR Y VGND
**
*.SEEDPROM
XM0 8 B VGND VNB sky130_fd_pr__nfet_01v8 L=0.15 W=0.74 m=1
XM1 Y A 8 VNB sky130_fd_pr__nfet_01v8 L=0.15 W=0.74 m=1
XM2 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1.12 m=1
XM3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1.12 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__model__pfet_highvoltage__example_55959141808420 2 3 4 5
**
XM0 5 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__hvsbt_nor 1 2 IN0 4 5
**
XM0 5 IN0 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
XM1 1 4 5 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
X2 2 IN0 4 6 5 sky130_fd_pr__model__pfet_highvoltage__example_55959141808421
X3 2 IN0 2 6 sky130_fd_pr__model__pfet_highvoltage__example_55959141808420
X4 2 4 5 6 sky130_fd_pr__model__pfet_highvoltage__example_55959141808420
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_559591418085 2 3 4 5
**
XM0 5 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_559591418089 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_559591418087 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__hvsbt_nand2 VGND VPWR IN0 IN1 OUT
**
X0 VPWR IN0 VPWR OUT sky130_fd_pr__pfet_01v8__example_559591418085
X1 VPWR IN0 VPWR OUT sky130_fd_pr__pfet_01v8__example_559591418085
X2 VPWR IN1 OUT VPWR sky130_fd_pr__pfet_01v8__example_559591418085
X3 VPWR IN1 OUT VPWR sky130_fd_pr__pfet_01v8__example_559591418085
X4 VGND IN0 6 sky130_fd_pr__nfet_01v8__example_559591418089
X5 VGND IN1 6 OUT sky130_fd_pr__nfet_01v8__example_559591418087
.ENDS
***************************************
.SUBCKT sky130_fd_io__nor2_1 VNB VPB A B VPWR Y VGND
**
*.SEEDPROM
XM0 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=0.15 W=0.74 m=1
XM1 VGND B Y VNB sky130_fd_pr__nfet_01v8 L=0.15 W=0.74 m=1
XM2 8 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1.12 m=1
XM3 Y B 8 VPB sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1.12 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_amux_decoder VSSD VCCD 5 6 7 ANALOG_SEL 9 10 11 12 AMUXBUSA_ON_N AMUXBUSA_ON 15 PU_ON_N 17 NMIDA_ON_N PU_ON 20 ANALOG_EN D_B
+ 23 PD_ON AMUXBUSB_ON_N PGA_AMX_VDDA_H_N 27 AMUXBUSB_ON PD_ON_N PGA_PAD_VDDIOQ_H_N PGB_AMX_VDDA_H_N 32 33 PGB_PAD_VDDIOQ_H_N NGA_PAD_VSWITCH_H 36 OUT ANALOG_POL NGB_PAD_VSWITCH_H 40 41 NGB_PAD_VSWITCH_H_N
+ NGA_PAD_VSWITCH_H_N PU_VDDIOQ_H_N PD_VSWITCH_H_N 46 NMIDA_VCCD_N
**
*.SEEDPROM
XM0 48 5 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 m=1
XM1 VSSD 6 48 VSSD sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 m=1
XM2 51 6 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 m=1
XM3 7 5 51 VSSD sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 m=1
XM4 VSSD 48 7 VSSD sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 m=1
XM5 49 5 48 VCCD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1.26 m=1
XM6 VCCD 6 49 VCCD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1.26 m=1
XM7 50 6 VCCD VCCD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1.26 m=1
XM8 VCCD 5 50 VCCD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1.26 m=1
XM9 50 48 7 VCCD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1.26 m=1
X10 VSSD VCCD sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X11 VSSD VCCD sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X15 VSSD VCCD 40 41 NGB_PAD_VSWITCH_H_N NGA_PAD_VSWITCH_H_N PGB_PAD_VDDIOQ_H_N PGA_PAD_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_nand5
X16 VSSD VCCD 57 15 NGB_PAD_VSWITCH_H_N NGA_PAD_VSWITCH_H_N PGB_PAD_VDDIOQ_H_N PGA_PAD_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_nand5
X17 VSSD VCCD 10 AMUXBUSB_ON_N 46 PD_VSWITCH_H_N PU_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_nand4
X18 VSSD VCCD 33 AMUXBUSA_ON_N NMIDA_VCCD_N PD_VSWITCH_H_N PU_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_nand4
X19 VSSD VCCD ANALOG_SEL VCCD 52 VSSD sky130_fd_io__inv_1
X20 VSSD VCCD 52 VCCD 9 VSSD sky130_fd_io__inv_1
X21 VSSD VCCD 10 VCCD 12 VSSD sky130_fd_io__inv_1
X22 VSSD VCCD AMUXBUSA_ON_N VCCD AMUXBUSA_ON VSSD sky130_fd_io__inv_1
X23 VSSD VCCD PU_ON VCCD PU_ON_N VSSD sky130_fd_io__inv_1
X24 VSSD VCCD ANALOG_EN VCCD 53 VSSD sky130_fd_io__inv_1
X25 VSSD VCCD PD_ON VCCD PD_ON_N VSSD sky130_fd_io__inv_1
X26 VSSD VCCD AMUXBUSB_ON_N VCCD AMUXBUSB_ON VSSD sky130_fd_io__inv_1
X27 VSSD VCCD 57 VCCD PU_ON VSSD sky130_fd_io__inv_1
X28 VSSD VCCD 33 VCCD 20 VSSD sky130_fd_io__inv_1
X29 VSSD VCCD 36 VCCD 5 VSSD sky130_fd_io__inv_1
X30 VSSD VCCD 58 VCCD 6 VSSD sky130_fd_io__inv_1
X31 VSSD VCCD OUT VCCD 36 VSSD sky130_fd_io__inv_1
X32 VSSD VCCD ANALOG_POL VCCD 58 VSSD sky130_fd_io__inv_1
X33 VSSD VCCD 40 VCCD PD_ON VSSD sky130_fd_io__inv_1
X34 VSSD VCCD 7 52 VCCD 11 VSSD sky130_fd_io__nand2_1
X35 VSSD VCCD 9 7 VCCD 54 VSSD sky130_fd_io__nand2_1
X36 VSSD VCCD 5 6 VCCD 55 VSSD sky130_fd_io__nand2_1
X37 VSSD VCCD 36 58 VCCD 56 VSSD sky130_fd_io__nand2_1
X38 VSSD VCCD NGA_PAD_VSWITCH_H 27 17 sky130_fd_io__hvsbt_nor
X39 VSSD VCCD NGB_PAD_VSWITCH_H 32 23 sky130_fd_io__hvsbt_nor
X40 VSSD VCCD 20 17 NMIDA_ON_N sky130_fd_io__hvsbt_nand2
X41 VSSD VCCD 12 23 D_B sky130_fd_io__hvsbt_nand2
X42 VSSD VCCD PGA_PAD_VDDIOQ_H_N PGA_AMX_VDDA_H_N 27 sky130_fd_io__hvsbt_nand2
X43 VSSD VCCD PGB_PAD_VDDIOQ_H_N PGB_AMX_VDDA_H_N 32 sky130_fd_io__hvsbt_nand2
X44 VSSD VCCD 53 54 VCCD 10 VSSD sky130_fd_io__nor2_1
X45 VSSD VCCD 53 55 VCCD 15 VSSD sky130_fd_io__nor2_1
X46 VSSD VCCD 53 56 VCCD 41 VSSD sky130_fd_io__nor2_1
X47 VSSD VCCD 53 11 VCCD 33 VSSD sky130_fd_io__nor2_1
*.CALIBRE WARNING OPEN Open circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_amux_ctl_logic VSSD VSSA VDDA VSWITCH VCCD 12 13 14 15 VDDIO_Q 17 PGA_AMX_VDDA_H_N NGB_PAD_VSWITCH_H NGA_PAD_VSWITCH_H AMUX_EN_VDDA_H_N PGB_AMX_VDDA_H_N 23 24 D_B 26
+ NMIDA_VCCD 28 ENABLE_VDDA_H ENABLE_VSWITCH_H 31 AMUX_EN_VDDIO_H_N 33 34 35 36 37 38 39 40 PGA_PAD_VDDIOQ_H_N PGB_PAD_VDDIOQ_H_N 43 44 45 46
+ 47 48 49 50 51 52 PD_CSD_VSWITCH_H 54 55 56 NGA_AMX_VSWITCH_H NGB_AMX_VSWITCH_H 59 60 61 62 PU_CSD_VDDIOQ_H_N 64 65 66
+ ANALOG_EN HLD_I_H_N HLD_I_H ANALOG_SEL 71 72 73 74 75 76 77 78 79 OUT ANALOG_POL 82 83 84 85 86
**
X0 VSSD VDDA sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X1 VSSD VCCD sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X2 VSSD VSSA VDDA VSWITCH VCCD VDDIO_Q 54 52 56 51 55 14 AMUX_EN_VDDA_H_N 17 89 61 AMUX_EN_VDDIO_H_N 62 65 PD_CSD_VSWITCH_H
+ PU_CSD_VDDIOQ_H_N PGA_AMX_VDDA_H_N PGB_AMX_VDDA_H_N 13 NGA_PAD_VSWITCH_H 35 34 NGA_AMX_VSWITCH_H NGB_AMX_VSWITCH_H NGB_PAD_VSWITCH_H 23 24 D_B 12 26 NMIDA_VCCD 43 15 60 49
+ 84 50 59 64 66 PGA_PAD_VDDIOQ_H_N PGB_PAD_VDDIOQ_H_N 40 33 45 39 38 46 47 37 36
+ sky130_fd_io__gpiov2_amux_drvr
X3 VSSA VSSD VSWITCH VDDA VDDIO_Q VCCD ENABLE_VDDA_H 15 31 ENABLE_VSWITCH_H AMUX_EN_VDDIO_H_N 28 91 90 88 HLD_I_H_N HLD_I_H AMUX_EN_VDDA_H_N 89 33
+ 34 ANALOG_EN
+ sky130_fd_io__gpiov2_amux_ls
X4 VSSD VCCD 85 72 74 ANALOG_SEL 71 83 92 76 40 39 48 46 73 26 47 75 ANALOG_EN 12
+ 77 36 45 PGA_AMX_VDDA_H_N 78 38 37 PGA_PAD_VDDIOQ_H_N PGB_AMX_VDDA_H_N 79 44 PGB_PAD_VDDIOQ_H_N NGA_PAD_VSWITCH_H 86 OUT ANALOG_POL NGB_PAD_VSWITCH_H 82 87 23
+ 35 PU_CSD_VDDIOQ_H_N 13 24 43
+ sky130_fd_io__gpiov2_amux_decoder
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_amux VSSD VSSIO_Q VSSA 4 5 6 7 VSWITCH VDDIO_Q VDDA HLD_I_H PAD VCCD 15 ENABLE_VDDA_H ENABLE_VSWITCH_H AMUXBUS_B AMUXBUS_A ANALOG_SEL ANALOG_EN
+ OUT ANALOG_POL HLD_I_H_N
**
XM0 36 27 VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
XM1 VSSIO_Q 27 36 VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
XM2 36 27 VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
XM3 VSSIO_Q 27 36 VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
XM4 36 27 VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
XM5 VSSIO_Q 27 36 VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
XM6 37 27 VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
XM7 VSSIO_Q 27 37 VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
XM8 37 27 VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
XM9 VSSIO_Q 27 37 VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
XM10 37 27 VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
XM11 VSSIO_Q 27 37 VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
XM12 37 27 VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
XM13 VSSIO_Q 27 37 VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
XM14 37 25 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 m=1
XM15 VDDIO_Q 25 37 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 m=1
XM16 37 25 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 m=1
XM17 VDDIO_Q 25 37 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 m=1
XM18 36 25 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 m=1
XM19 VDDIO_Q 25 36 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 m=1
XM20 36 25 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 m=1
X21 VSSA VSWITCH condiode m=1
X22 VSSA VSWITCH condiode m=1
X23 VSSA VSWITCH condiode m=1
X24 VSSIO_Q VDDA condiode m=1
X25 VSSA VDDA condiode m=1
X26 VSSIO_Q VDDA condiode m=1
X27 VSSD VDDA sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X28 VSSIO_Q VDDA sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X29 VSSA VDDA sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X30 VSSD VDDA sky130_fd_pr__model__parasitic__diode_ps2dn m=1
X31 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X33 VSSA 28 7 VSSA sky130_fd_pr__nfet_01v8__example_55959141808592
X34 VSSA 28 5 VSSA sky130_fd_pr__nfet_01v8__example_55959141808592
X35 VSSA 28 VSSA 4 sky130_fd_pr__nfet_01v8__example_55959141808592
X36 VSSA 28 VSSA 6 sky130_fd_pr__nfet_01v8__example_55959141808592
X37 VSSA HLD_I_H 4 VSSA sky130_fd_pr__nfet_01v8__example_55959141808592
X38 VSSA HLD_I_H 6 VSSA sky130_fd_pr__nfet_01v8__example_55959141808592
X39 VSSA HLD_I_H VSSA 7 sky130_fd_pr__nfet_01v8__example_55959141808592
X40 VSSA HLD_I_H VSSA 5 sky130_fd_pr__nfet_01v8__example_55959141808592
X41 VSSA 26 41 5 sky130_fd_pr__nfet_01v8__example_55959141808593
X42 VSSA 26 39 6 sky130_fd_pr__nfet_01v8__example_55959141808593
X43 VSSA 29 4 40 sky130_fd_pr__nfet_01v8__example_55959141808593
X44 VSSA 29 38 7 sky130_fd_pr__nfet_01v8__example_55959141808593
X52 PAD 30 sky130_fd_io__res75only_small
X53 31 32 sky130_fd_io__res75only_small
X54 PAD PAD sky130_fd_io__res75only_small
X55 PAD 31 sky130_fd_io__res75only_small
X56 PAD 33 sky130_fd_io__res75only_small
X57 PAD PAD sky130_fd_io__res75only_small
X58 33 34 sky130_fd_io__res75only_small
X59 PAD 35 sky130_fd_io__res75only_small
X60 PAD 36 sky130_fd_io__res75only_small
X61 PAD 37 sky130_fd_io__res75only_small
X62 VSSA 38 sky130_fd_io__res75only_small
X63 VSSA 39 sky130_fd_io__res75only_small
X64 VSSA 40 sky130_fd_io__res75only_small
X65 VSSA 41 sky130_fd_io__res75only_small
X66 VSSD 5 6 VDDIO_Q VDDA 77 15 65 45 30 35 AMUXBUS_B 32 32 34 34 sky130_fd_io__amux_switch_1v2b
X67 VSSD 4 7 VDDIO_Q VDDA 73 57 64 46 30 35 AMUXBUS_A 32 32 34 34 sky130_fd_io__amux_switch_1v2b
X76 VSSD VSSA VDDA VSWITCH VCCD 75 72 42 43 VDDIO_Q 44 57 45 46 47 15 99 48 26 78
+ 29 28 ENABLE_VDDA_H ENABLE_VSWITCH_H 52 68 51 58 74 67 89 54 53 49 73 77 81 96 50 79
+ 97 80 55 56 59 60 27 61 62 63 64 65 66 69 70 71 25 90 92 95
+ ANALOG_EN HLD_I_H_N HLD_I_H ANALOG_SEL 76 82 83 84 85 86 87 88 91 OUT ANALOG_POL 93 94 98 100 101
+ sky130_fd_io__gpiov2_amux_ctl_logic
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em2s_cdns_55959141808438 2 3
**
R0 2 4 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R1 4 3 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em1o_cdns_5595914180880 2 3 4
**
R0 2 3 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R1 5 4 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em1s_cdns_5595914180882 1 2
**
R0 1 3 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R1 3 2 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808620 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.25 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808430 2 3 4 5 6
**
*.SEEDPROM
XM0 5 3 4 2 sky130_fd_pr__pfet_01v8_hvt L=0.25 W=1 m=1
XM1 6 4 5 2 sky130_fd_pr__pfet_01v8_hvt L=0.25 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808116 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808622 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 m=1
XM1 1 2 3 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 m=1
XM2 3 2 1 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 m=1
XM3 1 2 3 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd__example_5595914180811
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_5595914180813 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808624 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808623 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=1 W=0.75 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_5595914180822 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.75 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__com_ctl_lsv2 VGND VCC_IO VPWR HLD_H_N SET_H RST_H IN OUT_H OUT_H_N
**
*.SEEDPROM
XM0 16 VPWR 14 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
XM1 17 VPWR 15 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
XM2 14 VPWR 16 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
XM3 15 VPWR 17 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
XM4 16 VPWR 14 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
XM5 17 VPWR 15 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
XM6 16 VPWR 14 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
XM7 15 VPWR 17 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
X8 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X9 VGND IN 12 sky130_fd_pr__nfet_01v8__example_55959141808620
X10 VGND 12 13 sky130_fd_pr__nfet_01v8__example_55959141808620
X11 VPWR IN 12 VPWR 13 sky130_fd_pr__pfet_01v8__example_55959141808430
X12 VGND HLD_H_N 15 10 sky130_fd_pr__nfet_01v8__example_55959141808116
X13 VGND SET_H VGND 10 sky130_fd_pr__nfet_01v8__example_55959141808116
X14 VGND RST_H VGND 11 sky130_fd_pr__nfet_01v8__example_55959141808116
X15 VGND HLD_H_N 16 11 sky130_fd_pr__nfet_01v8__example_55959141808116
X16 VGND 12 14 sky130_fd_pr__nfet_01v8__example_55959141808622
X17 VGND 13 17 sky130_fd_pr__nfet_01v8__example_55959141808622
X18 VCC_IO 11 OUT_H_N sky130_fd_pr__pfet_01v8__example_5595914180813
X19 VCC_IO 10 OUT_H sky130_fd_pr__pfet_01v8__example_5595914180813
X20 VGND 10 OUT_H sky130_fd_pr__nfet_01v8__example_55959141808624
X21 VGND 11 OUT_H_N sky130_fd_pr__nfet_01v8__example_55959141808624
X22 VGND 11 10 sky130_fd_pr__nfet_01v8__example_55959141808623
X23 VGND 10 11 sky130_fd_pr__nfet_01v8__example_55959141808623
X24 VCC_IO 11 10 sky130_fd_pr__pfet_01v8__example_5595914180822
X25 VCC_IO 10 11 sky130_fd_pr__pfet_01v8__example_5595914180822
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em1o_cdns_5595914180879 1 2
**
R0 1 3 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R1 4 2 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em1s_cdns_5595914180881 1 2
**
R0 1 3 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R1 3 2 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808383 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808382 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808423 1 2 3 4
**
XM0 1 2 4 1 sky130_fd_pr__nfet_01v8 L=0.25 W=1 m=1
XM1 2 3 1 1 sky130_fd_pr__nfet_01v8 L=0.25 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808428 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808424 1 2 3
**
XM0 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=1 W=0.75 m=1
XM1 2 3 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=1 W=0.75 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808429 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808427 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 m=1
XM1 1 2 3 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 m=1
XM2 3 2 1 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 m=1
XM3 1 2 3 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808426 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
XM1 3 2 4 1 sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808432 2 3 4
**
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd__example_55959141808102
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808431 2 3 4
**
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__via_pol1__example_55959141808394
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808380 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808435 2 3 4
**
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.75 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808433 2 3 4
**
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.75 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808379 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__com_ctl_ls_1v2 1 VCC_IO VPB VPWR HLD_H_N IN RST_H SET_H OUT_H_N OUT_H
**
*.SEEDPROM
X0 VPB IN 14 VPWR 13 sky130_fd_pr__pfet_01v8__example_55959141808430
X1 1 SET_H 12 sky130_fd_pr__nfet_01v8__example_55959141808383
X2 1 RST_H 11 sky130_fd_pr__nfet_01v8__example_55959141808382
X3 1 14 IN 13 sky130_fd_pr__nfet_01v8__example_55959141808423
X4 1 HLD_H_N 11 17 sky130_fd_pr__nfet_01v8__example_55959141808428
X5 1 12 11 sky130_fd_pr__nfet_01v8__example_55959141808424
X6 1 HLD_H_N 15 12 sky130_fd_pr__nfet_01v8__example_55959141808429
X7 1 13 16 sky130_fd_pr__nfet_01v8__example_55959141808427
X8 1 14 18 sky130_fd_pr__nfet_01v8__example_55959141808427
X9 1 VPWR 16 15 sky130_fd_pr__nfet_01v8__example_55959141808426
X10 1 VPWR 16 15 sky130_fd_pr__nfet_01v8__example_55959141808426
X11 1 VPWR 18 17 sky130_fd_pr__nfet_01v8__example_55959141808426
X12 1 VPWR 18 17 sky130_fd_pr__nfet_01v8__example_55959141808426
X13 VCC_IO 11 OUT_H_N sky130_fd_pr__pfet_01v8__example_55959141808432
X14 VCC_IO 12 OUT_H sky130_fd_pr__pfet_01v8__example_55959141808431
X16 1 12 OUT_H sky130_fd_pr__nfet_01v8__example_55959141808380
X17 VCC_IO 11 12 sky130_fd_pr__pfet_01v8__example_55959141808435
X18 VCC_IO 12 11 sky130_fd_pr__pfet_01v8__example_55959141808433
X19 1 11 OUT_H_N sky130_fd_pr__nfet_01v8__example_55959141808379
.ENDS
***************************************
.SUBCKT sky130_fd_io__com_ctl_ls_v2 1 VCC_IO VPB VPWR HLD_H_N IN RST_H SET_H OUT_H_N OUT_H
**
*.SEEDPROM
X0 1 VPB sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X1 VPB IN 14 VPWR 13 sky130_fd_pr__pfet_01v8__example_55959141808430
X2 1 SET_H 12 sky130_fd_pr__nfet_01v8__example_55959141808383
X3 1 RST_H 11 sky130_fd_pr__nfet_01v8__example_55959141808382
X4 1 14 IN 13 sky130_fd_pr__nfet_01v8__example_55959141808423
X5 1 HLD_H_N 11 17 sky130_fd_pr__nfet_01v8__example_55959141808428
X6 1 12 11 sky130_fd_pr__nfet_01v8__example_55959141808424
X7 1 HLD_H_N 15 12 sky130_fd_pr__nfet_01v8__example_55959141808429
X8 1 13 16 sky130_fd_pr__nfet_01v8__example_55959141808427
X9 1 14 18 sky130_fd_pr__nfet_01v8__example_55959141808427
X10 1 VPWR 16 15 sky130_fd_pr__nfet_01v8__example_55959141808426
X11 1 VPWR 16 15 sky130_fd_pr__nfet_01v8__example_55959141808426
X12 1 VPWR 18 17 sky130_fd_pr__nfet_01v8__example_55959141808426
X13 1 VPWR 18 17 sky130_fd_pr__nfet_01v8__example_55959141808426
X14 VCC_IO 11 OUT_H_N sky130_fd_pr__pfet_01v8__example_55959141808432
X15 VCC_IO 12 OUT_H sky130_fd_pr__pfet_01v8__example_55959141808431
X17 1 12 OUT_H sky130_fd_pr__nfet_01v8__example_55959141808380
X18 VCC_IO 11 12 sky130_fd_pr__pfet_01v8__example_55959141808435
X19 VCC_IO 12 11 sky130_fd_pr__pfet_01v8__example_55959141808433
X20 1 11 OUT_H_N sky130_fd_pr__nfet_01v8__example_55959141808379
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808617 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_01v8_hvt L=0.25 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__com_ctl_ls_en_1_v2 1 VCC_IO 3 VPWR HLD_H_N DM[1] RST_H SET_H OUT_H_N OUT_H
**
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VPB
X0 1 3 sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X1 1 SET_H 13 sky130_fd_pr__nfet_01v8__example_55959141808383
X2 1 RST_H 12 sky130_fd_pr__nfet_01v8__example_55959141808382
X3 1 15 DM[1] 14 sky130_fd_pr__nfet_01v8__example_55959141808423
X4 1 HLD_H_N 12 18 sky130_fd_pr__nfet_01v8__example_55959141808428
X5 1 13 12 sky130_fd_pr__nfet_01v8__example_55959141808424
X6 1 HLD_H_N 16 13 sky130_fd_pr__nfet_01v8__example_55959141808429
X7 1 14 17 sky130_fd_pr__nfet_01v8__example_55959141808427
X8 1 15 19 sky130_fd_pr__nfet_01v8__example_55959141808427
X9 1 VPWR 17 16 sky130_fd_pr__nfet_01v8__example_55959141808426
X10 1 VPWR 17 16 sky130_fd_pr__nfet_01v8__example_55959141808426
X11 1 VPWR 19 18 sky130_fd_pr__nfet_01v8__example_55959141808426
X12 1 VPWR 19 18 sky130_fd_pr__nfet_01v8__example_55959141808426
X13 VCC_IO 12 OUT_H_N sky130_fd_pr__pfet_01v8__example_55959141808432
X14 VCC_IO 13 OUT_H sky130_fd_pr__pfet_01v8__example_55959141808431
X16 1 13 OUT_H sky130_fd_pr__nfet_01v8__example_55959141808380
X17 VCC_IO 12 13 sky130_fd_pr__pfet_01v8__example_55959141808435
X18 VCC_IO 13 12 sky130_fd_pr__pfet_01v8__example_55959141808433
X19 1 12 OUT_H_N sky130_fd_pr__nfet_01v8__example_55959141808379
X20 3 DM[1] 15 sky130_fd_pr__pfet_01v8__example_55959141808617
X21 3 15 14 sky130_fd_pr__pfet_01v8__example_55959141808617
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_ctl_lsbank VGND VCC_IO VPWR IB_MODE_SEL HLD_I_H_N OD_I_H DM_H[1] DM_H_N[1] DM_H_N[0] DM_H[0] STARTUP_RST_H DM[0] INP_DIS STARTUP_ST_H INP_DIS_H_N DM_H_N[2] DM_H[2] DM[2] VTRIP_SEL_H_N VTRIP_SEL
+ IB_MODE_SEL_H IB_MODE_SEL_H_N DM[1]
**
*.SEEDPROM
X0 VGND VPWR sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X1 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X2 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
R3 OD_I_H 45 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R4 46 33 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
X5 32 OD_I_H sky130_fd_io__tk_em2s_cdns_55959141808438
X6 33 VGND sky130_fd_io__tk_em2s_cdns_55959141808438
X7 OD_I_H 34 35 sky130_fd_io__tk_em1o_cdns_5595914180880
X8 STARTUP_RST_H 36 37 sky130_fd_io__tk_em1o_cdns_5595914180880
X9 38 39 STARTUP_ST_H sky130_fd_io__tk_em1o_cdns_5595914180880
X10 OD_I_H 40 41 sky130_fd_io__tk_em1o_cdns_5595914180880
X11 OD_I_H 42 43 sky130_fd_io__tk_em1o_cdns_5595914180880
X12 VGND 44 32 sky130_fd_io__tk_em1o_cdns_5595914180880
X13 35 VGND sky130_fd_io__tk_em1s_cdns_5595914180882
X14 37 STARTUP_ST_H sky130_fd_io__tk_em1s_cdns_5595914180882
X15 STARTUP_RST_H 38 sky130_fd_io__tk_em1s_cdns_5595914180882
X16 41 VGND sky130_fd_io__tk_em1s_cdns_5595914180882
X17 VGND 43 sky130_fd_io__tk_em1s_cdns_5595914180882
X18 VGND VCC_IO VPWR HLD_I_H_N 33 32 IB_MODE_SEL IB_MODE_SEL_H IB_MODE_SEL_H_N sky130_fd_io__com_ctl_lsv2
X19 VGND 26 sky130_fd_io__tk_em1o_cdns_5595914180879
X20 STARTUP_ST_H 27 sky130_fd_io__tk_em1o_cdns_5595914180879
X21 28 STARTUP_RST_H sky130_fd_io__tk_em1o_cdns_5595914180879
X22 VGND 30 sky130_fd_io__tk_em1o_cdns_5595914180879
X23 VGND 31 sky130_fd_io__tk_em1o_cdns_5595914180879
X24 26 OD_I_H sky130_fd_io__tk_em1s_cdns_5595914180881
X25 27 STARTUP_RST_H sky130_fd_io__tk_em1s_cdns_5595914180881
X26 STARTUP_ST_H 28 sky130_fd_io__tk_em1s_cdns_5595914180881
X27 30 OD_I_H sky130_fd_io__tk_em1s_cdns_5595914180881
X28 OD_I_H 31 sky130_fd_io__tk_em1s_cdns_5595914180881
X29 VGND VCC_IO VPWR VPWR HLD_I_H_N VTRIP_SEL 31 43 VTRIP_SEL_H_N VTRIP_SEL_H sky130_fd_io__com_ctl_ls_1v2
X30 VGND VCC_IO VPWR VPWR HLD_I_H_N DM[0] 27 37 DM_H_N[0] DM_H[0] sky130_fd_io__com_ctl_ls_v2
X31 VGND VCC_IO VPWR VPWR HLD_I_H_N INP_DIS 28 38 INP_DIS_H_N INP_DIS_H sky130_fd_io__com_ctl_ls_v2
X32 VGND VCC_IO VPWR VPWR HLD_I_H_N DM[2] 30 41 DM_H_N[2] DM_H[2] sky130_fd_io__com_ctl_ls_v2
X33 VGND VCC_IO VPWR VPWR HLD_I_H_N DM[1] 26 35 DM_H_N[1] DM_H[1] sky130_fd_io__com_ctl_ls_en_1_v2
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em2s_cdns_55959141808652 2 3
**
R0 2 4 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R1 4 3 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em2o_cdns_55959141808653 2 3
**
R0 2 4 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R1 5 3 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_io__res250only_small PAD ROUT
**
R0 PAD 4 sky130_fd_pr__res_generic_po W=2 m=1 w=480000u l=45000u
R1 4 5 sky130_fd_pr__res_generic_po W=2 m=1 w=480000u l=45000u
R2 5 ROUT sky130_fd_pr__res_generic_po W=2 m=1 w=480000u l=45000u
R3 PAD 4 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R4 5 ROUT sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R5 PAD 4 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R6 5 ROUT sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_pr__via_pol1__example_5595914180854
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__via_pol1_centered__example_559591418080
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_5595914180850 1 2 3
**
XM0 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpio_pddrvr_weakv2 2 3 PD_H PAD
**
*.SEEDPROM
X0 2 3 sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X1 2 PD_H PAD sky130_fd_pr__nfet_01v8__example_5595914180850
X2 2 PD_H PAD sky130_fd_pr__nfet_01v8__example_5595914180850
X3 2 PD_H PAD sky130_fd_pr__nfet_01v8__example_5595914180850
X4 2 PD_H PAD sky130_fd_pr__nfet_01v8__example_5595914180850
X5 2 PD_H PAD sky130_fd_pr__nfet_01v8__example_5595914180850
X6 2 PD_H PAD sky130_fd_pr__nfet_01v8__example_5595914180850
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd__example_55959141808655
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808654 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM1 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM2 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
XM3 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__com_pudrvr_strong_slowv2 2 PU_H_N PAD
**
*.SEEDPROM
X0 2 PU_H_N PAD sky130_fd_pr__pfet_01v8__example_55959141808654
X1 2 PU_H_N PAD sky130_fd_pr__pfet_01v8__example_55959141808654
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_generic_po__example_5595914180864 2 3
**
R0 2 3 sky130_fd_pr__res_generic_po W=0.8 m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_5595914180862 2 3
**
R0 2 3 sky130_fd_pr__res_generic_po W=0.8 m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em1s_cdns_5595914180859 2 3
**
R0 2 4 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R1 4 3 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_5595914180863 2 3
**
R0 2 3 sky130_fd_pr__res_generic_po W=0.8 m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_io__com_res_weak RA 3 4 5 6 7 RB
**
R0 RA 3 sky130_fd_pr__res_generic_po W=0.8 m=1 w=480000u l=45000u
R1 11 4 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R2 12 5 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
X3 6 9 sky130_fd_pr__res_generic_po__example_5595914180864
X4 9 7 sky130_fd_pr__res_generic_po__example_5595914180864
X5 10 RB sky130_fd_pr__res_generic_po__example_5595914180864
X6 7 10 sky130_fd_pr__res_generic_po__example_5595914180864
X7 5 4 sky130_fd_pr__res_bent_po__example_5595914180862
X8 6 5 sky130_fd_pr__res_bent_po__example_5595914180862
X9 5 6 sky130_fd_io__tk_em1s_cdns_5595914180859
X10 6 9 sky130_fd_io__tk_em1s_cdns_5595914180859
X11 9 7 sky130_fd_io__tk_em1s_cdns_5595914180859
X12 10 RB sky130_fd_io__tk_em1s_cdns_5595914180859
X13 7 10 sky130_fd_io__tk_em1s_cdns_5595914180859
X14 4 3 sky130_fd_pr__res_bent_po__example_5595914180863
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd__example_5595914180848
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_5595914180849
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_generic_po__example_5595914180838 2 3
**
R0 2 3 sky130_fd_pr__res_generic_po W=0.5 m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpio_pddrvr_strong_slowv2 2 3 PD_H PAD
**
*.SEEDPROM
X0 2 3 sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X1 2 PD_H PAD sky130_fd_pr__nfet_01v8__example_5595914180850
X2 2 PD_H PAD sky130_fd_pr__nfet_01v8__example_5595914180850
X3 2 PD_H PAD sky130_fd_pr__nfet_01v8__example_5595914180850
X4 2 PD_H PAD sky130_fd_pr__nfet_01v8__example_5595914180850
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s__example_55959141808646
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808647 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
.ENDS
***************************************
.SUBCKT ICV_13
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpm1s2__example_55959141808649
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808648 1 2 3 4 5 6 7 8 9 10 11 12
**
XM0 12 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM1 1 2 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM2 12 3 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM3 1 3 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM4 12 3 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM5 1 4 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM6 12 4 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM7 1 4 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM8 12 5 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM9 1 5 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM10 12 5 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM11 1 6 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM12 12 7 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM13 1 7 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM14 12 7 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM15 1 8 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM16 12 8 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM17 1 8 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM18 12 8 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM19 1 8 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM20 12 8 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM21 1 9 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM22 12 10 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM23 1 11 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM24 12 11 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808651 1 2 3 4 5 6 7 8 9 10 11 12
**
XM0 12 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM1 1 2 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM2 12 3 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM3 1 3 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM4 12 3 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM5 1 4 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM6 12 4 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM7 1 4 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM8 12 5 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM9 1 5 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM10 12 5 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM11 1 6 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM12 12 7 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM13 1 7 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM14 12 7 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM15 1 8 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM16 12 8 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM17 1 8 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM18 12 8 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM19 1 8 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM20 12 8 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM21 1 9 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM22 12 10 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM23 1 11 12 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
XM24 12 11 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808650 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808645 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__nfet_con_diff_wo_abt_270v2 VSSIO VCC_IO 4 5 6 7 8 9 10 11 12 13 PAD
**
*.SEEDPROM
X0 VSSIO VCC_IO sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X3 VSSIO 4 PAD sky130_fd_pr__nfet_01v8__example_55959141808647
X4 VSSIO 13 PAD sky130_fd_pr__nfet_01v8__example_55959141808647
X5 VSSIO 13 PAD sky130_fd_pr__nfet_01v8__example_55959141808647
X32 VSSIO 4 5 6 7 8 9 10 11 12 13 PAD sky130_fd_pr__nfet_01v8__example_55959141808648
X33 VSSIO 4 5 6 7 8 9 10 11 12 13 PAD sky130_fd_pr__nfet_01v8__example_55959141808651
X34 VSSIO 4 PAD sky130_fd_pr__nfet_01v8__example_55959141808650
X35 VSSIO 4 PAD sky130_fd_pr__nfet_01v8__example_55959141808650
X36 VSSIO 4 PAD sky130_fd_pr__nfet_01v8__example_55959141808645
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd2__example_55959141808202
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808657 2 3 4
**
*.SEEDPROM
XM0 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
.ENDS
***************************************
.SUBCKT ICV_14
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpm1s2__example_55959141808659
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808658 2 3 4 5 6 7 8 9 10
**
*.SEEDPROM
XM0 10 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM1 2 3 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM2 10 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM3 2 3 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM4 10 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM5 2 3 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM6 10 4 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM7 2 4 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM8 10 4 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM9 2 4 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM10 10 4 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM11 2 4 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM12 10 4 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM13 2 4 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM14 10 4 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM15 2 5 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM16 10 5 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM17 2 5 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM18 10 6 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM19 2 6 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM20 10 6 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM21 2 7 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM22 10 7 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM23 2 7 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM24 10 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM25 2 8 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM26 10 9 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__pfet_con_diff_wo_abt_270v2 1 2 3 4 5 6 7 8 9 10
**
X0 1 2 sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X7 2 9 10 sky130_fd_pr__pfet_01v8__example_55959141808657
X8 2 9 10 sky130_fd_pr__pfet_01v8__example_55959141808657
X35 2 3 4 5 6 7 8 9 10 sky130_fd_pr__pfet_01v8__example_55959141808658
X36 2 3 4 5 6 7 8 9 10 sky130_fd_pr__pfet_01v8__example_55959141808658
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpio_pudrvr_strongv2 VNB TIE_HI_ESD VCC_IO PAD PU_H_N[2] PU_H_N[3]
**
X0 PU_H_N[2] 9 sky130_fd_io__tk_em2s_cdns_55959141808652
X1 PU_H_N[3] 10 sky130_fd_io__tk_em2s_cdns_55959141808652
X2 TIE_HI_ESD 11 sky130_fd_io__tk_em2s_cdns_55959141808652
X3 PU_H_N[3] 12 sky130_fd_io__tk_em2s_cdns_55959141808652
X4 TIE_HI_ESD 13 sky130_fd_io__tk_em2s_cdns_55959141808652
X5 TIE_HI_ESD 9 sky130_fd_io__tk_em2o_cdns_55959141808653
X6 PU_H_N[3] 9 sky130_fd_io__tk_em2o_cdns_55959141808653
X7 TIE_HI_ESD 10 sky130_fd_io__tk_em2o_cdns_55959141808653
X8 PU_H_N[2] 10 sky130_fd_io__tk_em2o_cdns_55959141808653
X9 PU_H_N[3] 11 sky130_fd_io__tk_em2o_cdns_55959141808653
X10 PU_H_N[2] 11 sky130_fd_io__tk_em2o_cdns_55959141808653
X11 TIE_HI_ESD 12 sky130_fd_io__tk_em2o_cdns_55959141808653
X12 PU_H_N[2] 12 sky130_fd_io__tk_em2o_cdns_55959141808653
X13 PU_H_N[3] 13 sky130_fd_io__tk_em2o_cdns_55959141808653
X14 PU_H_N[2] 13 sky130_fd_io__tk_em2o_cdns_55959141808653
X15 TIE_HI_ESD VCC_IO sky130_fd_pr__res_generic_po__example_5595914180838
X16 VNB VCC_IO PU_H_N[2] PU_H_N[3] 9 10 11 12 13 PAD sky130_fd_io__pfet_con_diff_wo_abt_270v2
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpio_odrvrv2 VGND VGND_IO VCC_IO TIE_LO_ESD PU_H_N[0] PD_H[2] PD_H[3] 14 PAD PD_H[1] PD_H[0] PU_H_N[1] PU_H_N[3] TIE_HI_ESD PU_H_N[2]
**
*.SEEDPROM
*.CALIBRE ISOLATED NETS: FORCE_HI_H_N VSSIO_AMX FORCE_LOVOL_H FORCE_LO_H
XM0 30 PU_H_N[0] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM1 VCC_IO PU_H_N[0] 30 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM2 30 PU_H_N[0] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM3 VCC_IO PU_H_N[0] 30 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
X4 VGND_IO VCC_IO condiode m=1
X5 VGND_IO VCC_IO condiode m=1
X6 VGND_IO VCC_IO condiode m=1
R7 26 27 sky130_fd_pr__res_generic_po W=2 m=1 w=480000u l=45000u
R8 27 28 sky130_fd_pr__res_generic_po W=2 m=1 w=480000u l=45000u
R9 28 29 sky130_fd_pr__res_generic_po W=2 m=1 w=480000u l=45000u
X10 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2dn m=1
X11 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
R12 27 43 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R13 43 28 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
X14 PD_H[3] 42 sky130_fd_io__tk_em2s_cdns_55959141808652
X15 PD_H[2] 41 sky130_fd_io__tk_em2s_cdns_55959141808652
X16 PD_H[3] 40 sky130_fd_io__tk_em2s_cdns_55959141808652
X17 PD_H[3] 39 sky130_fd_io__tk_em2s_cdns_55959141808652
X18 PD_H[3] 38 sky130_fd_io__tk_em2s_cdns_55959141808652
X19 PD_H[3] 37 sky130_fd_io__tk_em2s_cdns_55959141808652
X20 TIE_LO_ESD 36 sky130_fd_io__tk_em2s_cdns_55959141808652
X21 TIE_LO_ESD 42 sky130_fd_io__tk_em2o_cdns_55959141808653
X22 PD_H[2] 42 sky130_fd_io__tk_em2o_cdns_55959141808653
X23 PD_H[3] 41 sky130_fd_io__tk_em2o_cdns_55959141808653
X24 TIE_LO_ESD 41 sky130_fd_io__tk_em2o_cdns_55959141808653
X25 PD_H[2] 40 sky130_fd_io__tk_em2o_cdns_55959141808653
X26 TIE_LO_ESD 40 sky130_fd_io__tk_em2o_cdns_55959141808653
X27 PD_H[2] 39 sky130_fd_io__tk_em2o_cdns_55959141808653
X28 TIE_LO_ESD 39 sky130_fd_io__tk_em2o_cdns_55959141808653
X29 PD_H[2] 38 sky130_fd_io__tk_em2o_cdns_55959141808653
X30 TIE_LO_ESD 38 sky130_fd_io__tk_em2o_cdns_55959141808653
X31 PD_H[2] 37 sky130_fd_io__tk_em2o_cdns_55959141808653
X32 TIE_LO_ESD 37 sky130_fd_io__tk_em2o_cdns_55959141808653
X33 PD_H[2] 36 sky130_fd_io__tk_em2o_cdns_55959141808653
X34 PD_H[3] 36 sky130_fd_io__tk_em2o_cdns_55959141808653
X35 PAD 29 sky130_fd_io__res250only_small
X44 VGND_IO VCC_IO PD_H[0] 30 sky130_fd_io__gpio_pddrvr_weakv2
X45 VCC_IO PU_H_N[0] 30 sky130_fd_pr__pfet_01v8__example_55959141808654
X46 VCC_IO PU_H_N[1] 26 sky130_fd_io__com_pudrvr_strong_slowv2
X47 30 35 32 33 34 31 29 sky130_fd_io__com_res_weak
X53 TIE_LO_ESD VGND_IO sky130_fd_pr__res_generic_po__example_5595914180838
X54 VGND_IO VCC_IO PD_H[1] 26 sky130_fd_io__gpio_pddrvr_strong_slowv2
X55 VGND_IO VCC_IO 36 37 38 39 40 PD_H[2] PD_H[3] 14 41 42 PAD sky130_fd_io__nfet_con_diff_wo_abt_270v2
X56 VGND TIE_HI_ESD VCC_IO PAD PU_H_N[2] PU_H_N[3] sky130_fd_io__gpio_pudrvr_strongv2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__tpl1__example_55959141808151
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__tpl1__example_55959141808148
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__tpl1__example_55959141808150
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__tpl1__example_55959141808149
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1__example_55959141808158
**
.ENDS
***************************************
.SUBCKT sky130_fd_io__signal_5_sym_hv_local_5term NBODY NWELLRING GATE VGND IN 7
**
*.SEEDPROM
XM0 IN GATE VGND NBODY sky130_fd_pr__esd_nfet_g5v0d10v5 L=0.6 W=5.4 m=1
R1 NWELLRING 7 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R2 NBODY 8 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808555 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_buf_localesd VSSD VDDIO_Q VTRIP_SEL_H OUT_VT OUT_H IN_H
**
X0 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X1 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X2 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X3 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X4 IN_H OUT_H sky130_fd_io__res250only_small
X5 VSSD VDDIO_Q VSSD VSSD OUT_H 8 sky130_fd_io__signal_5_sym_hv_local_5term
X6 VSSD VDDIO_Q VSSD OUT_H VDDIO_Q 7 sky130_fd_io__signal_5_sym_hv_local_5term
X7 VSSD VTRIP_SEL_H OUT_VT OUT_H sky130_fd_pr__nfet_01v8__example_55959141808555
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd__example_55959141808517
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808533 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808230 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 m=1
XM1 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808604
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd2__example_55959141808518
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd__example_55959141808190
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808548 2 3 4 5
**
*.SEEDPROM
XM0 5 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd2__example_55959141808191
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808189 2 3 4 5
**
*.SEEDPROM
XM0 5 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM1 4 3 5 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808611
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808610 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM1 3 2 4 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM2 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM3 3 2 4 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM4 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_in_buf VSSD VDDIO_Q IN_H MODE_NORMAL_N IN_VT VTRIP_SEL_H_N OUT VTRIP_SEL_H
**
*.SEEDPROM
XM0 19 11 17 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM1 17 11 19 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM2 19 11 17 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM3 17 11 19 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM4 VSSD VTRIP_SEL_H_N IN_VT VSSD sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 m=1
XM5 18 11 17 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=1 m=1
XM6 17 11 18 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=1 m=1
XM7 18 11 17 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=1 m=1
XM8 17 11 18 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=1 m=1
XM9 VSSD IN_VT 17 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM10 VSSD IN_H 17 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM11 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM12 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM13 12 11 14 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
XM14 11 IN_H 16 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=5 m=1
XM15 15 IN_H 11 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=5 m=1
XM16 VDDIO_Q VDDIO_Q VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=5 m=1
X17 VSSD VDDIO_Q 20 10 sky130_fd_io__hvsbt_inv_x1
X20 VSSD VDDIO_Q VTRIP_SEL_H MODE_NORMAL_N 20 sky130_fd_io__hvsbt_nor
X25 VSSD 12 OUT_N VSSD sky130_fd_pr__nfet_01v8__example_55959141808533
X26 VSSD OUT_N VSSD OUT sky130_fd_pr__nfet_01v8__example_55959141808533
X27 VSSD MODE_NORMAL_N 12 sky130_fd_pr__nfet_01v8__example_55959141808230
X28 VSSD 11 12 sky130_fd_pr__nfet_01v8__example_55959141808230
X36 VDDIO_Q MODE_NORMAL_N VDDIO_Q 14 sky130_fd_pr__pfet_01v8__example_55959141808548
X37 VDDIO_Q 12 OUT_N VDDIO_Q sky130_fd_pr__pfet_01v8__example_55959141808548
X38 VDDIO_Q OUT_N VDDIO_Q OUT sky130_fd_pr__pfet_01v8__example_55959141808548
X39 VDDIO_Q MODE_NORMAL_N VDDIO_Q 16 sky130_fd_pr__pfet_01v8__example_55959141808189
X40 VDDIO_Q 10 15 VDDIO_Q sky130_fd_pr__pfet_01v8__example_55959141808189
X41 VDDIO_Q 10 VDDIO_Q 19 sky130_fd_pr__pfet_01v8__example_55959141808189
X42 VDDIO_Q MODE_NORMAL_N VDDIO_Q 18 sky130_fd_pr__pfet_01v8__example_55959141808189
X46 VSSD IN_H 11 17 sky130_fd_pr__nfet_01v8__example_55959141808610
X47 VSSD IN_H VSSD 17 sky130_fd_pr__nfet_01v8__example_55959141808610
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808550 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
XM1 3 2 4 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
XM2 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808607 1 2 3
**
XM0 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
XM1 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
XM2 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
XM3 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808528 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808600 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808481 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_ipath_hvls VSSD VDDIO_Q MODE_VCCHIB_N INB_VCCHIB MODE_VCCHIB MODE_NORMAL_N MODE_NORMAL IN_VDDIO IN_VCCHIB OUT
**
*.SEEDPROM
XM0 VDDIO_Q OUT_B OUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM1 OUT OUT_B VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM2 VDDIO_Q OUT_B OUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM3 OUT OUT_B VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM4 VDDIO_Q OUT_B OUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
X5 VSSD MODE_VCCHIB_N 11 VSSD sky130_fd_pr__nfet_01v8__example_55959141808533
X8 VDDIO_Q MODE_VCCHIB 15 OUT_B sky130_fd_pr__pfet_01v8__example_55959141808548
X9 VDDIO_Q MODE_NORMAL VDDIO_Q 15 sky130_fd_pr__pfet_01v8__example_55959141808548
X14 VDDIO_Q 13 16 OUT_B sky130_fd_pr__pfet_01v8__example_55959141808189
X15 VDDIO_Q MODE_VCCHIB_N 16 VDDIO_Q sky130_fd_pr__pfet_01v8__example_55959141808189
X16 VDDIO_Q MODE_NORMAL_N 17 VDDIO_Q sky130_fd_pr__pfet_01v8__example_55959141808189
X17 VDDIO_Q IN_VDDIO 17 OUT_B sky130_fd_pr__pfet_01v8__example_55959141808189
X18 VSSD INB_VCCHIB 18 11 sky130_fd_pr__nfet_01v8__example_55959141808550
X19 VSSD IN_VCCHIB 19 12 sky130_fd_pr__nfet_01v8__example_55959141808550
X20 VSSD OUT_B OUT VSSD sky130_fd_pr__nfet_01v8__example_55959141808550
X21 VSSD MODE_VCCHIB 18 sky130_fd_pr__nfet_01v8__example_55959141808607
X22 VSSD MODE_VCCHIB 19 sky130_fd_pr__nfet_01v8__example_55959141808607
X23 VSSD 13 OUT_B 20 sky130_fd_pr__nfet_01v8__example_55959141808528
X24 VSSD MODE_VCCHIB 20 VSSD sky130_fd_pr__nfet_01v8__example_55959141808528
X25 VSSD MODE_NORMAL 21 VSSD sky130_fd_pr__nfet_01v8__example_55959141808528
X26 VSSD IN_VDDIO OUT_B 21 sky130_fd_pr__nfet_01v8__example_55959141808528
X27 VSSD 12 VSSD 13 sky130_fd_pr__nfet_01v8__example_55959141808600
X28 VDDIO_Q 11 VDDIO_Q 12 sky130_fd_pr__pfet_01v8__example_55959141808481
X29 VDDIO_Q 12 11 VDDIO_Q sky130_fd_pr__pfet_01v8__example_55959141808481
X30 VDDIO_Q 12 VDDIO_Q 13 sky130_fd_pr__pfet_01v8__example_55959141808481
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808535 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM1 3 2 4 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808602 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_01v8 L=0.25 W=1 m=1
XM1 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.25 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_5595914180825 1 2 3
**
XM0 1 2 3 1 sky130_fd_pr__nfet_01v8 L=0.25 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808598 2 3 4 5
**
*.SEEDPROM
XM0 5 3 4 2 sky130_fd_pr__pfet_01v8 L=0.25 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808596 2 3 4 5
**
*.SEEDPROM
XM0 5 3 4 2 sky130_fd_pr__pfet_01v8 L=0.25 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_vcchib_in_buf VSSD VCCHIB MODE_VCCHIB_LV_N OUT_N IN_H OUT
**
*.SEEDPROM
XM0 VSSD OUT_N OUT VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=1 m=1
XM1 OUT OUT_N VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=1 m=1
XM2 VSSD OUT_N OUT VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=1 m=1
XM3 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=1 m=1
XM4 12 8 11 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=1 m=1
XM5 11 8 12 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=1 m=1
XM6 12 8 11 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=1 m=1
XM7 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM8 VCCHIB MODE_VCCHIB_LV_N 9 VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=5 m=1
XM9 9 MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=5 m=1
XM10 VCCHIB MODE_VCCHIB_LV_N 9 VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=5 m=1
XM11 7 8 10 VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=1 m=1
XM12 10 8 7 VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=1 m=1
XM13 8 IN_H 9 VCCHIB sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=5 m=1
XM14 9 IN_H 8 VCCHIB sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=5 m=1
X23 VSSD IN_H 12 8 sky130_fd_pr__nfet_01v8__example_55959141808535
X24 VSSD IN_H 12 VSSD sky130_fd_pr__nfet_01v8__example_55959141808535
X25 VSSD 8 7 sky130_fd_pr__nfet_01v8__example_55959141808602
X26 VSSD MODE_VCCHIB_LV_N 7 sky130_fd_pr__nfet_01v8__example_55959141808602
X27 VSSD 7 OUT_N sky130_fd_pr__nfet_01v8__example_5595914180825
X28 VCCHIB MODE_VCCHIB_LV_N 10 VCCHIB sky130_fd_pr__pfet_01v8__example_55959141808598
X29 VCCHIB MODE_VCCHIB_LV_N VCCHIB 11 sky130_fd_pr__pfet_01v8__example_55959141808596
X30 VCCHIB 7 VCCHIB OUT_N sky130_fd_pr__pfet_01v8__example_55959141808596
X31 VCCHIB OUT_N OUT VCCHIB sky130_fd_pr__pfet_01v8__example_55959141808596
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_inbuf_lvinv_x1 VGND VPWR IN OUT
**
*.SEEDPROM
XM0 VPWR IN OUT VPWR sky130_fd_pr__pfet_01v8_hvt L=0.25 W=3 m=1
X3 VGND IN OUT sky130_fd_pr__nfet_01v8__example_5595914180825
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808547 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_01v8 L=0.25 W=3 m=1
XM1 3 2 4 1 sky130_fd_pr__nfet_01v8 L=0.25 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd2__example_5595914180812
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808599 2 3 4 5
**
*.SEEDPROM
XM0 5 3 4 2 sky130_fd_pr__pfet_01v8 L=0.25 W=3 m=1
XM1 4 3 5 2 sky130_fd_pr__pfet_01v8 L=0.25 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808546 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_01v8 L=0.25 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_ipath_lvls VSSD VCCHIB MODE_NORMAL_LV IN_VDDIO 5 MODE_NORMAL_LV_N OUT_B MODE_VCCHIB_LV_N IN_VCCHIB MODE_VCCHIB_LV OUT
**
*.SEEDPROM
XM0 OUT OUT_B VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=3 m=1
XM1 VCCHIB OUT_B OUT VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=3 m=1
XM2 OUT OUT_B VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=3 m=1
XM3 VCCHIB OUT_B OUT VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=3 m=1
X6 VCCHIB IN_VDDIO VCCHIB 12 sky130_fd_pr__pfet_01v8__example_55959141808189
X7 VSSD IN_VDDIO 12 18 sky130_fd_pr__nfet_01v8__example_55959141808600
X8 VCCHIB MODE_NORMAL_LV OUT_B 13 sky130_fd_pr__pfet_01v8__example_55959141808598
X9 VCCHIB MODE_VCCHIB_LV 13 VCCHIB sky130_fd_pr__pfet_01v8__example_55959141808598
X10 VCCHIB MODE_NORMAL_LV VCCHIB 12 sky130_fd_pr__pfet_01v8__example_55959141808596
X11 VCCHIB 12 VCCHIB 5 sky130_fd_pr__pfet_01v8__example_55959141808596
X12 VSSD 5 16 OUT_B sky130_fd_pr__nfet_01v8__example_55959141808547
X13 VSSD MODE_NORMAL_LV 16 VSSD sky130_fd_pr__nfet_01v8__example_55959141808547
X14 VSSD OUT_B VSSD OUT sky130_fd_pr__nfet_01v8__example_55959141808547
X15 VSSD IN_VCCHIB 17 OUT_B sky130_fd_pr__nfet_01v8__example_55959141808547
X16 VSSD MODE_VCCHIB_LV 17 VSSD sky130_fd_pr__nfet_01v8__example_55959141808547
X20 VCCHIB 5 14 OUT_B sky130_fd_pr__pfet_01v8__example_55959141808599
X21 VCCHIB MODE_NORMAL_LV_N 14 VCCHIB sky130_fd_pr__pfet_01v8__example_55959141808599
X22 VCCHIB MODE_VCCHIB_LV_N 15 VCCHIB sky130_fd_pr__pfet_01v8__example_55959141808599
X23 VCCHIB IN_VCCHIB 15 OUT_B sky130_fd_pr__pfet_01v8__example_55959141808599
X24 VSSD MODE_NORMAL_LV 18 VSSD sky130_fd_pr__nfet_01v8__example_55959141808546
X25 VSSD 12 VSSD 5 sky130_fd_pr__nfet_01v8__example_55959141808546
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_ibuf_se VSSD VDDIO_Q VCCHIB MODE_NORMAL_N MODE_VCCHIB_N ENABLE_VDDIO_LV IN_H VTRIP_SEL_H VTRIP_SEL_H_N IN_VT IBUFMUX_OUT_H IBUFMUX_OUT 14
**
*.SEEDPROM
X0 VSSD VCCHIB sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X1 VSSD VCCHIB sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X2 VSSD VDDIO_Q MODE_NORMAL_N 15 sky130_fd_io__hvsbt_inv_x1
X3 VSSD VDDIO_Q MODE_VCCHIB_N 16 sky130_fd_io__hvsbt_inv_x1
X4 VSSD VCCHIB ENABLE_VDDIO_LV 16 17 sky130_fd_io__hvsbt_nand2
X5 VSSD VCCHIB ENABLE_VDDIO_LV 15 18 sky130_fd_io__hvsbt_nand2
X6 VSSD VDDIO_Q IN_H MODE_NORMAL_N IN_VT VTRIP_SEL_H_N 19 VTRIP_SEL_H sky130_fd_io__gpiov2_in_buf
X7 VSSD VDDIO_Q MODE_VCCHIB_N 21 16 MODE_NORMAL_N 15 19 20 IBUFMUX_OUT_H sky130_fd_io__gpiov2_ipath_hvls
X8 VSSD VCCHIB 17 21 IN_H 20 sky130_fd_io__gpiov2_vcchib_in_buf
X9 VSSD VCCHIB 17 22 sky130_fd_io__gpiov2_inbuf_lvinv_x1
X10 VSSD VCCHIB 18 23 sky130_fd_io__gpiov2_inbuf_lvinv_x1
X11 VSSD VCCHIB 23 19 14 18 24 17 20 22 IBUFMUX_OUT sky130_fd_io__gpiov2_ipath_lvls
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_ictl_logic VSSD VDDIO_Q DM_H_N[1] DM_H_N[0] DM_H_N[2] INP_DIS_H_N IB_MODE_SEL_H MODE_VCCHIB_N IB_MODE_SEL_H_N MODE_NORMAL_N TRIPSEL_I_H VTRIP_SEL_H_N TRIPSEL_I_H_N
**
*.SEEDPROM
X0 VSSD VDDIO_Q 14 16 sky130_fd_io__hvsbt_inv_x1
X1 VSSD VDDIO_Q INP_DIS_I_H INP_DIS_I_H_N sky130_fd_io__hvsbt_inv_x1
X2 VSSD VDDIO_Q TRIPSEL_I_H TRIPSEL_I_H_N sky130_fd_io__hvsbt_inv_x1
X3 VSSD VDDIO_Q VTRIP_SEL_H_N MODE_NORMAL_N TRIPSEL_I_H sky130_fd_io__hvsbt_nor
X4 VDDIO_Q DM_H_N[1] VDDIO_Q 14 sky130_fd_pr__pfet_01v8__example_559591418085
X5 VDDIO_Q DM_H_N[1] VDDIO_Q 14 sky130_fd_pr__pfet_01v8__example_559591418085
X6 VDDIO_Q DM_H_N[0] 14 VDDIO_Q sky130_fd_pr__pfet_01v8__example_559591418085
X7 VDDIO_Q DM_H_N[0] 14 VDDIO_Q sky130_fd_pr__pfet_01v8__example_559591418085
X8 VSSD DM_H_N[1] 15 sky130_fd_pr__nfet_01v8__example_559591418089
X9 VSSD DM_H_N[0] 15 14 sky130_fd_pr__nfet_01v8__example_559591418087
X10 VSSD VDDIO_Q DM_H_N[2] 16 17 sky130_fd_io__hvsbt_nand2
X11 VSSD VDDIO_Q 17 INP_DIS_H_N INP_DIS_I_H sky130_fd_io__hvsbt_nand2
X12 VSSD VDDIO_Q INP_DIS_I_H_N IB_MODE_SEL_H MODE_VCCHIB_N sky130_fd_io__hvsbt_nand2
X13 VSSD VDDIO_Q INP_DIS_I_H_N IB_MODE_SEL_H_N MODE_NORMAL_N sky130_fd_io__hvsbt_nand2
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_ipath VSSD VDDIO_Q ENABLE_VDDIO_LV DM_H_N[0] OUT_H MODE_VCCHIB_N PAD OUT VCCHIB DM_H_N[1] DM_H_N[2] INP_DIS_H_N IB_MODE_SEL_H IB_MODE_SEL_H_N VTRIP_SEL_H_N
**
*.SEEDPROM
X0 VSSD VDDIO_Q 22 21 19 PAD sky130_fd_io__gpiov2_buf_localesd
X1 VSSD VDDIO_Q VCCHIB 20 MODE_VCCHIB_N ENABLE_VDDIO_LV 19 22 23 21 OUT_H OUT 24 sky130_fd_io__gpiov2_ibuf_se
X2 VSSD VDDIO_Q DM_H_N[1] DM_H_N[0] DM_H_N[2] INP_DIS_H_N IB_MODE_SEL_H MODE_VCCHIB_N IB_MODE_SEL_H_N 20 22 VTRIP_SEL_H_N 23 sky130_fd_io__gpiov2_ictl_logic
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808314 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd2__example_55959141808143
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808362 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
XM1 3 2 4 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808364 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
XM1 3 2 4 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808360 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd__example_55959141808194
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808284 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808282 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em1o_cdns_55959141808289 2 3
**
R0 2 4 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R1 5 3 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em1s_cdns_55959141808288 1 2
**
R0 1 3 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R1 3 2 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_pr__via_pol1__example_55959141808272
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808283 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM1 1 2 3 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM2 3 2 1 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808287 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1.5 m=1
.ENDS
***************************************
.SUBCKT ICV_15 1 2 3 4 5
**
X0 1 2 4 sky130_fd_pr__nfet_01v8__example_55959141808287
X1 1 3 5 sky130_fd_pr__nfet_01v8__example_55959141808287
.ENDS
***************************************
.SUBCKT sky130_fd_pr__via_pol1__example_55959141808273
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__via_pol1__example_55959141808275
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_generic_po__example_55959141808285 1 2
**
R0 1 2 sky130_fd_pr__res_generic_po W=0.33 m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808281 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=0.42 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808644 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=0.42 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_generic_po__example_55959141808286 2 3
**
R0 2 3 sky130_fd_pr__res_generic_po W=0.33 m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_pr__via_pol1__example_55959141808294
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808304 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__via_pol1__example_55959141808295
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808307 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 m=1
XM1 3 2 4 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 m=1
XM2 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 m=1
XM3 3 2 4 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808315 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=1 m=1
XM1 1 2 3 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=1 m=1
XM2 3 2 1 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=1 m=1
XM3 1 2 3 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808313 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__feascom_pupredrvr_nbiasv2 VGND_IO VCC_IO EN_H NBIAS DRVHI_H PUEN_H 7 PU_H_N EN_H_N 10 11 12
**
XM0 VGND_IO DRVHI_H 16 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 m=1
XM1 20 14 19 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 m=1
XM2 13 DRVHI_H 20 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 m=1
XM3 15 VCC_IO VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=8 W=0.42 m=1
XM4 10 10 11 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 m=1
XM5 11 10 10 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 m=1
XM6 15 11 11 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 m=1
XM7 11 11 15 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 m=1
XM8 16 DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 m=1
XM9 VCC_IO DRVHI_H 16 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 m=1
XM10 18 PU_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=8 W=0.42 m=1
XM11 13 17 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
XM12 VCC_IO 17 13 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
XM13 13 17 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
XM14 VCC_IO 17 13 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
XM15 10 13 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM16 VCC_IO 13 10 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
R17 23 PU_H_N sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R18 23 14 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R19 25 14 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R20 26 17 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
X28 EN_H 27 14 sky130_fd_io__tk_em1o_cdns_5595914180880
X29 7 24 NBIAS sky130_fd_io__tk_em1o_cdns_5595914180880
X30 21 NBIAS sky130_fd_io__tk_em1s_cdns_5595914180882
X31 13 18 sky130_fd_io__tk_em1s_cdns_5595914180882
X32 NBIAS 22 sky130_fd_io__tk_em1s_cdns_5595914180881
X33 7 12 sky130_fd_io__tk_em1s_cdns_5595914180881
X36 VCC_IO 14 17 14 sky130_fd_pr__pfet_01v8__example_55959141808314
X42 VGND_IO EN_H VGND_IO 19 sky130_fd_pr__nfet_01v8__example_55959141808282
X43 VGND_IO 13 VGND_IO 21 sky130_fd_pr__nfet_01v8__example_55959141808281
X49 VGND_IO EN_H_N NBIAS VGND_IO sky130_fd_pr__nfet_01v8__example_55959141808304
X50 VGND_IO 16 NBIAS VGND_IO sky130_fd_pr__nfet_01v8__example_55959141808304
X51 VGND_IO 16 VGND_IO 15 sky130_fd_pr__nfet_01v8__example_55959141808304
X53 VGND_IO NBIAS 7 NBIAS sky130_fd_pr__nfet_01v8__example_55959141808307
X54 VGND_IO 7 VGND_IO 7 sky130_fd_pr__nfet_01v8__example_55959141808307
X55 VGND_IO 15 VGND_IO 12 sky130_fd_pr__nfet_01v8__example_55959141808307
X56 VCC_IO 13 NBIAS sky130_fd_pr__pfet_01v8__example_55959141808315
X57 VCC_IO 13 22 sky130_fd_pr__pfet_01v8__example_55959141808315
X58 VCC_IO DRVHI_H 13 sky130_fd_pr__pfet_01v8__example_55959141808313
X59 VCC_IO EN_H 13 sky130_fd_pr__pfet_01v8__example_55959141808313
X60 VCC_IO PUEN_H 17 sky130_fd_pr__pfet_01v8__example_55959141808313
X61 VCC_IO DRVHI_H 17 sky130_fd_pr__pfet_01v8__example_55959141808313
.ENDS
***************************************
.SUBCKT sky130_fd_pr__model__nfet_highvoltage__example_55959141808144 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpio_pupredrvr_strongv2 VGND_IO VCC_IO SLOW_H_N PUEN_H DRVHI_H PU_H_N[2] 7 PU_H_N[3] 9 10 11 12 13
**
XM0 23 14 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 m=1
XM1 14 SLOW_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 m=1
XM2 VCC_IO PUEN_H 14 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 m=1
XM3 23 14 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 m=1
X4 23 35 15 sky130_fd_io__tk_em1o_cdns_5595914180880
X5 23 36 21 sky130_fd_io__tk_em1o_cdns_5595914180880
X6 15 11 sky130_fd_io__tk_em1s_cdns_5595914180882
X7 17 PU_H_N[2] sky130_fd_io__tk_em1s_cdns_5595914180882
X8 21 11 sky130_fd_io__tk_em1s_cdns_5595914180882
X9 7 PU_H_N[3] sky130_fd_io__tk_em1s_cdns_5595914180882
X15 VCC_IO PUEN_H PU_H_N[2] sky130_fd_pr__pfet_01v8__example_55959141808284
X16 VCC_IO PUEN_H PU_H_N[3] sky130_fd_pr__pfet_01v8__example_55959141808284
X17 VGND_IO DRVHI_H 17 28 sky130_fd_pr__nfet_01v8__example_55959141808282
X18 VGND_IO DRVHI_H 17 29 sky130_fd_pr__nfet_01v8__example_55959141808282
X19 VGND_IO DRVHI_H 17 24 sky130_fd_pr__nfet_01v8__example_55959141808282
X20 VGND_IO DRVHI_H 17 25 sky130_fd_pr__nfet_01v8__example_55959141808282
X21 VGND_IO DRVHI_H 7 26 sky130_fd_pr__nfet_01v8__example_55959141808282
X22 VGND_IO DRVHI_H 7 27 sky130_fd_pr__nfet_01v8__example_55959141808282
X23 VGND_IO DRVHI_H 7 30 sky130_fd_pr__nfet_01v8__example_55959141808282
X24 VGND_IO DRVHI_H 7 31 sky130_fd_pr__nfet_01v8__example_55959141808282
X25 19 VGND_IO sky130_fd_io__tk_em1o_cdns_55959141808289
X26 20 21 sky130_fd_io__tk_em1o_cdns_55959141808289
X27 22 21 sky130_fd_io__tk_em1o_cdns_55959141808289
X28 19 21 sky130_fd_io__tk_em1s_cdns_55959141808288
X29 VGND_IO 20 sky130_fd_io__tk_em1s_cdns_55959141808288
X30 VGND_IO 22 sky130_fd_io__tk_em1s_cdns_55959141808288
X34 VCC_IO DRVHI_H PU_H_N[2] sky130_fd_pr__pfet_01v8__example_55959141808283
X35 VCC_IO DRVHI_H PU_H_N[3] sky130_fd_pr__pfet_01v8__example_55959141808283
X36 VGND_IO 15 15 24 28 ICV_15
X37 VGND_IO 15 15 25 29 ICV_15
X38 VGND_IO 21 19 30 26 ICV_15
X39 VGND_IO 22 20 31 27 ICV_15
X44 16 PU_H_N[2] sky130_fd_pr__res_generic_po__example_55959141808285
X45 18 PU_H_N[3] sky130_fd_pr__res_generic_po__example_55959141808285
X46 VGND_IO DRVHI_H 32 PU_H_N[2] sky130_fd_pr__nfet_01v8__example_55959141808281
X47 VGND_IO DRVHI_H 33 PU_H_N[3] sky130_fd_pr__nfet_01v8__example_55959141808281
X48 VGND_IO PUEN_H 32 sky130_fd_pr__nfet_01v8__example_55959141808644
X49 VGND_IO PUEN_H 33 sky130_fd_pr__nfet_01v8__example_55959141808644
X50 16 17 sky130_fd_pr__res_generic_po__example_55959141808286
X51 18 7 sky130_fd_pr__res_generic_po__example_55959141808286
X52 VGND_IO VCC_IO 23 11 DRVHI_H PUEN_H 9 PU_H_N[2] 14 13 12 10 sky130_fd_io__feascom_pupredrvr_nbiasv2
X53 VGND_IO SLOW_H_N 14 34 sky130_fd_pr__model__nfet_highvoltage__example_55959141808144
X54 VGND_IO PUEN_H VGND_IO 34 sky130_fd_pr__model__nfet_highvoltage__example_55959141808144
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808636 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__pfet_g5v0d10v5 L=2 W=0.42 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808630 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__pfet_g5v0d10v5 L=4 W=0.42 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808634 2 3 4 5
**
*.SEEDPROM
XM0 5 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__model__pfet_highvoltage__example_55959141808141 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808629 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__pfet_g5v0d10v5 L=1 W=0.42 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808631 1 2 3
**
XM0 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
XM1 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808354 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__pfet_g5v0d10v5 L=4 W=0.42 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808628 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808626 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
XM1 3 2 4 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_pdpredrvr_strong_nr2 VGND_IO VCC_IO I2C_MODE_H DRVLO_H_N EN_FAST_N[0] EN_FAST_N[1] PDEN_H_N PD_H PD_I2C_H
**
XM0 10 I2C_MODE_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
XM1 VCC_IO I2C_MODE_H 10 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
XM2 10 I2C_MODE_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
X3 VGND_IO I2C_MODE_H VGND_IO PD_H sky130_fd_pr__nfet_01v8__example_55959141808116
X4 VGND_IO PDEN_H_N VGND_IO PD_H sky130_fd_pr__nfet_01v8__example_55959141808116
X5 VGND_IO PDEN_H_N VGND_IO PD_I2C_H sky130_fd_pr__nfet_01v8__example_55959141808116
X10 VCC_IO PDEN_H_N VCC_IO 15 sky130_fd_pr__pfet_01v8__example_55959141808630
X11 VCC_IO DRVLO_H_N 15 PD_I2C_H sky130_fd_pr__pfet_01v8__example_55959141808630
X12 VCC_IO EN_FAST_N[1] VCC_IO 11 sky130_fd_pr__pfet_01v8__example_55959141808629
X13 VCC_IO DRVLO_H_N 11 PD_I2C_H sky130_fd_pr__pfet_01v8__example_55959141808629
X14 VCC_IO DRVLO_H_N 11 PD_I2C_H sky130_fd_pr__pfet_01v8__example_55959141808629
X15 VGND_IO DRVLO_H_N PD_H sky130_fd_pr__nfet_01v8__example_55959141808631
X16 VGND_IO DRVLO_H_N PD_I2C_H sky130_fd_pr__nfet_01v8__example_55959141808631
X17 VCC_IO PDEN_H_N 14 16 sky130_fd_pr__pfet_01v8__example_55959141808354
X18 VCC_IO PDEN_H_N 10 16 sky130_fd_pr__pfet_01v8__example_55959141808354
X19 VCC_IO DRVLO_H_N 14 PD_H sky130_fd_pr__pfet_01v8__example_55959141808354
X20 VCC_IO EN_FAST_N[0] 10 12 sky130_fd_pr__pfet_01v8__example_55959141808628
X21 VCC_IO EN_FAST_N[1] 10 13 sky130_fd_pr__pfet_01v8__example_55959141808628
X22 VCC_IO DRVLO_H_N PD_H 12 sky130_fd_pr__pfet_01v8__example_55959141808626
X23 VCC_IO DRVLO_H_N PD_H 13 sky130_fd_pr__pfet_01v8__example_55959141808626
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_5595914180888 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808344 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808346 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM1 3 2 4 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM2 4 2 3 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM3 3 2 4 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__via_pol1__example_55959141808321
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808343 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM1 3 2 4 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM2 4 2 3 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM3 3 2 4 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM4 4 2 3 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM5 3 2 4 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM6 4 2 3 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM7 3 2 4 1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808329 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808330 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__via_pol1__example_55959141808322
**
.ENDS
***************************************
.SUBCKT sky130_fd_io__com_pdpredrvr_pbiasv2 VGND_IO VCC_IO PD_H DRVLO_H_N PDEN_H_N EN_H_N EN_H 9 PBIAS 11 12 13 14 15
**
XM0 23 17 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 m=1
XM1 VGND_IO 17 23 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 m=1
XM2 PBIAS 17 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 m=1
XM3 VGND_IO 17 PBIAS VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 m=1
XM4 VGND_IO PD_H 14 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=4 W=0.42 m=1
XM5 24 PD_H 14 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=4 W=0.42 m=1
XM6 VGND_IO PDEN_H_N 18 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 m=1
XM7 20 17 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=0.42 m=1
XM8 21 DRVLO_H_N 17 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
XM9 19 DRVLO_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 m=1
XM10 22 16 21 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
XM11 VCC_IO EN_H_N 22 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
XM12 VCC_IO DRVLO_H_N 19 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 m=1
XM13 11 VGND_IO VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=8 W=0.42 m=1
R14 25 16 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R15 26 18 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R16 16 27 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R17 28 EN_H_N sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
X18 16 PD_H sky130_fd_io__tk_em1s_cdns_5595914180882
X19 23 PBIAS sky130_fd_io__tk_em1s_cdns_5595914180882
X20 PBIAS 9 sky130_fd_io__tk_em1o_cdns_5595914180879
X21 9 15 sky130_fd_io__tk_em1s_cdns_5595914180881
X24 24 17 sky130_fd_io__tk_em1s_cdns_55959141808288
X25 PBIAS 20 sky130_fd_io__tk_em1s_cdns_55959141808288
X29 VGND_IO 16 18 16 sky130_fd_pr__nfet_01v8__example_55959141808304
X30 VCC_IO EN_H PBIAS sky130_fd_pr__pfet_01v8__example_55959141808344
X31 VCC_IO 19 11 sky130_fd_pr__pfet_01v8__example_55959141808344
X32 VCC_IO 19 PBIAS sky130_fd_pr__pfet_01v8__example_55959141808344
X33 VCC_IO 12 13 12 sky130_fd_pr__pfet_01v8__example_55959141808346
X34 VCC_IO 13 13 11 sky130_fd_pr__pfet_01v8__example_55959141808346
X38 VCC_IO 9 VCC_IO 9 sky130_fd_pr__pfet_01v8__example_55959141808343
X39 VCC_IO PBIAS 9 PBIAS sky130_fd_pr__pfet_01v8__example_55959141808343
X40 VCC_IO 11 VCC_IO 15 sky130_fd_pr__pfet_01v8__example_55959141808343
X41 VGND_IO DRVLO_H_N 18 sky130_fd_pr__nfet_01v8__example_55959141808329
X42 VGND_IO DRVLO_H_N 17 sky130_fd_pr__nfet_01v8__example_55959141808329
X43 VGND_IO EN_H_N 17 sky130_fd_pr__nfet_01v8__example_55959141808329
X44 VGND_IO DRVLO_H_N 19 sky130_fd_pr__nfet_01v8__example_55959141808329
X45 VGND_IO 17 12 sky130_fd_pr__nfet_01v8__example_55959141808330
X46 VGND_IO 18 17 sky130_fd_pr__nfet_01v8__example_55959141808330
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_pdpredrvr_strong VGND_IO VGND VCC_IO PD_H[4] I2C_MODE_H_N PDEN_H_N 7 PD_H[3] DRVLO_H_N SLOW_H 11 12 13 14 15 16 17 PD_H[2]
**
*.SEEDPROM
XM0 VGND PD_H[4] 26 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 m=1
XM1 22 PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 m=1
XM2 VGND_IO 21 22 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 m=1
XM3 27 22 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 m=1
XM4 VGND_IO 7 PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
XM5 PD_H[3] 7 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
XM6 VGND_IO 7 PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
XM7 PD_H[3] 7 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
XM8 VGND_IO 7 PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
XM9 PD_H[3] PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
XM10 VGND_IO PDEN_H_N PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
XM11 VCC_IO PD_H[4] 26 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
XM12 27 22 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 m=1
XM13 VCC_IO 23 28 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 m=1
XM14 28 23 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 m=1
XM15 PD_H[3] 7 29 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 m=1
XM16 29 7 PD_H[3] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 m=1
X17 VCC_IO I2C_MODE_H_N 20 sky130_fd_pr__model__pfet_highvoltage__example_55959141808371
X18 VCC_IO I2C_MODE_H_N 20 sky130_fd_pr__model__pfet_highvoltage__example_55959141808371
X19 VGND I2C_MODE_H_N 20 sky130_fd_pr__model__nfet_highvoltage__example_55959141808369
X20 VGND VCC_IO 35 21 sky130_fd_io__hvsbt_inv_x1
X21 VGND VCC_IO 36 23 sky130_fd_io__hvsbt_inv_x1
X31 VGND VCC_IO I2C_MODE_H_N SLOW_H 35 sky130_fd_io__hvsbt_nand2
X32 VGND VCC_IO 20 SLOW_H 36 sky130_fd_io__hvsbt_nand2
X33 27 38 37 sky130_fd_io__tk_em1o_cdns_5595914180880
X34 27 39 24 sky130_fd_io__tk_em1o_cdns_5595914180880
X35 25 40 24 sky130_fd_io__tk_em1o_cdns_5595914180880
X36 37 11 sky130_fd_io__tk_em1s_cdns_5595914180882
X37 24 11 sky130_fd_io__tk_em1s_cdns_5595914180882
X38 25 VCC_IO sky130_fd_io__tk_em1s_cdns_5595914180882
X43 VCC_IO 7 30 PD_H[3] sky130_fd_pr__pfet_01v8__example_55959141808481
X44 VCC_IO 7 31 PD_H[3] sky130_fd_pr__pfet_01v8__example_55959141808481
X45 VCC_IO 24 VCC_IO 31 sky130_fd_pr__pfet_01v8__example_55959141808481
X46 VCC_IO 25 VCC_IO 30 sky130_fd_pr__pfet_01v8__example_55959141808481
X47 VCC_IO 7 32 PD_H[3] sky130_fd_pr__pfet_01v8__example_55959141808636
X48 VCC_IO 7 33 PD_H[3] sky130_fd_pr__pfet_01v8__example_55959141808636
X49 VCC_IO PDEN_H_N 28 33 sky130_fd_pr__pfet_01v8__example_55959141808636
X50 VCC_IO PDEN_H_N VCC_IO 32 sky130_fd_pr__pfet_01v8__example_55959141808630
X51 VCC_IO 24 28 29 sky130_fd_pr__pfet_01v8__example_55959141808634
X52 VCC_IO 25 28 29 sky130_fd_pr__pfet_01v8__example_55959141808634
X53 VCC_IO PDEN_H_N 22 34 sky130_fd_pr__model__pfet_highvoltage__example_55959141808141
X54 VCC_IO 21 VCC_IO 34 sky130_fd_pr__model__pfet_highvoltage__example_55959141808141
X55 VCC_IO 20 DRVLO_H_N 7 sky130_fd_pr__pfet_01v8__example_55959141808628
X56 VCC_IO I2C_MODE_H_N 26 7 sky130_fd_pr__pfet_01v8__example_55959141808628
X57 VGND_IO VCC_IO 23 DRVLO_H_N 11 11 PDEN_H_N PD_H[2] PD_H[4] sky130_fd_io__gpiov2_pdpredrvr_strong_nr2
X58 VGND_IO 20 7 26 sky130_fd_pr__nfet_01v8__example_5595914180888
X59 VGND_IO I2C_MODE_H_N 7 DRVLO_H_N sky130_fd_pr__nfet_01v8__example_5595914180888
X60 VGND_IO VCC_IO PD_H[4] DRVLO_H_N PDEN_H_N 27 22 13 11 17 16 15 12 14 sky130_fd_io__com_pdpredrvr_pbiasv2
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_obpredrvr VGND VGND_IO VCC_IO DRVHI_H PUEN_H[0] DRVLO_H_N PDEN_H_N[0] PDEN_H_N[1] PUEN_H[1] PD_H[0] PU_H_N[1] PU_H_N[0] 13 PD_H[1] 15 16 17 18 19 PU_H_N[2]
+ 21 22 23 24 25 26 27 28 PD_H[3] SLOW_H_N PU_H_N[3] I2C_MODE_H_N SLOW_H PD_H[2] PD_H[4] 36
**
*.SEEDPROM
XM0 PU_H_N[0] DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM1 VCC_IO DRVHI_H PU_H_N[0] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM2 37 DRVLO_H_N PD_H[0] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 m=1
XM3 VCC_IO PDEN_H_N[0] 37 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 m=1
XM4 37 PDEN_H_N[0] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 m=1
XM5 VCC_IO DRVHI_H PU_H_N[1] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
XM6 PU_H_N[1] DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
XM7 VCC_IO DRVHI_H PU_H_N[1] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
X8 VGND_IO VCC_IO condiode m=1
X9 VGND_IO VCC_IO sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X10 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2dn m=1
X19 VCC_IO PUEN_H[1] VCC_IO PU_H_N[1] sky130_fd_pr__pfet_01v8__example_55959141808314
X23 VGND_IO DRVHI_H 13 PU_H_N[1] sky130_fd_pr__nfet_01v8__example_55959141808362
X24 VGND_IO PUEN_H[1] 13 VGND_IO sky130_fd_pr__nfet_01v8__example_55959141808362
X25 VCC_IO PDEN_H_N[1] 38 VCC_IO sky130_fd_pr__pfet_01v8__example_55959141808364
X26 VCC_IO DRVLO_H_N 38 PD_H[1] sky130_fd_pr__pfet_01v8__example_55959141808364
X27 VGND_IO DRVHI_H 39 PU_H_N[0] sky130_fd_pr__nfet_01v8__example_55959141808360
X28 VGND_IO PUEN_H[0] VGND_IO 39 sky130_fd_pr__nfet_01v8__example_55959141808360
X29 VGND_IO DRVLO_H_N VGND_IO PD_H[0] sky130_fd_pr__nfet_01v8__example_55959141808360
X30 VGND_IO PDEN_H_N[0] VGND_IO PD_H[0] sky130_fd_pr__nfet_01v8__example_55959141808360
X31 VGND_IO PDEN_H_N[1] VGND_IO PD_H[1] sky130_fd_pr__nfet_01v8__example_55959141808360
X32 VGND_IO DRVLO_H_N VGND_IO PD_H[1] sky130_fd_pr__nfet_01v8__example_55959141808360
X35 VCC_IO PUEN_H[0] PU_H_N[0] sky130_fd_pr__pfet_01v8__example_55959141808284
X36 VGND_IO VCC_IO SLOW_H_N PUEN_H[1] DRVHI_H PU_H_N[2] 21 PU_H_N[3] 15 16 17 18 19 sky130_fd_io__gpio_pupredrvr_strongv2
X37 VGND_IO VGND VCC_IO PD_H[4] I2C_MODE_H_N PDEN_H_N[1] 36 PD_H[3] DRVLO_H_N SLOW_H 22 28 27 26 24 25 23 PD_H[2] sky130_fd_io__gpiov2_pdpredrvr_strong
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808417 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808416 2 3 4 5
**
*.SEEDPROM
XM0 5 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
.ENDS
***************************************
.SUBCKT ICV_16 2 3 4 5
**
*.SEEDPROM
X0 2 3 2 4 sky130_fd_pr__pfet_01v8__example_55959141808416
X1 2 3 2 5 sky130_fd_pr__pfet_01v8__example_55959141808416
.ENDS
***************************************
.SUBCKT sky130_fd_io__com_ctl_ls_octl SET_H VCC_IO VPB 4 HLD_H_N IN RST_H OUT_H_N OUT_H
**
*.SEEDPROM
X0 SET_H VPB sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X1 VPB IN 4 VPB 12 sky130_fd_pr__pfet_01v8__example_55959141808430
X2 SET_H SET_H 11 sky130_fd_pr__nfet_01v8__example_55959141808383
X3 SET_H RST_H 10 sky130_fd_pr__nfet_01v8__example_55959141808382
X4 SET_H 4 IN 12 sky130_fd_pr__nfet_01v8__example_55959141808423
X5 SET_H HLD_H_N 10 15 sky130_fd_pr__nfet_01v8__example_55959141808428
X6 SET_H 11 10 sky130_fd_pr__nfet_01v8__example_55959141808424
X7 SET_H HLD_H_N 13 11 sky130_fd_pr__nfet_01v8__example_55959141808429
X8 SET_H 12 14 sky130_fd_pr__nfet_01v8__example_55959141808427
X9 SET_H 4 16 sky130_fd_pr__nfet_01v8__example_55959141808427
X10 SET_H VPB 14 13 sky130_fd_pr__nfet_01v8__example_55959141808426
X11 SET_H VPB 14 13 sky130_fd_pr__nfet_01v8__example_55959141808426
X12 SET_H VPB 16 15 sky130_fd_pr__nfet_01v8__example_55959141808426
X13 SET_H VPB 16 15 sky130_fd_pr__nfet_01v8__example_55959141808426
X14 VCC_IO 10 OUT_H_N sky130_fd_pr__pfet_01v8__example_55959141808432
X15 VCC_IO 11 OUT_H sky130_fd_pr__pfet_01v8__example_55959141808431
X17 SET_H 11 OUT_H sky130_fd_pr__nfet_01v8__example_55959141808380
X18 VCC_IO 10 11 sky130_fd_pr__pfet_01v8__example_55959141808435
X19 VCC_IO 11 10 sky130_fd_pr__pfet_01v8__example_55959141808433
X20 SET_H 10 OUT_H_N sky130_fd_pr__nfet_01v8__example_55959141808379
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_octl VGND VCC_IO DM_H[2] DM_H[0] 6 DM_H[1] 8 DM_H_N[1] DM_H_N[2] DM_H_N[0] 12 13 PDEN_H_N[0] PDEN_H_N[1] VPWR SLOW_H SLOW_H_N HLD_I_H_N SLOW OD_H
**
*.SEEDPROM
X0 VGND VCC_IO 37 45 sky130_fd_io__hvsbt_inv_x1
X1 VGND VCC_IO 39 46 sky130_fd_io__hvsbt_inv_x1
X2 VGND VCC_IO 44 47 sky130_fd_io__hvsbt_inv_x1
X3 VGND VCC_IO 45 48 sky130_fd_io__hvsbt_inv_x1
X4 VGND VCC_IO 43 49 sky130_fd_io__hvsbt_inv_x1
X5 VGND VCC_IO 48 12 sky130_fd_io__hvsbt_inv_x2
X6 VGND VCC_IO 49 13 sky130_fd_io__hvsbt_inv_x2
X7 VGND VCC_IO 46 PDEN_H_N[0] sky130_fd_io__hvsbt_inv_x2
X8 VGND VCC_IO 47 PDEN_H_N[1] sky130_fd_io__hvsbt_inv_x2
X9 VGND VCC_IO DM_H[1] DM_H[0] 35 sky130_fd_io__hvsbt_nor
X10 VGND VCC_IO DM_H_N[2] DM_H_N[1] 36 sky130_fd_io__hvsbt_nor
X11 VGND VCC_IO 26 DM_H_N[1] 43 sky130_fd_io__hvsbt_nor
X12 VGND VCC_IO DM_H[2] 35 8 sky130_fd_io__hvsbt_nand2
X13 VGND VCC_IO PUEN_2OR1_H VCC_IO 37 sky130_fd_io__hvsbt_nand2
X14 VGND VCC_IO 36 DM_H_N[0] 40 sky130_fd_io__hvsbt_nand2
X15 VGND VCC_IO DM_H[1] DM_H[0] 39 sky130_fd_io__hvsbt_nand2
X16 VGND VCC_IO DM_H_N[2] DM_H_N[1] 41 sky130_fd_io__hvsbt_nand2
X17 VGND VCC_IO 42 40 PUEN_2OR1_H sky130_fd_io__hvsbt_nand2
X18 VGND VCC_IO 28 DM_H[0] 42 sky130_fd_io__hvsbt_nand2
X19 VGND VCC_IO DM_H_N[0] 41 44 sky130_fd_io__hvsbt_nand2
X20 VGND DM_H[2] VGND 23 sky130_fd_pr__nfet_01v8__example_55959141808417
X21 VGND DM_H[2] VGND 24 sky130_fd_pr__nfet_01v8__example_55959141808417
X22 VGND DM_H[2] VGND 31 sky130_fd_pr__nfet_01v8__example_55959141808417
X23 VGND DM_H[2] VGND 32 sky130_fd_pr__nfet_01v8__example_55959141808417
X24 VGND DM_H[0] 31 26 sky130_fd_pr__nfet_01v8__example_55959141808417
X25 VGND DM_H[1] 32 28 sky130_fd_pr__nfet_01v8__example_55959141808417
X26 VGND 6 33 26 sky130_fd_pr__nfet_01v8__example_55959141808417
X27 VGND 22 34 28 sky130_fd_pr__nfet_01v8__example_55959141808417
X28 VGND 23 VGND 33 sky130_fd_pr__nfet_01v8__example_55959141808417
X29 VGND 24 VGND 34 sky130_fd_pr__nfet_01v8__example_55959141808417
X30 VGND DM_H[0] VGND 6 sky130_fd_pr__nfet_01v8__example_55959141808417
X31 VGND DM_H[1] VGND 22 sky130_fd_pr__nfet_01v8__example_55959141808417
X32 VCC_IO 6 25 26 sky130_fd_pr__pfet_01v8__example_55959141808416
X33 VCC_IO 6 25 26 sky130_fd_pr__pfet_01v8__example_55959141808416
X34 VCC_IO 22 27 28 sky130_fd_pr__pfet_01v8__example_55959141808416
X35 VCC_IO 22 27 28 sky130_fd_pr__pfet_01v8__example_55959141808416
X36 VCC_IO 23 29 26 sky130_fd_pr__pfet_01v8__example_55959141808416
X37 VCC_IO 23 29 26 sky130_fd_pr__pfet_01v8__example_55959141808416
X38 VCC_IO 24 30 28 sky130_fd_pr__pfet_01v8__example_55959141808416
X39 VCC_IO 24 30 28 sky130_fd_pr__pfet_01v8__example_55959141808416
X40 VCC_IO DM_H[2] 25 23 ICV_16
X41 VCC_IO DM_H[2] 25 23 ICV_16
X42 VCC_IO DM_H[2] 27 24 ICV_16
X43 VCC_IO DM_H[2] 27 24 ICV_16
X44 VCC_IO DM_H[0] 6 29 ICV_16
X45 VCC_IO DM_H[0] 6 29 ICV_16
X46 VCC_IO DM_H[1] 22 30 ICV_16
X47 VCC_IO DM_H[1] 22 30 ICV_16
X48 VGND VCC_IO VPWR 50 HLD_I_H_N SLOW OD_H SLOW_H_N SLOW_H sky130_fd_io__com_ctl_ls_octl
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808389 2 3 4 5
**
*.SEEDPROM
XM0 2 3 5 2 sky130_fd_pr__pfet_01v8_hvt L=0.25 W=3 m=1
XM1 3 4 2 2 sky130_fd_pr__pfet_01v8_hvt L=0.25 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808375 1 2 3 4
**
XM0 4 2 1 1 sky130_fd_pr__nfet_01v8 L=0.25 W=1 m=1
XM1 1 2 4 1 sky130_fd_pr__nfet_01v8 L=0.25 W=1 m=1
XM2 2 3 1 1 sky130_fd_pr__nfet_01v8 L=0.25 W=1 m=1
XM3 1 3 2 1 sky130_fd_pr__nfet_01v8 L=0.25 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808387 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808388 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 m=1
XM1 1 2 3 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 m=1
.ENDS
***************************************
.SUBCKT ICV_17 1 2 3 4 5 6
**
X0 1 2 4 5 sky130_fd_pr__nfet_01v8__example_55959141808387
X1 1 3 6 sky130_fd_pr__nfet_01v8__example_55959141808388
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808376 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808377 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808386 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
XM1 3 2 4 1 sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__tpl1__example_55959141808374
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808384 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808381 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808392 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808393 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808391 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808390 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpio_dat_lsv2 VGND VCC_IO VPWR_KA 4 RST_H SET_H HLD_H_N IN OUT_H OUT_H_N
**
*.SEEDPROM
X0 VGND RST_H 4 sky130_fd_pr__nfet_01v8__example_55959141808383
X1 VGND SET_H 11 sky130_fd_pr__nfet_01v8__example_55959141808382
X2 VGND 4 OUT_H_N sky130_fd_pr__nfet_01v8__example_55959141808380
X3 VGND 11 OUT_H sky130_fd_pr__nfet_01v8__example_55959141808379
X6 VPWR_KA 13 IN 12 sky130_fd_pr__pfet_01v8__example_55959141808389
X7 VGND 13 IN 12 sky130_fd_pr__nfet_01v8__example_55959141808375
X8 VGND VPWR_KA 12 16 17 15 ICV_17
X9 VGND VPWR_KA 12 16 17 15 ICV_17
X10 VGND VPWR_KA 12 16 17 15 ICV_17
X11 VGND VPWR_KA 12 16 17 15 ICV_17
X12 VGND VPWR_KA 13 16 17 17 ICV_17
X13 VGND VPWR_KA 13 16 17 17 ICV_17
X14 VGND VPWR_KA 13 16 17 17 ICV_17
X15 VGND VPWR_KA 13 16 17 17 ICV_17
X16 VGND HLD_H_N 4 16 sky130_fd_pr__nfet_01v8__example_55959141808376
X17 VGND HLD_H_N 14 11 sky130_fd_pr__nfet_01v8__example_55959141808377
X18 VGND VPWR_KA 14 15 sky130_fd_pr__nfet_01v8__example_55959141808386
X19 VGND VPWR_KA 14 15 sky130_fd_pr__nfet_01v8__example_55959141808386
X20 VGND VPWR_KA 14 15 sky130_fd_pr__nfet_01v8__example_55959141808386
X21 VGND VPWR_KA 14 15 sky130_fd_pr__nfet_01v8__example_55959141808386
X23 VGND 4 11 sky130_fd_pr__nfet_01v8__example_55959141808384
X24 VGND 11 4 sky130_fd_pr__nfet_01v8__example_55959141808381
X25 VCC_IO 11 OUT_H sky130_fd_pr__pfet_01v8__example_55959141808392
X26 VCC_IO 4 OUT_H_N sky130_fd_pr__pfet_01v8__example_55959141808393
X27 VCC_IO 11 4 sky130_fd_pr__pfet_01v8__example_55959141808391
X28 VCC_IO 4 11 sky130_fd_pr__pfet_01v8__example_55959141808390
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpio_dat_ls_1v2 VGND VCC_IO VPWR_KA RST_H SET_H HLD_H_N IN OUT_H OUT_H_N
**
*.SEEDPROM
X0 VGND RST_H 11 sky130_fd_pr__nfet_01v8__example_55959141808383
X1 VGND SET_H 10 sky130_fd_pr__nfet_01v8__example_55959141808382
X2 VGND 11 OUT_H_N sky130_fd_pr__nfet_01v8__example_55959141808380
X3 VGND 10 OUT_H sky130_fd_pr__nfet_01v8__example_55959141808379
X6 VPWR_KA 13 IN 12 sky130_fd_pr__pfet_01v8__example_55959141808389
X7 VGND 13 IN 12 sky130_fd_pr__nfet_01v8__example_55959141808375
X8 VGND VPWR_KA 12 16 17 15 ICV_17
X9 VGND VPWR_KA 12 16 17 15 ICV_17
X10 VGND VPWR_KA 12 16 17 15 ICV_17
X11 VGND VPWR_KA 12 16 17 15 ICV_17
X12 VGND VPWR_KA 13 16 17 17 ICV_17
X13 VGND VPWR_KA 13 16 17 17 ICV_17
X14 VGND VPWR_KA 13 16 17 17 ICV_17
X15 VGND VPWR_KA 13 16 17 17 ICV_17
X16 VGND HLD_H_N 11 16 sky130_fd_pr__nfet_01v8__example_55959141808376
X17 VGND HLD_H_N 14 10 sky130_fd_pr__nfet_01v8__example_55959141808377
X18 VGND VPWR_KA 14 15 sky130_fd_pr__nfet_01v8__example_55959141808386
X19 VGND VPWR_KA 14 15 sky130_fd_pr__nfet_01v8__example_55959141808386
X20 VGND VPWR_KA 14 15 sky130_fd_pr__nfet_01v8__example_55959141808386
X21 VGND VPWR_KA 14 15 sky130_fd_pr__nfet_01v8__example_55959141808386
X23 VGND 11 10 sky130_fd_pr__nfet_01v8__example_55959141808384
X24 VGND 10 11 sky130_fd_pr__nfet_01v8__example_55959141808381
X25 VCC_IO 10 OUT_H sky130_fd_pr__pfet_01v8__example_55959141808392
X26 VCC_IO 11 OUT_H_N sky130_fd_pr__pfet_01v8__example_55959141808393
X27 VCC_IO 10 11 sky130_fd_pr__pfet_01v8__example_55959141808391
X28 VCC_IO 11 10 sky130_fd_pr__pfet_01v8__example_55959141808390
.ENDS
***************************************
.SUBCKT sky130_fd_pr__tpl1__example_55959141808625
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808406 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
XM1 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__via_pol1__example_55959141808396
**
.ENDS
***************************************
.SUBCKT ICV_18
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808404 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
XM1 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
XM2 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
XM3 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
XM4 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
XM5 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
.ENDS
***************************************
.SUBCKT ICV_19
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808409 2 3 4 5
**
*.SEEDPROM
XM0 5 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__com_cclat VGND VCC_IO OE_H_N PU_DIS_H DRVLO_H_N DRVHI_H PD_DIS_H
**
*.SEEDPROM
XM0 12 8 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
XM1 15 8 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
XM2 VGND 8 15 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
XM3 15 8 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
XM4 VGND 8 15 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 m=1
XM5 DRVHI_H 10 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM6 VCC_IO 10 DRVHI_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM7 DRVHI_H 10 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM8 VCC_IO 10 DRVHI_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM9 DRVHI_H 10 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM10 VCC_IO 10 DRVHI_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM11 DRVLO_H_N 11 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM12 VCC_IO 11 DRVLO_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM13 DRVLO_H_N 11 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM14 VCC_IO 11 DRVLO_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM15 DRVLO_H_N 11 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM16 VCC_IO 11 DRVLO_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM17 13 12 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM18 VCC_IO 12 13 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM19 13 12 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM20 VCC_IO 12 13 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM21 13 12 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM22 VCC_IO 12 13 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM23 13 12 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
XM24 VCC_IO 12 13 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 m=1
X32 VGND OE_H_N VGND 8 sky130_fd_pr__nfet_01v8__example_55959141808429
X38 VGND DRVLO_H_N 16 15 sky130_fd_pr__nfet_01v8__example_55959141808362
X39 VGND 9 16 10 sky130_fd_pr__nfet_01v8__example_55959141808362
X40 VGND PU_DIS_H VGND 9 sky130_fd_pr__nfet_01v8__example_55959141808360
X50 VCC_IO DRVHI_H 14 13 sky130_fd_pr__pfet_01v8__example_55959141808346
X51 VCC_IO PD_DIS_H 14 11 sky130_fd_pr__pfet_01v8__example_55959141808346
X54 VGND 12 11 sky130_fd_pr__nfet_01v8__example_55959141808406
X55 VGND DRVHI_H 11 sky130_fd_pr__nfet_01v8__example_55959141808406
X56 VGND PD_DIS_H 11 sky130_fd_pr__nfet_01v8__example_55959141808406
X62 VGND 11 DRVLO_H_N sky130_fd_pr__nfet_01v8__example_55959141808404
X63 VGND 10 DRVHI_H sky130_fd_pr__nfet_01v8__example_55959141808404
X68 VCC_IO OE_H_N VCC_IO 8 sky130_fd_pr__pfet_01v8__example_55959141808409
X69 VCC_IO 8 VCC_IO 12 sky130_fd_pr__pfet_01v8__example_55959141808409
X70 VCC_IO PU_DIS_H 9 VCC_IO sky130_fd_pr__pfet_01v8__example_55959141808409
X71 VCC_IO 8 10 VCC_IO sky130_fd_pr__pfet_01v8__example_55959141808409
X72 VCC_IO 9 VCC_IO 10 sky130_fd_pr__pfet_01v8__example_55959141808409
X73 VCC_IO DRVLO_H_N VCC_IO 10 sky130_fd_pr__pfet_01v8__example_55959141808409
.ENDS
***************************************
.SUBCKT sky130_fd_io__com_opath_datoev2 VGND VCC_IO VPWR_KA HLD_I_OVR_H OD_H 6 OE_N DRVHI_H DRVLO_H_N OUT
**
*.SEEDPROM
X0 VGND VPWR_KA sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X1 VGND VCC_IO VPWR_KA 11 VGND OD_H HLD_I_OVR_H OE_N 12 OE_H sky130_fd_io__gpio_dat_lsv2
X2 VGND VCC_IO VPWR_KA VGND OD_H HLD_I_OVR_H OUT 6 13 sky130_fd_io__gpio_dat_ls_1v2
X5 VGND VCC_IO 12 13 DRVLO_H_N DRVHI_H 6 sky130_fd_io__com_cclat
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_octl_dat VGND VGND_IO VCC_IO 5 OD_H 7 8 9 10 11 12 13 14 15 16 17 PU_H_N[2] 19 PU_H_N[0] PD_H[0]
+ 22 PD_H[1] PU_H_N[1] PD_H[3] DM_H[0] DM_H[1] DM_H[2] PU_H_N[3] PD_H[2] PD_H[4] VPWR DM_H_N[1] HLD_I_H_N SLOW VPWR_KA OE_N HLD_I_OVR_H DM_H_N[0] DM_H_N[2] OUT
+ 42
**
*.SEEDPROM
X0 VGND VGND_IO VCC_IO DRVHI_H 44 DRVLO_H_N 51 50 49 PD_H[0] PU_H_N[1] PU_H_N[0] 5 PD_H[1] 11 12 14 15 17 PU_H_N[2]
+ 19 7 8 9 10 13 16 22 PD_H[3] SLOW_H_N PU_H_N[3] 52 46 PD_H[2] PD_H[4] 42
+ sky130_fd_io__gpiov2_obpredrvr
X1 VGND VCC_IO DM_H[2] DM_H[0] 43 DM_H[1] 52 DM_H_N[1] DM_H_N[2] DM_H_N[0] 49 44 51 50 VPWR 46 SLOW_H_N HLD_I_H_N SLOW OD_H sky130_fd_io__gpiov2_octl
X2 VGND VCC_IO VPWR_KA HLD_I_OVR_H OD_H 47 OE_N DRVHI_H DRVLO_H_N OUT sky130_fd_io__com_opath_datoev2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__model__pfet_highvoltage__example_55959141808616 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
XM1 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
XM2 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
XM3 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__hvsbt_inv_x4 1 2 IN OUT
**
*.SEEDPROM
XM0 OUT IN 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
XM1 1 IN OUT 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
XM2 OUT IN 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
XM3 1 IN OUT 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
X4 2 IN OUT sky130_fd_pr__model__pfet_highvoltage__example_55959141808616
X5 2 IN OUT sky130_fd_pr__model__pfet_highvoltage__example_55959141808616
.ENDS
***************************************
.SUBCKT sky130_fd_io__com_ctl_ls SET_H VCC_IO VPB VPWR HLD_H_N IN RST_H OUT_H
**
*.SEEDPROM
X0 SET_H VPB sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X1 VPB IN 12 VPWR 11 sky130_fd_pr__pfet_01v8__example_55959141808430
X2 SET_H SET_H 10 sky130_fd_pr__nfet_01v8__example_55959141808383
X3 SET_H RST_H 9 sky130_fd_pr__nfet_01v8__example_55959141808382
X4 SET_H 12 IN 11 sky130_fd_pr__nfet_01v8__example_55959141808423
X5 SET_H HLD_H_N 9 16 sky130_fd_pr__nfet_01v8__example_55959141808428
X6 SET_H 10 9 sky130_fd_pr__nfet_01v8__example_55959141808424
X7 SET_H HLD_H_N 13 10 sky130_fd_pr__nfet_01v8__example_55959141808429
X8 SET_H 11 15 sky130_fd_pr__nfet_01v8__example_55959141808427
X9 SET_H 12 17 sky130_fd_pr__nfet_01v8__example_55959141808427
X10 SET_H VPWR 15 13 sky130_fd_pr__nfet_01v8__example_55959141808426
X11 SET_H VPWR 15 13 sky130_fd_pr__nfet_01v8__example_55959141808426
X12 SET_H VPWR 17 16 sky130_fd_pr__nfet_01v8__example_55959141808426
X13 SET_H VPWR 17 16 sky130_fd_pr__nfet_01v8__example_55959141808426
X14 VCC_IO 9 OUT_H_N sky130_fd_pr__pfet_01v8__example_55959141808432
X15 VCC_IO 10 OUT_H sky130_fd_pr__pfet_01v8__example_55959141808431
X17 SET_H 10 OUT_H sky130_fd_pr__nfet_01v8__example_55959141808380
X18 VCC_IO 9 10 sky130_fd_pr__pfet_01v8__example_55959141808435
X19 VCC_IO 10 9 sky130_fd_pr__pfet_01v8__example_55959141808433
X20 SET_H 9 OUT_H_N sky130_fd_pr__nfet_01v8__example_55959141808379
.ENDS
***************************************
.SUBCKT sky130_fd_pr__model__pfet_highvoltage__example_55959141808614 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
XM1 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
XM2 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
XM3 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
XM4 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
XM5 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
XM6 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
XM7 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__model__nfet_highvoltage__example_55959141808613 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
XM1 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
XM2 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
XM3 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
XM4 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
XM5 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
XM6 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
XM7 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__com_ctl_hldv2 VGND VCC_IO 3 4 5 OD_I_H HLD_I_H HLD_OVR HLD_I_H_N VPWR
**
*.SEEDPROM
R0 HLD_I_H 11 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R1 15 HLD_I_H_N sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R2 HLD_I_H_N 16 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
X3 VGND VCC_IO 3 12 sky130_fd_io__hvsbt_inv_x1
X4 VGND VCC_IO 13 14 sky130_fd_io__hvsbt_inv_x1
X5 VGND VCC_IO 12 17 sky130_fd_io__hvsbt_inv_x1
X6 VGND VCC_IO OD_I_H 18 5 sky130_fd_io__hvsbt_nor
X7 VGND VCC_IO 14 19 18 sky130_fd_io__hvsbt_nor
X8 VGND VCC_IO 3 4 13 sky130_fd_io__hvsbt_nand2
X9 VGND VCC_IO 14 11 sky130_fd_io__hvsbt_inv_x4
X10 VGND VCC_IO 17 OD_I_H sky130_fd_io__hvsbt_inv_x4
X11 VGND VCC_IO VPWR VPWR 14 HLD_OVR 12 19 sky130_fd_io__com_ctl_ls
X12 VCC_IO 11 15 sky130_fd_pr__model__pfet_highvoltage__example_55959141808614
X13 VCC_IO 11 15 sky130_fd_pr__model__pfet_highvoltage__example_55959141808614
X14 VCC_IO 11 16 sky130_fd_pr__model__pfet_highvoltage__example_55959141808614
X15 VCC_IO 11 16 sky130_fd_pr__model__pfet_highvoltage__example_55959141808614
X16 VGND 11 15 sky130_fd_pr__model__nfet_highvoltage__example_55959141808613
X17 VGND 11 16 sky130_fd_pr__model__nfet_highvoltage__example_55959141808613
.ENDS
***************************************
.SUBCKT sky130_ef_io__gpiov2_pad_wrapped VSSD VSSA VSSIO VSSIO_Q VDDIO VDDIO_Q PAD PAD_A_ESD_0_H IB_MODE_SEL ENABLE_INP_H ENABLE_H VDDA VCCD OE_N ENABLE_VDDA_H VTRIP_SEL VCCHIB ENABLE_VSWITCH_H OUT HLD_OVR
+ DM[2] ANALOG_SEL HLD_H_N ANALOG_EN INP_DIS ANALOG_POL DM[0] DM[1] SLOW IN ENABLE_VDDIO TIE_LO_ESD VSWITCH AMUXBUS_A AMUXBUS_B
**
X0 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X1 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X2 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X3 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X4 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X5 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw m=1
R6 PAD_A_NOESD_H PAD sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R7 PAD_A_NOESD_H PAD sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R8 PAD_A_NOESD_H PAD sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
X9 PAD_A_ESD_1_H 41 sky130_fd_io__res75only_small
X10 41 PAD sky130_fd_io__res75only_small
X11 42 PAD sky130_fd_io__res75only_small
X12 PAD_A_ESD_0_H 42 sky130_fd_io__res75only_small
X13 VSSD VDDIO_Q 57 59 sky130_fd_io__hvsbt_inv_x1
X14 VSSD VDDIO_Q ENABLE_INP_H ENABLE_H 60 sky130_fd_io__hvsbt_nor
X15 VSSD VDDIO_Q 58 ENABLE_INP_H 57 sky130_fd_io__hvsbt_nand2
X16 VSSD VSSIO_Q VSSA 37 36 38 39 VSWITCH VDDIO_Q VDDA 74 PAD VCCD 86 ENABLE_VDDA_H ENABLE_VSWITCH_H AMUXBUS_B AMUXBUS_A ANALOG_SEL ANALOG_EN
+ OUT ANALOG_POL 73
+ sky130_fd_io__gpiov2_amux
X17 VSSD VDDIO_Q VCCD IB_MODE_SEL 73 58 82 81 63 79 60 DM[0] INP_DIS 59 78 75 76 DM[2] 72 VTRIP_SEL
+ 68 69 DM[1]
+ sky130_fd_io__gpiov2_ctl_lsbank
X18 VSSD VSSIO VDDIO TIE_LO_ESD 64 77 62 87 PAD 66 65 67 83 TIE_HI_ESD 55 sky130_fd_io__gpio_odrvrv2
X19 VSSD VDDIO_Q ENABLE_VDDIO 63 IN_H 70 PAD IN VCCHIB 81 75 78 68 69 72 sky130_fd_io__gpiov2_ipath
X20 VSSD VSSIO VDDIO 43 58 44 45 46 47 48 49 50 51 52 54 53 55 56 64 65
+ 61 66 67 62 79 82 76 83 77 87 VCCD 81 73 SLOW VCCHIB OE_N 71 63 75 OUT
+ 88
+ sky130_fd_io__gpiov2_octl_dat
X21 VSSD VDDIO_Q ENABLE_H HLD_H_N 71 58 74 HLD_OVR 73 VCCD sky130_fd_io__com_ctl_hldv2
.ENDS
***************************************
.SUBCKT sky130_ef_io__vssio_hvc_clamped_pad VSSD VDDIO VSSIO 12
**
*.CALIBRE ISOLATED NETS: VCCHIB VCCD VDDA VSWITCH VSSA AMUXBUS_B AMUXBUS_A VDDIO_Q
X0 VSSD VSSIO VDDIO VDDIO VSSIO 12 sky130_fd_io__top_ground_hvc_wpad
*.CALIBRE WARNING SHORT Short circuit(s) detected by extraction in this cell. See extraction report for details.
*.CALIBRE WARNING OPEN Open circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT sky130_ef_io__vssd_lvc_clamped_pad VSSD VSSIO VCCD VDDIO 13
**
*.CALIBRE ISOLATED NETS: VCCHIB VDDA VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
X0 VSSD VSSD VSSD VCCD VDDIO VCCD VSSIO VSSD 13 sky130_fd_io__top_ground_lvc_wpad
*.CALIBRE WARNING OPEN Open circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 2 3
**
R0 2 4 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R1 5 3 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_p_em1c_cdns_55959141808753 2
**
R0 2 3 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R1 2 4 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT ICV_20 2 3
**
X0 2 3 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X1 2 sky130_fd_io__xres_p_em1c_cdns_55959141808753
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_generic_nd__example_55959141808754 2 3
**
*.SEEDPROM
R0 2 3 sky130_fd_pr__res_generic_nd L=14 W=0.5 m=1
.ENDS
***************************************
.SUBCKT ICV_21 2 3 4 5
**
*.SEEDPROM
X0 2 3 sky130_fd_pr__res_generic_nd__example_55959141808754
X1 4 5 sky130_fd_pr__res_generic_nd__example_55959141808754
.ENDS
***************************************
.SUBCKT ICV_22 2 3 4 5 6 7 8 9
**
*.SEEDPROM
X0 4 2 3 5 ICV_21
X1 8 6 7 9 ICV_21
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758 2 3
**
R0 2 4 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R1 5 3 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1c_cdns_55959141808760 2
**
R0 2 3 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R1 2 4 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1c_cdns_55959141808761 2
**
R0 2 3 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R1 2 4 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd__example_55959141808338
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd2__example_55959141808337
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_23
**
.ENDS
***************************************
.SUBCKT ICV_24
**
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759 1
**
R0 1 2 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R1 1 3 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT ICV_25 2 3 4
**
X0 2 3 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X1 4 sky130_fd_io__xres_p_em1c_cdns_55959141808753
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1o_cdns_55959141808756 1 2
**
R0 2 3 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
R1 4 1 sky130_fd_pr__res_generic_po m=1 w=480000u l=45000u
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_generic_nd__example_55959141808755 2 3
**
*.SEEDPROM
R0 2 3 sky130_fd_pr__res_generic_nd L=47 W=0.5 m=1
.ENDS
***************************************
.SUBCKT ICV_26 2 3 4
**
*.SEEDPROM
X0 2 3 sky130_fd_pr__res_generic_nd__example_55959141808754
X1 4 2 sky130_fd_pr__res_generic_nd__example_55959141808755
.ENDS
***************************************
.SUBCKT ICV_27 2 3
**
*.SEEDPROM
X0 2 2 sky130_fd_pr__res_generic_nd__example_55959141808754
X1 2 3 sky130_fd_pr__res_generic_nd__example_55959141808755
.ENDS
***************************************
.SUBCKT ICV_28 2 3 4 5 6
**
*.SEEDPROM
X0 3 4 2 ICV_26
X1 5 6 ICV_27
.ENDS
***************************************
.SUBCKT ICV_29 2 3 4 5 6 7 8 9 10 11
**
*.SEEDPROM
X0 2 4 6 5 3 ICV_28
X1 7 9 11 10 8 ICV_28
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres2v2_rcfilter_lpfv2 1 VCC_IO 3 4 5 6 7 8 9 10 11 12 13 IN
**
XM0 1 3 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 m=1
XM1 1 4 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 m=1
XM2 1 5 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 m=1
XM3 1 6 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 m=1
XM4 1 7 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 m=1
XM5 1 8 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 m=1
XM6 1 9 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 m=1
XM7 1 10 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 m=1
XM8 1 11 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 m=1
XM9 1 11 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 m=1
XM10 1 12 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 m=1
XM11 1 13 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 m=1
XM12 VCC_IO 3 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 m=1
XM13 VCC_IO 4 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 m=1
XM14 VCC_IO 5 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 m=1
XM15 VCC_IO 6 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 m=1
XM16 VCC_IO 7 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 m=1
XM17 VCC_IO 8 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 m=1
XM18 VCC_IO 9 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 m=1
XM19 VCC_IO 10 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 m=1
XM20 VCC_IO 11 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 m=1
XM21 VCC_IO 11 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 m=1
XM22 VCC_IO 12 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 m=1
XM23 VCC_IO 13 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 m=1
X24 1 8 sky130_fd_pr__diode_pw2nd_05v5 m=1
X25 1 1 sky130_fd_pr__diode_pw2nd_05v5 m=1
X26 1 7 sky130_fd_pr__diode_pw2nd_05v5 m=1
X27 1 1 sky130_fd_pr__diode_pw2nd_05v5 m=1
X28 1 6 sky130_fd_pr__diode_pw2nd_05v5 m=1
X29 1 1 sky130_fd_pr__diode_pw2nd_05v5 m=1
X30 1 5 sky130_fd_pr__diode_pw2nd_05v5 m=1
X31 1 1 sky130_fd_pr__diode_pw2nd_05v5 m=1
X32 1 4 sky130_fd_pr__diode_pw2nd_05v5 m=1
X33 1 3 sky130_fd_pr__diode_pw2nd_05v5 m=1
X34 1 3 sky130_fd_pr__diode_pw2nd_05v5 m=1
X35 1 9 sky130_fd_pr__diode_pw2nd_05v5 m=1
X36 1 15 sky130_fd_pr__diode_pw2nd_05v5 m=1
X37 1 15 sky130_fd_pr__diode_pw2nd_05v5 m=1
X38 1 16 sky130_fd_pr__diode_pw2nd_05v5 m=1
X39 1 16 sky130_fd_pr__diode_pw2nd_05v5 m=1
X40 1 17 sky130_fd_pr__diode_pw2nd_05v5 m=1
X41 1 17 sky130_fd_pr__diode_pw2nd_05v5 m=1
X42 1 18 sky130_fd_pr__diode_pw2nd_05v5 m=1
X43 1 18 sky130_fd_pr__diode_pw2nd_05v5 m=1
X44 1 19 sky130_fd_pr__diode_pw2nd_05v5 m=1
X45 1 19 sky130_fd_pr__diode_pw2nd_05v5 m=1
X46 1 20 sky130_fd_pr__diode_pw2nd_05v5 m=1
X47 1 20 sky130_fd_pr__diode_pw2nd_05v5 m=1
X48 1 21 sky130_fd_pr__diode_pw2nd_05v5 m=1
X49 1 1 sky130_fd_pr__diode_pw2nd_05v5 m=1
X50 1 22 sky130_fd_pr__diode_pw2nd_05v5 m=1
X51 1 1 sky130_fd_pr__diode_pw2nd_05v5 m=1
X52 1 23 sky130_fd_pr__diode_pw2nd_05v5 m=1
X53 1 1 sky130_fd_pr__diode_pw2nd_05v5 m=1
X54 1 24 sky130_fd_pr__diode_pw2nd_05v5 m=1
X55 1 1 sky130_fd_pr__diode_pw2nd_05v5 m=1
X56 1 25 sky130_fd_pr__diode_pw2nd_05v5 m=1
X57 1 3 sky130_fd_pr__diode_pw2nd_05v5 m=1
X58 1 26 sky130_fd_pr__diode_pw2nd_05v5 m=1
X59 1 9 sky130_fd_pr__diode_pw2nd_05v5 m=1
X60 1 15 sky130_fd_pr__diode_pw2nd_05v5 m=1
X61 1 27 sky130_fd_pr__diode_pw2nd_05v5 m=1
X62 1 16 sky130_fd_pr__diode_pw2nd_05v5 m=1
X63 1 28 sky130_fd_pr__diode_pw2nd_05v5 m=1
X64 1 17 sky130_fd_pr__diode_pw2nd_05v5 m=1
X65 1 29 sky130_fd_pr__diode_pw2nd_05v5 m=1
X66 1 18 sky130_fd_pr__diode_pw2nd_05v5 m=1
X67 1 30 sky130_fd_pr__diode_pw2nd_05v5 m=1
X68 1 19 sky130_fd_pr__diode_pw2nd_05v5 m=1
X69 1 31 sky130_fd_pr__diode_pw2nd_05v5 m=1
X70 1 20 sky130_fd_pr__diode_pw2nd_05v5 m=1
X71 1 32 sky130_fd_pr__diode_pw2nd_05v5 m=1
X72 1 33 sky130_fd_pr__diode_pw2nd_05v5 m=1
X73 1 33 sky130_fd_pr__diode_pw2nd_05v5 m=1
X74 1 34 sky130_fd_pr__diode_pw2nd_05v5 m=1
X75 1 34 sky130_fd_pr__diode_pw2nd_05v5 m=1
X76 1 35 sky130_fd_pr__diode_pw2nd_05v5 m=1
X77 1 35 sky130_fd_pr__diode_pw2nd_05v5 m=1
X78 1 36 sky130_fd_pr__diode_pw2nd_05v5 m=1
X79 1 36 sky130_fd_pr__diode_pw2nd_05v5 m=1
X80 1 37 sky130_fd_pr__diode_pw2nd_05v5 m=1
X81 1 37 sky130_fd_pr__diode_pw2nd_05v5 m=1
X82 1 38 sky130_fd_pr__diode_pw2nd_05v5 m=1
X83 1 38 sky130_fd_pr__diode_pw2nd_05v5 m=1
X84 1 IN sky130_fd_pr__diode_pw2nd_05v5 m=1
X85 1 13 sky130_fd_pr__diode_pw2nd_05v5 m=1
X86 1 13 sky130_fd_pr__diode_pw2nd_05v5 m=1
X87 1 12 sky130_fd_pr__diode_pw2nd_05v5 m=1
X88 1 12 sky130_fd_pr__diode_pw2nd_05v5 m=1
X89 1 11 sky130_fd_pr__diode_pw2nd_05v5 m=1
X90 1 11 sky130_fd_pr__diode_pw2nd_05v5 m=1
X91 1 11 sky130_fd_pr__diode_pw2nd_05v5 m=1
X92 1 11 sky130_fd_pr__diode_pw2nd_05v5 m=1
X93 1 10 sky130_fd_pr__diode_pw2nd_05v5 m=1
X94 1 10 sky130_fd_pr__diode_pw2nd_05v5 m=1
X95 1 9 sky130_fd_pr__diode_pw2nd_05v5 m=1
X96 1 38 sky130_fd_pr__diode_pw2nd_05v5 m=1
X97 1 39 sky130_fd_pr__diode_pw2nd_05v5 m=1
X98 1 37 sky130_fd_pr__diode_pw2nd_05v5 m=1
X99 1 40 sky130_fd_pr__diode_pw2nd_05v5 m=1
X100 1 36 sky130_fd_pr__diode_pw2nd_05v5 m=1
X101 1 41 sky130_fd_pr__diode_pw2nd_05v5 m=1
X102 1 35 sky130_fd_pr__diode_pw2nd_05v5 m=1
X103 1 42 sky130_fd_pr__diode_pw2nd_05v5 m=1
X104 1 34 sky130_fd_pr__diode_pw2nd_05v5 m=1
X105 1 43 sky130_fd_pr__diode_pw2nd_05v5 m=1
X106 1 33 sky130_fd_pr__diode_pw2nd_05v5 m=1
X107 1 44 sky130_fd_pr__diode_pw2nd_05v5 m=1
X108 1 45 sky130_fd_pr__diode_pw2nd_05v5 m=1
X109 1 10 sky130_fd_pr__diode_pw2nd_05v5 m=1
X110 1 46 sky130_fd_pr__diode_pw2nd_05v5 m=1
X111 1 11 sky130_fd_pr__diode_pw2nd_05v5 m=1
X112 1 47 sky130_fd_pr__diode_pw2nd_05v5 m=1
X113 1 11 sky130_fd_pr__diode_pw2nd_05v5 m=1
X114 1 48 sky130_fd_pr__diode_pw2nd_05v5 m=1
X115 1 12 sky130_fd_pr__diode_pw2nd_05v5 m=1
X116 1 49 sky130_fd_pr__diode_pw2nd_05v5 m=1
X117 1 13 sky130_fd_pr__diode_pw2nd_05v5 m=1
X118 1 50 sky130_fd_pr__diode_pw2nd_05v5 m=1
X119 1 IN sky130_fd_pr__diode_pw2nd_05v5 m=1
X120 1 44 sky130_fd_pr__diode_pw2nd_05v5 m=1
X121 1 33 sky130_fd_pr__diode_pw2nd_05v5 m=1
X122 1 43 sky130_fd_pr__diode_pw2nd_05v5 m=1
X123 1 34 sky130_fd_pr__diode_pw2nd_05v5 m=1
X124 1 42 sky130_fd_pr__diode_pw2nd_05v5 m=1
X125 1 35 sky130_fd_pr__diode_pw2nd_05v5 m=1
X126 1 41 sky130_fd_pr__diode_pw2nd_05v5 m=1
X127 1 36 sky130_fd_pr__diode_pw2nd_05v5 m=1
X128 1 40 sky130_fd_pr__diode_pw2nd_05v5 m=1
X129 1 37 sky130_fd_pr__diode_pw2nd_05v5 m=1
X130 1 39 sky130_fd_pr__diode_pw2nd_05v5 m=1
X131 1 38 sky130_fd_pr__diode_pw2nd_05v5 m=1
X132 1 IN sky130_fd_pr__diode_pw2nd_05v5 m=1
X133 1 50 sky130_fd_pr__diode_pw2nd_05v5 m=1
X134 1 13 sky130_fd_pr__diode_pw2nd_05v5 m=1
X135 1 49 sky130_fd_pr__diode_pw2nd_05v5 m=1
X136 1 12 sky130_fd_pr__diode_pw2nd_05v5 m=1
X137 1 48 sky130_fd_pr__diode_pw2nd_05v5 m=1
X138 1 11 sky130_fd_pr__diode_pw2nd_05v5 m=1
X139 1 47 sky130_fd_pr__diode_pw2nd_05v5 m=1
X140 1 11 sky130_fd_pr__diode_pw2nd_05v5 m=1
X141 1 46 sky130_fd_pr__diode_pw2nd_05v5 m=1
X142 1 10 sky130_fd_pr__diode_pw2nd_05v5 m=1
X143 1 45 sky130_fd_pr__diode_pw2nd_05v5 m=1
X144 1 VCC_IO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X164 20 32 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X165 8 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X166 7 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X167 6 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X168 5 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X169 3 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X170 9 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X171 12 49 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X172 11 47 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X173 9 45 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X174 15 sky130_fd_io__xres_p_em1c_cdns_55959141808753
X175 IN sky130_fd_io__xres_p_em1c_cdns_55959141808753
X176 12 sky130_fd_io__xres_p_em1c_cdns_55959141808753
X177 11 sky130_fd_io__xres_p_em1c_cdns_55959141808753
X178 33 44 ICV_20
X179 34 43 ICV_20
X180 35 42 ICV_20
X181 36 41 ICV_20
X182 37 40 ICV_20
X183 38 39 ICV_20
X184 13 50 ICV_20
X185 11 48 ICV_20
X186 10 46 ICV_20
X187 34 43 34 34 33 44 33 33 ICV_22
X188 36 41 36 36 35 42 35 35 ICV_22
X189 38 39 38 38 37 40 37 37 ICV_22
X190 12 13 49 13 13 IN 50 IN ICV_22
X191 11 11 47 11 11 12 48 12 ICV_22
X192 9 10 45 10 10 11 46 11 ICV_22
X193 1 7 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758
X194 1 6 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758
X195 1 5 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758
X196 1 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758
X197 13 12 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758
X198 12 11 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758
X199 11 10 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758
X200 10 9 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758
X201 3 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808760
X202 11 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808760
X203 9 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808761
X204 4 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808761
X218 1 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759
X219 1 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759
X220 1 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759
X221 1 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759
X222 8 21 1 ICV_25
X223 7 22 1 ICV_25
X224 6 23 1 ICV_25
X225 5 24 1 ICV_25
X226 4 25 3 ICV_25
X227 3 26 9 ICV_25
X228 15 27 16 ICV_25
X229 16 28 17 ICV_25
X230 17 29 18 ICV_25
X231 18 30 19 ICV_25
X232 19 31 20 ICV_25
X233 1 9 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808756
X234 1 3 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808756
X235 32 20 IN ICV_26
X236 15 45 ICV_27
X237 13 31 19 20 50 ICV_28
X238 38 39 21 1 8 37 40 22 1 7 ICV_29
X239 36 41 23 1 6 35 42 24 1 5 ICV_29
X240 34 43 25 3 4 33 44 26 9 3 ICV_29
X241 10 46 27 16 15 11 47 28 17 16 ICV_29
X242 11 48 29 18 17 12 49 30 19 18 ICV_29
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_55959141808243
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808723 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_55959141808719
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808720 2 3 4 5
**
*.SEEDPROM
XM0 5 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=1 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_5595914180829
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808767 2 3 4 5
**
*.SEEDPROM
XM0 5 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_tie_r_out_esd A B
**
X0 A B sky130_fd_pr__res_generic_po__example_5595914180838
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_55959141808765
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808764 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808779 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808777 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_5595914180827
**
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808778 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
XM1 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808784 2 3 4
**
*.SEEDPROM
XM0 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=1 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808783 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd__example_55959141808782
**
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808786 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808787 2 3 4 5
**
*.SEEDPROM
XM0 5 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpio_buf_localesdv2 VGND VCC_IO VTRIP_SEL_H OUT_H 5
**
X0 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X1 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X2 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X3 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X4 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X5 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X6 5 OUT_H sky130_fd_io__res250only_small
X7 VGND VCC_IO VGND VGND OUT_VT 8 sky130_fd_io__signal_5_sym_hv_local_5term
X8 VGND VCC_IO VGND VGND OUT_H 10 sky130_fd_io__signal_5_sym_hv_local_5term
X9 VGND VCC_IO VGND OUT_VT VCC_IO 7 sky130_fd_io__signal_5_sym_hv_local_5term
X10 VGND VCC_IO VGND OUT_H VCC_IO 9 sky130_fd_io__signal_5_sym_hv_local_5term
X11 VGND VTRIP_SEL_H OUT_VT OUT_H sky130_fd_pr__nfet_01v8__example_55959141808555
.ENDS
***************************************
.SUBCKT sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2 1 2 VCC_IO 4 5 6 7 8 9 10 11 12 13 14
**
X0 1 VCC_IO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X1 2 VCC_IO sky130_fd_pr__model__parasitic__diode_pw2dn m=1
X2 1 VCC_IO sky130_fd_pr__model__parasitic__diode_ps2dn m=1
X5 2 4 14 sky130_fd_pr__nfet_01v8__example_55959141808647
X6 2 13 14 sky130_fd_pr__nfet_01v8__example_55959141808647
X7 2 13 14 sky130_fd_pr__nfet_01v8__example_55959141808647
X34 2 4 5 6 7 8 9 10 11 12 13 14 sky130_fd_pr__nfet_01v8__example_55959141808648
X35 2 4 5 6 7 8 9 10 11 12 13 14 sky130_fd_pr__nfet_01v8__example_55959141808651
X36 2 4 14 sky130_fd_pr__nfet_01v8__example_55959141808650
X37 2 4 14 sky130_fd_pr__nfet_01v8__example_55959141808650
X38 2 4 14 sky130_fd_pr__nfet_01v8__example_55959141808645
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpio_pddrvr_strong_xres4v2 1 TIE_LO_ESD 3 VCC_IO PD_H[2] PD_H[3] 7 8
**
X0 3 VCC_IO condiode m=1
X1 TIE_LO_ESD 7 sky130_fd_io__tk_em2s_cdns_55959141808652
X2 PD_H[2] 15 sky130_fd_io__tk_em2s_cdns_55959141808652
X3 PD_H[2] 14 sky130_fd_io__tk_em2s_cdns_55959141808652
X4 PD_H[3] 13 sky130_fd_io__tk_em2s_cdns_55959141808652
X5 PD_H[3] 12 sky130_fd_io__tk_em2s_cdns_55959141808652
X6 PD_H[3] 11 sky130_fd_io__tk_em2s_cdns_55959141808652
X7 PD_H[3] 10 sky130_fd_io__tk_em2s_cdns_55959141808652
X8 TIE_LO_ESD 9 sky130_fd_io__tk_em2s_cdns_55959141808652
X9 PD_H[3] 7 sky130_fd_io__tk_em2o_cdns_55959141808653
X10 PD_H[2] 7 sky130_fd_io__tk_em2o_cdns_55959141808653
X11 PD_H[3] 15 sky130_fd_io__tk_em2o_cdns_55959141808653
X12 TIE_LO_ESD 15 sky130_fd_io__tk_em2o_cdns_55959141808653
X13 PD_H[3] 14 sky130_fd_io__tk_em2o_cdns_55959141808653
X14 TIE_LO_ESD 14 sky130_fd_io__tk_em2o_cdns_55959141808653
X15 PD_H[2] 13 sky130_fd_io__tk_em2o_cdns_55959141808653
X16 TIE_LO_ESD 13 sky130_fd_io__tk_em2o_cdns_55959141808653
X17 PD_H[2] 12 sky130_fd_io__tk_em2o_cdns_55959141808653
X18 TIE_LO_ESD 12 sky130_fd_io__tk_em2o_cdns_55959141808653
X19 PD_H[2] 11 sky130_fd_io__tk_em2o_cdns_55959141808653
X20 TIE_LO_ESD 11 sky130_fd_io__tk_em2o_cdns_55959141808653
X21 PD_H[2] 10 sky130_fd_io__tk_em2o_cdns_55959141808653
X22 TIE_LO_ESD 10 sky130_fd_io__tk_em2o_cdns_55959141808653
X23 PD_H[2] 9 sky130_fd_io__tk_em2o_cdns_55959141808653
X24 PD_H[3] 9 sky130_fd_io__tk_em2o_cdns_55959141808653
X25 TIE_LO_ESD 3 sky130_fd_pr__res_generic_po__example_5595914180838
X26 1 3 VCC_IO 9 10 11 12 13 PD_H[2] PD_H[3] 14 15 7 8 sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2
.ENDS
***************************************
.SUBCKT sky130_fd_io__top_xres4v2 VSSD VDDIO VCCHIB VDDIO_Q ENABLE_H EN_VDDIO_SIG_H INP_SEL_H PAD PULLUP_H ENABLE_VDDIO DISABLE_PULLUP_H PAD_A_ESD_H VSSIO FILT_IN_H XRES_H_N TIE_WEAK_HI_H
**
*.CALIBRE ISOLATED NETS: VCCD VDDA VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q
R0 54 50 sky130_fd_pr__res_generic_nd__hv L=1077.19 W=0.29 m=1
XM1 61 37 59 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM2 59 37 61 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM3 61 37 59 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM4 59 37 61 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM5 VSSD 30 59 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM6 59 30 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM7 37 30 59 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM8 59 30 37 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM9 59 37 55 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 m=1
XM10 VSSD 31 51 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 m=1
XM11 51 31 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 m=1
XM12 VSSD 31 51 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 m=1
XM13 VSSD 40 60 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=1 W=0.42 m=1
XM14 40 43 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 m=1
XM15 24 34 58 VSSD sky130_fd_pr__nfet_05v0_nvt L=0.9 W=10 m=1
XM16 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_05v0_nvt L=0.9 W=10 m=1
XM17 50 30 37 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM18 VDDIO_Q 31 51 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
XM19 51 31 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
XM20 VDDIO_Q 31 51 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
XM21 VDDIO_Q 32 31 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
XM22 40 43 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 m=1
XM23 52 40 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=1 W=0.42 m=1
XM24 29 42 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM25 VDDIO 42 29 VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM26 29 42 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
XM27 VDDIO 42 29 VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 m=1
R28 44 26 sky130_fd_pr__res_generic_po W=0.4 m=1 w=480000u l=45000u
R29 28 29 sky130_fd_pr__res_generic_po W=0.8 m=1 w=480000u l=45000u
X30 VSSD 54 sky130_fd_pr__diode_pw2nd_11v0 m=1
X31 VSSD 50 sky130_fd_pr__diode_pw2nd_11v0 m=1
X32 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X33 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X34 VSSD VCCHIB sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X35 VSSD 24 sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X36 VSSD 25 sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X37 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X38 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X39 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X40 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X41 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X42 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X43 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X44 VSSD VCCHIB sky130_fd_pr__model__parasitic__diode_ps2nw m=1
X45 VSSD VDDIO_Q 63 34 sky130_fd_io__hvsbt_inv_x1
X46 VSSD VDDIO_Q 40 70 sky130_fd_io__hvsbt_inv_x1
X47 VSSD VDDIO 69 42 sky130_fd_io__hvsbt_inv_x2
X48 VSSD VDDIO DISABLE_PULLUP_H 69 sky130_fd_io__hvsbt_inv_x2
X49 VSSD VDDIO_Q INP_SEL_H 39 sky130_fd_io__hvsbt_inv_x2
X50 VSSD VDDIO_Q EN_VDDIO_SIG_H 35 sky130_fd_io__hvsbt_inv_x2
X55 VSSD VCCHIB ENABLE_VDDIO VCCHIB 36 VSSD sky130_fd_io__inv_1
X56 VSSD VDDIO_Q 35 ENABLE_H 63 sky130_fd_io__hvsbt_nand2
X57 27 45 sky130_fd_io__tk_em2s_cdns_55959141808652
X58 27 46 sky130_fd_io__tk_em2s_cdns_55959141808652
X59 27 47 sky130_fd_io__tk_em2s_cdns_55959141808652
X60 27 48 sky130_fd_io__tk_em2s_cdns_55959141808652
X61 27 49 sky130_fd_io__tk_em2s_cdns_55959141808652
X62 27 45 sky130_fd_io__tk_em2o_cdns_55959141808653
X63 27 45 sky130_fd_io__tk_em2o_cdns_55959141808653
X64 27 46 sky130_fd_io__tk_em2o_cdns_55959141808653
X65 27 46 sky130_fd_io__tk_em2o_cdns_55959141808653
X66 27 47 sky130_fd_io__tk_em2o_cdns_55959141808653
X67 27 47 sky130_fd_io__tk_em2o_cdns_55959141808653
X68 27 48 sky130_fd_io__tk_em2o_cdns_55959141808653
X69 27 48 sky130_fd_io__tk_em2o_cdns_55959141808653
X70 27 49 sky130_fd_io__tk_em2o_cdns_55959141808653
X71 27 49 sky130_fd_io__tk_em2o_cdns_55959141808653
X72 PAD PAD_A_ESD_H sky130_fd_io__res250only_small
X73 TIE_WEAK_HI_H 74 sky130_fd_io__res250only_small
X74 64 PULLUP_H sky130_fd_pr__res_generic_po__example_5595914180864
X75 66 64 sky130_fd_pr__res_generic_po__example_5595914180864
X76 67 66 sky130_fd_pr__res_generic_po__example_5595914180864
X77 62 67 sky130_fd_pr__res_generic_po__example_5595914180864
X78 65 62 sky130_fd_pr__res_bent_po__example_5595914180862
X79 68 65 sky130_fd_pr__res_bent_po__example_5595914180862
X80 64 PULLUP_H sky130_fd_io__tk_em1s_cdns_5595914180859
X81 66 64 sky130_fd_io__tk_em1s_cdns_5595914180859
X82 67 66 sky130_fd_io__tk_em1s_cdns_5595914180859
X83 62 67 sky130_fd_io__tk_em1s_cdns_5595914180859
X84 68 28 sky130_fd_pr__res_bent_po__example_5595914180863
X85 VDDIO 71 72 73 75 76 74 sky130_fd_io__com_res_weak
X93 27 VDDIO sky130_fd_pr__res_generic_po__example_5595914180838
X100 VDDIO 49 PAD sky130_fd_pr__pfet_01v8__example_55959141808657
X101 VDDIO 49 PAD sky130_fd_pr__pfet_01v8__example_55959141808657
X128 VDDIO 27 27 45 46 47 48 49 PAD sky130_fd_pr__pfet_01v8__example_55959141808658
X129 VDDIO 27 27 45 46 47 48 49 PAD sky130_fd_pr__pfet_01v8__example_55959141808658
X130 68 65 sky130_fd_io__tk_em1o_cdns_55959141808289
X131 65 62 sky130_fd_io__tk_em1s_cdns_55959141808288
X132 VSSD VDDIO_Q 70 XRES_H_N sky130_fd_io__hvsbt_inv_x4
X133 VSSD VDDIO_Q 70 XRES_H_N sky130_fd_io__hvsbt_inv_x4
X134 VSSD VDDIO_Q 77 41 78 79 80 81 82 83 84 85 86 88 sky130_fd_io__xres2v2_rcfilter_lpfv2
X140 VSSD 41 VSSD 60 sky130_fd_pr__nfet_01v8__example_55959141808723
X141 VSSD 41 60 43 sky130_fd_pr__nfet_01v8__example_55959141808723
X148 VDDIO_Q 41 VDDIO_Q 52 sky130_fd_pr__pfet_01v8__example_55959141808720
X149 VDDIO_Q 41 52 43 sky130_fd_pr__pfet_01v8__example_55959141808720
X153 VDDIO_Q INP_SEL_H 51 88 sky130_fd_pr__pfet_01v8__example_55959141808767
X154 VDDIO_Q 39 88 FILT_IN_H sky130_fd_pr__pfet_01v8__example_55959141808767
X155 VSSIO TIE_LO_ESD sky130_fd_io__tk_tie_r_out_esd
X156 VDDIO TIE_HI_ESD sky130_fd_io__tk_tie_r_out_esd
X157 VSSD 39 51 88 sky130_fd_pr__nfet_01v8__example_55959141808764
X158 VSSD INP_SEL_H 88 FILT_IN_H sky130_fd_pr__nfet_01v8__example_55959141808764
X159 VSSD 30 61 56 sky130_fd_pr__nfet_01v8__example_55959141808779
X160 VSSD 34 57 25 sky130_fd_pr__nfet_01v8__example_55959141808779
X161 VSSD 32 31 sky130_fd_pr__nfet_01v8__example_55959141808777
X162 VSSD 37 38 sky130_fd_pr__nfet_01v8__example_55959141808777
X163 VSSD ENABLE_H 53 sky130_fd_pr__nfet_01v8__example_55959141808777
X175 VSSD 38 33 sky130_fd_pr__nfet_01v8__example_55959141808778
X176 VSSD 37 32 sky130_fd_pr__nfet_01v8__example_55959141808778
X177 24 24 24 sky130_fd_pr__pfet_01v8__example_55959141808784
X178 24 30 37 sky130_fd_pr__pfet_01v8__example_55959141808784
X179 VDDIO_Q 32 33 sky130_fd_pr__pfet_01v8__example_55959141808783
X180 VDDIO_Q 33 32 sky130_fd_pr__pfet_01v8__example_55959141808783
X183 VDDIO_Q ENABLE_H 53 sky130_fd_pr__pfet_01v8__example_55959141808786
X184 VDDIO_Q 34 54 sky130_fd_pr__pfet_01v8__example_55959141808786
X185 VDDIO_Q 35 55 sky130_fd_pr__pfet_01v8__example_55959141808786
X186 VDDIO_Q EN_VDDIO_SIG_H 56 sky130_fd_pr__pfet_01v8__example_55959141808786
X187 VCCHIB 36 57 sky130_fd_pr__pfet_01v8__example_55959141808786
X188 VCCHIB 36 58 sky130_fd_pr__pfet_01v8__example_55959141808786
X189 VDDIO_Q 34 26 sky130_fd_pr__pfet_01v8__example_55959141808786
X190 VDDIO_Q 35 54 50 sky130_fd_pr__pfet_01v8__example_55959141808787
X191 25 37 38 25 sky130_fd_pr__pfet_01v8__example_55959141808787
X192 VDDIO_Q 37 44 38 sky130_fd_pr__pfet_01v8__example_55959141808787
X193 VDDIO_Q 35 26 44 sky130_fd_pr__pfet_01v8__example_55959141808787
X194 VSSD VDDIO VSSD 30 PAD sky130_fd_io__gpio_buf_localesdv2
X195 VSSD 91 VSSIO VDDIO 91 91 87 PAD sky130_fd_io__gpio_pddrvr_strong_xres4v2
.ENDS
***************************************
.SUBCKT sky130_ef_io__vddio_hvc_clamped_pad VSSD VSSIO VDDIO 12
**
*.CALIBRE ISOLATED NETS: VCCHIB VCCD VDDA VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q
X0 VSSD VSSIO VDDIO VDDIO VDDIO 12 sky130_fd_io__top_power_hvc_wpadv2
*.CALIBRE WARNING SHORT Short circuit(s) detected by extraction in this cell. See extraction report for details.
*.CALIBRE WARNING OPEN Open circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT sky130_ef_io__vccd_lvc_clamped_pad VSSD VSSIO VCCD VDDIO 13
**
*.CALIBRE ISOLATED NETS: VCCHIB VDDA VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
X0 VSSD VSSD VSSD VCCD VDDIO VCCD VSSIO VCCD 13 sky130_fd_io__top_power_lvc_wpad
*.CALIBRE WARNING OPEN Open circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT chip_io vssd porb_h vssio vccd vddio vssa flash_io0_ieb_core flash_io0_oeb_core flash_io1_ieb_core vssa1 vdda1 mprj_io_oeb[37] mprj_io_ib_mode_sel[37] mprj_io_vtrip_sel[37] mprj_io_out[37] mprj_io_holdover[37] mprj_io_dm[113] mprj_io_analog_sel[37] mprj_io_hldh_n[37] mprj_io_enh[37]
+ mprj_io_inp_dis[37] mprj_io_analog_pol[37] mprj_io_dm[111] mprj_io_analog_en[37] mprj_io_dm[112] mprj_analog_io[30] mprj_io_slow_sel[37] mprj_io_in[37] mprj_io_oeb[36] mprj_io_ib_mode_sel[36] mprj_io_vtrip_sel[36] mprj_io_out[36] mprj_io_holdover[36] mprj_io_dm[110] mprj_io_analog_sel[36] mprj_io_hldh_n[36] mprj_io_enh[36] mprj_io_inp_dis[36] mprj_io_analog_pol[36] mprj_io_dm[108]
+ mprj_io_analog_en[36] mprj_io_dm[109] mprj_analog_io[29] mprj_io_slow_sel[36] mprj_io_in[36] mprj_io_oeb[35] mprj_io_ib_mode_sel[35] mprj_io_vtrip_sel[35] mprj_io_out[35] mprj_io_holdover[35] mprj_io_dm[107] mprj_io_analog_sel[35] mprj_io_hldh_n[35] mprj_io_enh[35] mprj_io_inp_dis[35] mprj_io_analog_pol[35] mprj_io_dm[105] mprj_io_analog_en[35] mprj_io_dm[106] mprj_analog_io[28]
+ mprj_io_slow_sel[35] mprj_io_in[35] mprj_io_oeb[34] mprj_io_ib_mode_sel[34] mprj_io_vtrip_sel[34] mprj_io_out[34] mprj_io_holdover[34] mprj_io_dm[104] mprj_io_analog_sel[34] mprj_io_hldh_n[34] mprj_io_enh[34] mprj_io_inp_dis[34] mprj_io_analog_pol[34] mprj_io_dm[102] mprj_io_analog_en[34] mprj_io_dm[103] mprj_analog_io[27] mprj_io_slow_sel[34] mprj_io_in[34] mprj_io_oeb[33]
+ mprj_io_ib_mode_sel[33] mprj_io_vtrip_sel[33] mprj_io_out[33] mprj_io_holdover[33] mprj_io_dm[101] mprj_io_analog_sel[33] mprj_io_hldh_n[33] mprj_io_enh[33] mprj_io_inp_dis[33] mprj_io_analog_pol[33] mprj_io_dm[99] mprj_io_analog_en[33] mprj_io_dm[100] mprj_analog_io[26] mprj_io_slow_sel[33] mprj_io_in[33] mprj_io_oeb[32] mprj_io_ib_mode_sel[32] mprj_io_vtrip_sel[32] mprj_io_out[32]
+ mprj_io_holdover[32] mprj_io_dm[98] mprj_io_analog_sel[32] mprj_io_hldh_n[32] mprj_io_enh[32] mprj_io_inp_dis[32] mprj_io_analog_pol[32] mprj_io_dm[96] mprj_io_analog_en[32] mprj_io_dm[97] mprj_analog_io[25] mprj_io_slow_sel[32] mprj_io_in[32] mprj_io_oeb[31] mprj_io_ib_mode_sel[31] mprj_io_vtrip_sel[31] mprj_io_out[31] mprj_io_holdover[31] mprj_io_dm[95] mprj_io_analog_sel[31]
+ mprj_io_hldh_n[31] mprj_io_enh[31] mprj_io_inp_dis[31] mprj_io_analog_pol[31] mprj_io_dm[93] mprj_io_analog_en[31] mprj_io_dm[94] mprj_analog_io[24] mprj_io_slow_sel[31] mprj_io_in[31] mprj_io_oeb[30] mprj_io_ib_mode_sel[30] mprj_io_vtrip_sel[30] mprj_io_out[30] mprj_io_holdover[30] mprj_io_dm[92] mprj_io_analog_sel[30] mprj_io_hldh_n[30] mprj_io_enh[30] mprj_io_inp_dis[30]
+ mprj_io_analog_pol[30] mprj_io_dm[90] mprj_io_analog_en[30] mprj_io_dm[91] mprj_analog_io[23] mprj_io_slow_sel[30] mprj_io_in[30] mprj_io_oeb[29] mprj_io_ib_mode_sel[29] mprj_io_vtrip_sel[29] mprj_io_out[29] mprj_io_holdover[29] mprj_io_dm[89] mprj_io_analog_sel[29] mprj_io_hldh_n[29] mprj_io_enh[29] mprj_io_inp_dis[29] mprj_io_analog_pol[29] mprj_io_dm[87] mprj_io_analog_en[29]
+ mprj_io_dm[88] mprj_analog_io[22] mprj_io_slow_sel[29] mprj_io_in[29] mprj_io_oeb[28] mprj_io_ib_mode_sel[28] mprj_io_vtrip_sel[28] mprj_io_out[28] mprj_io_holdover[28] mprj_io_dm[86] mprj_io_analog_sel[28] mprj_io_hldh_n[28] mprj_io_enh[28] mprj_io_inp_dis[28] mprj_io_analog_pol[28] mprj_io_dm[84] mprj_io_analog_en[28] mprj_io_dm[85] mprj_analog_io[21] mprj_io_slow_sel[28]
+ mprj_io_in[28] mprj_io_oeb[27] mprj_io_ib_mode_sel[27] mprj_io_vtrip_sel[27] mprj_io_out[27] mprj_io_holdover[27] mprj_io_dm[83] mprj_io_analog_sel[27] mprj_io_hldh_n[27] mprj_io_enh[27] mprj_io_inp_dis[27] mprj_io_analog_pol[27] mprj_io_dm[81] mprj_io_analog_en[27] mprj_io_dm[82] mprj_analog_io[20] mprj_io_slow_sel[27] mprj_io_in[27] mprj_io_oeb[26] mprj_io_ib_mode_sel[26]
+ mprj_io_vtrip_sel[26] mprj_io_out[26] mprj_io_holdover[26] mprj_io_dm[80] mprj_io_analog_sel[26] mprj_io_hldh_n[26] mprj_io_enh[26] mprj_io_inp_dis[26] mprj_io_analog_pol[26] mprj_io_dm[78] mprj_io_analog_en[26] mprj_io_dm[79] mprj_analog_io[19] mprj_io_slow_sel[26] mprj_io_in[26] mprj_io_oeb[25] mprj_io_ib_mode_sel[25] mprj_io_vtrip_sel[25] mprj_io_out[25] mprj_io_holdover[25]
+ mprj_io_dm[77] mprj_io_analog_sel[25] mprj_io_hldh_n[25] mprj_io_enh[25] mprj_io_inp_dis[25] mprj_io_analog_pol[25] mprj_io_dm[75] mprj_io_analog_en[25] mprj_io_dm[76] mprj_analog_io[18] mprj_io_slow_sel[25] mprj_io_in[25] mprj_io_oeb[24] mprj_io_ib_mode_sel[24] mprj_io_vtrip_sel[24] mprj_io_out[24] mprj_io_holdover[24] mprj_io_dm[74] mprj_io_analog_sel[24] mprj_io_hldh_n[24]
+ mprj_io_enh[24] mprj_io_inp_dis[24] mprj_io_analog_pol[24] mprj_io_dm[72] mprj_io_analog_en[24] mprj_io_dm[73] mprj_analog_io[17] mprj_io_slow_sel[24] mprj_io_in[24] mprj_io_oeb[23] mprj_io_ib_mode_sel[23] mprj_io_vtrip_sel[23] mprj_io_out[23] mprj_io_holdover[23] mprj_io_dm[71] mprj_io_analog_sel[23] mprj_io_hldh_n[23] mprj_io_enh[23] mprj_io_inp_dis[23] mprj_io_analog_pol[23]
+ mprj_io_dm[69] mprj_io_analog_en[23] mprj_io_dm[70] mprj_analog_io[16] mprj_io_slow_sel[23] mprj_io_in[23] mprj_io_oeb[22] mprj_io_ib_mode_sel[22] mprj_io_vtrip_sel[22] mprj_io_out[22] mprj_io_holdover[22] mprj_io_dm[68] mprj_io_analog_sel[22] mprj_io_hldh_n[22] mprj_io_enh[22] mprj_io_inp_dis[22] mprj_io_analog_pol[22] mprj_io_dm[66] mprj_io_analog_en[22] mprj_io_dm[67]
+ mprj_analog_io[15] mprj_io_slow_sel[22] resetb_core_h mprj_io_in[22] mprj_io_oeb[21] mprj_io_ib_mode_sel[21] mprj_io_vtrip_sel[21] mprj_io_out[21] mprj_io_holdover[21] mprj_io_dm[65] mprj_io_analog_sel[21] mprj_io_hldh_n[21] mprj_io_enh[21] mprj_io_inp_dis[21] clock_core mprj_io_analog_pol[21] mprj_io_dm[63] mprj_io_analog_en[21] mprj_io_dm[64] mprj_analog_io[14]
+ mprj_io_slow_sel[21] mprj_io_in[21] por mprj_io_oeb[20] mprj_io_ib_mode_sel[20] mprj_io_vtrip_sel[20] mprj_io_out[20] mprj_io_holdover[20] mprj_io_dm[62] mprj_io_analog_sel[20] mprj_io_hldh_n[20] mprj_io_enh[20] mprj_io_inp_dis[20] mprj_io_analog_pol[20] mprj_io_dm[60] mprj_io_analog_en[20] mprj_io_dm[61] mprj_analog_io[13] mprj_io_slow_sel[20] mprj_io_in[20]
+ mprj_io_oeb[19] mprj_io_ib_mode_sel[19] mprj_io_vtrip_sel[19] mprj_io_out[19] mprj_io_holdover[19] mprj_io_dm[59] mprj_io_analog_sel[19] mprj_io_hldh_n[19] mprj_io_enh[19] mprj_io_inp_dis[19] mprj_io_analog_pol[19] mprj_io_dm[57] mprj_io_analog_en[19] mprj_io_dm[58] mprj_analog_io[12] mprj_io_slow_sel[19] mprj_io_in[19] flash_csb_ieb_core flash_csb_core flash_csb_oeb_core
+ flash_clk_ieb_core flash_clk_core flash_clk_oeb_core mprj_io_oeb[18] mprj_io_ib_mode_sel[18] mprj_io_vtrip_sel[18] mprj_io_out[18] mprj_io_holdover[18] mprj_io_dm[56] mprj_io_analog_sel[18] mprj_io_hldh_n[18] mprj_io_enh[18] mprj_io_inp_dis[18] mprj_io_analog_pol[18] mprj_io_dm[54] mprj_io_analog_en[18] mprj_io_dm[55] mprj_analog_io[11] mprj_io_slow_sel[18] mprj_io_in[18]
+ flash_io0_di_core flash_io0_do_core flash_io1_di_core flash_io1_oeb_core flash_io1_do_core mprj_io_oeb[17] mprj_io_ib_mode_sel[17] mprj_io_vtrip_sel[17] mprj_io_out[17] mprj_io_holdover[17] mprj_io_dm[53] mprj_io_analog_sel[17] mprj_io_hldh_n[17] mprj_io_enh[17] mprj_io_inp_dis[17] mprj_io_analog_pol[17] mprj_io_dm[51] mprj_io_analog_en[17] mprj_io_dm[52] mprj_analog_io[10]
+ mprj_io_slow_sel[17] mprj_io_in[17] gpio_in_core gpio_mode1_core gpio_mode0_core gpio_inenb_core mprj_io_oeb[16] mprj_io_ib_mode_sel[16] gpio_out_core mprj_io_vtrip_sel[16] mprj_io_out[16] mprj_io_holdover[16] gpio_outenb_core mprj_io_dm[50] mprj_io_analog_sel[16] mprj_io_hldh_n[16] mprj_io_enh[16] mprj_io_inp_dis[16] mprj_io_analog_pol[16] mprj_io_dm[48]
+ mprj_io_analog_en[16] mprj_io_dm[49] mprj_analog_io[9] mprj_io_slow_sel[16] mprj_io_in[16] mprj_io_oeb[15] mprj_io_ib_mode_sel[15] mprj_io_vtrip_sel[15] mprj_io_out[15] mprj_io_holdover[15] mprj_io_dm[47] mprj_io_analog_sel[15] mprj_io_hldh_n[15] mprj_io_enh[15] mprj_io_inp_dis[15] mprj_io_analog_pol[15] mprj_io_dm[45] mprj_io_analog_en[15] mprj_io_dm[46] mprj_analog_io[8]
+ mprj_io_slow_sel[15] mprj_io_in[15] mprj_io_in[0] mprj_io_slow_sel[0] mprj_io_dm[1] mprj_io_analog_en[0] mprj_io_dm[0] mprj_io_analog_pol[0] mprj_io_inp_dis[0] mprj_io_enh[0] mprj_io_hldh_n[0] mprj_io_analog_sel[0] mprj_io_dm[2] mprj_io_holdover[0] mprj_io_out[0] mprj_io_vtrip_sel[0] mprj_io_ib_mode_sel[0] mprj_io_oeb[0] mprj_io_in[1] mprj_io_slow_sel[1]
+ mprj_io_dm[4] mprj_io_analog_en[1] mprj_io_dm[3] mprj_io_analog_pol[1] mprj_io_inp_dis[1] mprj_io_enh[1] mprj_io_hldh_n[1] mprj_io_analog_sel[1] mprj_io_dm[5] mprj_io_holdover[1] mprj_io_out[1] mprj_io_vtrip_sel[1] mprj_io_ib_mode_sel[1] mprj_io_oeb[1] mprj_io_in[2] mprj_io_slow_sel[2] mprj_io_dm[7] mprj_io_analog_en[2] mprj_io_dm[6] mprj_io_analog_pol[2]
+ mprj_io_inp_dis[2] mprj_io_enh[2] mprj_io_hldh_n[2] mprj_io_analog_sel[2] mprj_io_dm[8] mprj_io_holdover[2] mprj_io_out[2] mprj_io_vtrip_sel[2] mprj_io_ib_mode_sel[2] mprj_io_oeb[2] mprj_io_in[3] mprj_io_slow_sel[3] mprj_io_dm[10] mprj_io_analog_en[3] mprj_io_dm[9] mprj_io_analog_pol[3] mprj_io_inp_dis[3] mprj_io_enh[3] mprj_io_hldh_n[3] mprj_io_analog_sel[3]
+ mprj_io_dm[11] mprj_io_holdover[3] mprj_io_out[3] mprj_io_vtrip_sel[3] mprj_io_ib_mode_sel[3] mprj_io_oeb[3] mprj_io_in[4] mprj_io_slow_sel[4] mprj_io_dm[13] mprj_io_analog_en[4] mprj_io_dm[12] mprj_io_analog_pol[4] mprj_io_inp_dis[4] mprj_io_enh[4] mprj_io_hldh_n[4] mprj_io_analog_sel[4] mprj_io_dm[14] mprj_io_holdover[4] mprj_io_out[4] mprj_io_vtrip_sel[4]
+ mprj_io_ib_mode_sel[4] mprj_io_oeb[4] mprj_io_in[5] mprj_io_slow_sel[5] mprj_io_dm[16] mprj_io_analog_en[5] mprj_io_dm[15] mprj_io_analog_pol[5] mprj_io_inp_dis[5] mprj_io_enh[5] mprj_io_hldh_n[5] mprj_io_analog_sel[5] mprj_io_dm[17] mprj_io_holdover[5] mprj_io_out[5] mprj_io_vtrip_sel[5] mprj_io_ib_mode_sel[5] mprj_io_oeb[5] mprj_io_in[6] mprj_io_slow_sel[6]
+ mprj_io_dm[19] mprj_io_analog_en[6] mprj_io_dm[18] mprj_io_analog_pol[6] mprj_io_inp_dis[6] mprj_io_enh[6] mprj_io_hldh_n[6] mprj_io_analog_sel[6] mprj_io_dm[20] mprj_io_holdover[6] mprj_io_out[6] mprj_io_vtrip_sel[6] mprj_io_ib_mode_sel[6] mprj_io_oeb[6] mprj_io_in[7] mprj_io_slow_sel[7] mprj_analog_io[0] mprj_io_dm[22] mprj_io_analog_en[7] mprj_io_dm[21]
+ mprj_io_analog_pol[7] mprj_io_inp_dis[7] mprj_io_enh[7] mprj_io_hldh_n[7] mprj_io_analog_sel[7] mprj_io_dm[23] mprj_io_holdover[7] mprj_io_out[7] mprj_io_vtrip_sel[7] mprj_io_ib_mode_sel[7] mprj_io_oeb[7] mprj_io_in[8] mprj_io_slow_sel[8] mprj_analog_io[1] mprj_io_dm[25] mprj_io_analog_en[8] mprj_io_dm[24] mprj_io_analog_pol[8] mprj_io_inp_dis[8] mprj_io_enh[8]
+ mprj_io_hldh_n[8] mprj_io_analog_sel[8] mprj_io_dm[26] mprj_io_holdover[8] mprj_io_out[8] mprj_io_vtrip_sel[8] mprj_io_ib_mode_sel[8] mprj_io_oeb[8] mprj_io_in[9] mprj_io_slow_sel[9] mprj_analog_io[2] mprj_io_dm[28] mprj_io_analog_en[9] mprj_io_dm[27] mprj_io_analog_pol[9] mprj_io_inp_dis[9] mprj_io_enh[9] mprj_io_hldh_n[9] mprj_io_analog_sel[9] mprj_io_dm[29]
+ mprj_io_holdover[9] mprj_io_out[9] mprj_io_vtrip_sel[9] mprj_io_ib_mode_sel[9] mprj_io_oeb[9] mprj_io_in[10] mprj_io_slow_sel[10] mprj_analog_io[3] mprj_io_dm[31] mprj_io_analog_en[10] mprj_io_dm[30] mprj_io_analog_pol[10] mprj_io_inp_dis[10] mprj_io_enh[10] mprj_io_hldh_n[10] mprj_io_analog_sel[10] mprj_io_dm[32] mprj_io_holdover[10] mprj_io_out[10] mprj_io_vtrip_sel[10]
+ mprj_io_ib_mode_sel[10] mprj_io_oeb[10] mprj_io_in[11] mprj_io_slow_sel[11] mprj_analog_io[4] mprj_io_dm[34] mprj_io_analog_en[11] mprj_io_dm[33] mprj_io_analog_pol[11] mprj_io_inp_dis[11] mprj_io_enh[11] mprj_io_hldh_n[11] mprj_io_analog_sel[11] mprj_io_dm[35] mprj_io_holdover[11] mprj_io_out[11] mprj_io_vtrip_sel[11] mprj_io_ib_mode_sel[11] mprj_io_oeb[11] mprj_io_in[12]
+ mprj_io_slow_sel[12] mprj_analog_io[5] mprj_io_dm[37] mprj_io_analog_en[12] mprj_io_dm[36] mprj_io_analog_pol[12] mprj_io_inp_dis[12] mprj_io_enh[12] mprj_io_hldh_n[12] mprj_io_analog_sel[12] mprj_io_dm[38] mprj_io_holdover[12] mprj_io_out[12] mprj_io_vtrip_sel[12] mprj_io_ib_mode_sel[12] mprj_io_oeb[12] mprj_io_in[13] mprj_io_slow_sel[13] mprj_analog_io[6] mprj_io_dm[40]
+ mprj_io_analog_en[13] mprj_io_dm[39] mprj_io_analog_pol[13] mprj_io_inp_dis[13] mprj_io_enh[13] mprj_io_hldh_n[13] mprj_io_analog_sel[13] mprj_io_dm[41] mprj_io_holdover[13] mprj_io_out[13] mprj_io_vtrip_sel[13] mprj_io_ib_mode_sel[13] mprj_io_oeb[13] mprj_io_in[14] mprj_io_slow_sel[14] mprj_analog_io[7] mprj_io_dm[43] mprj_io_analog_en[14] mprj_io_dm[42] mprj_io_analog_pol[14]
+ mprj_io_inp_dis[14] mprj_io_enh[14] mprj_io_hldh_n[14] mprj_io_analog_sel[14] mprj_io_dm[44] mprj_io_holdover[14] mprj_io_out[14] mprj_io_vtrip_sel[14] mprj_io_ib_mode_sel[14] mprj_io_oeb[14] vssa2 vdda2 vccd2 vdda vccd1 738 vssd2 740 mprj_io[37] mprj_io[36]
+ mprj_io[35] mprj_io[34] mprj_io[33] mprj_io[32] mprj_io[31] mprj_io[30] mprj_io[29] mprj_io[28] mprj_io[27] mprj_io[26] mprj_io[25] mprj_io[24] 755 756 757 mprj_io[23] 759 mprj_io[22] resetb mprj_io[21]
+ clock mprj_io[20] 765 mprj_io[19] flash_csb 768 flash_clk mprj_io[18] flash_io0 flash_io1 mprj_io[17] gpio mprj_io[16] 776 777 778 mprj_io[15] vssd1 781 mprj_io[0]
+ mprj_io[1] mprj_io[2] mprj_io[3] mprj_io[4] mprj_io[5] mprj_io[6] mprj_io[7] mprj_io[8] mprj_io[9] mprj_io[10] mprj_io[11] mprj_io[12] mprj_io[13] mprj_io[14] 797
**
X0 vssd vssa2 vddio vdda2 756 sky130_ef_io__vdda_hvc_clamped_pad
X1 vssd vssa vddio vdda 778 sky130_ef_io__vdda_hvc_clamped_pad
X2 vssd vssa1 vddio vdda1 798 sky130_ef_io__vdda_hvc_clamped_pad
X3 vssd vssa1 vddio vdda1 797 sky130_ef_io__vdda_hvc_clamped_pad
X4 vssd vddio vssa2 vdda2 757 sky130_ef_io__vssa_hvc_clamped_pad
X5 vssd vddio vssa vdda 759 sky130_ef_io__vssa_hvc_clamped_pad
X6 vssd vddio vssa1 vdda1 777 sky130_ef_io__vssa_hvc_clamped_pad
X7 vssd vddio vssa1 vdda1 799 sky130_ef_io__vssa_hvc_clamped_pad
X8 vssd vssa2 vssio vccd2 vddio 740 sky130_ef_io__vccd_lvc_clamped2_pad
X9 vssd vssa1 vssio vccd1 vddio 781 sky130_ef_io__vccd_lvc_clamped2_pad
X10 vssd vssa2 vssio vccd2 vddio vssd2 sky130_ef_io__vssd_lvc_clamped2_pad
X11 vssd vssa1 vssio vccd1 vddio vssd1 sky130_ef_io__vssd_lvc_clamped2_pad
X12 vssd vssa2 vssio vssio vddio vddio mprj_io[37] mprj_analog_io[30] mprj_io_ib_mode_sel[37] 3 mprj_io_enh[37] vdda2 vccd2 mprj_io_oeb[37] porb_h mprj_io_vtrip_sel[37] vccd vssio mprj_io_out[37] mprj_io_holdover[37]
+ mprj_io_dm[113] mprj_io_analog_sel[37] mprj_io_hldh_n[37] mprj_io_analog_en[37] mprj_io_inp_dis[37] mprj_io_analog_pol[37] mprj_io_dm[111] mprj_io_dm[112] mprj_io_slow_sel[37] mprj_io_in[37] vccd 3 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X13 vssd vssa2 vssio vssio vddio vddio mprj_io[36] mprj_analog_io[29] mprj_io_ib_mode_sel[36] 4 mprj_io_enh[36] vdda2 vccd2 mprj_io_oeb[36] porb_h mprj_io_vtrip_sel[36] vccd vssio mprj_io_out[36] mprj_io_holdover[36]
+ mprj_io_dm[110] mprj_io_analog_sel[36] mprj_io_hldh_n[36] mprj_io_analog_en[36] mprj_io_inp_dis[36] mprj_io_analog_pol[36] mprj_io_dm[108] mprj_io_dm[109] mprj_io_slow_sel[36] mprj_io_in[36] vccd 4 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X14 vssd vssa2 vssio vssio vddio vddio mprj_io[35] mprj_analog_io[28] mprj_io_ib_mode_sel[35] 5 mprj_io_enh[35] vdda2 vccd2 mprj_io_oeb[35] porb_h mprj_io_vtrip_sel[35] vccd vssio mprj_io_out[35] mprj_io_holdover[35]
+ mprj_io_dm[107] mprj_io_analog_sel[35] mprj_io_hldh_n[35] mprj_io_analog_en[35] mprj_io_inp_dis[35] mprj_io_analog_pol[35] mprj_io_dm[105] mprj_io_dm[106] mprj_io_slow_sel[35] mprj_io_in[35] vccd 5 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X15 vssd vssa2 vssio vssio vddio vddio mprj_io[34] mprj_analog_io[27] mprj_io_ib_mode_sel[34] 6 mprj_io_enh[34] vdda2 vccd2 mprj_io_oeb[34] porb_h mprj_io_vtrip_sel[34] vccd vssio mprj_io_out[34] mprj_io_holdover[34]
+ mprj_io_dm[104] mprj_io_analog_sel[34] mprj_io_hldh_n[34] mprj_io_analog_en[34] mprj_io_inp_dis[34] mprj_io_analog_pol[34] mprj_io_dm[102] mprj_io_dm[103] mprj_io_slow_sel[34] mprj_io_in[34] vccd 6 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X16 vssd vssa2 vssio vssio vddio vddio mprj_io[33] mprj_analog_io[26] mprj_io_ib_mode_sel[33] 7 mprj_io_enh[33] vdda2 vccd2 mprj_io_oeb[33] porb_h mprj_io_vtrip_sel[33] vccd vssio mprj_io_out[33] mprj_io_holdover[33]
+ mprj_io_dm[101] mprj_io_analog_sel[33] mprj_io_hldh_n[33] mprj_io_analog_en[33] mprj_io_inp_dis[33] mprj_io_analog_pol[33] mprj_io_dm[99] mprj_io_dm[100] mprj_io_slow_sel[33] mprj_io_in[33] vccd 7 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X17 vssd vssa2 vssio vssio vddio vddio mprj_io[32] mprj_analog_io[25] mprj_io_ib_mode_sel[32] 8 mprj_io_enh[32] vdda2 vccd2 mprj_io_oeb[32] porb_h mprj_io_vtrip_sel[32] vccd vssio mprj_io_out[32] mprj_io_holdover[32]
+ mprj_io_dm[98] mprj_io_analog_sel[32] mprj_io_hldh_n[32] mprj_io_analog_en[32] mprj_io_inp_dis[32] mprj_io_analog_pol[32] mprj_io_dm[96] mprj_io_dm[97] mprj_io_slow_sel[32] mprj_io_in[32] vccd 8 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X18 vssd vssa2 vssio vssio vddio vddio mprj_io[31] mprj_analog_io[24] mprj_io_ib_mode_sel[31] 9 mprj_io_enh[31] vdda2 vccd2 mprj_io_oeb[31] porb_h mprj_io_vtrip_sel[31] vccd vssio mprj_io_out[31] mprj_io_holdover[31]
+ mprj_io_dm[95] mprj_io_analog_sel[31] mprj_io_hldh_n[31] mprj_io_analog_en[31] mprj_io_inp_dis[31] mprj_io_analog_pol[31] mprj_io_dm[93] mprj_io_dm[94] mprj_io_slow_sel[31] mprj_io_in[31] vccd 9 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X19 vssd vssa2 vssio vssio vddio vddio mprj_io[30] mprj_analog_io[23] mprj_io_ib_mode_sel[30] 10 mprj_io_enh[30] vdda2 vccd2 mprj_io_oeb[30] porb_h mprj_io_vtrip_sel[30] vccd vssio mprj_io_out[30] mprj_io_holdover[30]
+ mprj_io_dm[92] mprj_io_analog_sel[30] mprj_io_hldh_n[30] mprj_io_analog_en[30] mprj_io_inp_dis[30] mprj_io_analog_pol[30] mprj_io_dm[90] mprj_io_dm[91] mprj_io_slow_sel[30] mprj_io_in[30] vccd 10 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X20 vssd vssa2 vssio vssio vddio vddio mprj_io[29] mprj_analog_io[22] mprj_io_ib_mode_sel[29] 11 mprj_io_enh[29] vdda2 vccd2 mprj_io_oeb[29] porb_h mprj_io_vtrip_sel[29] vccd vssio mprj_io_out[29] mprj_io_holdover[29]
+ mprj_io_dm[89] mprj_io_analog_sel[29] mprj_io_hldh_n[29] mprj_io_analog_en[29] mprj_io_inp_dis[29] mprj_io_analog_pol[29] mprj_io_dm[87] mprj_io_dm[88] mprj_io_slow_sel[29] mprj_io_in[29] vccd 11 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X21 vssd vssa2 vssio vssio vddio vddio mprj_io[28] mprj_analog_io[21] mprj_io_ib_mode_sel[28] 12 mprj_io_enh[28] vdda2 vccd2 mprj_io_oeb[28] porb_h mprj_io_vtrip_sel[28] vccd vssio mprj_io_out[28] mprj_io_holdover[28]
+ mprj_io_dm[86] mprj_io_analog_sel[28] mprj_io_hldh_n[28] mprj_io_analog_en[28] mprj_io_inp_dis[28] mprj_io_analog_pol[28] mprj_io_dm[84] mprj_io_dm[85] mprj_io_slow_sel[28] mprj_io_in[28] vccd 12 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X22 vssd vssa2 vssio vssio vddio vddio mprj_io[27] mprj_analog_io[20] mprj_io_ib_mode_sel[27] 13 mprj_io_enh[27] vdda2 vccd2 mprj_io_oeb[27] porb_h mprj_io_vtrip_sel[27] vccd vssio mprj_io_out[27] mprj_io_holdover[27]
+ mprj_io_dm[83] mprj_io_analog_sel[27] mprj_io_hldh_n[27] mprj_io_analog_en[27] mprj_io_inp_dis[27] mprj_io_analog_pol[27] mprj_io_dm[81] mprj_io_dm[82] mprj_io_slow_sel[27] mprj_io_in[27] vccd 13 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X23 vssd vssa2 vssio vssio vddio vddio mprj_io[26] mprj_analog_io[19] mprj_io_ib_mode_sel[26] 14 mprj_io_enh[26] vdda2 vccd2 mprj_io_oeb[26] porb_h mprj_io_vtrip_sel[26] vccd vssio mprj_io_out[26] mprj_io_holdover[26]
+ mprj_io_dm[80] mprj_io_analog_sel[26] mprj_io_hldh_n[26] mprj_io_analog_en[26] mprj_io_inp_dis[26] mprj_io_analog_pol[26] mprj_io_dm[78] mprj_io_dm[79] mprj_io_slow_sel[26] mprj_io_in[26] vccd 14 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X24 vssd vssa2 vssio vssio vddio vddio mprj_io[25] mprj_analog_io[18] mprj_io_ib_mode_sel[25] 15 mprj_io_enh[25] vdda2 vccd2 mprj_io_oeb[25] porb_h mprj_io_vtrip_sel[25] vccd vssio mprj_io_out[25] mprj_io_holdover[25]
+ mprj_io_dm[77] mprj_io_analog_sel[25] mprj_io_hldh_n[25] mprj_io_analog_en[25] mprj_io_inp_dis[25] mprj_io_analog_pol[25] mprj_io_dm[75] mprj_io_dm[76] mprj_io_slow_sel[25] mprj_io_in[25] vccd 15 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X25 vssd vssa2 vssio vssio vddio vddio mprj_io[24] mprj_analog_io[17] mprj_io_ib_mode_sel[24] 18 mprj_io_enh[24] vdda2 vccd2 mprj_io_oeb[24] porb_h mprj_io_vtrip_sel[24] vccd vssio mprj_io_out[24] mprj_io_holdover[24]
+ mprj_io_dm[74] mprj_io_analog_sel[24] mprj_io_hldh_n[24] mprj_io_analog_en[24] mprj_io_inp_dis[24] mprj_io_analog_pol[24] mprj_io_dm[72] mprj_io_dm[73] mprj_io_slow_sel[24] mprj_io_in[24] vccd 18 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X26 vssd vssa2 vssio vssio vddio vddio mprj_io[23] mprj_analog_io[16] mprj_io_ib_mode_sel[23] 20 mprj_io_enh[23] vdda2 vccd2 mprj_io_oeb[23] porb_h mprj_io_vtrip_sel[23] vccd vssio mprj_io_out[23] mprj_io_holdover[23]
+ mprj_io_dm[71] mprj_io_analog_sel[23] mprj_io_hldh_n[23] mprj_io_analog_en[23] mprj_io_inp_dis[23] mprj_io_analog_pol[23] mprj_io_dm[69] mprj_io_dm[70] mprj_io_slow_sel[23] mprj_io_in[23] vccd 20 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X27 vssd vssa2 vssio vssio vddio vddio mprj_io[22] mprj_analog_io[15] mprj_io_ib_mode_sel[22] 22 mprj_io_enh[22] vdda2 vccd2 mprj_io_oeb[22] porb_h mprj_io_vtrip_sel[22] vccd vssio mprj_io_out[22] mprj_io_holdover[22]
+ mprj_io_dm[68] mprj_io_analog_sel[22] mprj_io_hldh_n[22] mprj_io_analog_en[22] mprj_io_inp_dis[22] mprj_io_analog_pol[22] mprj_io_dm[66] mprj_io_dm[67] mprj_io_slow_sel[22] mprj_io_in[22] vccd 22 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X28 vssd vssa2 vssio vssio vddio vddio mprj_io[21] mprj_analog_io[14] mprj_io_ib_mode_sel[21] 25 mprj_io_enh[21] vdda2 vccd2 mprj_io_oeb[21] porb_h mprj_io_vtrip_sel[21] vccd vssio mprj_io_out[21] mprj_io_holdover[21]
+ mprj_io_dm[65] mprj_io_analog_sel[21] mprj_io_hldh_n[21] mprj_io_analog_en[21] mprj_io_inp_dis[21] mprj_io_analog_pol[21] mprj_io_dm[63] mprj_io_dm[64] mprj_io_slow_sel[21] mprj_io_in[21] vccd 25 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X29 vssd vssa vssio vssio vddio vddio clock 716 vssd 24 porb_h vdda vccd vccd porb_h vssd vccd vssa vssd vssd
+ vssd vssd vddio vssd por vssd vccd vssd vssd clock_core vccd 24 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X30 vssd vssa2 vssio vssio vddio vddio mprj_io[20] mprj_analog_io[13] mprj_io_ib_mode_sel[20] 26 mprj_io_enh[20] vdda2 vccd2 mprj_io_oeb[20] porb_h mprj_io_vtrip_sel[20] vccd vssio mprj_io_out[20] mprj_io_holdover[20]
+ mprj_io_dm[62] mprj_io_analog_sel[20] mprj_io_hldh_n[20] mprj_io_analog_en[20] mprj_io_inp_dis[20] mprj_io_analog_pol[20] mprj_io_dm[60] mprj_io_dm[61] mprj_io_slow_sel[20] mprj_io_in[20] vccd 26 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X31 vssd vssa2 vssio vssio vddio vddio mprj_io[19] mprj_analog_io[12] mprj_io_ib_mode_sel[19] 27 mprj_io_enh[19] vdda2 vccd2 mprj_io_oeb[19] porb_h mprj_io_vtrip_sel[19] vccd vssio mprj_io_out[19] mprj_io_holdover[19]
+ mprj_io_dm[59] mprj_io_analog_sel[19] mprj_io_hldh_n[19] mprj_io_analog_en[19] mprj_io_inp_dis[19] mprj_io_analog_pol[19] mprj_io_dm[57] mprj_io_dm[58] mprj_io_slow_sel[19] mprj_io_in[19] vccd 27 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X32 vssd vssa vssio vssio vddio vddio flash_csb 717 vssd 28 porb_h vdda vccd flash_csb_oeb_core porb_h vssd vccd vssa flash_csb_core vssd
+ vccd vssd vddio vssd flash_csb_ieb_core vssd vssd vccd vssd 718 vccd 28 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X33 vssd vssa vssio vssio vddio vddio flash_clk 719 vssd 29 porb_h vdda vccd flash_clk_oeb_core porb_h vssd vccd vssa flash_clk_core vssd
+ vccd vssd vddio vssd flash_clk_ieb_core vssd vssd vccd vssd 720 vccd 29 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X34 vssd vssa2 vssio vssio vddio vddio mprj_io[18] mprj_analog_io[11] mprj_io_ib_mode_sel[18] 30 mprj_io_enh[18] vdda2 vccd2 mprj_io_oeb[18] porb_h mprj_io_vtrip_sel[18] vccd vssio mprj_io_out[18] mprj_io_holdover[18]
+ mprj_io_dm[56] mprj_io_analog_sel[18] mprj_io_hldh_n[18] mprj_io_analog_en[18] mprj_io_inp_dis[18] mprj_io_analog_pol[18] mprj_io_dm[54] mprj_io_dm[55] mprj_io_slow_sel[18] mprj_io_in[18] vccd 30 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X35 vssd vssa vssio vssio vddio vddio flash_io0 721 vssd 31 porb_h vdda vccd flash_io0_oeb_core porb_h vssd vccd vssa flash_io0_do_core vssd
+ flash_io0_ieb_core vssd vddio vssd flash_io0_ieb_core vssd flash_io0_oeb_core flash_io0_ieb_core vssd flash_io0_di_core vccd 31 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X36 vssd vssa vssio vssio vddio vddio flash_io1 722 vssd 34 porb_h vdda vccd flash_io1_oeb_core porb_h vssd vccd vssa flash_io1_do_core vssd
+ flash_io1_ieb_core vssd vddio vssd flash_io1_ieb_core vssd flash_io1_oeb_core flash_io1_ieb_core vssd flash_io1_di_core vccd 34 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X37 vssd vssa1 vssio vssio vddio vddio mprj_io[17] mprj_analog_io[10] mprj_io_ib_mode_sel[17] 36 mprj_io_enh[17] vdda1 vccd1 mprj_io_oeb[17] porb_h mprj_io_vtrip_sel[17] vccd vssio mprj_io_out[17] mprj_io_holdover[17]
+ mprj_io_dm[53] mprj_io_analog_sel[17] mprj_io_hldh_n[17] mprj_io_analog_en[17] mprj_io_inp_dis[17] mprj_io_analog_pol[17] mprj_io_dm[51] mprj_io_dm[52] mprj_io_slow_sel[17] mprj_io_in[17] vccd 36 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X38 vssd vssa vssio vssio vddio vddio gpio 723 vssd 37 porb_h vdda vccd gpio_outenb_core porb_h vssd vccd vssa gpio_out_core vssd
+ gpio_mode1_core vssd vddio vssd gpio_inenb_core vssd gpio_mode0_core gpio_mode1_core vssd gpio_in_core vccd 37 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X39 vssd vssa1 vssio vssio vddio vddio mprj_io[16] mprj_analog_io[9] mprj_io_ib_mode_sel[16] 38 mprj_io_enh[16] vdda1 vccd1 mprj_io_oeb[16] porb_h mprj_io_vtrip_sel[16] vccd vssio mprj_io_out[16] mprj_io_holdover[16]
+ mprj_io_dm[50] mprj_io_analog_sel[16] mprj_io_hldh_n[16] mprj_io_analog_en[16] mprj_io_inp_dis[16] mprj_io_analog_pol[16] mprj_io_dm[48] mprj_io_dm[49] mprj_io_slow_sel[16] mprj_io_in[16] vccd 38 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X40 vssd vssa1 vssio vssio vddio vddio mprj_io[15] mprj_analog_io[8] mprj_io_ib_mode_sel[15] 39 mprj_io_enh[15] vdda1 vccd1 mprj_io_oeb[15] porb_h mprj_io_vtrip_sel[15] vccd vssio mprj_io_out[15] mprj_io_holdover[15]
+ mprj_io_dm[47] mprj_io_analog_sel[15] mprj_io_hldh_n[15] mprj_io_analog_en[15] mprj_io_inp_dis[15] mprj_io_analog_pol[15] mprj_io_dm[45] mprj_io_dm[46] mprj_io_slow_sel[15] mprj_io_in[15] vccd 39 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X41 vssd vssa1 vssio vssio vddio vddio mprj_io[0] 724 mprj_io_ib_mode_sel[0] 457 mprj_io_enh[0] vdda1 vccd1 mprj_io_oeb[0] porb_h mprj_io_vtrip_sel[0] vccd vssio mprj_io_out[0] mprj_io_holdover[0]
+ mprj_io_dm[2] mprj_io_analog_sel[0] mprj_io_hldh_n[0] mprj_io_analog_en[0] mprj_io_inp_dis[0] mprj_io_analog_pol[0] mprj_io_dm[0] mprj_io_dm[1] mprj_io_slow_sel[0] mprj_io_in[0] vccd 457 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X42 vssd vssa1 vssio vssio vddio vddio mprj_io[1] 725 mprj_io_ib_mode_sel[1] 458 mprj_io_enh[1] vdda1 vccd1 mprj_io_oeb[1] porb_h mprj_io_vtrip_sel[1] vccd vssio mprj_io_out[1] mprj_io_holdover[1]
+ mprj_io_dm[5] mprj_io_analog_sel[1] mprj_io_hldh_n[1] mprj_io_analog_en[1] mprj_io_inp_dis[1] mprj_io_analog_pol[1] mprj_io_dm[3] mprj_io_dm[4] mprj_io_slow_sel[1] mprj_io_in[1] vccd 458 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X43 vssd vssa1 vssio vssio vddio vddio mprj_io[2] 726 mprj_io_ib_mode_sel[2] 463 mprj_io_enh[2] vdda1 vccd1 mprj_io_oeb[2] porb_h mprj_io_vtrip_sel[2] vccd vssio mprj_io_out[2] mprj_io_holdover[2]
+ mprj_io_dm[8] mprj_io_analog_sel[2] mprj_io_hldh_n[2] mprj_io_analog_en[2] mprj_io_inp_dis[2] mprj_io_analog_pol[2] mprj_io_dm[6] mprj_io_dm[7] mprj_io_slow_sel[2] mprj_io_in[2] vccd 463 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X44 vssd vssa1 vssio vssio vddio vddio mprj_io[3] 727 mprj_io_ib_mode_sel[3] 459 mprj_io_enh[3] vdda1 vccd1 mprj_io_oeb[3] porb_h mprj_io_vtrip_sel[3] vccd vssio mprj_io_out[3] mprj_io_holdover[3]
+ mprj_io_dm[11] mprj_io_analog_sel[3] mprj_io_hldh_n[3] mprj_io_analog_en[3] mprj_io_inp_dis[3] mprj_io_analog_pol[3] mprj_io_dm[9] mprj_io_dm[10] mprj_io_slow_sel[3] mprj_io_in[3] vccd 459 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X45 vssd vssa1 vssio vssio vddio vddio mprj_io[4] 728 mprj_io_ib_mode_sel[4] 460 mprj_io_enh[4] vdda1 vccd1 mprj_io_oeb[4] porb_h mprj_io_vtrip_sel[4] vccd vssio mprj_io_out[4] mprj_io_holdover[4]
+ mprj_io_dm[14] mprj_io_analog_sel[4] mprj_io_hldh_n[4] mprj_io_analog_en[4] mprj_io_inp_dis[4] mprj_io_analog_pol[4] mprj_io_dm[12] mprj_io_dm[13] mprj_io_slow_sel[4] mprj_io_in[4] vccd 460 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X46 vssd vssa1 vssio vssio vddio vddio mprj_io[5] 729 mprj_io_ib_mode_sel[5] 461 mprj_io_enh[5] vdda1 vccd1 mprj_io_oeb[5] porb_h mprj_io_vtrip_sel[5] vccd vssio mprj_io_out[5] mprj_io_holdover[5]
+ mprj_io_dm[17] mprj_io_analog_sel[5] mprj_io_hldh_n[5] mprj_io_analog_en[5] mprj_io_inp_dis[5] mprj_io_analog_pol[5] mprj_io_dm[15] mprj_io_dm[16] mprj_io_slow_sel[5] mprj_io_in[5] vccd 461 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X47 vssd vssa1 vssio vssio vddio vddio mprj_io[6] 730 mprj_io_ib_mode_sel[6] 462 mprj_io_enh[6] vdda1 vccd1 mprj_io_oeb[6] porb_h mprj_io_vtrip_sel[6] vccd vssio mprj_io_out[6] mprj_io_holdover[6]
+ mprj_io_dm[20] mprj_io_analog_sel[6] mprj_io_hldh_n[6] mprj_io_analog_en[6] mprj_io_inp_dis[6] mprj_io_analog_pol[6] mprj_io_dm[18] mprj_io_dm[19] mprj_io_slow_sel[6] mprj_io_in[6] vccd 462 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X48 vssd vssa1 vssio vssio vddio vddio mprj_io[7] mprj_analog_io[0] mprj_io_ib_mode_sel[7] 464 mprj_io_enh[7] vdda1 vccd1 mprj_io_oeb[7] porb_h mprj_io_vtrip_sel[7] vccd vssio mprj_io_out[7] mprj_io_holdover[7]
+ mprj_io_dm[23] mprj_io_analog_sel[7] mprj_io_hldh_n[7] mprj_io_analog_en[7] mprj_io_inp_dis[7] mprj_io_analog_pol[7] mprj_io_dm[21] mprj_io_dm[22] mprj_io_slow_sel[7] mprj_io_in[7] vccd 464 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X49 vssd vssa1 vssio vssio vddio vddio mprj_io[8] mprj_analog_io[1] mprj_io_ib_mode_sel[8] 42 mprj_io_enh[8] vdda1 vccd1 mprj_io_oeb[8] porb_h mprj_io_vtrip_sel[8] vccd vssio mprj_io_out[8] mprj_io_holdover[8]
+ mprj_io_dm[26] mprj_io_analog_sel[8] mprj_io_hldh_n[8] mprj_io_analog_en[8] mprj_io_inp_dis[8] mprj_io_analog_pol[8] mprj_io_dm[24] mprj_io_dm[25] mprj_io_slow_sel[8] mprj_io_in[8] vccd 42 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X50 vssd vssa1 vssio vssio vddio vddio mprj_io[9] mprj_analog_io[2] mprj_io_ib_mode_sel[9] 43 mprj_io_enh[9] vdda1 vccd1 mprj_io_oeb[9] porb_h mprj_io_vtrip_sel[9] vccd vssio mprj_io_out[9] mprj_io_holdover[9]
+ mprj_io_dm[29] mprj_io_analog_sel[9] mprj_io_hldh_n[9] mprj_io_analog_en[9] mprj_io_inp_dis[9] mprj_io_analog_pol[9] mprj_io_dm[27] mprj_io_dm[28] mprj_io_slow_sel[9] mprj_io_in[9] vccd 43 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X51 vssd vssa1 vssio vssio vddio vddio mprj_io[10] mprj_analog_io[3] mprj_io_ib_mode_sel[10] 715 mprj_io_enh[10] vdda1 vccd1 mprj_io_oeb[10] porb_h mprj_io_vtrip_sel[10] vccd vssio mprj_io_out[10] mprj_io_holdover[10]
+ mprj_io_dm[32] mprj_io_analog_sel[10] mprj_io_hldh_n[10] mprj_io_analog_en[10] mprj_io_inp_dis[10] mprj_io_analog_pol[10] mprj_io_dm[30] mprj_io_dm[31] mprj_io_slow_sel[10] mprj_io_in[10] vccd 715 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X52 vssd vssa1 vssio vssio vddio vddio mprj_io[11] mprj_analog_io[4] mprj_io_ib_mode_sel[11] 465 mprj_io_enh[11] vdda1 vccd1 mprj_io_oeb[11] porb_h mprj_io_vtrip_sel[11] vccd vssio mprj_io_out[11] mprj_io_holdover[11]
+ mprj_io_dm[35] mprj_io_analog_sel[11] mprj_io_hldh_n[11] mprj_io_analog_en[11] mprj_io_inp_dis[11] mprj_io_analog_pol[11] mprj_io_dm[33] mprj_io_dm[34] mprj_io_slow_sel[11] mprj_io_in[11] vccd 465 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X53 vssd vssa1 vssio vssio vddio vddio mprj_io[12] mprj_analog_io[5] mprj_io_ib_mode_sel[12] 44 mprj_io_enh[12] vdda1 vccd1 mprj_io_oeb[12] porb_h mprj_io_vtrip_sel[12] vccd vssio mprj_io_out[12] mprj_io_holdover[12]
+ mprj_io_dm[38] mprj_io_analog_sel[12] mprj_io_hldh_n[12] mprj_io_analog_en[12] mprj_io_inp_dis[12] mprj_io_analog_pol[12] mprj_io_dm[36] mprj_io_dm[37] mprj_io_slow_sel[12] mprj_io_in[12] vccd 44 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X54 vssd vssa1 vssio vssio vddio vddio mprj_io[13] mprj_analog_io[6] mprj_io_ib_mode_sel[13] 45 mprj_io_enh[13] vdda1 vccd1 mprj_io_oeb[13] porb_h mprj_io_vtrip_sel[13] vccd vssio mprj_io_out[13] mprj_io_holdover[13]
+ mprj_io_dm[41] mprj_io_analog_sel[13] mprj_io_hldh_n[13] mprj_io_analog_en[13] mprj_io_inp_dis[13] mprj_io_analog_pol[13] mprj_io_dm[39] mprj_io_dm[40] mprj_io_slow_sel[13] mprj_io_in[13] vccd 45 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X55 vssd vssa1 vssio vssio vddio vddio mprj_io[14] mprj_analog_io[7] mprj_io_ib_mode_sel[14] 466 mprj_io_enh[14] vdda1 vccd1 mprj_io_oeb[14] porb_h mprj_io_vtrip_sel[14] vccd vssio mprj_io_out[14] mprj_io_holdover[14]
+ mprj_io_dm[44] mprj_io_analog_sel[14] mprj_io_hldh_n[14] mprj_io_analog_en[14] mprj_io_inp_dis[14] mprj_io_analog_pol[14] mprj_io_dm[42] mprj_io_dm[43] mprj_io_slow_sel[14] mprj_io_in[14] vccd 466 vddio 736 737
+ sky130_ef_io__gpiov2_pad_wrapped
X56 vssd vddio vssio 768 sky130_ef_io__vssio_hvc_clamped_pad
X57 vssd vddio vssio 776 sky130_ef_io__vssio_hvc_clamped_pad
X58 vssd vssio vccd vddio 765 sky130_ef_io__vssd_lvc_clamped_pad
X59 vssd vddio vccd vddio porb_h vssio vssio resetb vssio vccd vssio 23 vssio vssio resetb_core_h 23 sky130_fd_io__top_xres4v2
X60 vssd vssio vddio 755 sky130_ef_io__vddio_hvc_clamped_pad
X61 vssd vssio vddio 800 sky130_ef_io__vddio_hvc_clamped_pad
X62 vssd vssio vccd vddio 738 sky130_ef_io__vccd_lvc_clamped_pad
*.CALIBRE WARNING SHORT Short circuit(s) detected by extraction in this cell. See extraction report for details.
*.CALIBRE WARNING OPEN Open circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
