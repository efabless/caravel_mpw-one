magic
tech sky130A
magscale 12 1
timestamp 1598777870
<< metal5 >>
rect 0 20 15 75
rect 30 20 45 75
rect 0 10 45 20
rect 5 5 45 10
rect 10 0 45 5
rect 25 -15 45 0
rect 0 -20 45 -15
rect 0 -25 40 -20
rect 0 -30 35 -25
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
