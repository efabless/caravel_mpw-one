magic
tech sky130A
magscale 1 2
timestamp 1625664533
<< error_s >>
rect 145464 39289 145492 39299
rect 145436 39285 145492 39289
rect 145436 39271 145489 39285
rect 144523 39241 144579 39269
rect 144623 39261 144653 39269
rect 144523 39233 144551 39241
rect 144571 39233 144579 39241
rect 144597 39241 144653 39261
rect 145436 39261 145442 39271
rect 145436 39247 145461 39261
rect 145464 39247 145489 39271
rect 145436 39243 145464 39247
rect 145502 39242 145558 39247
rect 144523 39215 144571 39233
rect 144597 39215 144625 39241
rect 144523 39213 144625 39215
rect 145433 39219 145558 39242
rect 145433 39214 145489 39219
rect 144551 39205 144599 39213
rect 144543 39187 144599 39205
rect 145461 39191 145525 39214
rect 145530 39191 145558 39219
rect 144543 39159 144571 39187
rect 145461 39186 145489 39191
rect 145497 39163 145530 39178
rect 145497 39150 145553 39163
rect 145525 39122 145553 39150
rect 145571 39150 145627 39178
rect 145571 39135 145591 39150
rect 145599 39135 145627 39150
rect 145591 39122 145627 39135
rect 145573 39084 145591 39085
rect 141748 39020 141804 39048
rect 141847 39039 143068 39077
rect 143128 39039 144423 39077
rect 145601 39056 145619 39085
rect 141748 39011 141776 39020
rect 141784 39011 141804 39020
rect 141822 39020 141878 39039
rect 141748 38992 141784 39011
rect 141822 38992 141850 39020
rect 141682 38954 141738 38982
rect 141776 38969 141812 38982
rect 141684 38934 141712 38954
rect 141736 38934 141738 38954
rect 141684 38928 141738 38934
rect 141756 38954 141812 38969
rect 141684 38926 141736 38928
rect 141756 38926 141784 38954
rect 143002 38377 143122 38433
rect 143375 38390 143448 38433
rect 143328 38377 143448 38390
rect 142946 38373 143122 38377
rect 142946 38360 143066 38373
rect 143079 38360 143122 38373
rect 143315 38373 143448 38377
rect 142946 38317 143079 38360
rect 143315 38330 143392 38373
rect 142946 38300 143006 38317
rect 143019 38313 143079 38317
rect 143272 38317 143392 38330
rect 143019 38300 143066 38313
rect 142946 38257 143019 38300
rect 143272 38257 143332 38317
rect 145505 38178 145561 38188
rect 145601 38178 145635 38188
rect 145505 38148 145567 38178
rect 145579 38160 145635 38178
rect 145579 38148 145607 38160
rect 145465 38136 145607 38148
rect 145465 38132 145533 38136
rect 145539 38132 145607 38136
rect 145465 38120 145521 38132
rect 145539 38120 145595 38132
rect 145465 38108 145493 38120
rect 145501 38108 145521 38120
rect 145533 38108 145567 38120
rect 145465 38092 145501 38108
rect 145539 38092 145567 38108
rect 145493 38080 145529 38082
rect 145473 38054 145529 38080
rect 141813 37971 141933 38031
rect 145473 38026 145501 38054
rect 141813 37911 141820 37971
rect 141873 37911 141933 37971
rect 141656 37805 141684 37811
rect 141736 37795 141748 37811
rect 141684 37783 141748 37795
rect 141692 37767 141748 37783
rect 141684 37755 141720 37767
rect 141692 37739 141720 37755
rect 141594 36821 141629 36832
rect 141573 36804 141629 36821
rect 141573 36776 141601 36804
rect 145874 36711 145936 36743
rect 145874 36683 145994 36711
rect 145934 36623 145994 36683
rect 145418 34371 145470 34398
rect 145418 34343 145470 34370
rect 145318 33775 145374 33782
rect 145318 33737 145375 33775
rect 145273 33733 145403 33737
rect 145273 33710 145346 33733
rect 145347 33710 145403 33733
rect 145273 33709 145403 33710
rect 145296 33704 145376 33709
rect 145296 33682 145375 33704
rect 145296 33681 145348 33682
rect 145964 33624 146084 33684
rect 146155 33639 146230 33684
rect 145964 33609 146024 33624
rect 146027 33609 146084 33624
rect 146110 33624 146230 33639
rect 145964 33564 146027 33609
rect 146110 33564 146170 33624
rect 145821 33481 145941 33541
rect 146024 33489 146087 33541
rect 145821 33459 145881 33481
rect 145889 33459 145941 33481
rect 145967 33481 146087 33489
rect 145821 33424 145889 33459
rect 145967 33424 146027 33481
rect 145704 33421 146027 33424
rect 145704 33364 145824 33421
rect 145885 33369 145970 33421
rect 145721 33339 145824 33364
rect 145850 33364 145970 33369
rect 145721 33321 145769 33339
rect 145704 33304 145769 33321
rect 145850 33320 145910 33364
rect 145777 33304 145910 33320
rect 145777 33261 145866 33304
rect 145746 33260 145866 33261
rect 145746 33200 145806 33260
rect 133422 26450 133502 26500
rect 133422 26440 133542 26450
rect 133482 26380 133542 26440
rect 133889 26293 134009 26353
rect 133889 26270 133942 26293
rect 133949 26270 134009 26293
rect 133679 26210 133742 26243
rect 133942 26233 134009 26270
rect 133679 26183 133799 26210
rect 133739 26123 133799 26183
rect 133869 26000 133952 26053
rect 133869 25993 133989 26000
rect 133929 25933 133989 25993
rect 134062 25820 134132 25860
rect 134062 25800 134182 25820
rect 134122 25740 134182 25800
rect 134304 25584 134368 25618
rect 134304 25558 134424 25584
rect 134364 25520 134424 25558
rect 134402 25498 134424 25520
<< metal1 >>
rect 675426 875711 675482 875717
rect 671564 875655 671570 875711
rect 671626 875655 675426 875711
rect 675426 875649 675482 875655
rect 675465 875067 675521 875073
rect 671266 875011 671272 875067
rect 671328 875011 675465 875067
rect 675465 875005 675521 875011
rect 675437 872031 675493 872037
rect 671159 871975 671165 872031
rect 671221 871975 675437 872031
rect 675437 871969 675493 871975
rect 675471 871387 675527 871393
rect 671575 871331 671581 871387
rect 671637 871331 675471 871387
rect 675471 871325 675527 871331
rect 675419 870743 675475 870749
rect 673645 870687 673651 870743
rect 673707 870687 675419 870743
rect 675419 870681 675475 870687
rect 675434 864579 675490 864585
rect 671364 864523 671370 864579
rect 671426 864523 675434 864579
rect 675434 864517 675490 864523
rect 673652 862683 673658 862735
rect 673710 862683 675505 862735
rect 675557 862683 675563 862735
rect 42068 800067 42074 800123
rect 42130 800067 43597 800123
rect 43653 800067 43659 800123
rect 42068 798223 42074 798279
rect 42130 798223 43904 798279
rect 43960 798223 43966 798279
rect 42068 792055 42074 792111
rect 42130 792055 43594 792111
rect 43650 792055 43656 792111
rect 42068 791413 42074 791469
rect 42130 791413 43697 791469
rect 43753 791413 43759 791469
rect 42068 790771 42074 790827
rect 42130 790771 44111 790827
rect 44167 790771 44173 790827
rect 42068 787733 42074 787789
rect 42130 787733 44006 787789
rect 44062 787733 44068 787789
rect 42068 787087 42074 787143
rect 42130 787087 43693 787143
rect 43749 787087 43755 787143
rect 675426 786511 675482 786517
rect 671564 786455 671570 786511
rect 671626 786455 675426 786511
rect 675426 786449 675482 786455
rect 675465 785867 675521 785873
rect 671266 785811 671272 785867
rect 671328 785811 675465 785867
rect 675465 785805 675521 785811
rect 675437 782831 675493 782837
rect 671159 782775 671165 782831
rect 671221 782775 675437 782831
rect 675437 782769 675493 782775
rect 675471 782187 675527 782193
rect 671575 782131 671581 782187
rect 671637 782131 675471 782187
rect 675471 782125 675527 782131
rect 675419 781543 675475 781549
rect 673645 781487 673651 781543
rect 673707 781487 675419 781543
rect 675419 781481 675475 781487
rect 675434 775379 675490 775385
rect 671364 775323 671370 775379
rect 671426 775323 675434 775379
rect 675434 775317 675490 775323
rect 673652 773483 673658 773535
rect 673710 773483 675505 773535
rect 675557 773483 675563 773535
rect 41945 756467 41951 756523
rect 42007 756467 43597 756523
rect 43653 756467 43659 756523
rect 42068 755023 42074 755079
rect 42130 755023 43904 755079
rect 43960 755023 43966 755079
rect 42068 748855 42074 748911
rect 42130 748855 43594 748911
rect 43650 748855 43656 748911
rect 42068 748213 42074 748269
rect 42130 748213 43697 748269
rect 43753 748213 43759 748269
rect 42068 747571 42074 747627
rect 42130 747571 44111 747627
rect 44167 747571 44173 747627
rect 42068 744533 42074 744589
rect 42130 744533 44006 744589
rect 44062 744533 44068 744589
rect 42068 743887 42074 743943
rect 42130 743887 43693 743943
rect 43749 743887 43755 743943
rect 675426 741511 675482 741517
rect 671564 741455 671570 741511
rect 671626 741455 675426 741511
rect 675426 741449 675482 741455
rect 675465 740867 675521 740873
rect 671266 740811 671272 740867
rect 671328 740811 675465 740867
rect 675465 740805 675521 740811
rect 675437 737831 675493 737837
rect 671159 737775 671165 737831
rect 671221 737775 675437 737831
rect 675437 737769 675493 737775
rect 675471 737187 675527 737193
rect 671575 737131 671581 737187
rect 671637 737131 675471 737187
rect 675471 737125 675527 737131
rect 675419 736543 675475 736549
rect 674045 736487 674051 736543
rect 674107 736487 675419 736543
rect 675419 736481 675475 736487
rect 675434 730379 675490 730385
rect 671364 730323 671370 730379
rect 671426 730323 675434 730379
rect 675434 730317 675490 730323
rect 674052 728483 674058 728535
rect 674110 728483 675505 728535
rect 675557 728483 675563 728535
rect 42131 714045 42137 714101
rect 42193 714045 44223 714101
rect 44279 714045 44285 714101
rect 42068 711823 42074 711879
rect 42130 711823 43904 711879
rect 43960 711823 43966 711879
rect 42068 705655 42074 705711
rect 42130 705655 44228 705711
rect 44284 705655 44290 705711
rect 42068 705013 42074 705069
rect 42130 705013 43697 705069
rect 43753 705013 43759 705069
rect 42068 704371 42074 704427
rect 42130 704371 44111 704427
rect 44167 704371 44173 704427
rect 42068 701333 42074 701389
rect 42130 701333 44006 701389
rect 44062 701333 44068 701389
rect 42068 700687 42074 700743
rect 42130 700687 43693 700743
rect 43749 700687 43755 700743
rect 675426 696511 675482 696517
rect 671564 696455 671570 696511
rect 671626 696455 675426 696511
rect 675426 696449 675482 696455
rect 675465 695867 675521 695873
rect 671266 695811 671272 695867
rect 671328 695811 675465 695867
rect 675465 695805 675521 695811
rect 675437 692831 675493 692837
rect 671159 692775 671165 692831
rect 671221 692775 675437 692831
rect 675437 692769 675493 692775
rect 675471 692187 675527 692193
rect 671575 692131 671581 692187
rect 671637 692131 675471 692187
rect 675471 692125 675527 692131
rect 675419 691543 675475 691549
rect 674045 691487 674051 691543
rect 674107 691487 675419 691543
rect 675419 691481 675475 691487
rect 675434 685379 675490 685385
rect 671364 685323 671370 685379
rect 671426 685323 675434 685379
rect 675434 685317 675490 685323
rect 674052 683483 674058 683535
rect 674110 683483 675505 683535
rect 675557 683483 675563 683535
rect 41963 670067 41969 670123
rect 42025 670067 43597 670123
rect 43653 670067 43659 670123
rect 42068 668623 42074 668679
rect 42130 668623 43904 668679
rect 43960 668623 43966 668679
rect 42068 662455 42074 662511
rect 42130 662455 43594 662511
rect 43650 662455 43656 662511
rect 42068 661813 42074 661869
rect 42130 661813 43697 661869
rect 43753 661813 43759 661869
rect 42068 661171 42074 661227
rect 42130 661171 44111 661227
rect 44167 661171 44173 661227
rect 42068 658133 42074 658189
rect 42130 658133 44006 658189
rect 44062 658133 44068 658189
rect 42068 657487 42074 657543
rect 42130 657487 43693 657543
rect 43749 657487 43755 657543
rect 675426 651311 675482 651317
rect 671564 651255 671570 651311
rect 671626 651255 675426 651311
rect 675426 651249 675482 651255
rect 675465 650667 675521 650673
rect 671266 650611 671272 650667
rect 671328 650611 675465 650667
rect 675465 650605 675521 650611
rect 675437 647631 675493 647637
rect 671159 647575 671165 647631
rect 671221 647575 675437 647631
rect 675437 647569 675493 647575
rect 675471 646987 675527 646993
rect 671575 646931 671581 646987
rect 671637 646931 675471 646987
rect 675471 646925 675527 646931
rect 675419 646343 675475 646349
rect 673645 646287 673651 646343
rect 673707 646287 675419 646343
rect 675419 646281 675475 646287
rect 675434 640179 675490 640185
rect 671364 640123 671370 640179
rect 671426 640123 675434 640179
rect 675434 640117 675490 640123
rect 673652 638283 673658 638335
rect 673710 638283 675505 638335
rect 675557 638283 675563 638335
rect 42068 627267 42074 627323
rect 42130 627267 43597 627323
rect 43653 627267 43659 627323
rect 42068 625623 42074 625679
rect 42130 625623 43904 625679
rect 43960 625623 43966 625679
rect 42068 619255 42074 619311
rect 42130 619255 43594 619311
rect 43650 619255 43656 619311
rect 42068 618613 42074 618669
rect 42130 618613 43697 618669
rect 43753 618613 43759 618669
rect 42068 617971 42074 618027
rect 42130 617971 44111 618027
rect 44167 617971 44173 618027
rect 42068 614933 42074 614989
rect 42130 614933 44006 614989
rect 44062 614933 44068 614989
rect 42068 614287 42074 614343
rect 42130 614287 43693 614343
rect 43749 614287 43755 614343
rect 675426 606311 675482 606317
rect 671564 606255 671570 606311
rect 671626 606255 675426 606311
rect 675426 606249 675482 606255
rect 675465 605667 675521 605673
rect 671266 605611 671272 605667
rect 671328 605611 675465 605667
rect 675465 605605 675521 605611
rect 675437 602631 675493 602637
rect 671159 602575 671165 602631
rect 671221 602575 675437 602631
rect 675437 602569 675493 602575
rect 675471 601987 675527 601993
rect 675133 601952 675471 601987
rect 671575 601896 671581 601952
rect 671637 601931 675471 601952
rect 671637 601896 675189 601931
rect 675471 601925 675527 601931
rect 675419 601343 675475 601349
rect 674015 601287 674021 601343
rect 674077 601287 675419 601343
rect 675419 601281 675475 601287
rect 675434 595179 675490 595185
rect 671364 595123 671370 595179
rect 671426 595123 675434 595179
rect 675434 595117 675490 595123
rect 674022 593283 674028 593335
rect 674080 593283 675505 593335
rect 675557 593283 675563 593335
rect 42068 584067 42074 584123
rect 42130 584067 43217 584123
rect 43273 584067 43279 584123
rect 42099 582479 42105 582482
rect 42098 582426 42105 582479
rect 42161 582479 42167 582482
rect 42161 582426 43904 582479
rect 42098 582423 43904 582426
rect 43960 582423 43966 582479
rect 42068 576055 42074 576111
rect 42130 576055 43214 576111
rect 43270 576055 43276 576111
rect 42068 575413 42074 575469
rect 42130 575413 43697 575469
rect 43753 575413 43759 575469
rect 42068 574771 42074 574827
rect 42130 574771 44111 574827
rect 44167 574771 44173 574827
rect 42068 571733 42074 571789
rect 42130 571733 44006 571789
rect 44062 571733 44068 571789
rect 42068 571087 42074 571143
rect 42130 571087 43693 571143
rect 43749 571087 43755 571143
rect 675426 561111 675482 561117
rect 671564 561055 671570 561111
rect 671626 561055 675426 561111
rect 675426 561049 675482 561055
rect 675465 560467 675521 560473
rect 671266 560411 671272 560467
rect 671328 560411 675465 560467
rect 675465 560405 675521 560411
rect 675437 557431 675493 557437
rect 671159 557375 671165 557431
rect 671221 557375 675437 557431
rect 675437 557369 675493 557375
rect 675471 556787 675527 556793
rect 671575 556731 671581 556787
rect 671637 556731 675471 556787
rect 675471 556725 675527 556731
rect 675419 556143 675475 556149
rect 673245 556087 673251 556143
rect 673307 556087 675419 556143
rect 675419 556081 675475 556087
rect 675434 549979 675490 549985
rect 671364 549923 671370 549979
rect 671426 549923 675434 549979
rect 675434 549917 675490 549923
rect 673252 548083 673258 548135
rect 673310 548083 675505 548135
rect 675557 548083 675563 548135
rect 42068 540867 42074 540923
rect 42130 540867 43197 540923
rect 43253 540867 43259 540923
rect 42068 539023 42074 539079
rect 42130 539023 43904 539079
rect 43960 539023 43966 539079
rect 42068 532855 42074 532911
rect 42130 532855 43194 532911
rect 43250 532855 43256 532911
rect 42068 532213 42074 532269
rect 42130 532213 43697 532269
rect 43753 532213 43759 532269
rect 42068 531571 42074 531627
rect 42130 531571 44111 531627
rect 44167 531571 44173 531627
rect 42068 528533 42074 528589
rect 42130 528533 44006 528589
rect 44062 528533 44068 528589
rect 42068 527887 42074 527943
rect 42130 527887 43693 527943
rect 43749 527887 43755 527943
rect 42068 413267 42074 413323
rect 42130 413267 43597 413323
rect 43653 413267 43659 413323
rect 42068 411423 42074 411479
rect 42130 411423 43904 411479
rect 43960 411423 43966 411479
rect 42068 405255 42074 405311
rect 42130 405255 43594 405311
rect 43650 405255 43656 405311
rect 42068 404613 42074 404669
rect 42130 404613 43697 404669
rect 43753 404613 43759 404669
rect 42068 403971 42074 404027
rect 42130 403971 44111 404027
rect 44167 403971 44173 404027
rect 42068 400933 42074 400989
rect 42130 400933 44006 400989
rect 44062 400933 44068 400989
rect 42068 400287 42074 400343
rect 42130 400287 43693 400343
rect 43749 400287 43755 400343
rect 675426 383911 675482 383917
rect 671564 383855 671570 383911
rect 671626 383855 675426 383911
rect 675426 383849 675482 383855
rect 675465 383267 675521 383273
rect 671266 383211 671272 383267
rect 671328 383211 675465 383267
rect 675465 383205 675521 383211
rect 675437 380231 675493 380237
rect 671159 380175 671165 380231
rect 671221 380175 675437 380231
rect 675437 380169 675493 380175
rect 675471 379587 675527 379593
rect 671575 379531 671581 379587
rect 671637 379531 675471 379587
rect 675471 379525 675527 379531
rect 675419 378943 675475 378949
rect 673645 378887 673651 378943
rect 673707 378887 675419 378943
rect 675419 378881 675475 378887
rect 675434 372779 675490 372785
rect 671364 372723 671370 372779
rect 671426 372723 675434 372779
rect 675434 372717 675490 372723
rect 673652 370883 673658 370935
rect 673710 370883 675505 370935
rect 675557 370883 675563 370935
rect 42068 370067 42074 370123
rect 42130 370067 43597 370123
rect 43653 370067 43659 370123
rect 42068 368223 42074 368279
rect 42130 368223 43904 368279
rect 43960 368223 43966 368279
rect 42068 362055 42074 362111
rect 42130 362055 43594 362111
rect 43650 362055 43656 362111
rect 42068 361413 42074 361469
rect 42130 361413 43697 361469
rect 43753 361413 43759 361469
rect 42068 360771 42074 360827
rect 42130 360771 44111 360827
rect 44167 360771 44173 360827
rect 42068 357733 42074 357789
rect 42130 357733 44006 357789
rect 44062 357733 44068 357789
rect 42068 357087 42074 357143
rect 42130 357087 43693 357143
rect 43749 357087 43755 357143
rect 675426 338711 675482 338717
rect 671564 338655 671570 338711
rect 671626 338655 675426 338711
rect 675426 338649 675482 338655
rect 675465 338067 675521 338073
rect 671266 338011 671272 338067
rect 671328 338011 675465 338067
rect 675465 338005 675521 338011
rect 675437 335031 675493 335037
rect 671159 334975 671165 335031
rect 671221 334975 675437 335031
rect 675437 334969 675493 334975
rect 675471 334387 675527 334393
rect 671575 334331 671581 334387
rect 671637 334331 675471 334387
rect 675471 334325 675527 334331
rect 675419 333743 675475 333749
rect 673645 333687 673651 333743
rect 673707 333687 675419 333743
rect 675419 333681 675475 333687
rect 675434 327579 675490 327585
rect 671364 327523 671370 327579
rect 671426 327523 675434 327579
rect 675434 327517 675490 327523
rect 42068 326867 42074 326923
rect 42130 326867 43597 326923
rect 43653 326867 43659 326923
rect 673652 325683 673658 325735
rect 673710 325683 675505 325735
rect 675557 325683 675563 325735
rect 42068 325023 42074 325079
rect 42130 325023 43904 325079
rect 43960 325023 43966 325079
rect 42068 318855 42074 318911
rect 42130 318855 43594 318911
rect 43650 318855 43656 318911
rect 42068 318213 42074 318269
rect 42130 318213 43697 318269
rect 43753 318213 43759 318269
rect 42068 317571 42074 317627
rect 42130 317571 44111 317627
rect 44167 317571 44173 317627
rect 42068 314533 42074 314589
rect 42130 314533 44006 314589
rect 44062 314533 44068 314589
rect 42068 313887 42074 313943
rect 42130 313887 43693 313943
rect 43749 313887 43755 313943
rect 675426 293711 675482 293717
rect 671564 293655 671570 293711
rect 671626 293655 675426 293711
rect 675426 293649 675482 293655
rect 675465 293067 675521 293073
rect 671266 293011 671272 293067
rect 671328 293011 675465 293067
rect 675465 293005 675521 293011
rect 675437 290031 675493 290037
rect 671159 289975 671165 290031
rect 671221 289975 675437 290031
rect 675437 289969 675493 289975
rect 675471 289387 675527 289393
rect 671575 289331 671581 289387
rect 671637 289331 675471 289387
rect 675471 289325 675527 289331
rect 675419 288743 675475 288749
rect 673645 288687 673651 288743
rect 673707 288687 675419 288743
rect 675419 288681 675475 288687
rect 42068 283667 42074 283723
rect 42130 283667 43597 283723
rect 43653 283667 43659 283723
rect 675434 282579 675490 282585
rect 671364 282523 671370 282579
rect 671426 282523 675434 282579
rect 675434 282517 675490 282523
rect 42068 281823 42074 281879
rect 42130 281823 43904 281879
rect 43960 281823 43966 281879
rect 673652 280683 673658 280735
rect 673710 280683 675505 280735
rect 675557 280683 675563 280735
rect 42068 275655 42074 275711
rect 42130 275655 43594 275711
rect 43650 275655 43656 275711
rect 42068 275013 42074 275069
rect 42130 275013 43697 275069
rect 43753 275013 43759 275069
rect 42068 274371 42074 274427
rect 42130 274371 44111 274427
rect 44167 274371 44173 274427
rect 42068 271333 42074 271389
rect 42130 271333 44006 271389
rect 44062 271333 44068 271389
rect 42068 270687 42074 270743
rect 42130 270687 43693 270743
rect 43749 270687 43755 270743
rect 675426 248711 675482 248717
rect 671564 248655 671570 248711
rect 671626 248655 675426 248711
rect 675426 248649 675482 248655
rect 675465 248067 675521 248073
rect 671266 248011 671272 248067
rect 671328 248011 675465 248067
rect 675465 248005 675521 248011
rect 675437 245031 675493 245037
rect 671159 244975 671165 245031
rect 671221 244975 675437 245031
rect 675437 244969 675493 244975
rect 675471 244387 675527 244393
rect 671575 244331 671581 244387
rect 671637 244331 675471 244387
rect 675471 244325 675527 244331
rect 675419 243743 675475 243749
rect 673645 243687 673651 243743
rect 673707 243687 675419 243743
rect 675419 243681 675475 243687
rect 42068 240467 42074 240523
rect 42130 240467 43597 240523
rect 43653 240467 43659 240523
rect 42068 238623 42074 238679
rect 42130 238623 43904 238679
rect 43960 238623 43966 238679
rect 675434 237579 675490 237585
rect 671364 237523 671370 237579
rect 671426 237523 675434 237579
rect 675434 237517 675490 237523
rect 673652 235683 673658 235735
rect 673710 235683 675505 235735
rect 675557 235683 675563 235735
rect 42068 232455 42074 232511
rect 42130 232455 43594 232511
rect 43650 232455 43656 232511
rect 42068 231813 42074 231869
rect 42130 231813 43697 231869
rect 43753 231813 43759 231869
rect 42068 231171 42074 231227
rect 42130 231171 44111 231227
rect 44167 231171 44173 231227
rect 42068 228133 42074 228189
rect 42130 228133 44006 228189
rect 44062 228133 44068 228189
rect 42068 227487 42074 227543
rect 42130 227487 43693 227543
rect 43749 227487 43755 227543
rect 675426 203511 675482 203517
rect 671564 203455 671570 203511
rect 671626 203455 675426 203511
rect 675426 203449 675482 203455
rect 675465 202867 675521 202873
rect 671266 202811 671272 202867
rect 671328 202811 675465 202867
rect 675465 202805 675521 202811
rect 675437 199831 675493 199837
rect 671159 199775 671165 199831
rect 671221 199775 675437 199831
rect 675437 199769 675493 199775
rect 675471 199187 675527 199193
rect 671575 199131 671581 199187
rect 671637 199131 675471 199187
rect 675471 199125 675527 199131
rect 675419 198543 675475 198549
rect 673645 198487 673651 198543
rect 673707 198487 675419 198543
rect 675419 198481 675475 198487
rect 42068 197267 42074 197323
rect 42130 197267 43597 197323
rect 43653 197267 43659 197323
rect 42068 195423 42074 195479
rect 42130 195423 43904 195479
rect 43960 195423 43966 195479
rect 675434 192379 675490 192385
rect 671364 192323 671370 192379
rect 671426 192323 675434 192379
rect 675434 192317 675490 192323
rect 673652 190483 673658 190535
rect 673710 190483 675505 190535
rect 675557 190483 675563 190535
rect 42068 189255 42074 189311
rect 42130 189255 43594 189311
rect 43650 189255 43656 189311
rect 42068 188613 42074 188669
rect 42130 188613 43697 188669
rect 43753 188613 43759 188669
rect 42068 187971 42074 188027
rect 42130 187971 44111 188027
rect 44167 187971 44173 188027
rect 42068 184933 42074 184989
rect 42130 184933 44006 184989
rect 44062 184933 44068 184989
rect 43693 181266 43699 181278
rect 41414 181238 43699 181266
rect 41414 177471 41442 181238
rect 43693 181226 43699 181238
rect 43751 181226 43757 181278
rect 43904 181079 43910 181080
rect 41624 181029 43910 181079
rect 41624 177703 41674 181029
rect 43904 181028 43910 181029
rect 43962 181079 43968 181080
rect 43962 181029 43977 181079
rect 43962 181028 43968 181029
rect 44006 180979 44012 180980
rect 41724 180929 44012 180979
rect 41724 177803 41774 180929
rect 44006 180928 44012 180929
rect 44064 180979 44070 180980
rect 44064 180929 44086 180979
rect 44064 180928 44070 180929
rect 44104 180879 44110 180880
rect 41824 180829 44110 180879
rect 41824 177903 41874 180829
rect 44104 180828 44110 180829
rect 44162 180879 44168 180880
rect 44162 180829 44183 180879
rect 44162 180828 44168 180829
rect 41824 177853 42474 177903
rect 41724 177753 42374 177803
rect 41624 177653 42274 177703
rect 41414 177443 42042 177471
rect 42014 41861 42042 177443
rect 42224 69987 42274 177653
rect 42210 69967 42296 69987
rect 42210 69441 42216 69967
rect 42289 69441 42296 69967
rect 42210 69425 42296 69441
rect 42224 42134 42274 69425
rect 42324 42550 42374 177753
rect 42424 112755 42474 177853
rect 675426 158511 675482 158517
rect 671564 158455 671570 158511
rect 671626 158455 675426 158511
rect 675426 158449 675482 158455
rect 675465 157867 675521 157873
rect 671266 157811 671272 157867
rect 671328 157811 675465 157867
rect 675465 157805 675521 157811
rect 675437 154831 675493 154837
rect 671159 154775 671165 154831
rect 671221 154775 675437 154831
rect 675437 154769 675493 154775
rect 675471 154187 675527 154193
rect 671575 154131 671581 154187
rect 671637 154131 675471 154187
rect 675471 154125 675527 154131
rect 675419 153543 675475 153549
rect 673645 153487 673651 153543
rect 673707 153487 675419 153543
rect 675419 153481 675475 153487
rect 675434 147379 675490 147385
rect 671364 147323 671370 147379
rect 671426 147323 675434 147379
rect 675434 147317 675490 147323
rect 673652 145483 673658 145535
rect 673710 145483 675505 145535
rect 675557 145483 675563 145535
rect 675426 113311 675482 113317
rect 671564 113255 671570 113311
rect 671626 113255 675426 113311
rect 675426 113249 675482 113255
rect 42414 112734 42519 112755
rect 42414 112371 42428 112734
rect 42510 112371 42519 112734
rect 675465 112667 675521 112673
rect 671266 112611 671272 112667
rect 671328 112611 675465 112667
rect 675465 112605 675521 112611
rect 42414 112354 42519 112371
rect 42321 42544 42374 42550
rect 42321 42406 42374 42412
rect 42324 42395 42374 42406
rect 42424 42334 42474 112354
rect 675437 109631 675493 109637
rect 671159 109575 671165 109631
rect 671221 109575 675437 109631
rect 675437 109569 675493 109575
rect 675471 108987 675527 108993
rect 671575 108931 671581 108987
rect 671637 108931 675471 108987
rect 675471 108925 675527 108931
rect 675419 108343 675475 108349
rect 673645 108287 673651 108343
rect 673707 108287 675419 108343
rect 675419 108281 675475 108287
rect 675434 102179 675490 102185
rect 671364 102123 671370 102179
rect 671426 102123 675434 102179
rect 675434 102117 675490 102123
rect 673652 100283 673658 100335
rect 673710 100283 675505 100335
rect 675557 100283 675563 100335
rect 571321 42961 571764 42984
rect 467043 42754 467099 42760
rect 411009 42744 419695 42748
rect 411009 42692 411046 42744
rect 411040 42685 411046 42692
rect 411105 42692 419695 42744
rect 419751 42692 419757 42748
rect 464000 42698 464006 42754
rect 464062 42698 467043 42754
rect 467099 42698 470169 42754
rect 470225 42698 470231 42754
rect 467043 42692 467099 42698
rect 411105 42685 411111 42692
rect 518798 42671 518804 42723
rect 518856 42711 518862 42723
rect 524946 42711 524952 42723
rect 518856 42683 524952 42711
rect 518856 42671 518862 42683
rect 524946 42671 524952 42683
rect 525004 42671 525010 42723
rect 409204 42597 409210 42653
rect 409266 42597 412243 42653
rect 412299 42649 415444 42653
rect 412299 42597 415371 42649
rect 415365 42593 415371 42597
rect 415427 42597 415444 42649
rect 571321 42637 571346 42961
rect 415427 42593 415433 42597
rect 465839 42564 465845 42620
rect 465901 42564 474495 42620
rect 474551 42564 474557 42620
rect 505902 42601 571346 42637
rect 571737 42637 571764 42961
rect 571737 42601 671271 42637
rect 505902 42585 671271 42601
rect 671323 42585 671329 42637
rect 295280 42550 295286 42555
rect 295276 42508 295286 42550
rect 295280 42503 295286 42508
rect 295338 42550 295344 42555
rect 303284 42550 303290 42555
rect 295338 42508 303290 42550
rect 295338 42503 295344 42508
rect 303284 42503 303290 42508
rect 303342 42503 303348 42555
rect 350080 42550 350086 42555
rect 350076 42508 350086 42550
rect 350080 42503 350086 42508
rect 350138 42550 350144 42555
rect 358084 42550 358090 42555
rect 350138 42508 358090 42550
rect 350138 42503 350144 42508
rect 358084 42503 358090 42508
rect 358142 42503 358148 42555
rect 404880 42550 404886 42555
rect 404876 42508 404886 42550
rect 404880 42503 404886 42508
rect 404938 42550 404944 42555
rect 412884 42550 412890 42555
rect 404938 42508 412890 42550
rect 404938 42503 404944 42508
rect 412884 42503 412890 42508
rect 412942 42503 412948 42555
rect 505902 42464 505954 42585
rect 571321 42583 571764 42585
rect 523776 42508 523782 42509
rect 42527 42412 42582 42464
rect 42734 42412 140996 42464
rect 141048 42412 142570 42464
rect 142622 42412 143075 42464
rect 143127 42412 143432 42464
rect 143484 42412 144602 42464
rect 144654 42412 505954 42464
rect 506084 42458 523782 42508
rect 195976 42334 195982 42335
rect 42424 42284 195982 42334
rect 195976 42283 195982 42284
rect 196034 42334 196040 42335
rect 304576 42334 304582 42335
rect 196034 42284 304582 42334
rect 196034 42283 196040 42284
rect 304576 42283 304582 42284
rect 304634 42334 304640 42335
rect 359376 42334 359382 42335
rect 304634 42284 359382 42334
rect 304634 42283 304640 42284
rect 359376 42283 359382 42284
rect 359434 42334 359440 42335
rect 414176 42334 414182 42335
rect 359434 42284 414182 42334
rect 359434 42283 359440 42284
rect 414176 42283 414182 42284
rect 414234 42334 414240 42335
rect 468976 42334 468982 42335
rect 414234 42284 468982 42334
rect 414234 42283 414240 42284
rect 468976 42283 468982 42284
rect 469034 42334 469040 42335
rect 506084 42334 506134 42458
rect 523776 42457 523782 42458
rect 523834 42508 523840 42509
rect 671160 42508 671166 42509
rect 523834 42458 671166 42508
rect 523834 42457 523840 42458
rect 671160 42457 671166 42458
rect 671218 42508 671224 42509
rect 671218 42458 671236 42508
rect 671218 42457 671224 42458
rect 526810 42408 526816 42409
rect 469034 42284 506134 42334
rect 506184 42358 526816 42408
rect 469034 42283 469040 42284
rect 90863 42239 91094 42245
rect 90863 42234 90872 42239
rect 90846 42184 90872 42234
rect 90863 42183 90872 42184
rect 91085 42234 91094 42239
rect 199016 42234 199022 42235
rect 91085 42184 199022 42234
rect 91085 42183 91094 42184
rect 199016 42183 199022 42184
rect 199074 42234 199080 42235
rect 307610 42234 307616 42235
rect 199074 42184 307616 42234
rect 199074 42183 199080 42184
rect 307610 42183 307616 42184
rect 307668 42234 307674 42235
rect 362410 42234 362416 42235
rect 307668 42184 362416 42234
rect 307668 42183 307674 42184
rect 362410 42183 362416 42184
rect 362468 42234 362474 42235
rect 417210 42234 417216 42235
rect 362468 42184 417216 42234
rect 362468 42183 362474 42184
rect 417210 42183 417216 42184
rect 417268 42234 417274 42235
rect 472010 42234 472016 42235
rect 417268 42184 472016 42234
rect 417268 42183 417274 42184
rect 472010 42183 472016 42184
rect 472068 42234 472074 42235
rect 506184 42234 506234 42358
rect 526810 42357 526816 42358
rect 526868 42408 526874 42409
rect 526868 42358 526888 42408
rect 526868 42357 526874 42358
rect 516320 42308 516326 42309
rect 472068 42184 506234 42234
rect 506284 42258 516326 42308
rect 472068 42183 472074 42184
rect 90863 42174 91094 42183
rect 145847 42134 145853 42136
rect 42224 42084 145853 42134
rect 145847 42082 145853 42084
rect 145907 42134 145913 42136
rect 188520 42134 188526 42135
rect 145907 42084 188526 42134
rect 145907 42082 145913 42084
rect 188520 42083 188526 42084
rect 188578 42134 188584 42135
rect 192840 42134 192846 42135
rect 188578 42084 192846 42134
rect 188578 42083 188584 42084
rect 192840 42083 192846 42084
rect 192898 42134 192904 42135
rect 201486 42134 201492 42135
rect 192898 42084 201492 42134
rect 192898 42083 192904 42084
rect 201486 42083 201492 42084
rect 201544 42134 201550 42135
rect 297120 42134 297126 42135
rect 201544 42084 297126 42134
rect 201544 42083 201550 42084
rect 297120 42083 297126 42084
rect 297178 42134 297184 42135
rect 351920 42134 351926 42135
rect 297178 42132 351926 42134
rect 297178 42084 299607 42132
rect 297178 42083 297184 42084
rect 299601 42076 299607 42084
rect 299663 42130 351926 42132
rect 299663 42084 305771 42130
rect 299663 42076 299669 42084
rect 305765 42074 305771 42084
rect 305827 42084 351926 42130
rect 305827 42074 305833 42084
rect 351920 42083 351926 42084
rect 351978 42134 351984 42135
rect 360565 42134 360571 42139
rect 351978 42084 354407 42134
rect 351978 42083 351984 42084
rect 354401 42078 354407 42084
rect 354463 42084 360571 42134
rect 354463 42078 354469 42084
rect 360565 42083 360571 42084
rect 360627 42134 360633 42139
rect 406720 42134 406726 42135
rect 360627 42084 406726 42134
rect 360627 42083 360633 42084
rect 406720 42083 406726 42084
rect 406778 42134 406784 42135
rect 461520 42134 461526 42135
rect 406778 42084 461526 42134
rect 406778 42083 406784 42084
rect 461520 42083 461526 42084
rect 461578 42134 461584 42135
rect 506284 42134 506334 42258
rect 516320 42257 516326 42258
rect 516378 42308 516384 42309
rect 671360 42308 671366 42309
rect 516378 42258 671366 42308
rect 516378 42257 516384 42258
rect 671360 42257 671366 42258
rect 671418 42308 671424 42309
rect 671418 42258 671432 42308
rect 671418 42257 671424 42258
rect 516962 42208 516968 42209
rect 461578 42084 506334 42134
rect 506384 42158 516968 42208
rect 461578 42083 461584 42084
rect 189162 42034 189168 42035
rect 189160 41984 189168 42034
rect 189162 41983 189168 41984
rect 189220 42034 189226 42035
rect 191004 42034 191010 42035
rect 189220 41984 191010 42034
rect 189220 41983 189226 41984
rect 191004 41983 191010 41984
rect 191062 42034 191068 42035
rect 192194 42034 192200 42035
rect 191062 41984 192200 42034
rect 191062 41983 191068 41984
rect 192194 41983 192200 41984
rect 192252 42034 192258 42035
rect 193494 42034 193500 42035
rect 192252 41984 193500 42034
rect 192252 41983 192258 41984
rect 193494 41983 193500 41984
rect 193552 42034 193558 42035
rect 196518 42034 196524 42035
rect 193552 41984 196524 42034
rect 193552 41983 193558 41984
rect 196518 41983 196524 41984
rect 196576 42034 196582 42035
rect 197170 42034 197176 42035
rect 196576 41984 197176 42034
rect 196576 41983 196582 41984
rect 197170 41983 197176 41984
rect 197228 42034 197234 42035
rect 197810 42034 197816 42035
rect 197228 41984 197816 42034
rect 197228 41983 197234 41984
rect 197810 41983 197816 41984
rect 197868 42034 197874 42035
rect 198368 42034 198374 42035
rect 197868 41984 198374 42034
rect 197868 41983 197874 41984
rect 198368 41983 198374 41984
rect 198426 42034 198432 42035
rect 200208 42034 200214 42035
rect 198426 41984 200214 42034
rect 198426 41983 198432 41984
rect 200208 41983 200214 41984
rect 200266 42034 200272 42035
rect 200846 42034 200852 42035
rect 200266 41984 200852 42034
rect 200266 41983 200272 41984
rect 200846 41983 200852 41984
rect 200904 42034 200910 42035
rect 253613 42034 253827 42043
rect 297762 42034 297768 42035
rect 200904 41984 253622 42034
rect 200904 41983 200910 41984
rect 253613 41962 253622 41984
rect 253815 41984 297768 42034
rect 253815 41962 253827 41984
rect 297762 41983 297768 41984
rect 297820 42034 297826 42035
rect 300794 42034 300800 42035
rect 297820 41984 300800 42034
rect 297820 41983 297826 41984
rect 300794 41983 300800 41984
rect 300852 42034 300858 42035
rect 302094 42034 302100 42035
rect 300852 42033 302100 42034
rect 300852 41984 301447 42033
rect 300852 41983 300858 41984
rect 301441 41977 301447 41984
rect 301503 41984 302100 42033
rect 301503 41977 301509 41984
rect 302094 41983 302100 41984
rect 302152 42034 302158 42035
rect 305118 42034 305124 42035
rect 302152 41984 305124 42034
rect 302152 41983 302158 41984
rect 305118 41983 305124 41984
rect 305176 42034 305182 42035
rect 306410 42034 306416 42035
rect 305176 41984 306416 42034
rect 305176 41983 305182 41984
rect 306410 41983 306416 41984
rect 306468 42034 306474 42035
rect 308808 42034 308814 42035
rect 306468 41984 308814 42034
rect 306468 41983 306474 41984
rect 308808 41983 308814 41984
rect 308866 42034 308872 42035
rect 309446 42034 309452 42035
rect 308866 41984 309452 42034
rect 308866 41983 308872 41984
rect 309446 41983 309452 41984
rect 309504 42034 309510 42035
rect 352562 42034 352568 42035
rect 309504 41984 352568 42034
rect 309504 41983 309510 41984
rect 352562 41983 352568 41984
rect 352620 42034 352626 42035
rect 355594 42034 355600 42035
rect 352620 41984 355600 42034
rect 352620 41983 352626 41984
rect 355594 41983 355600 41984
rect 355652 42034 355658 42035
rect 356894 42034 356900 42035
rect 355652 42030 356900 42034
rect 355652 41984 356247 42030
rect 355652 41983 355658 41984
rect 356241 41974 356247 41984
rect 356303 41984 356900 42030
rect 356303 41974 356309 41984
rect 356894 41983 356900 41984
rect 356952 42034 356958 42035
rect 359918 42034 359924 42035
rect 356952 41984 359924 42034
rect 356952 41983 356958 41984
rect 359918 41983 359924 41984
rect 359976 42034 359982 42035
rect 361210 42034 361216 42035
rect 359976 41984 361216 42034
rect 359976 41983 359982 41984
rect 361210 41983 361216 41984
rect 361268 42034 361274 42035
rect 363608 42034 363614 42035
rect 361268 41984 363614 42034
rect 361268 41983 361274 41984
rect 363608 41983 363614 41984
rect 363666 42034 363672 42035
rect 364246 42034 364252 42035
rect 363666 41984 364252 42034
rect 363666 41983 363672 41984
rect 364246 41983 364252 41984
rect 364304 42034 364310 42035
rect 407362 42034 407368 42035
rect 364304 41984 407368 42034
rect 364304 41983 364310 41984
rect 407362 41983 407368 41984
rect 407420 42034 407426 42035
rect 410394 42034 410400 42035
rect 407420 41984 410400 42034
rect 407420 41983 407426 41984
rect 410394 41983 410400 41984
rect 410452 42034 410458 42035
rect 411694 42034 411700 42035
rect 410452 41984 411700 42034
rect 410452 41983 410458 41984
rect 411694 41983 411700 41984
rect 411752 42034 411758 42035
rect 414718 42034 414724 42035
rect 411752 41984 414724 42034
rect 411752 41983 411758 41984
rect 414718 41983 414724 41984
rect 414776 42034 414782 42035
rect 416010 42034 416016 42035
rect 414776 41984 416016 42034
rect 414776 41983 414782 41984
rect 416010 41983 416016 41984
rect 416068 42034 416074 42035
rect 418408 42034 418414 42035
rect 416068 41984 418414 42034
rect 416068 41983 416074 41984
rect 418408 41983 418414 41984
rect 418466 42034 418472 42035
rect 419046 42034 419052 42035
rect 418466 41984 419052 42034
rect 418466 41983 418472 41984
rect 419046 41983 419052 41984
rect 419104 42034 419110 42035
rect 462162 42034 462168 42035
rect 419104 41984 462168 42034
rect 419104 41983 419110 41984
rect 462162 41983 462168 41984
rect 462220 42034 462226 42035
rect 465194 42034 465200 42035
rect 462220 41984 465200 42034
rect 462220 41983 462226 41984
rect 465194 41983 465200 41984
rect 465252 42034 465258 42035
rect 466494 42034 466500 42035
rect 465252 41984 466500 42034
rect 465252 41983 465258 41984
rect 466494 41983 466500 41984
rect 466552 42034 466558 42035
rect 469518 42034 469524 42035
rect 466552 41984 469524 42034
rect 466552 41983 466558 41984
rect 469518 41983 469524 41984
rect 469576 42034 469582 42035
rect 470810 42034 470816 42035
rect 469576 41984 470816 42034
rect 469576 41983 469582 41984
rect 470810 41983 470816 41984
rect 470868 42034 470874 42035
rect 473208 42034 473214 42035
rect 470868 41984 473214 42034
rect 470868 41983 470874 41984
rect 473208 41983 473214 41984
rect 473266 42034 473272 42035
rect 473846 42034 473852 42035
rect 473266 41984 473852 42034
rect 473266 41983 473272 41984
rect 473846 41983 473852 41984
rect 473904 42034 473910 42035
rect 506384 42034 506434 42158
rect 516962 42157 516968 42158
rect 517020 42208 517026 42209
rect 519994 42208 520000 42209
rect 517020 42158 520000 42208
rect 517020 42157 517026 42158
rect 519994 42157 520000 42158
rect 520052 42208 520058 42209
rect 521294 42208 521300 42209
rect 520052 42158 521300 42208
rect 520052 42157 520058 42158
rect 521294 42157 521300 42158
rect 521352 42208 521358 42209
rect 524318 42208 524324 42209
rect 521352 42158 524324 42208
rect 521352 42157 521358 42158
rect 524318 42157 524324 42158
rect 524376 42208 524382 42209
rect 525610 42208 525616 42209
rect 524376 42158 525616 42208
rect 524376 42157 524382 42158
rect 525610 42157 525616 42158
rect 525668 42208 525674 42209
rect 528008 42208 528014 42209
rect 525668 42158 528014 42208
rect 525668 42157 525674 42158
rect 528008 42157 528014 42158
rect 528066 42208 528072 42209
rect 528646 42208 528652 42209
rect 528066 42158 528652 42208
rect 528066 42157 528072 42158
rect 528646 42157 528652 42158
rect 528704 42208 528710 42209
rect 528704 42158 528736 42208
rect 528704 42157 528710 42158
rect 514480 42114 514486 42119
rect 514476 42072 514486 42114
rect 514480 42067 514486 42072
rect 514538 42114 514544 42119
rect 522484 42114 522490 42119
rect 514538 42072 522490 42114
rect 514538 42067 514544 42072
rect 522484 42067 522490 42072
rect 522542 42067 522548 42119
rect 671563 42095 671569 42107
rect 636516 42067 671569 42095
rect 473904 41984 506434 42034
rect 473904 41983 473910 41984
rect 253613 41951 253827 41962
rect 186680 41940 186686 41945
rect 186676 41898 186686 41940
rect 186680 41893 186686 41898
rect 186738 41940 186744 41945
rect 194684 41940 194690 41945
rect 186738 41898 194690 41940
rect 186738 41893 186744 41898
rect 194684 41893 194690 41898
rect 194742 41893 194748 41945
rect 459680 41940 459686 41945
rect 459676 41898 459686 41940
rect 459680 41893 459686 41898
rect 459738 41940 459744 41945
rect 467684 41940 467690 41945
rect 459738 41898 467690 41940
rect 459738 41893 459744 41898
rect 467684 41893 467690 41898
rect 467742 41893 467748 41945
rect 195325 41861 195331 41887
rect 42014 41833 145091 41861
rect 145085 41809 145091 41833
rect 145143 41833 195331 41861
rect 145143 41809 145149 41833
rect 195325 41831 195331 41833
rect 195387 41861 195393 41887
rect 199649 41861 199655 41887
rect 195387 41833 199655 41861
rect 195387 41831 195393 41833
rect 199649 41831 199655 41833
rect 199711 41861 199717 41887
rect 303925 41861 303931 41871
rect 199711 41833 303931 41861
rect 199711 41831 199717 41833
rect 303925 41815 303931 41833
rect 303987 41861 303993 41871
rect 308249 41861 308255 41873
rect 303987 41833 308255 41861
rect 303987 41815 303993 41833
rect 308249 41817 308255 41833
rect 308311 41861 308317 41873
rect 358725 41861 358731 41871
rect 308311 41833 358731 41861
rect 308311 41817 308317 41833
rect 358725 41815 358731 41833
rect 358787 41861 358793 41871
rect 363049 41861 363055 41873
rect 358787 41833 363055 41861
rect 358787 41815 358793 41833
rect 363049 41817 363055 41833
rect 363111 41861 363117 41873
rect 413525 41861 413531 41871
rect 363111 41833 413531 41861
rect 363111 41817 363117 41833
rect 413525 41815 413531 41833
rect 413587 41861 413593 41871
rect 417849 41861 417855 41873
rect 413587 41833 417855 41861
rect 413587 41815 413593 41833
rect 417849 41817 417855 41833
rect 417911 41861 417917 41873
rect 468325 41861 468331 41875
rect 417911 41833 468331 41861
rect 417911 41817 417917 41833
rect 468325 41819 468331 41833
rect 468387 41861 468393 41875
rect 472649 41861 472655 41876
rect 468387 41833 472655 41861
rect 468387 41819 468393 41833
rect 472649 41820 472655 41833
rect 472711 41861 472717 41876
rect 523125 41861 523131 41873
rect 472711 41833 523131 41861
rect 472711 41820 472717 41833
rect 523125 41817 523131 41833
rect 523187 41861 523193 41873
rect 527449 41861 527455 41871
rect 523187 41833 527455 41861
rect 523187 41817 523193 41833
rect 527449 41815 527455 41833
rect 527511 41861 527517 41871
rect 636516 41861 636544 42067
rect 671563 42055 671569 42067
rect 671621 42055 671627 42107
rect 527511 41833 636544 41861
rect 527511 41815 527517 41833
rect 132992 40176 132998 40228
rect 133050 40221 133056 40228
rect 143919 40221 143925 40228
rect 133050 40183 143925 40221
rect 133050 40176 133056 40183
rect 143919 40176 143925 40183
rect 143977 40176 143983 40228
rect 142570 40122 142622 40128
rect 142570 40064 142622 40070
rect 142573 39946 142619 40064
<< via1 >>
rect 671570 875655 671626 875711
rect 675426 875655 675482 875711
rect 671272 875011 671328 875067
rect 675465 875011 675521 875067
rect 671165 871975 671221 872031
rect 675437 871975 675493 872031
rect 671581 871331 671637 871387
rect 675471 871331 675527 871387
rect 673651 870687 673707 870743
rect 675419 870687 675475 870743
rect 671370 864523 671426 864579
rect 675434 864523 675490 864579
rect 673658 862683 673710 862735
rect 675505 862683 675557 862735
rect 42074 800067 42130 800123
rect 43597 800067 43653 800123
rect 42074 798223 42130 798279
rect 43904 798223 43960 798279
rect 42074 792055 42130 792111
rect 43594 792055 43650 792111
rect 42074 791413 42130 791469
rect 43697 791413 43753 791469
rect 42074 790771 42130 790827
rect 44111 790771 44167 790827
rect 42074 787733 42130 787789
rect 44006 787733 44062 787789
rect 42074 787087 42130 787143
rect 43693 787087 43749 787143
rect 671570 786455 671626 786511
rect 675426 786455 675482 786511
rect 671272 785811 671328 785867
rect 675465 785811 675521 785867
rect 671165 782775 671221 782831
rect 675437 782775 675493 782831
rect 671581 782131 671637 782187
rect 675471 782131 675527 782187
rect 673651 781487 673707 781543
rect 675419 781487 675475 781543
rect 671370 775323 671426 775379
rect 675434 775323 675490 775379
rect 673658 773483 673710 773535
rect 675505 773483 675557 773535
rect 41951 756467 42007 756523
rect 43597 756467 43653 756523
rect 42074 755023 42130 755079
rect 43904 755023 43960 755079
rect 42074 748855 42130 748911
rect 43594 748855 43650 748911
rect 42074 748213 42130 748269
rect 43697 748213 43753 748269
rect 42074 747571 42130 747627
rect 44111 747571 44167 747627
rect 42074 744533 42130 744589
rect 44006 744533 44062 744589
rect 42074 743887 42130 743943
rect 43693 743887 43749 743943
rect 671570 741455 671626 741511
rect 675426 741455 675482 741511
rect 671272 740811 671328 740867
rect 675465 740811 675521 740867
rect 671165 737775 671221 737831
rect 675437 737775 675493 737831
rect 671581 737131 671637 737187
rect 675471 737131 675527 737187
rect 674051 736487 674107 736543
rect 675419 736487 675475 736543
rect 671370 730323 671426 730379
rect 675434 730323 675490 730379
rect 674058 728483 674110 728535
rect 675505 728483 675557 728535
rect 42137 714045 42193 714101
rect 44223 714045 44279 714101
rect 42074 711823 42130 711879
rect 43904 711823 43960 711879
rect 42074 705655 42130 705711
rect 44228 705655 44284 705711
rect 42074 705013 42130 705069
rect 43697 705013 43753 705069
rect 42074 704371 42130 704427
rect 44111 704371 44167 704427
rect 42074 701333 42130 701389
rect 44006 701333 44062 701389
rect 42074 700687 42130 700743
rect 43693 700687 43749 700743
rect 671570 696455 671626 696511
rect 675426 696455 675482 696511
rect 671272 695811 671328 695867
rect 675465 695811 675521 695867
rect 671165 692775 671221 692831
rect 675437 692775 675493 692831
rect 671581 692131 671637 692187
rect 675471 692131 675527 692187
rect 674051 691487 674107 691543
rect 675419 691487 675475 691543
rect 671370 685323 671426 685379
rect 675434 685323 675490 685379
rect 674058 683483 674110 683535
rect 675505 683483 675557 683535
rect 41969 670067 42025 670123
rect 43597 670067 43653 670123
rect 42074 668623 42130 668679
rect 43904 668623 43960 668679
rect 42074 662455 42130 662511
rect 43594 662455 43650 662511
rect 42074 661813 42130 661869
rect 43697 661813 43753 661869
rect 42074 661171 42130 661227
rect 44111 661171 44167 661227
rect 42074 658133 42130 658189
rect 44006 658133 44062 658189
rect 42074 657487 42130 657543
rect 43693 657487 43749 657543
rect 671570 651255 671626 651311
rect 675426 651255 675482 651311
rect 671272 650611 671328 650667
rect 675465 650611 675521 650667
rect 671165 647575 671221 647631
rect 675437 647575 675493 647631
rect 671581 646931 671637 646987
rect 675471 646931 675527 646987
rect 673651 646287 673707 646343
rect 675419 646287 675475 646343
rect 671370 640123 671426 640179
rect 675434 640123 675490 640179
rect 673658 638283 673710 638335
rect 675505 638283 675557 638335
rect 42074 627267 42130 627323
rect 43597 627267 43653 627323
rect 42074 625623 42130 625679
rect 43904 625623 43960 625679
rect 42074 619255 42130 619311
rect 43594 619255 43650 619311
rect 42074 618613 42130 618669
rect 43697 618613 43753 618669
rect 42074 617971 42130 618027
rect 44111 617971 44167 618027
rect 42074 614933 42130 614989
rect 44006 614933 44062 614989
rect 42074 614287 42130 614343
rect 43693 614287 43749 614343
rect 671570 606255 671626 606311
rect 675426 606255 675482 606311
rect 671272 605611 671328 605667
rect 675465 605611 675521 605667
rect 671165 602575 671221 602631
rect 675437 602575 675493 602631
rect 671581 601896 671637 601952
rect 675471 601931 675527 601987
rect 674021 601287 674077 601343
rect 675419 601287 675475 601343
rect 671370 595123 671426 595179
rect 675434 595123 675490 595179
rect 674028 593283 674080 593335
rect 675505 593283 675557 593335
rect 42074 584067 42130 584123
rect 43217 584067 43273 584123
rect 42105 582426 42161 582482
rect 43904 582423 43960 582479
rect 42074 576055 42130 576111
rect 43214 576055 43270 576111
rect 42074 575413 42130 575469
rect 43697 575413 43753 575469
rect 42074 574771 42130 574827
rect 44111 574771 44167 574827
rect 42074 571733 42130 571789
rect 44006 571733 44062 571789
rect 42074 571087 42130 571143
rect 43693 571087 43749 571143
rect 671570 561055 671626 561111
rect 675426 561055 675482 561111
rect 671272 560411 671328 560467
rect 675465 560411 675521 560467
rect 671165 557375 671221 557431
rect 675437 557375 675493 557431
rect 671581 556731 671637 556787
rect 675471 556731 675527 556787
rect 673251 556087 673307 556143
rect 675419 556087 675475 556143
rect 671370 549923 671426 549979
rect 675434 549923 675490 549979
rect 673258 548083 673310 548135
rect 675505 548083 675557 548135
rect 42074 540867 42130 540923
rect 43197 540867 43253 540923
rect 42074 539023 42130 539079
rect 43904 539023 43960 539079
rect 42074 532855 42130 532911
rect 43194 532855 43250 532911
rect 42074 532213 42130 532269
rect 43697 532213 43753 532269
rect 42074 531571 42130 531627
rect 44111 531571 44167 531627
rect 42074 528533 42130 528589
rect 44006 528533 44062 528589
rect 42074 527887 42130 527943
rect 43693 527887 43749 527943
rect 42074 413267 42130 413323
rect 43597 413267 43653 413323
rect 42074 411423 42130 411479
rect 43904 411423 43960 411479
rect 42074 405255 42130 405311
rect 43594 405255 43650 405311
rect 42074 404613 42130 404669
rect 43697 404613 43753 404669
rect 42074 403971 42130 404027
rect 44111 403971 44167 404027
rect 42074 400933 42130 400989
rect 44006 400933 44062 400989
rect 42074 400287 42130 400343
rect 43693 400287 43749 400343
rect 671570 383855 671626 383911
rect 675426 383855 675482 383911
rect 671272 383211 671328 383267
rect 675465 383211 675521 383267
rect 671165 380175 671221 380231
rect 675437 380175 675493 380231
rect 671581 379531 671637 379587
rect 675471 379531 675527 379587
rect 673651 378887 673707 378943
rect 675419 378887 675475 378943
rect 671370 372723 671426 372779
rect 675434 372723 675490 372779
rect 673658 370883 673710 370935
rect 675505 370883 675557 370935
rect 42074 370067 42130 370123
rect 43597 370067 43653 370123
rect 42074 368223 42130 368279
rect 43904 368223 43960 368279
rect 42074 362055 42130 362111
rect 43594 362055 43650 362111
rect 42074 361413 42130 361469
rect 43697 361413 43753 361469
rect 42074 360771 42130 360827
rect 44111 360771 44167 360827
rect 42074 357733 42130 357789
rect 44006 357733 44062 357789
rect 42074 357087 42130 357143
rect 43693 357087 43749 357143
rect 671570 338655 671626 338711
rect 675426 338655 675482 338711
rect 671272 338011 671328 338067
rect 675465 338011 675521 338067
rect 671165 334975 671221 335031
rect 675437 334975 675493 335031
rect 671581 334331 671637 334387
rect 675471 334331 675527 334387
rect 673651 333687 673707 333743
rect 675419 333687 675475 333743
rect 671370 327523 671426 327579
rect 675434 327523 675490 327579
rect 42074 326867 42130 326923
rect 43597 326867 43653 326923
rect 673658 325683 673710 325735
rect 675505 325683 675557 325735
rect 42074 325023 42130 325079
rect 43904 325023 43960 325079
rect 42074 318855 42130 318911
rect 43594 318855 43650 318911
rect 42074 318213 42130 318269
rect 43697 318213 43753 318269
rect 42074 317571 42130 317627
rect 44111 317571 44167 317627
rect 42074 314533 42130 314589
rect 44006 314533 44062 314589
rect 42074 313887 42130 313943
rect 43693 313887 43749 313943
rect 671570 293655 671626 293711
rect 675426 293655 675482 293711
rect 671272 293011 671328 293067
rect 675465 293011 675521 293067
rect 671165 289975 671221 290031
rect 675437 289975 675493 290031
rect 671581 289331 671637 289387
rect 675471 289331 675527 289387
rect 673651 288687 673707 288743
rect 675419 288687 675475 288743
rect 42074 283667 42130 283723
rect 43597 283667 43653 283723
rect 671370 282523 671426 282579
rect 675434 282523 675490 282579
rect 42074 281823 42130 281879
rect 43904 281823 43960 281879
rect 673658 280683 673710 280735
rect 675505 280683 675557 280735
rect 42074 275655 42130 275711
rect 43594 275655 43650 275711
rect 42074 275013 42130 275069
rect 43697 275013 43753 275069
rect 42074 274371 42130 274427
rect 44111 274371 44167 274427
rect 42074 271333 42130 271389
rect 44006 271333 44062 271389
rect 42074 270687 42130 270743
rect 43693 270687 43749 270743
rect 671570 248655 671626 248711
rect 675426 248655 675482 248711
rect 671272 248011 671328 248067
rect 675465 248011 675521 248067
rect 671165 244975 671221 245031
rect 675437 244975 675493 245031
rect 671581 244331 671637 244387
rect 675471 244331 675527 244387
rect 673651 243687 673707 243743
rect 675419 243687 675475 243743
rect 42074 240467 42130 240523
rect 43597 240467 43653 240523
rect 42074 238623 42130 238679
rect 43904 238623 43960 238679
rect 671370 237523 671426 237579
rect 675434 237523 675490 237579
rect 673658 235683 673710 235735
rect 675505 235683 675557 235735
rect 42074 232455 42130 232511
rect 43594 232455 43650 232511
rect 42074 231813 42130 231869
rect 43697 231813 43753 231869
rect 42074 231171 42130 231227
rect 44111 231171 44167 231227
rect 42074 228133 42130 228189
rect 44006 228133 44062 228189
rect 42074 227487 42130 227543
rect 43693 227487 43749 227543
rect 671570 203455 671626 203511
rect 675426 203455 675482 203511
rect 671272 202811 671328 202867
rect 675465 202811 675521 202867
rect 671165 199775 671221 199831
rect 675437 199775 675493 199831
rect 671581 199131 671637 199187
rect 675471 199131 675527 199187
rect 673651 198487 673707 198543
rect 675419 198487 675475 198543
rect 42074 197267 42130 197323
rect 43597 197267 43653 197323
rect 42074 195423 42130 195479
rect 43904 195423 43960 195479
rect 671370 192323 671426 192379
rect 675434 192323 675490 192379
rect 673658 190483 673710 190535
rect 675505 190483 675557 190535
rect 42074 189255 42130 189311
rect 43594 189255 43650 189311
rect 42074 188613 42130 188669
rect 43697 188613 43753 188669
rect 42074 187971 42130 188027
rect 44111 187971 44167 188027
rect 42074 184933 42130 184989
rect 44006 184933 44062 184989
rect 43699 181226 43751 181278
rect 43910 181028 43962 181080
rect 44012 180928 44064 180980
rect 44110 180828 44162 180880
rect 42216 69441 42289 69967
rect 671570 158455 671626 158511
rect 675426 158455 675482 158511
rect 671272 157811 671328 157867
rect 675465 157811 675521 157867
rect 671165 154775 671221 154831
rect 675437 154775 675493 154831
rect 671581 154131 671637 154187
rect 675471 154131 675527 154187
rect 673651 153487 673707 153543
rect 675419 153487 675475 153543
rect 671370 147323 671426 147379
rect 675434 147323 675490 147379
rect 673658 145483 673710 145535
rect 675505 145483 675557 145535
rect 671570 113255 671626 113311
rect 675426 113255 675482 113311
rect 42428 112371 42510 112734
rect 671272 112611 671328 112667
rect 675465 112611 675521 112667
rect 42321 42412 42374 42544
rect 671165 109575 671221 109631
rect 675437 109575 675493 109631
rect 671581 108931 671637 108987
rect 675471 108931 675527 108987
rect 673651 108287 673707 108343
rect 675419 108287 675475 108343
rect 671370 102123 671426 102179
rect 675434 102123 675490 102179
rect 673658 100283 673710 100335
rect 675505 100283 675557 100335
rect 411046 42685 411105 42744
rect 419695 42692 419751 42748
rect 464006 42698 464062 42754
rect 467043 42698 467099 42754
rect 470169 42698 470225 42754
rect 518804 42671 518856 42723
rect 524952 42671 525004 42723
rect 409210 42597 409266 42653
rect 412243 42597 412299 42653
rect 415371 42593 415427 42649
rect 465845 42564 465901 42620
rect 474495 42564 474551 42620
rect 571346 42601 571737 42961
rect 671271 42585 671323 42637
rect 295286 42503 295338 42555
rect 303290 42503 303342 42555
rect 350086 42503 350138 42555
rect 358090 42503 358142 42555
rect 404886 42503 404938 42555
rect 412890 42503 412942 42555
rect 42582 42412 42734 42464
rect 140996 42412 141048 42464
rect 142570 42412 142622 42464
rect 143075 42412 143127 42464
rect 143432 42412 143484 42464
rect 144602 42412 144654 42464
rect 195982 42283 196034 42335
rect 304582 42283 304634 42335
rect 359382 42283 359434 42335
rect 414182 42283 414234 42335
rect 468982 42283 469034 42335
rect 523782 42457 523834 42509
rect 671166 42457 671218 42509
rect 90872 42183 91085 42239
rect 199022 42183 199074 42235
rect 307616 42183 307668 42235
rect 362416 42183 362468 42235
rect 417216 42183 417268 42235
rect 472016 42183 472068 42235
rect 526816 42357 526868 42409
rect 145853 42082 145907 42136
rect 188526 42083 188578 42135
rect 192846 42083 192898 42135
rect 201492 42083 201544 42135
rect 297126 42083 297178 42135
rect 299607 42076 299663 42132
rect 305771 42074 305827 42130
rect 351926 42083 351978 42135
rect 354407 42078 354463 42134
rect 360571 42083 360627 42139
rect 406726 42083 406778 42135
rect 461526 42083 461578 42135
rect 516326 42257 516378 42309
rect 671366 42257 671418 42309
rect 189168 41983 189220 42035
rect 191010 41983 191062 42035
rect 192200 41983 192252 42035
rect 193500 41983 193552 42035
rect 196524 41983 196576 42035
rect 197176 41983 197228 42035
rect 197816 41983 197868 42035
rect 198374 41983 198426 42035
rect 200214 41983 200266 42035
rect 200852 41983 200904 42035
rect 253622 41962 253815 42034
rect 297768 41983 297820 42035
rect 300800 41983 300852 42035
rect 301447 41977 301503 42033
rect 302100 41983 302152 42035
rect 305124 41983 305176 42035
rect 306416 41983 306468 42035
rect 308814 41983 308866 42035
rect 309452 41983 309504 42035
rect 352568 41983 352620 42035
rect 355600 41983 355652 42035
rect 356247 41974 356303 42030
rect 356900 41983 356952 42035
rect 359924 41983 359976 42035
rect 361216 41983 361268 42035
rect 363614 41983 363666 42035
rect 364252 41983 364304 42035
rect 407368 41983 407420 42035
rect 410400 41983 410452 42035
rect 411700 41983 411752 42035
rect 414724 41983 414776 42035
rect 416016 41983 416068 42035
rect 418414 41983 418466 42035
rect 419052 41983 419104 42035
rect 462168 41983 462220 42035
rect 465200 41983 465252 42035
rect 466500 41983 466552 42035
rect 469524 41983 469576 42035
rect 470816 41983 470868 42035
rect 473214 41983 473266 42035
rect 473852 41983 473904 42035
rect 516968 42157 517020 42209
rect 520000 42157 520052 42209
rect 521300 42157 521352 42209
rect 524324 42157 524376 42209
rect 525616 42157 525668 42209
rect 528014 42157 528066 42209
rect 528652 42157 528704 42209
rect 514486 42067 514538 42119
rect 522490 42067 522542 42119
rect 186686 41893 186738 41945
rect 194690 41893 194742 41945
rect 459686 41893 459738 41945
rect 467690 41893 467742 41945
rect 145091 41809 145143 41861
rect 195331 41831 195387 41887
rect 199655 41831 199711 41887
rect 303931 41815 303987 41871
rect 308255 41817 308311 41873
rect 358731 41815 358787 41871
rect 363055 41817 363111 41873
rect 413531 41815 413587 41871
rect 417855 41817 417911 41873
rect 468331 41819 468387 41875
rect 472655 41820 472711 41876
rect 523131 41817 523187 41873
rect 527455 41815 527511 41871
rect 671569 42055 671621 42107
rect 132998 40176 133050 40228
rect 143925 40176 143977 40228
rect 142570 40070 142622 40122
<< metal2 >>
rect 230499 997600 235279 998010
rect 240478 997600 245258 1002732
rect 283099 997600 287879 998010
rect 293078 997600 297858 1002732
rect 384899 997600 389679 998010
rect 394878 997600 399658 1002732
rect 675407 878047 675887 878103
rect 675407 877495 675887 877551
rect 675407 876851 675887 876907
rect 675407 876207 675887 876263
rect 671576 875717 671614 875747
rect 671570 875711 671626 875717
rect 675407 875655 675426 875711
rect 675482 875655 675517 875711
rect 671570 875649 671626 875655
rect 671266 875073 671316 875102
rect 671266 875067 671328 875073
rect 671266 875011 671272 875067
rect 671266 875005 671328 875011
rect 671166 872037 671216 872055
rect 671161 872031 671221 872037
rect 671161 871975 671165 872031
rect 671161 871969 671221 871975
rect 43594 800129 43650 800144
rect 42074 800125 42130 800129
rect 41989 800123 42193 800125
rect 41989 800121 42074 800123
rect 41982 800117 42074 800121
rect 41970 800067 42074 800117
rect 42130 800067 42193 800123
rect 41970 800061 42193 800067
rect 43594 800123 43653 800129
rect 43594 800067 43597 800123
rect 43594 800061 43653 800067
rect 41713 799417 42193 799473
rect 42074 798281 42130 798285
rect 41989 798279 42193 798281
rect 41989 798277 42074 798279
rect 41980 798223 42074 798277
rect 42130 798223 42193 798279
rect 41980 798221 42193 798223
rect 42074 798217 42130 798221
rect 41713 797577 42193 797633
rect 41713 796933 42193 796989
rect 41713 795737 42193 795793
rect 41713 795093 42193 795149
rect 41713 794541 42193 794597
rect 41713 793897 42193 793953
rect 41713 793253 42193 793309
rect 41713 792701 42193 792757
rect 42074 792113 42130 792117
rect 41851 792111 42193 792113
rect 41851 792057 42074 792111
rect 41880 792055 42074 792057
rect 42130 792055 42193 792111
rect 41880 792053 42193 792055
rect 43594 792111 43650 800061
rect 43912 798285 43962 798355
rect 43904 798279 43962 798285
rect 43960 798223 43962 798279
rect 43904 798217 43962 798223
rect 42074 792049 42130 792053
rect 43594 792049 43650 792055
rect 43706 791475 43745 791509
rect 42074 791469 42130 791475
rect 43697 791469 43753 791475
rect 42031 791413 42074 791469
rect 42130 791413 42193 791469
rect 42031 791411 42193 791413
rect 42074 791407 42130 791411
rect 43697 791407 43753 791413
rect 42074 790827 42130 790833
rect 42029 790771 42074 790827
rect 42130 790771 42193 790827
rect 42029 790769 42193 790771
rect 42074 790765 42130 790769
rect 41713 790217 42193 790273
rect 41713 789573 42193 789629
rect 41713 788929 42193 788985
rect 41713 788377 42193 788433
rect 42074 787789 42130 787795
rect 42024 787733 42074 787789
rect 42130 787733 42193 787789
rect 42074 787727 42130 787733
rect 43706 787149 43745 791407
rect 42074 787145 42130 787149
rect 42008 787143 42193 787145
rect 42008 787089 42074 787143
rect 42017 787087 42074 787089
rect 42130 787087 42193 787143
rect 43693 787143 43749 787149
rect 42074 787081 42130 787087
rect 43693 787081 43749 787087
rect 41713 786537 42193 786593
rect 41713 785893 42193 785949
rect 41713 785249 42193 785305
rect 41713 784697 42193 784753
rect 41951 756523 42007 756881
rect 41951 756461 42007 756467
rect 43594 756529 43650 756544
rect 43594 756523 43653 756529
rect 43594 756467 43597 756523
rect 43594 756461 43653 756467
rect 41713 756217 42193 756273
rect 42074 755081 42130 755085
rect 41989 755079 42193 755081
rect 41989 755077 42074 755079
rect 41980 755023 42074 755077
rect 42130 755023 42193 755079
rect 41980 755021 42193 755023
rect 42074 755017 42130 755021
rect 41713 754377 42193 754433
rect 41713 753733 42193 753789
rect 41713 752537 42193 752593
rect 41713 751893 42193 751949
rect 41713 751341 42193 751397
rect 41713 750697 42193 750753
rect 41713 750053 42193 750109
rect 41713 749501 42193 749557
rect 42074 748913 42130 748917
rect 41851 748911 42193 748913
rect 41851 748857 42074 748911
rect 41880 748855 42074 748857
rect 42130 748855 42193 748911
rect 41880 748853 42193 748855
rect 43594 748911 43650 756461
rect 42074 748849 42130 748853
rect 43594 748849 43650 748855
rect 43706 748275 43745 787081
rect 43912 755085 43962 798217
rect 44112 790833 44162 790885
rect 44111 790827 44167 790833
rect 44111 790765 44167 790771
rect 44012 787795 44062 787820
rect 44006 787789 44062 787795
rect 44006 787727 44062 787733
rect 43904 755079 43962 755085
rect 43960 755023 43962 755079
rect 43904 755017 43962 755023
rect 42074 748269 42130 748275
rect 43697 748269 43753 748275
rect 42031 748213 42074 748269
rect 42130 748213 42193 748269
rect 42031 748211 42193 748213
rect 42074 748207 42130 748211
rect 43697 748207 43753 748213
rect 42074 747627 42130 747633
rect 42029 747571 42074 747627
rect 42130 747571 42193 747627
rect 42029 747569 42193 747571
rect 42074 747565 42130 747569
rect 41713 747017 42193 747073
rect 41713 746373 42193 746429
rect 41713 745729 42193 745785
rect 41713 745177 42193 745233
rect 42074 744589 42130 744595
rect 42024 744533 42074 744589
rect 42130 744533 42193 744589
rect 42074 744527 42130 744533
rect 43706 743949 43745 748207
rect 42074 743945 42130 743949
rect 42008 743943 42193 743945
rect 42008 743889 42074 743943
rect 42017 743887 42074 743889
rect 42130 743887 42193 743943
rect 43693 743943 43749 743949
rect 42074 743881 42130 743887
rect 43693 743881 43749 743887
rect 41713 743337 42193 743393
rect 41713 742693 42193 742749
rect 41713 742049 42193 742105
rect 41713 741497 42193 741553
rect 42137 714101 42193 714107
rect 42137 713717 42193 714045
rect 41967 713661 42193 713717
rect 41713 713017 42193 713073
rect 42074 711881 42130 711885
rect 41989 711879 42193 711881
rect 41989 711877 42074 711879
rect 41980 711823 42074 711877
rect 42130 711823 42193 711879
rect 41980 711821 42193 711823
rect 42074 711817 42130 711821
rect 41713 711177 42193 711233
rect 41713 710533 42193 710589
rect 41713 709337 42193 709393
rect 41713 708693 42193 708749
rect 41713 708141 42193 708197
rect 41713 707497 42193 707553
rect 41713 706853 42193 706909
rect 41713 706301 42193 706357
rect 42074 705713 42130 705717
rect 41851 705711 42193 705713
rect 41851 705657 42074 705711
rect 41880 705655 42074 705657
rect 42130 705655 42193 705711
rect 41880 705653 42193 705655
rect 42074 705649 42130 705653
rect 43706 705075 43745 743881
rect 43912 711885 43962 755017
rect 44012 744595 44062 787727
rect 44112 747633 44162 790765
rect 671166 782837 671216 871969
rect 671266 785873 671316 875005
rect 671576 871393 671614 875649
rect 675407 875011 675465 875067
rect 675521 875011 675591 875067
rect 675407 874367 675887 874423
rect 675407 873815 675887 873871
rect 675407 873171 675887 873227
rect 675407 872527 675887 872583
rect 675407 871975 675437 872031
rect 675493 871975 675566 872031
rect 671576 871387 671637 871393
rect 671576 871331 671581 871387
rect 675407 871331 675471 871387
rect 675527 871331 675573 871387
rect 671576 871325 671637 871331
rect 671366 864585 671416 864602
rect 671366 864579 671426 864585
rect 671366 864523 671370 864579
rect 671366 864517 671426 864523
rect 671266 785867 671328 785873
rect 671266 785811 671272 785867
rect 671266 785805 671328 785811
rect 671161 782831 671221 782837
rect 671161 782775 671165 782831
rect 671161 782769 671221 782775
rect 44111 747627 44167 747633
rect 44111 747565 44167 747571
rect 44006 744589 44062 744595
rect 44006 744527 44062 744533
rect 43904 711879 43962 711885
rect 43960 711823 43962 711879
rect 43904 711817 43962 711823
rect 42074 705069 42130 705075
rect 43697 705069 43753 705075
rect 42031 705013 42074 705069
rect 42130 705013 42193 705069
rect 42031 705011 42193 705013
rect 42074 705007 42130 705011
rect 43697 705007 43753 705013
rect 42074 704427 42130 704433
rect 42029 704371 42074 704427
rect 42130 704371 42193 704427
rect 42029 704369 42193 704371
rect 42074 704365 42130 704369
rect 41713 703817 42193 703873
rect 41713 703173 42193 703229
rect 41713 702529 42193 702585
rect 41713 701977 42193 702033
rect 42074 701389 42130 701395
rect 42024 701333 42074 701389
rect 42130 701333 42193 701389
rect 42074 701327 42130 701333
rect 43706 700749 43745 705007
rect 42074 700745 42130 700749
rect 42008 700743 42193 700745
rect 42008 700689 42074 700743
rect 42017 700687 42074 700689
rect 42130 700687 42193 700743
rect 43693 700743 43749 700749
rect 42074 700681 42130 700687
rect 43693 700681 43749 700687
rect 41713 700137 42193 700193
rect 41713 699493 42193 699549
rect 41713 698849 42193 698905
rect 41713 698297 42193 698353
rect 41969 670123 42025 670509
rect 41969 670061 42025 670067
rect 43594 670129 43650 670144
rect 43594 670123 43653 670129
rect 43594 670067 43597 670123
rect 43594 670061 43653 670067
rect 41713 669817 42193 669873
rect 42074 668681 42130 668685
rect 41989 668679 42193 668681
rect 41989 668677 42074 668679
rect 41980 668623 42074 668677
rect 42130 668623 42193 668679
rect 41980 668621 42193 668623
rect 42074 668617 42130 668621
rect 41713 667977 42193 668033
rect 41713 667333 42193 667389
rect 41713 666137 42193 666193
rect 41713 665493 42193 665549
rect 41713 664941 42193 664997
rect 41713 664297 42193 664353
rect 41713 663653 42193 663709
rect 41713 663101 42193 663157
rect 42074 662513 42130 662517
rect 41851 662511 42193 662513
rect 41851 662457 42074 662511
rect 41880 662455 42074 662457
rect 42130 662455 42193 662511
rect 41880 662453 42193 662455
rect 43594 662511 43650 670061
rect 42074 662449 42130 662453
rect 43594 662449 43650 662455
rect 43706 661875 43745 700681
rect 43912 668685 43962 711817
rect 44012 701395 44062 744527
rect 44112 704433 44162 747565
rect 671166 737837 671216 782769
rect 671266 740873 671316 785805
rect 671366 775385 671416 864517
rect 671576 786517 671614 871325
rect 673658 870749 673714 870768
rect 673651 870743 673714 870749
rect 673707 870687 673714 870743
rect 675407 870687 675419 870743
rect 675475 870687 675490 870743
rect 673651 870681 673714 870687
rect 673658 862735 673714 870681
rect 675407 870043 675887 870099
rect 675407 869491 675887 869547
rect 675407 868847 675887 868903
rect 675407 868203 675887 868259
rect 675407 867651 675887 867707
rect 675407 867007 675887 867063
rect 675407 865811 675887 865867
rect 675407 865167 675887 865223
rect 675407 864523 675434 864579
rect 675490 864523 675513 864579
rect 675407 863327 675887 863383
rect 675505 862739 675557 862741
rect 673710 862683 673714 862735
rect 675425 862735 675580 862739
rect 675425 862683 675505 862735
rect 675557 862683 675580 862735
rect 673658 862677 673714 862683
rect 675505 862677 675557 862683
rect 675407 788847 675887 788903
rect 675407 788295 675887 788351
rect 675407 787651 675887 787707
rect 675407 787007 675887 787063
rect 671570 786511 671626 786517
rect 675407 786455 675426 786511
rect 675482 786455 675517 786511
rect 671570 786449 671626 786455
rect 671576 782193 671614 786449
rect 675407 785811 675465 785867
rect 675521 785811 675591 785867
rect 675407 785167 675887 785223
rect 675407 784615 675887 784671
rect 675407 783971 675887 784027
rect 675407 783327 675887 783383
rect 675407 782775 675437 782831
rect 675493 782775 675566 782831
rect 671576 782187 671637 782193
rect 671576 782131 671581 782187
rect 675407 782131 675471 782187
rect 675527 782131 675573 782187
rect 671576 782125 671637 782131
rect 671366 775379 671426 775385
rect 671366 775323 671370 775379
rect 671366 775317 671426 775323
rect 671266 740867 671328 740873
rect 671266 740811 671272 740867
rect 671266 740805 671328 740811
rect 671161 737831 671221 737837
rect 671161 737775 671165 737831
rect 671161 737769 671221 737775
rect 44223 714101 44279 714107
rect 44223 705717 44279 714045
rect 44223 705711 44284 705717
rect 44223 705655 44228 705711
rect 44223 705649 44284 705655
rect 44223 705648 44279 705649
rect 44111 704427 44167 704433
rect 44111 704365 44167 704371
rect 44006 701389 44062 701395
rect 44006 701327 44062 701333
rect 43904 668679 43962 668685
rect 43960 668623 43962 668679
rect 43904 668617 43962 668623
rect 42074 661869 42130 661875
rect 43697 661869 43753 661875
rect 42031 661813 42074 661869
rect 42130 661813 42193 661869
rect 42031 661811 42193 661813
rect 42074 661807 42130 661811
rect 43697 661807 43753 661813
rect 42074 661227 42130 661233
rect 42029 661171 42074 661227
rect 42130 661171 42193 661227
rect 42029 661169 42193 661171
rect 42074 661165 42130 661169
rect 41713 660617 42193 660673
rect 41713 659973 42193 660029
rect 41713 659329 42193 659385
rect 41713 658777 42193 658833
rect 42074 658189 42130 658195
rect 42024 658133 42074 658189
rect 42130 658133 42193 658189
rect 42074 658127 42130 658133
rect 43706 657549 43745 661807
rect 42074 657545 42130 657549
rect 42008 657543 42193 657545
rect 42008 657489 42074 657543
rect 42017 657487 42074 657489
rect 42130 657487 42193 657543
rect 43693 657543 43749 657549
rect 42074 657481 42130 657487
rect 43693 657481 43749 657487
rect 41713 656937 42193 656993
rect 41713 656293 42193 656349
rect 41713 655649 42193 655705
rect 41713 655097 42193 655153
rect 43594 627329 43650 627344
rect 42074 627325 42130 627329
rect 41989 627323 42193 627325
rect 41989 627321 42074 627323
rect 41982 627317 42074 627321
rect 41970 627267 42074 627317
rect 42130 627267 42193 627323
rect 41970 627261 42193 627267
rect 43594 627323 43653 627329
rect 43594 627267 43597 627323
rect 43594 627261 43653 627267
rect 41713 626617 42193 626673
rect 42069 625685 42125 625691
rect 42069 625681 42130 625685
rect 42058 625679 42143 625681
rect 42058 625623 42074 625679
rect 42130 625623 42143 625679
rect 42058 625621 42143 625623
rect 42069 625617 42130 625621
rect 42069 625421 42125 625617
rect 41713 624777 42193 624833
rect 41713 624133 42193 624189
rect 41713 622937 42193 622993
rect 41713 622293 42193 622349
rect 41713 621741 42193 621797
rect 41713 621097 42193 621153
rect 41713 620453 42193 620509
rect 41713 619901 42193 619957
rect 42074 619313 42130 619317
rect 41851 619311 42193 619313
rect 41851 619257 42074 619311
rect 41880 619255 42074 619257
rect 42130 619255 42193 619311
rect 41880 619253 42193 619255
rect 43594 619311 43650 627261
rect 42074 619249 42130 619253
rect 43594 619249 43650 619255
rect 43706 618675 43745 657481
rect 43912 625685 43962 668617
rect 44012 658195 44062 701327
rect 44112 661233 44162 704365
rect 671166 692837 671216 737769
rect 671266 695873 671316 740805
rect 671366 730385 671416 775317
rect 671576 741517 671614 782125
rect 673658 781549 673714 781568
rect 673651 781543 673714 781549
rect 673707 781487 673714 781543
rect 675407 781487 675419 781543
rect 675475 781487 675490 781543
rect 673651 781481 673714 781487
rect 673658 773535 673714 781481
rect 675407 780843 675887 780899
rect 675407 780291 675887 780347
rect 675407 779647 675887 779703
rect 675407 779003 675887 779059
rect 675407 778451 675887 778507
rect 675407 777807 675887 777863
rect 675407 776611 675887 776667
rect 675407 775967 675887 776023
rect 675407 775323 675434 775379
rect 675490 775323 675513 775379
rect 675407 774127 675887 774183
rect 675505 773539 675557 773541
rect 673710 773483 673714 773535
rect 675425 773535 675580 773539
rect 675425 773483 675505 773535
rect 675557 773483 675580 773535
rect 673658 773477 673714 773483
rect 675505 773477 675557 773483
rect 675407 743847 675887 743903
rect 675407 743295 675887 743351
rect 675407 742651 675887 742707
rect 675407 742007 675887 742063
rect 671570 741511 671626 741517
rect 675407 741455 675426 741511
rect 675482 741455 675517 741511
rect 671570 741449 671626 741455
rect 671576 737193 671614 741449
rect 675407 740811 675465 740867
rect 675521 740811 675591 740867
rect 675407 740167 675887 740223
rect 675407 739615 675887 739671
rect 675407 738971 675887 739027
rect 675407 738327 675887 738383
rect 675407 737775 675437 737831
rect 675493 737775 675566 737831
rect 671576 737187 671637 737193
rect 671576 737131 671581 737187
rect 675407 737131 675471 737187
rect 675527 737131 675573 737187
rect 671576 737125 671637 737131
rect 671366 730379 671426 730385
rect 671366 730323 671370 730379
rect 671366 730317 671426 730323
rect 671266 695867 671328 695873
rect 671266 695811 671272 695867
rect 671266 695805 671328 695811
rect 671161 692831 671221 692837
rect 671161 692775 671165 692831
rect 671161 692769 671221 692775
rect 44111 661227 44167 661233
rect 44111 661165 44167 661171
rect 44006 658189 44062 658195
rect 44006 658127 44062 658133
rect 43904 625679 43962 625685
rect 43960 625623 43962 625679
rect 43904 625617 43962 625623
rect 42074 618669 42130 618675
rect 43697 618669 43753 618675
rect 42031 618613 42074 618669
rect 42130 618613 42193 618669
rect 42031 618611 42193 618613
rect 42074 618607 42130 618611
rect 43697 618607 43753 618613
rect 42074 618027 42130 618033
rect 42029 617971 42074 618027
rect 42130 617971 42193 618027
rect 42029 617969 42193 617971
rect 42074 617965 42130 617969
rect 41713 617417 42193 617473
rect 41713 616773 42193 616829
rect 41713 616129 42193 616185
rect 41713 615577 42193 615633
rect 42074 614989 42130 614995
rect 42024 614933 42074 614989
rect 42130 614933 42193 614989
rect 42074 614927 42130 614933
rect 43706 614349 43745 618607
rect 42074 614345 42130 614349
rect 42008 614343 42193 614345
rect 42008 614289 42074 614343
rect 42017 614287 42074 614289
rect 42130 614287 42193 614343
rect 43693 614343 43749 614349
rect 42074 614281 42130 614287
rect 43693 614281 43749 614287
rect 41713 613737 42193 613793
rect 41713 613093 42193 613149
rect 41713 612449 42193 612505
rect 41713 611897 42193 611953
rect 43214 584129 43270 584144
rect 42074 584125 42130 584129
rect 41989 584123 42193 584125
rect 41989 584121 42074 584123
rect 41982 584117 42074 584121
rect 41970 584067 42074 584117
rect 42130 584067 42193 584123
rect 41970 584061 42193 584067
rect 43214 584123 43273 584129
rect 43214 584067 43217 584123
rect 43214 584061 43273 584067
rect 41713 583417 42193 583473
rect 42105 582482 42161 582488
rect 42105 582221 42161 582426
rect 41713 581577 42193 581633
rect 41713 580933 42193 580989
rect 41713 579737 42193 579793
rect 41713 579093 42193 579149
rect 41713 578541 42193 578597
rect 41713 577897 42193 577953
rect 41713 577253 42193 577309
rect 41713 576701 42193 576757
rect 42074 576113 42130 576117
rect 41851 576111 42193 576113
rect 41851 576057 42074 576111
rect 41880 576055 42074 576057
rect 42130 576055 42193 576111
rect 41880 576053 42193 576055
rect 43214 576111 43270 584061
rect 42074 576049 42130 576053
rect 43214 576049 43270 576055
rect 43706 575475 43745 614281
rect 43912 582485 43962 625617
rect 44012 614995 44062 658127
rect 44112 618033 44162 661165
rect 671166 647637 671216 692769
rect 671266 650673 671316 695805
rect 671366 685385 671416 730317
rect 671576 696517 671614 737125
rect 674058 736549 674114 736568
rect 674051 736543 674114 736549
rect 674107 736487 674114 736543
rect 675407 736487 675419 736543
rect 675475 736487 675490 736543
rect 674051 736481 674114 736487
rect 674058 728535 674114 736481
rect 675407 735843 675887 735899
rect 675407 735291 675887 735347
rect 675407 734647 675887 734703
rect 675407 734003 675887 734059
rect 675407 733451 675887 733507
rect 675407 732807 675887 732863
rect 675407 731611 675887 731667
rect 675407 730967 675887 731023
rect 675407 730323 675434 730379
rect 675490 730323 675513 730379
rect 675407 729127 675887 729183
rect 675505 728539 675557 728541
rect 674110 728483 674114 728535
rect 675425 728535 675580 728539
rect 675425 728483 675505 728535
rect 675557 728483 675580 728535
rect 674058 728477 674114 728483
rect 675505 728477 675557 728483
rect 675407 698847 675887 698903
rect 675407 698295 675887 698351
rect 675407 697651 675887 697707
rect 675407 697007 675887 697063
rect 671570 696511 671626 696517
rect 675407 696455 675426 696511
rect 675482 696455 675517 696511
rect 671570 696449 671626 696455
rect 671576 692193 671614 696449
rect 675407 695811 675465 695867
rect 675521 695811 675591 695867
rect 675407 695167 675887 695223
rect 675407 694615 675887 694671
rect 675407 693971 675887 694027
rect 675407 693327 675887 693383
rect 675407 692775 675437 692831
rect 675493 692775 675566 692831
rect 671576 692187 671637 692193
rect 671576 692131 671581 692187
rect 675407 692131 675471 692187
rect 675527 692131 675573 692187
rect 671576 692125 671637 692131
rect 671366 685379 671426 685385
rect 671366 685323 671370 685379
rect 671366 685317 671426 685323
rect 671266 650667 671328 650673
rect 671266 650611 671272 650667
rect 671266 650605 671328 650611
rect 671161 647631 671221 647637
rect 671161 647575 671165 647631
rect 671161 647569 671221 647575
rect 44111 618027 44167 618033
rect 44111 617965 44167 617971
rect 44006 614989 44062 614995
rect 44006 614927 44062 614933
rect 43904 582479 43962 582485
rect 43960 582423 43962 582479
rect 43904 582417 43962 582423
rect 42074 575469 42130 575475
rect 43697 575469 43753 575475
rect 42031 575413 42074 575469
rect 42130 575413 42193 575469
rect 42031 575411 42193 575413
rect 42074 575407 42130 575411
rect 43697 575407 43753 575413
rect 42074 574827 42130 574833
rect 42029 574771 42074 574827
rect 42130 574771 42193 574827
rect 42029 574769 42193 574771
rect 42074 574765 42130 574769
rect 41713 574217 42193 574273
rect 41713 573573 42193 573629
rect 41713 572929 42193 572985
rect 41713 572377 42193 572433
rect 42074 571789 42130 571795
rect 42024 571733 42074 571789
rect 42130 571733 42193 571789
rect 42074 571727 42130 571733
rect 43706 571149 43745 575407
rect 42074 571145 42130 571149
rect 42008 571143 42193 571145
rect 42008 571089 42074 571143
rect 42017 571087 42074 571089
rect 42130 571087 42193 571143
rect 43693 571143 43749 571149
rect 42074 571081 42130 571087
rect 43693 571081 43749 571087
rect 41713 570537 42193 570593
rect 41713 569893 42193 569949
rect 41713 569249 42193 569305
rect 41713 568697 42193 568753
rect 43194 540929 43250 540944
rect 42074 540925 42130 540929
rect 41989 540923 42193 540925
rect 41989 540921 42074 540923
rect 41982 540917 42074 540921
rect 41970 540867 42074 540917
rect 42130 540867 42193 540923
rect 41970 540861 42193 540867
rect 43194 540923 43253 540929
rect 43194 540867 43197 540923
rect 43194 540861 43253 540867
rect 41713 540217 42193 540273
rect 42074 539081 42130 539085
rect 41989 539079 42193 539081
rect 41989 539077 42074 539079
rect 41980 539023 42074 539077
rect 42130 539023 42193 539079
rect 41980 539021 42193 539023
rect 42074 539017 42130 539021
rect 41713 538377 42193 538433
rect 41713 537733 42193 537789
rect 41713 536537 42193 536593
rect 41713 535893 42193 535949
rect 41713 535341 42193 535397
rect 41713 534697 42193 534753
rect 41713 534053 42193 534109
rect 41713 533501 42193 533557
rect 42074 532913 42130 532917
rect 41851 532911 42193 532913
rect 41851 532857 42074 532911
rect 41880 532855 42074 532857
rect 42130 532855 42193 532911
rect 41880 532853 42193 532855
rect 43194 532911 43250 540861
rect 42074 532849 42130 532853
rect 43194 532849 43250 532855
rect 43706 532275 43745 571081
rect 43912 539085 43962 582417
rect 44012 571795 44062 614927
rect 44112 574833 44162 617965
rect 671166 602637 671216 647569
rect 671266 605673 671316 650605
rect 671366 640185 671416 685317
rect 671576 651317 671614 692125
rect 674058 691549 674114 691568
rect 674051 691543 674114 691549
rect 674107 691487 674114 691543
rect 675407 691487 675419 691543
rect 675475 691487 675490 691543
rect 674051 691481 674114 691487
rect 674058 683535 674114 691481
rect 675407 690843 675887 690899
rect 675407 690291 675887 690347
rect 675407 689647 675887 689703
rect 675407 689003 675887 689059
rect 675407 688451 675887 688507
rect 675407 687807 675887 687863
rect 675407 686611 675887 686667
rect 675407 685967 675887 686023
rect 675407 685323 675434 685379
rect 675490 685323 675513 685379
rect 675407 684127 675887 684183
rect 675505 683539 675557 683541
rect 674110 683483 674114 683535
rect 675425 683535 675580 683539
rect 675425 683483 675505 683535
rect 675557 683483 675580 683535
rect 674058 683477 674114 683483
rect 675505 683477 675557 683483
rect 675407 653647 675887 653703
rect 675407 653095 675887 653151
rect 675407 652451 675887 652507
rect 675407 651807 675887 651863
rect 671570 651311 671626 651317
rect 675407 651255 675426 651311
rect 675482 651255 675517 651311
rect 671570 651249 671626 651255
rect 671576 646993 671614 651249
rect 675407 650611 675465 650667
rect 675521 650611 675591 650667
rect 675407 649967 675887 650023
rect 675407 649415 675887 649471
rect 675407 648771 675887 648827
rect 675407 648127 675887 648183
rect 675407 647575 675437 647631
rect 675493 647575 675566 647631
rect 671576 646987 671637 646993
rect 671576 646931 671581 646987
rect 675407 646931 675471 646987
rect 675527 646931 675573 646987
rect 671576 646925 671637 646931
rect 671366 640179 671426 640185
rect 671366 640123 671370 640179
rect 671366 640117 671426 640123
rect 671266 605667 671328 605673
rect 671266 605611 671272 605667
rect 671266 605605 671328 605611
rect 671161 602631 671221 602637
rect 671161 602575 671165 602631
rect 671161 602569 671221 602575
rect 44111 574827 44167 574833
rect 44111 574765 44167 574771
rect 44006 571789 44062 571795
rect 44006 571727 44062 571733
rect 43904 539079 43962 539085
rect 43960 539023 43962 539079
rect 43904 539017 43962 539023
rect 42074 532269 42130 532275
rect 43697 532269 43753 532275
rect 42031 532213 42074 532269
rect 42130 532213 42193 532269
rect 42031 532211 42193 532213
rect 42074 532207 42130 532211
rect 43697 532207 43753 532213
rect 42074 531627 42130 531633
rect 42029 531571 42074 531627
rect 42130 531571 42193 531627
rect 42029 531569 42193 531571
rect 42074 531565 42130 531569
rect 41713 531017 42193 531073
rect 41713 530373 42193 530429
rect 41713 529729 42193 529785
rect 41713 529177 42193 529233
rect 42074 528589 42130 528595
rect 42024 528533 42074 528589
rect 42130 528533 42193 528589
rect 42074 528527 42130 528533
rect 43706 527949 43745 532207
rect 42074 527945 42130 527949
rect 42008 527943 42193 527945
rect 42008 527889 42074 527943
rect 42017 527887 42074 527889
rect 42130 527887 42193 527943
rect 43693 527943 43749 527949
rect 42074 527881 42130 527887
rect 43693 527881 43749 527887
rect 41713 527337 42193 527393
rect 41713 526693 42193 526749
rect 41713 526049 42193 526105
rect 41713 525497 42193 525553
rect 43594 413329 43650 413344
rect 42074 413325 42130 413329
rect 41989 413323 42193 413325
rect 41989 413321 42074 413323
rect 41982 413317 42074 413321
rect 41970 413267 42074 413317
rect 42130 413267 42193 413323
rect 41970 413261 42193 413267
rect 43594 413323 43653 413329
rect 43594 413267 43597 413323
rect 43594 413261 43653 413267
rect 41713 412617 42193 412673
rect 42074 411481 42130 411485
rect 41989 411479 42193 411481
rect 41989 411477 42074 411479
rect 41980 411423 42074 411477
rect 42130 411423 42193 411479
rect 41980 411421 42193 411423
rect 42074 411417 42130 411421
rect 41713 410777 42193 410833
rect 41713 410133 42193 410189
rect 41713 408937 42193 408993
rect 41713 408293 42193 408349
rect 41713 407741 42193 407797
rect 41713 407097 42193 407153
rect 41713 406453 42193 406509
rect 41713 405901 42193 405957
rect 42074 405313 42130 405317
rect 41851 405311 42193 405313
rect 41851 405257 42074 405311
rect 41880 405255 42074 405257
rect 42130 405255 42193 405311
rect 41880 405253 42193 405255
rect 43594 405311 43650 413261
rect 42074 405249 42130 405253
rect 43594 405249 43650 405255
rect 43706 404675 43745 527881
rect 43912 411485 43962 539017
rect 44012 528595 44062 571727
rect 44112 531633 44162 574765
rect 671166 557437 671216 602569
rect 671266 560473 671316 605605
rect 671366 595185 671416 640117
rect 671576 606317 671614 646925
rect 673658 646349 673714 646368
rect 673651 646343 673714 646349
rect 673707 646287 673714 646343
rect 675407 646287 675419 646343
rect 675475 646287 675490 646343
rect 673651 646281 673714 646287
rect 673658 638335 673714 646281
rect 675407 645643 675887 645699
rect 675407 645091 675887 645147
rect 675407 644447 675887 644503
rect 675407 643803 675887 643859
rect 675407 643251 675887 643307
rect 675407 642607 675887 642663
rect 675407 641411 675887 641467
rect 675407 640767 675887 640823
rect 675407 640123 675434 640179
rect 675490 640123 675513 640179
rect 675407 638927 675887 638983
rect 675505 638339 675557 638341
rect 673710 638283 673714 638335
rect 675425 638335 675580 638339
rect 675425 638283 675505 638335
rect 675557 638283 675580 638335
rect 673658 638277 673714 638283
rect 675505 638277 675557 638283
rect 675407 608647 675887 608703
rect 675407 608095 675887 608151
rect 675407 607451 675887 607507
rect 675407 606807 675887 606863
rect 671570 606311 671626 606317
rect 675407 606255 675426 606311
rect 675482 606255 675517 606311
rect 671570 606249 671626 606255
rect 671576 601958 671614 606249
rect 675407 605611 675465 605667
rect 675521 605611 675591 605667
rect 675407 604967 675887 605023
rect 675407 604415 675887 604471
rect 675407 603771 675887 603827
rect 675407 603127 675887 603183
rect 675407 602575 675437 602631
rect 675493 602575 675566 602631
rect 671576 601952 671637 601958
rect 671576 601896 671581 601952
rect 675407 601931 675471 601987
rect 675527 601931 675573 601987
rect 671576 601890 671637 601896
rect 671366 595179 671426 595185
rect 671366 595123 671370 595179
rect 671366 595117 671426 595123
rect 671266 560467 671328 560473
rect 671266 560411 671272 560467
rect 671266 560405 671328 560411
rect 671161 557431 671221 557437
rect 671161 557375 671165 557431
rect 671161 557369 671221 557375
rect 44111 531627 44167 531633
rect 44111 531565 44167 531571
rect 44006 528589 44062 528595
rect 44006 528527 44062 528533
rect 43904 411479 43962 411485
rect 43960 411423 43962 411479
rect 43904 411417 43962 411423
rect 42074 404669 42130 404675
rect 43697 404669 43753 404675
rect 42031 404613 42074 404669
rect 42130 404613 42193 404669
rect 42031 404611 42193 404613
rect 42074 404607 42130 404611
rect 43697 404607 43753 404613
rect 42074 404027 42130 404033
rect 42029 403971 42074 404027
rect 42130 403971 42193 404027
rect 42029 403969 42193 403971
rect 42074 403965 42130 403969
rect 41713 403417 42193 403473
rect 41713 402773 42193 402829
rect 41713 402129 42193 402185
rect 41713 401577 42193 401633
rect 42074 400989 42130 400995
rect 42024 400933 42074 400989
rect 42130 400933 42193 400989
rect 42074 400927 42130 400933
rect 43706 400349 43745 404607
rect 42074 400345 42130 400349
rect 42008 400343 42193 400345
rect 42008 400289 42074 400343
rect 42017 400287 42074 400289
rect 42130 400287 42193 400343
rect 43693 400343 43749 400349
rect 42074 400281 42130 400287
rect 43693 400281 43749 400287
rect 41713 399737 42193 399793
rect 41713 399093 42193 399149
rect 41713 398449 42193 398505
rect 41713 397897 42193 397953
rect 43594 370129 43650 370144
rect 42074 370125 42130 370129
rect 41989 370123 42193 370125
rect 41989 370121 42074 370123
rect 41982 370117 42074 370121
rect 41970 370067 42074 370117
rect 42130 370067 42193 370123
rect 41970 370061 42193 370067
rect 43594 370123 43653 370129
rect 43594 370067 43597 370123
rect 43594 370061 43653 370067
rect 41713 369417 42193 369473
rect 42074 368281 42130 368285
rect 41989 368279 42193 368281
rect 41989 368277 42074 368279
rect 41980 368223 42074 368277
rect 42130 368223 42193 368279
rect 41980 368221 42193 368223
rect 42074 368217 42130 368221
rect 41713 367577 42193 367633
rect 41713 366933 42193 366989
rect 41713 365737 42193 365793
rect 41713 365093 42193 365149
rect 41713 364541 42193 364597
rect 41713 363897 42193 363953
rect 41713 363253 42193 363309
rect 41713 362701 42193 362757
rect 42074 362113 42130 362117
rect 41851 362111 42193 362113
rect 41851 362057 42074 362111
rect 41880 362055 42074 362057
rect 42130 362055 42193 362111
rect 41880 362053 42193 362055
rect 43594 362111 43650 370061
rect 42074 362049 42130 362053
rect 43594 362049 43650 362055
rect 43706 361475 43745 400281
rect 43912 368285 43962 411417
rect 44012 400995 44062 528527
rect 44112 404033 44162 531565
rect 44111 404027 44167 404033
rect 44111 403965 44167 403971
rect 44006 400989 44062 400995
rect 44006 400927 44062 400933
rect 43904 368279 43962 368285
rect 43960 368223 43962 368279
rect 43904 368217 43962 368223
rect 42074 361469 42130 361475
rect 43697 361469 43753 361475
rect 42031 361413 42074 361469
rect 42130 361413 42193 361469
rect 42031 361411 42193 361413
rect 42074 361407 42130 361411
rect 43697 361407 43753 361413
rect 42074 360827 42130 360833
rect 42029 360771 42074 360827
rect 42130 360771 42193 360827
rect 42029 360769 42193 360771
rect 42074 360765 42130 360769
rect 41713 360217 42193 360273
rect 41713 359573 42193 359629
rect 41713 358929 42193 358985
rect 41713 358377 42193 358433
rect 42074 357789 42130 357795
rect 42024 357733 42074 357789
rect 42130 357733 42193 357789
rect 42074 357727 42130 357733
rect 43706 357149 43745 361407
rect 42074 357145 42130 357149
rect 42008 357143 42193 357145
rect 42008 357089 42074 357143
rect 42017 357087 42074 357089
rect 42130 357087 42193 357143
rect 43693 357143 43749 357149
rect 42074 357081 42130 357087
rect 43693 357081 43749 357087
rect 41713 356537 42193 356593
rect 41713 355893 42193 355949
rect 41713 355249 42193 355305
rect 41713 354697 42193 354753
rect 43594 326929 43650 326944
rect 42074 326925 42130 326929
rect 41989 326923 42193 326925
rect 41989 326921 42074 326923
rect 41982 326917 42074 326921
rect 41970 326867 42074 326917
rect 42130 326867 42193 326923
rect 41970 326861 42193 326867
rect 43594 326923 43653 326929
rect 43594 326867 43597 326923
rect 43594 326861 43653 326867
rect 41713 326217 42193 326273
rect 42074 325081 42130 325085
rect 41989 325079 42193 325081
rect 41989 325077 42074 325079
rect 41980 325023 42074 325077
rect 42130 325023 42193 325079
rect 41980 325021 42193 325023
rect 42074 325017 42130 325021
rect 41713 324377 42193 324433
rect 41713 323733 42193 323789
rect 41713 322537 42193 322593
rect 41713 321893 42193 321949
rect 41713 321341 42193 321397
rect 41713 320697 42193 320753
rect 41713 320053 42193 320109
rect 41713 319501 42193 319557
rect 42074 318913 42130 318917
rect 41851 318911 42193 318913
rect 41851 318857 42074 318911
rect 41880 318855 42074 318857
rect 42130 318855 42193 318911
rect 41880 318853 42193 318855
rect 43594 318911 43650 326861
rect 42074 318849 42130 318853
rect 43594 318849 43650 318855
rect 43706 318275 43745 357081
rect 43912 325085 43962 368217
rect 44012 357795 44062 400927
rect 44112 360833 44162 403965
rect 671166 380237 671216 557369
rect 671266 383273 671316 560405
rect 671366 549985 671416 595117
rect 671576 561117 671614 601890
rect 674028 601349 674081 601368
rect 674021 601343 674081 601349
rect 674077 601287 674081 601343
rect 675407 601287 675419 601343
rect 675475 601287 675490 601343
rect 674021 601281 674081 601287
rect 674028 593335 674081 601281
rect 675407 600643 675887 600699
rect 675407 600091 675887 600147
rect 675407 599447 675887 599503
rect 675407 598803 675887 598859
rect 675407 598251 675887 598307
rect 675407 597607 675887 597663
rect 675407 596411 675887 596467
rect 675407 595767 675887 595823
rect 675407 595123 675434 595179
rect 675490 595123 675513 595179
rect 675407 593927 675887 593983
rect 675505 593339 675557 593341
rect 674080 593283 674081 593335
rect 675425 593335 675580 593339
rect 675425 593283 675505 593335
rect 675557 593283 675580 593335
rect 674028 593277 674081 593283
rect 675505 593277 675557 593283
rect 675407 563447 675887 563503
rect 675407 562895 675887 562951
rect 675407 562251 675887 562307
rect 675407 561607 675887 561663
rect 671570 561111 671626 561117
rect 675407 561055 675426 561111
rect 675482 561055 675517 561111
rect 671570 561049 671626 561055
rect 671576 556793 671614 561049
rect 675407 560411 675465 560467
rect 675521 560411 675591 560467
rect 675407 559767 675887 559823
rect 675407 559215 675887 559271
rect 675407 558571 675887 558627
rect 675407 557927 675887 557983
rect 675407 557375 675437 557431
rect 675493 557375 675566 557431
rect 671576 556787 671637 556793
rect 671576 556731 671581 556787
rect 675407 556731 675471 556787
rect 675527 556731 675573 556787
rect 671576 556725 671637 556731
rect 671366 549979 671426 549985
rect 671366 549923 671370 549979
rect 671366 549917 671426 549923
rect 671266 383267 671328 383273
rect 671266 383211 671272 383267
rect 671266 383205 671328 383211
rect 671161 380231 671221 380237
rect 671161 380175 671165 380231
rect 671161 380169 671221 380175
rect 44111 360827 44167 360833
rect 44111 360765 44167 360771
rect 44006 357789 44062 357795
rect 44006 357727 44062 357733
rect 43904 325079 43962 325085
rect 43960 325023 43962 325079
rect 43904 325017 43962 325023
rect 42074 318269 42130 318275
rect 43697 318269 43753 318275
rect 42031 318213 42074 318269
rect 42130 318213 42193 318269
rect 42031 318211 42193 318213
rect 42074 318207 42130 318211
rect 43697 318207 43753 318213
rect 42074 317627 42130 317633
rect 42029 317571 42074 317627
rect 42130 317571 42193 317627
rect 42029 317569 42193 317571
rect 42074 317565 42130 317569
rect 41713 317017 42193 317073
rect 41713 316373 42193 316429
rect 41713 315729 42193 315785
rect 41713 315177 42193 315233
rect 42074 314589 42130 314595
rect 42024 314533 42074 314589
rect 42130 314533 42193 314589
rect 42074 314527 42130 314533
rect 43706 313949 43745 318207
rect 42074 313945 42130 313949
rect 42008 313943 42193 313945
rect 42008 313889 42074 313943
rect 42017 313887 42074 313889
rect 42130 313887 42193 313943
rect 43693 313943 43749 313949
rect 42074 313881 42130 313887
rect 43693 313881 43749 313887
rect 41713 313337 42193 313393
rect 41713 312693 42193 312749
rect 41713 312049 42193 312105
rect 41713 311497 42193 311553
rect 43594 283729 43650 283744
rect 42074 283725 42130 283729
rect 41989 283723 42193 283725
rect 41989 283721 42074 283723
rect 41982 283717 42074 283721
rect 41970 283667 42074 283717
rect 42130 283667 42193 283723
rect 41970 283661 42193 283667
rect 43594 283723 43653 283729
rect 43594 283667 43597 283723
rect 43594 283661 43653 283667
rect 41713 283017 42193 283073
rect 42074 281881 42130 281885
rect 41989 281879 42193 281881
rect 41989 281877 42074 281879
rect 41980 281823 42074 281877
rect 42130 281823 42193 281879
rect 41980 281821 42193 281823
rect 42074 281817 42130 281821
rect 41713 281177 42193 281233
rect 41713 280533 42193 280589
rect 41713 279337 42193 279393
rect 41713 278693 42193 278749
rect 41713 278141 42193 278197
rect 41713 277497 42193 277553
rect 41713 276853 42193 276909
rect 41713 276301 42193 276357
rect 42074 275713 42130 275717
rect 41851 275711 42193 275713
rect 41851 275657 42074 275711
rect 41880 275655 42074 275657
rect 42130 275655 42193 275711
rect 41880 275653 42193 275655
rect 43594 275711 43650 283661
rect 42074 275649 42130 275653
rect 43594 275649 43650 275655
rect 43706 275075 43745 313881
rect 43912 281885 43962 325017
rect 44012 314595 44062 357727
rect 44112 317633 44162 360765
rect 671166 335037 671216 380169
rect 671266 338073 671316 383205
rect 671366 372785 671416 549917
rect 671576 383917 671614 556725
rect 673258 556149 673314 556168
rect 673251 556143 673314 556149
rect 673307 556087 673314 556143
rect 675407 556087 675419 556143
rect 675475 556087 675490 556143
rect 673251 556081 673314 556087
rect 673258 548135 673314 556081
rect 675407 555443 675887 555499
rect 675407 554891 675887 554947
rect 675407 554247 675887 554303
rect 675407 553603 675887 553659
rect 675407 553051 675887 553107
rect 675407 552407 675887 552463
rect 675407 551211 675887 551267
rect 675407 550567 675887 550623
rect 675407 549923 675434 549979
rect 675490 549923 675513 549979
rect 675407 548727 675887 548783
rect 675505 548139 675557 548141
rect 673310 548083 673314 548135
rect 675425 548135 675580 548139
rect 675425 548083 675505 548135
rect 675557 548083 675580 548135
rect 673258 548077 673314 548083
rect 675505 548077 675557 548083
rect 675407 386247 675887 386303
rect 675407 385695 675887 385751
rect 675407 385051 675887 385107
rect 675407 384407 675887 384463
rect 671570 383911 671626 383917
rect 675407 383855 675426 383911
rect 675482 383855 675517 383911
rect 671570 383849 671626 383855
rect 671576 379593 671614 383849
rect 675407 383211 675465 383267
rect 675521 383211 675591 383267
rect 675407 382567 675887 382623
rect 675407 382015 675887 382071
rect 675407 381371 675887 381427
rect 675407 380727 675887 380783
rect 675407 380175 675437 380231
rect 675493 380175 675566 380231
rect 671576 379587 671637 379593
rect 671576 379531 671581 379587
rect 675407 379531 675471 379587
rect 675527 379531 675573 379587
rect 671576 379525 671637 379531
rect 671366 372779 671426 372785
rect 671366 372723 671370 372779
rect 671366 372717 671426 372723
rect 671266 338067 671328 338073
rect 671266 338011 671272 338067
rect 671266 338005 671328 338011
rect 671161 335031 671221 335037
rect 671161 334975 671165 335031
rect 671161 334969 671221 334975
rect 44111 317627 44167 317633
rect 44111 317565 44167 317571
rect 44006 314589 44062 314595
rect 44006 314527 44062 314533
rect 43904 281879 43962 281885
rect 43960 281823 43962 281879
rect 43904 281817 43962 281823
rect 42074 275069 42130 275075
rect 43697 275069 43753 275075
rect 42031 275013 42074 275069
rect 42130 275013 42193 275069
rect 42031 275011 42193 275013
rect 42074 275007 42130 275011
rect 43697 275007 43753 275013
rect 42074 274427 42130 274433
rect 42029 274371 42074 274427
rect 42130 274371 42193 274427
rect 42029 274369 42193 274371
rect 42074 274365 42130 274369
rect 41713 273817 42193 273873
rect 41713 273173 42193 273229
rect 41713 272529 42193 272585
rect 41713 271977 42193 272033
rect 42074 271389 42130 271395
rect 42024 271333 42074 271389
rect 42130 271333 42193 271389
rect 42074 271327 42130 271333
rect 43706 270749 43745 275007
rect 42074 270745 42130 270749
rect 42008 270743 42193 270745
rect 42008 270689 42074 270743
rect 42017 270687 42074 270689
rect 42130 270687 42193 270743
rect 43693 270743 43749 270749
rect 42074 270681 42130 270687
rect 43693 270681 43749 270687
rect 41713 270137 42193 270193
rect 41713 269493 42193 269549
rect 41713 268849 42193 268905
rect 41713 268297 42193 268353
rect 43594 240529 43650 240544
rect 42074 240525 42130 240529
rect 41989 240523 42193 240525
rect 41989 240521 42074 240523
rect 41982 240517 42074 240521
rect 41970 240467 42074 240517
rect 42130 240467 42193 240523
rect 41970 240461 42193 240467
rect 43594 240523 43653 240529
rect 43594 240467 43597 240523
rect 43594 240461 43653 240467
rect 41713 239817 42193 239873
rect 42074 238681 42130 238685
rect 41989 238679 42193 238681
rect 41989 238677 42074 238679
rect 41980 238623 42074 238677
rect 42130 238623 42193 238679
rect 41980 238621 42193 238623
rect 42074 238617 42130 238621
rect 41713 237977 42193 238033
rect 41713 236137 42193 236193
rect 41713 234941 42193 234997
rect 41713 234297 42193 234353
rect 41713 233653 42193 233709
rect 41713 233101 42193 233157
rect 42074 232513 42130 232517
rect 41851 232511 42193 232513
rect 41851 232457 42074 232511
rect 41880 232455 42074 232457
rect 42130 232455 42193 232511
rect 41880 232453 42193 232455
rect 43594 232511 43650 240461
rect 42074 232449 42130 232453
rect 43594 232449 43650 232455
rect 43706 231875 43745 270681
rect 43912 238685 43962 281817
rect 44012 271395 44062 314527
rect 44112 274433 44162 317565
rect 671166 290037 671216 334969
rect 671266 293073 671316 338005
rect 671366 327585 671416 372717
rect 671576 338717 671614 379525
rect 673658 378949 673714 378968
rect 673651 378943 673714 378949
rect 673707 378887 673714 378943
rect 675407 378887 675419 378943
rect 675475 378887 675490 378943
rect 673651 378881 673714 378887
rect 673658 370935 673714 378881
rect 675407 378243 675887 378299
rect 675407 377691 675887 377747
rect 675407 377047 675887 377103
rect 675407 376403 675887 376459
rect 675407 375207 675887 375263
rect 675407 373367 675887 373423
rect 675407 372723 675434 372779
rect 675490 372723 675513 372779
rect 675407 371527 675887 371583
rect 675505 370939 675557 370941
rect 673710 370883 673714 370935
rect 675425 370935 675580 370939
rect 675425 370883 675505 370935
rect 675557 370883 675580 370935
rect 673658 370877 673714 370883
rect 675505 370877 675557 370883
rect 675407 341047 675887 341103
rect 675407 340495 675887 340551
rect 675407 339851 675887 339907
rect 675407 339207 675887 339263
rect 671570 338711 671626 338717
rect 675407 338655 675426 338711
rect 675482 338655 675517 338711
rect 671570 338649 671626 338655
rect 671576 334393 671614 338649
rect 675407 338011 675465 338067
rect 675521 338011 675591 338067
rect 675407 337367 675887 337423
rect 675407 336815 675887 336871
rect 675407 336171 675887 336227
rect 675407 335527 675887 335583
rect 675407 334975 675437 335031
rect 675493 334975 675566 335031
rect 671576 334387 671637 334393
rect 671576 334331 671581 334387
rect 675407 334331 675471 334387
rect 675527 334331 675573 334387
rect 671576 334325 671637 334331
rect 671366 327579 671426 327585
rect 671366 327523 671370 327579
rect 671366 327517 671426 327523
rect 671266 293067 671328 293073
rect 671266 293011 671272 293067
rect 671266 293005 671328 293011
rect 671161 290031 671221 290037
rect 671161 289975 671165 290031
rect 671161 289969 671221 289975
rect 44111 274427 44167 274433
rect 44111 274365 44167 274371
rect 44006 271389 44062 271395
rect 44006 271327 44062 271333
rect 43904 238679 43962 238685
rect 43960 238623 43962 238679
rect 43904 238617 43962 238623
rect 42074 231869 42130 231875
rect 43697 231869 43753 231875
rect 42031 231813 42074 231869
rect 42130 231813 42193 231869
rect 42031 231811 42193 231813
rect 42074 231807 42130 231811
rect 43697 231807 43753 231813
rect 42074 231227 42130 231233
rect 42029 231171 42074 231227
rect 42130 231171 42193 231227
rect 42029 231169 42193 231171
rect 42074 231165 42130 231169
rect 41713 230617 42193 230673
rect 41713 229973 42193 230029
rect 41713 229329 42193 229385
rect 41713 228777 42193 228833
rect 42074 228189 42130 228195
rect 42024 228133 42074 228189
rect 42130 228133 42193 228189
rect 42074 228127 42130 228133
rect 43706 227549 43745 231807
rect 42074 227543 42130 227549
rect 43693 227543 43749 227549
rect 42017 227487 42074 227543
rect 42130 227487 42193 227543
rect 42074 227481 42130 227487
rect 43693 227481 43749 227487
rect 41713 226937 42193 226993
rect 41713 226293 42193 226349
rect 41713 225649 42193 225705
rect 41713 225097 42193 225153
rect 43594 197329 43650 197344
rect 42074 197325 42130 197329
rect 41989 197323 42193 197325
rect 41989 197321 42074 197323
rect 41982 197267 42074 197321
rect 42130 197267 42193 197323
rect 41982 197265 42193 197267
rect 43594 197323 43653 197329
rect 43594 197267 43597 197323
rect 42074 197261 42130 197265
rect 43594 197261 43653 197267
rect 41713 196617 42193 196673
rect 42074 195481 42130 195485
rect 41989 195479 42193 195481
rect 41989 195423 42074 195479
rect 42130 195423 42193 195479
rect 41989 195421 42193 195423
rect 42074 195417 42130 195421
rect 41713 194777 42193 194833
rect 41713 192937 42193 192993
rect 41713 191741 42193 191797
rect 41713 191097 42193 191153
rect 41713 190453 42193 190509
rect 41713 189901 42193 189957
rect 42074 189311 42130 189317
rect 43594 189311 43650 197261
rect 41987 189309 42074 189311
rect 41880 189255 42074 189309
rect 42130 189255 42193 189311
rect 41880 189253 42193 189255
rect 42074 189249 42130 189253
rect 43594 189249 43650 189255
rect 43706 188675 43745 227481
rect 43912 195485 43962 238617
rect 44012 228195 44062 271327
rect 44112 231233 44162 274365
rect 671166 245037 671216 289969
rect 671266 248073 671316 293005
rect 671366 282585 671416 327517
rect 671576 293717 671614 334325
rect 673658 333749 673714 333768
rect 673651 333743 673714 333749
rect 673707 333687 673714 333743
rect 675407 333687 675419 333743
rect 675475 333687 675490 333743
rect 673651 333681 673714 333687
rect 673658 325735 673714 333681
rect 675407 333043 675887 333099
rect 675407 332491 675887 332547
rect 675407 331847 675887 331903
rect 675407 331203 675887 331259
rect 675407 330007 675887 330063
rect 675407 328167 675887 328223
rect 675407 327523 675434 327579
rect 675490 327523 675513 327579
rect 675407 326327 675887 326383
rect 675505 325739 675557 325741
rect 673710 325683 673714 325735
rect 675425 325735 675580 325739
rect 675425 325683 675505 325735
rect 675557 325683 675580 325735
rect 673658 325677 673714 325683
rect 675505 325677 675557 325683
rect 675407 296047 675887 296103
rect 675407 295495 675887 295551
rect 675407 294851 675887 294907
rect 675407 294207 675887 294263
rect 671570 293711 671626 293717
rect 675407 293655 675426 293711
rect 675482 293655 675517 293711
rect 671570 293649 671626 293655
rect 671576 289393 671614 293649
rect 675407 293011 675465 293067
rect 675521 293011 675591 293067
rect 675407 292367 675887 292423
rect 675407 291815 675887 291871
rect 675407 291171 675887 291227
rect 675407 290527 675887 290583
rect 675407 289975 675437 290031
rect 675493 289975 675566 290031
rect 671576 289387 671637 289393
rect 671576 289331 671581 289387
rect 675407 289331 675471 289387
rect 675527 289331 675573 289387
rect 671576 289325 671637 289331
rect 671366 282579 671426 282585
rect 671366 282523 671370 282579
rect 671366 282517 671426 282523
rect 671266 248067 671328 248073
rect 671266 248011 671272 248067
rect 671266 248005 671328 248011
rect 671161 245031 671221 245037
rect 671161 244975 671165 245031
rect 671161 244969 671221 244975
rect 44111 231227 44167 231233
rect 44111 231165 44167 231171
rect 44006 228189 44062 228195
rect 44006 228127 44062 228133
rect 43904 195479 43962 195485
rect 43960 195423 43962 195479
rect 43904 195417 43962 195423
rect 42074 188669 42130 188675
rect 43697 188669 43753 188675
rect 41987 188667 42074 188669
rect 41880 188613 42074 188667
rect 42130 188613 42193 188669
rect 41880 188611 42193 188613
rect 42074 188607 42130 188611
rect 43697 188607 43753 188613
rect 42074 188027 42130 188033
rect 41987 187971 42074 188027
rect 42130 187971 42193 188027
rect 42074 187965 42130 187971
rect 41713 187417 42193 187473
rect 41713 186773 42193 186829
rect 41713 186129 42193 186185
rect 41713 185577 42193 185633
rect 42074 184989 42130 184995
rect 42074 184927 42130 184933
rect 43706 184345 43745 188607
rect 42137 184289 43745 184345
rect 41713 183737 42193 183793
rect 41713 183093 42193 183149
rect 41713 182449 42193 182505
rect 41713 181897 42193 181953
rect 43706 181284 43745 184289
rect 43699 181278 43751 181284
rect 43699 181220 43751 181226
rect 43912 181086 43962 195417
rect 44012 184995 44062 228127
rect 44112 188033 44162 231165
rect 671166 199837 671216 244969
rect 671266 202873 671316 248005
rect 671366 237585 671416 282517
rect 671576 248717 671614 289325
rect 673658 288749 673714 288768
rect 673651 288743 673714 288749
rect 673707 288687 673714 288743
rect 675407 288687 675419 288743
rect 675475 288687 675490 288743
rect 673651 288681 673714 288687
rect 673658 280735 673714 288681
rect 675407 288043 675887 288099
rect 675407 287491 675887 287547
rect 675407 286847 675887 286903
rect 675407 286203 675887 286259
rect 675407 285007 675887 285063
rect 675407 283167 675887 283223
rect 675407 282523 675434 282579
rect 675490 282523 675513 282579
rect 675407 281327 675887 281383
rect 675505 280739 675557 280741
rect 673710 280683 673714 280735
rect 675425 280735 675580 280739
rect 675425 280683 675505 280735
rect 675557 280683 675580 280735
rect 673658 280677 673714 280683
rect 675505 280677 675557 280683
rect 675407 251047 675887 251103
rect 675407 250495 675887 250551
rect 675407 249851 675887 249907
rect 675407 249207 675887 249263
rect 671570 248711 671626 248717
rect 675407 248655 675426 248711
rect 675482 248655 675517 248711
rect 671570 248649 671626 248655
rect 671576 244393 671614 248649
rect 675407 248011 675465 248067
rect 675521 248011 675591 248067
rect 675407 247367 675887 247423
rect 675407 246815 675887 246871
rect 675407 246171 675887 246227
rect 675407 245527 675887 245583
rect 675407 244975 675437 245031
rect 675493 244975 675566 245031
rect 671576 244387 671637 244393
rect 671576 244331 671581 244387
rect 675407 244331 675471 244387
rect 675527 244331 675573 244387
rect 671576 244325 671637 244331
rect 671366 237579 671426 237585
rect 671366 237523 671370 237579
rect 671366 237517 671426 237523
rect 671266 202867 671328 202873
rect 671266 202811 671272 202867
rect 671266 202805 671328 202811
rect 671161 199831 671221 199837
rect 671161 199775 671165 199831
rect 671161 199769 671221 199775
rect 44111 188027 44167 188033
rect 44111 187965 44167 187971
rect 44006 184989 44062 184995
rect 44006 184927 44062 184933
rect 43910 181080 43962 181086
rect 43910 181022 43962 181028
rect 43912 181018 43962 181022
rect 44012 180986 44062 184927
rect 44012 180980 44064 180986
rect 44012 180922 44064 180928
rect 44012 180907 44062 180922
rect 44112 180886 44162 187965
rect 44110 180880 44162 180886
rect 44110 180822 44162 180828
rect 44112 180808 44162 180822
rect 671166 154837 671216 199769
rect 671266 157873 671316 202805
rect 671366 192385 671416 237517
rect 671576 203517 671614 244325
rect 673658 243749 673714 243768
rect 673651 243743 673714 243749
rect 673707 243687 673714 243743
rect 675407 243687 675419 243743
rect 675475 243687 675490 243743
rect 673651 243681 673714 243687
rect 673658 235735 673714 243681
rect 675407 243043 675887 243099
rect 675407 242491 675887 242547
rect 675407 241847 675887 241903
rect 675407 241203 675887 241259
rect 675407 240007 675887 240063
rect 675407 238167 675887 238223
rect 675407 237523 675434 237579
rect 675490 237523 675513 237579
rect 675407 236327 675887 236383
rect 675505 235739 675557 235741
rect 673710 235683 673714 235735
rect 675425 235735 675580 235739
rect 675425 235683 675505 235735
rect 675557 235683 675580 235735
rect 673658 235677 673714 235683
rect 675505 235677 675557 235683
rect 675407 205847 675887 205903
rect 675407 205295 675887 205351
rect 675407 204651 675887 204707
rect 675407 204007 675887 204063
rect 671570 203511 671626 203517
rect 675407 203455 675426 203511
rect 675482 203455 675517 203511
rect 671570 203449 671626 203455
rect 671576 199193 671614 203449
rect 675407 202811 675465 202867
rect 675521 202811 675591 202867
rect 675407 202167 675887 202223
rect 675407 201615 675887 201671
rect 675407 200971 675887 201027
rect 675407 200327 675887 200383
rect 675407 199775 675437 199831
rect 675493 199775 675566 199831
rect 671576 199187 671637 199193
rect 671576 199131 671581 199187
rect 675407 199131 675471 199187
rect 675527 199131 675573 199187
rect 671576 199125 671637 199131
rect 671366 192379 671426 192385
rect 671366 192323 671370 192379
rect 671366 192317 671426 192323
rect 671266 157867 671328 157873
rect 671266 157811 671272 157867
rect 671266 157805 671328 157811
rect 671161 154831 671221 154837
rect 671161 154775 671165 154831
rect 671161 154769 671221 154775
rect 42414 112734 42519 112755
rect 42414 112371 42428 112734
rect 42510 112371 42519 112734
rect 42414 112354 42519 112371
rect 671166 109637 671216 154769
rect 671266 112673 671316 157805
rect 671366 147385 671416 192317
rect 671576 158517 671614 199125
rect 673658 198549 673714 198568
rect 673651 198543 673714 198549
rect 673707 198487 673714 198543
rect 675407 198487 675419 198543
rect 675475 198487 675490 198543
rect 673651 198481 673714 198487
rect 673658 190535 673714 198481
rect 675407 197843 675887 197899
rect 675407 197291 675887 197347
rect 675407 196647 675887 196703
rect 675407 196003 675887 196059
rect 675407 194807 675887 194863
rect 675407 192967 675887 193023
rect 675407 192323 675434 192379
rect 675490 192323 675513 192379
rect 675407 191127 675887 191183
rect 675505 190539 675557 190541
rect 673710 190483 673714 190535
rect 675425 190535 675580 190539
rect 675425 190483 675505 190535
rect 675557 190483 675580 190535
rect 673658 190477 673714 190483
rect 675505 190477 675557 190483
rect 675407 160847 675887 160903
rect 675407 160295 675887 160351
rect 675407 159651 675887 159707
rect 675407 159007 675887 159063
rect 671570 158511 671626 158517
rect 675407 158455 675426 158511
rect 675482 158455 675517 158511
rect 671570 158449 671626 158455
rect 671576 154193 671614 158449
rect 675407 157811 675465 157867
rect 675521 157811 675591 157867
rect 675407 157167 675887 157223
rect 675407 156615 675887 156671
rect 675407 155971 675887 156027
rect 675407 155327 675887 155383
rect 675407 154775 675437 154831
rect 675493 154775 675566 154831
rect 671576 154187 671637 154193
rect 671576 154131 671581 154187
rect 675407 154131 675471 154187
rect 675527 154131 675573 154187
rect 671576 154125 671637 154131
rect 671366 147379 671426 147385
rect 671366 147323 671370 147379
rect 671366 147317 671426 147323
rect 671266 112667 671328 112673
rect 671266 112611 671272 112667
rect 671266 112605 671328 112611
rect 671161 109631 671221 109637
rect 671161 109575 671165 109631
rect 671161 109569 671221 109575
rect 42210 69967 42296 69987
rect 42210 69441 42216 69967
rect 42289 69441 42296 69967
rect 42210 69425 42296 69441
rect 571321 42961 571764 42984
rect 464007 42760 464063 42768
rect 464006 42754 464063 42760
rect 470169 42758 470225 42760
rect 470169 42754 470227 42758
rect 411046 42744 411105 42750
rect 409207 42659 409263 42672
rect 409207 42653 409266 42659
rect 409207 42597 409210 42653
rect 409207 42591 409266 42597
rect 295283 42555 295339 42568
rect 42315 42412 42321 42544
rect 42374 42464 42381 42544
rect 295283 42503 295286 42555
rect 295338 42503 295339 42555
rect 42582 42464 42734 42470
rect 42374 42412 42582 42464
rect 42582 42406 42734 42412
rect 140996 42464 141048 42470
rect 90863 42239 91094 42245
rect 90863 42183 90872 42239
rect 91085 42183 91094 42239
rect 90863 42174 91094 42183
rect 133004 40234 133052 40238
rect 132998 40228 133052 40234
rect 133050 40176 133052 40228
rect 132998 40170 133052 40176
rect 133004 39978 133052 40170
rect 140996 39942 141048 42412
rect 142570 42464 142622 42500
rect 143075 42469 143127 42470
rect 142570 40122 142622 42412
rect 143068 42464 143128 42469
rect 143068 42412 143075 42464
rect 143127 42412 143128 42464
rect 142564 40070 142570 40122
rect 142622 40070 142628 40122
rect 143068 39940 143128 42412
rect 143429 42464 143485 42484
rect 143429 42412 143432 42464
rect 143484 42412 143485 42464
rect 143429 40320 143485 42412
rect 144601 42464 144655 42483
rect 144601 42412 144602 42464
rect 144654 42412 144655 42464
rect 143420 40264 143429 40320
rect 143485 40264 143494 40320
rect 143925 40228 143977 40234
rect 143925 40170 143977 40176
rect 143932 39980 143970 40170
rect 144601 39971 144655 42412
rect 195975 42341 196031 42368
rect 195975 42335 196034 42341
rect 195975 42283 195982 42335
rect 195975 42277 196034 42283
rect 145853 42136 145907 42142
rect 145091 41861 145143 41867
rect 145091 39706 145143 41809
rect 145853 39981 145907 42082
rect 186686 41945 186738 41951
rect 186686 41887 186738 41893
rect 187327 41713 187383 42193
rect 188526 42135 188578 42141
rect 188526 42077 188578 42083
rect 192846 42135 192898 42141
rect 192846 42077 192898 42083
rect 189168 42035 189220 42041
rect 189168 41977 189220 41983
rect 191010 42035 191062 42041
rect 191010 41977 191062 41983
rect 192200 42035 192252 42041
rect 192200 41977 192252 41983
rect 193500 42035 193552 42041
rect 193500 41977 193552 41983
rect 194043 41713 194099 42193
rect 194690 41945 194742 41950
rect 194690 41887 194742 41893
rect 195331 41887 195387 42199
rect 195975 42136 196031 42277
rect 199011 42241 199067 42264
rect 199011 42235 199074 42241
rect 199011 42183 199022 42235
rect 199011 42177 199074 42183
rect 199011 42130 199067 42177
rect 196524 42035 196576 42041
rect 196524 41977 196576 41983
rect 197176 42035 197228 42041
rect 197176 41977 197228 41983
rect 197816 42035 197868 42041
rect 197816 41977 197868 41983
rect 198374 42035 198426 42041
rect 198374 41977 198426 41983
rect 195331 41825 195387 41831
rect 199655 41887 199711 42198
rect 201492 42135 201544 42141
rect 295283 42129 295339 42503
rect 303287 42555 303343 42568
rect 303287 42503 303290 42555
rect 303342 42503 303343 42555
rect 297123 42135 297179 42179
rect 201492 42077 201544 42083
rect 297123 42083 297126 42135
rect 297178 42083 297179 42135
rect 299607 42132 299663 42138
rect 297123 42056 297179 42083
rect 200214 42035 200266 42041
rect 200214 41977 200266 41983
rect 200852 42035 200904 42041
rect 200852 41977 200904 41983
rect 253613 42034 253827 42043
rect 253613 41962 253622 42034
rect 253815 41962 253827 42034
rect 297767 42035 297823 42086
rect 297767 41983 297768 42035
rect 297820 41983 297823 42035
rect 297767 41963 297823 41983
rect 253613 41951 253827 41962
rect 299607 41929 299663 42076
rect 300803 42041 300859 42075
rect 300800 42035 300859 42041
rect 302091 42041 302147 42081
rect 300852 41983 300859 42035
rect 300800 41977 300859 41983
rect 300803 41952 300859 41977
rect 301447 42033 301503 42039
rect 301447 41905 301503 41977
rect 302091 42035 302152 42041
rect 302091 41983 302100 42035
rect 302091 41977 302152 41983
rect 302091 41958 302147 41977
rect 199655 41825 199711 41831
rect 302643 41713 302699 42193
rect 303287 42137 303343 42503
rect 350083 42555 350139 42568
rect 350083 42503 350086 42555
rect 350138 42503 350139 42555
rect 304575 42341 304631 42363
rect 304575 42335 304634 42341
rect 304575 42283 304582 42335
rect 304575 42277 304634 42283
rect 304575 42113 304631 42277
rect 307611 42242 307668 42246
rect 307610 42235 307668 42242
rect 305771 42130 305827 42136
rect 305127 42041 305183 42064
rect 305124 42035 305183 42041
rect 305176 41983 305183 42035
rect 305124 41977 305183 41983
rect 305127 41960 305183 41977
rect 303931 41871 303987 41899
rect 305771 41894 305827 42074
rect 306415 42035 306471 42064
rect 306415 41983 306416 42035
rect 306468 41983 306471 42035
rect 306415 41960 306471 41983
rect 303931 41800 303987 41815
rect 306967 41713 307023 42193
rect 307610 42183 307616 42235
rect 307610 42176 307668 42183
rect 307611 42161 307667 42176
rect 308807 42041 308863 42056
rect 308807 42035 308866 42041
rect 308807 41983 308814 42035
rect 308807 41977 308866 41983
rect 309451 42035 309507 42072
rect 309451 41983 309452 42035
rect 309504 41983 309507 42035
rect 308807 41952 308863 41977
rect 309451 41968 309507 41983
rect 308255 41873 308311 41907
rect 308255 41803 308311 41817
rect 310095 41713 310151 42193
rect 350083 42129 350139 42503
rect 358087 42555 358143 42568
rect 358087 42503 358090 42555
rect 358142 42503 358143 42555
rect 351923 42135 351979 42179
rect 351923 42083 351926 42135
rect 351978 42083 351979 42135
rect 354407 42134 354463 42140
rect 351923 42056 351979 42083
rect 352567 42035 352623 42086
rect 352567 41983 352568 42035
rect 352620 41983 352623 42035
rect 352567 41963 352623 41983
rect 354407 41934 354463 42078
rect 355603 42041 355659 42075
rect 355600 42035 355659 42041
rect 356891 42041 356947 42081
rect 355652 41983 355659 42035
rect 355600 41977 355659 41983
rect 355603 41952 355659 41977
rect 356247 42030 356303 42036
rect 356247 41915 356303 41974
rect 356891 42035 356952 42041
rect 356891 41983 356900 42035
rect 356891 41977 356952 41983
rect 356891 41958 356947 41977
rect 357443 41713 357499 42193
rect 358087 42137 358143 42503
rect 404883 42555 404939 42568
rect 404883 42503 404886 42555
rect 404938 42503 404939 42555
rect 359375 42341 359431 42363
rect 359375 42335 359434 42341
rect 359375 42283 359382 42335
rect 359375 42277 359434 42283
rect 359375 42120 359431 42277
rect 362411 42242 362468 42246
rect 362410 42235 362468 42242
rect 360571 42139 360627 42145
rect 359927 42041 359983 42064
rect 359924 42035 359983 42041
rect 359976 41983 359983 42035
rect 359924 41977 359983 41983
rect 359927 41960 359983 41977
rect 360571 41913 360627 42083
rect 361215 42035 361271 42064
rect 361215 41983 361216 42035
rect 361268 41983 361271 42035
rect 361215 41960 361271 41983
rect 358731 41871 358787 41891
rect 358731 41800 358787 41815
rect 361767 41713 361823 42193
rect 362410 42183 362416 42235
rect 362410 42176 362468 42183
rect 362411 42161 362467 42176
rect 363607 42041 363663 42056
rect 363607 42035 363666 42041
rect 363607 41983 363614 42035
rect 363607 41977 363666 41983
rect 364251 42035 364307 42072
rect 364251 41983 364252 42035
rect 364304 41983 364307 42035
rect 363607 41952 363663 41977
rect 364251 41968 364307 41983
rect 363055 41873 363111 41907
rect 363055 41803 363111 41817
rect 364895 41713 364951 42193
rect 404883 42127 404939 42503
rect 405527 41713 405583 42193
rect 406726 42135 406778 42141
rect 406726 42077 406778 42083
rect 407368 42035 407420 42041
rect 407368 41977 407420 41983
rect 409207 41944 409263 42591
rect 410400 42035 410452 42041
rect 411046 42031 411105 42685
rect 419695 42748 419751 42754
rect 464062 42698 464063 42754
rect 467037 42698 467043 42754
rect 467099 42698 467105 42754
rect 470225 42698 470227 42754
rect 518816 42729 518844 42747
rect 464006 42692 464063 42698
rect 412243 42653 412299 42678
rect 411700 42035 411752 42041
rect 410400 41977 410452 41983
rect 411700 41977 411752 41983
rect 412243 41713 412299 42597
rect 415371 42649 415427 42667
rect 412887 42555 412943 42568
rect 412887 42503 412890 42555
rect 412942 42503 412943 42555
rect 412887 42125 412943 42503
rect 414175 42341 414231 42368
rect 414175 42335 414234 42341
rect 414175 42283 414182 42335
rect 414175 42277 414234 42283
rect 413531 41871 413587 42194
rect 414175 42136 414231 42277
rect 415371 42132 415427 42593
rect 417211 42242 417268 42246
rect 417210 42235 417268 42242
rect 414724 42035 414776 42041
rect 414724 41977 414776 41983
rect 416016 42035 416068 42041
rect 416016 41977 416068 41983
rect 413531 41809 413587 41815
rect 416567 41713 416623 42193
rect 417210 42183 417216 42235
rect 417210 42176 417268 42183
rect 417211 42130 417267 42176
rect 417855 41873 417911 42193
rect 418414 42035 418466 42041
rect 418414 41977 418466 41983
rect 419052 42035 419104 42041
rect 419052 41977 419104 41983
rect 417855 41811 417911 41817
rect 419695 41713 419751 42692
rect 459686 41945 459738 41951
rect 459686 41887 459738 41893
rect 460327 41713 460383 42193
rect 461526 42135 461578 42141
rect 464007 42120 464063 42692
rect 465847 42626 465903 42634
rect 465845 42620 465903 42626
rect 465901 42564 465903 42620
rect 465845 42558 465903 42564
rect 465847 42127 465903 42558
rect 461526 42077 461578 42083
rect 462168 42035 462220 42041
rect 462168 41977 462220 41983
rect 465200 42035 465252 42041
rect 465200 41977 465252 41983
rect 466500 42035 466552 42041
rect 466500 41977 466552 41983
rect 467043 41713 467099 42698
rect 470169 42692 470227 42698
rect 468975 42341 469031 42368
rect 468975 42335 469034 42341
rect 468975 42283 468982 42335
rect 468975 42277 469034 42283
rect 467690 41945 467742 41950
rect 467690 41887 467742 41893
rect 468331 41875 468387 42199
rect 468975 42136 469031 42277
rect 470171 42120 470227 42692
rect 518804 42723 518856 42729
rect 518804 42665 518856 42671
rect 524952 42723 525004 42729
rect 524952 42665 525004 42671
rect 474495 42620 474551 42626
rect 472011 42242 472068 42246
rect 472010 42235 472068 42242
rect 469524 42035 469576 42041
rect 469524 41977 469576 41983
rect 470816 42035 470868 42041
rect 470816 41977 470868 41983
rect 468331 41813 468387 41819
rect 471367 41713 471423 42193
rect 472010 42183 472016 42235
rect 472010 42176 472068 42183
rect 472011 42130 472067 42176
rect 472655 41876 472711 42195
rect 473214 42035 473266 42041
rect 473214 41977 473266 41983
rect 473852 42035 473904 42041
rect 473852 41977 473904 41983
rect 472655 41814 472711 41820
rect 474495 41713 474551 42564
rect 516323 42309 516379 42322
rect 516323 42257 516326 42309
rect 516378 42257 516379 42309
rect 514486 42119 514538 42125
rect 514486 42061 514538 42067
rect 515127 41713 515183 42193
rect 516323 42094 516379 42257
rect 516968 42209 517020 42215
rect 516968 42151 517020 42157
rect 518816 42016 518844 42665
rect 523775 42515 523831 42542
rect 523775 42509 523834 42515
rect 523775 42457 523782 42509
rect 523775 42451 523834 42457
rect 520000 42209 520052 42215
rect 521300 42209 521352 42215
rect 520000 42151 520052 42157
rect 520647 41713 520703 42193
rect 521300 42151 521352 42157
rect 521843 41713 521899 42193
rect 522490 42119 522542 42124
rect 522490 42061 522542 42067
rect 523131 41873 523187 42197
rect 523775 42120 523831 42451
rect 524324 42209 524376 42215
rect 524324 42151 524376 42157
rect 524964 42195 524992 42665
rect 571321 42601 571346 42961
rect 571737 42601 571764 42961
rect 571321 42583 571764 42601
rect 671166 42515 671216 109569
rect 671266 42643 671316 112605
rect 671366 102185 671416 147317
rect 671576 113317 671614 154125
rect 673658 153549 673714 153568
rect 673651 153543 673714 153549
rect 673707 153487 673714 153543
rect 675407 153487 675419 153543
rect 675475 153487 675490 153543
rect 673651 153481 673714 153487
rect 673658 145535 673714 153481
rect 675407 152843 675887 152899
rect 675407 152291 675887 152347
rect 675407 151647 675887 151703
rect 675407 151003 675887 151059
rect 675407 149807 675887 149863
rect 675407 147967 675887 148023
rect 675407 147323 675434 147379
rect 675490 147323 675513 147379
rect 675407 146127 675887 146183
rect 675505 145539 675557 145541
rect 673710 145483 673714 145535
rect 675425 145535 675580 145539
rect 675425 145483 675505 145535
rect 675557 145483 675580 145535
rect 673658 145477 673714 145483
rect 675505 145477 675557 145483
rect 675407 115647 675887 115703
rect 675407 115095 675887 115151
rect 675407 114451 675887 114507
rect 675407 113807 675887 113863
rect 671570 113311 671626 113317
rect 675420 113255 675426 113311
rect 675482 113255 675554 113311
rect 671570 113249 671626 113255
rect 671576 108993 671614 113249
rect 675459 112611 675465 112667
rect 675521 112611 675609 112667
rect 675407 111967 675887 112023
rect 675407 111415 675887 111471
rect 675407 110771 675887 110827
rect 675407 110127 675887 110183
rect 675431 109575 675437 109631
rect 675493 109575 675561 109631
rect 671576 108987 671637 108993
rect 671576 108931 671581 108987
rect 675465 108931 675471 108987
rect 675527 108931 675595 108987
rect 671576 108925 671637 108931
rect 671366 102179 671426 102185
rect 671366 102123 671370 102179
rect 671366 102117 671426 102123
rect 671266 42637 671323 42643
rect 671266 42585 671271 42637
rect 671266 42579 671323 42585
rect 671266 42570 671316 42579
rect 671166 42509 671218 42515
rect 671166 42451 671218 42457
rect 671166 42431 671216 42451
rect 526811 42416 526868 42420
rect 526810 42409 526868 42416
rect 526810 42357 526816 42409
rect 526810 42350 526868 42357
rect 525616 42209 525668 42215
rect 524964 42102 525027 42195
rect 525616 42151 525668 42157
rect 523131 41811 523187 41817
rect 524971 41713 525027 42102
rect 526167 41713 526223 42193
rect 526811 42112 526867 42350
rect 671366 42315 671416 102117
rect 671366 42309 671418 42315
rect 671366 42251 671418 42257
rect 671366 42243 671416 42251
rect 528014 42209 528066 42215
rect 527455 41871 527511 42201
rect 528014 42151 528066 42157
rect 528652 42209 528704 42215
rect 528652 42151 528704 42157
rect 527455 41809 527511 41815
rect 529295 41713 529351 42193
rect 671576 42113 671614 108925
rect 673658 108349 673714 108368
rect 673651 108343 673714 108349
rect 673707 108287 673714 108343
rect 675413 108287 675419 108343
rect 675475 108287 675602 108343
rect 673651 108281 673714 108287
rect 673658 100335 673714 108281
rect 675407 107643 675887 107699
rect 675407 107091 675887 107147
rect 675407 106447 675887 106503
rect 675407 105803 675887 105859
rect 675407 104607 675887 104663
rect 675407 102767 675887 102823
rect 675428 102123 675434 102179
rect 675490 102123 675592 102179
rect 675407 100927 675887 100983
rect 673710 100283 673714 100335
rect 673658 100277 673714 100283
rect 675505 100335 675557 100341
rect 675505 100277 675557 100283
rect 671569 42107 671621 42113
rect 671569 42049 671621 42055
<< via2 >>
rect 42428 112371 42510 112734
rect 42216 69441 42289 69967
rect 90872 42183 91085 42239
rect 143429 40264 143485 40320
rect 253622 41962 253815 42034
rect 571346 42601 571737 42961
<< metal3 >>
rect 82144 997600 87144 1014070
rect 133544 997600 138544 1014070
rect 184944 997600 189944 1014070
rect 240478 997600 254800 1000736
rect 293078 997600 307400 1000736
rect 394878 997600 409200 1000736
rect 478744 997600 483744 1014070
rect 530144 997600 535144 1014070
rect 631944 997600 636944 1014070
rect 23530 960144 40000 965144
rect 677600 956656 694070 961656
rect 678000 469900 685920 474700
rect 31680 440900 39600 445700
rect 42414 112734 42519 112755
rect 42414 112725 42428 112734
rect 39977 112380 42428 112725
rect 42414 112371 42428 112380
rect 42510 112371 42519 112734
rect 42414 112354 42519 112371
rect 42210 69967 42296 69987
rect 42210 69966 42216 69967
rect 39580 69441 42216 69966
rect 42289 69441 42296 69967
rect 42210 69425 42296 69441
rect 571321 42961 571764 42984
rect 571321 42601 571346 42961
rect 571737 42601 571764 42961
rect 571321 42583 571764 42601
rect 90866 42245 91092 42384
rect 90863 42239 91094 42245
rect 90863 42183 90872 42239
rect 91085 42183 91094 42239
rect 90863 42174 91094 42183
rect 90866 39940 91092 42174
rect 253613 42034 253827 42043
rect 253613 41962 253622 42034
rect 253815 41962 253827 42034
rect 143424 40320 143490 40325
rect 143424 40264 143429 40320
rect 143485 40264 143490 40320
rect 141667 38031 141813 39999
rect 143424 39971 143490 40264
rect 253613 39600 253827 41962
rect 571393 39973 571692 42583
<< metal4 >>
rect 679377 459800 680307 460054
rect 680587 459800 681277 459992
rect 688881 459800 688947 474800
rect 7 455645 4843 456093
rect 28653 440800 28719 455800
rect 32933 455546 33623 455800
rect 36323 455607 37013 455799
rect 37293 455546 38223 455800
rect 38503 455546 39593 455800
rect 41663 44090 43230 67615
rect 41663 42523 78849 44090
rect 132600 36323 132792 37013
rect 132600 30762 132868 31674
rect 132600 28653 147600 28719
<< metal5 >>
rect 78610 1018624 90778 1030788
rect 130010 1018624 142178 1030788
rect 181410 1018624 193578 1030788
rect 231810 1018624 243978 1030788
rect 284410 1018624 296578 1030788
rect 334810 1018624 346978 1030788
rect 386210 1018624 398378 1030788
rect 475210 1018624 487378 1030788
rect 526610 1018624 538778 1030788
rect 577010 1018624 589178 1030788
rect 628410 1018624 640578 1030788
rect 6811 956610 18975 968778
rect 698624 953022 710788 965190
rect 6167 914054 19619 924934
rect 697980 909666 711432 920546
rect 6811 871210 18975 883378
rect 698512 863640 711002 876160
rect 6811 829010 18975 841178
rect 698624 819822 710788 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710788 517390
rect 6811 484410 18975 496578
rect 697980 461866 711432 472746
rect 6167 442854 19619 453734
rect 698624 417022 710788 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 28653 125200 30453 125266
rect 31983 125200 32632 125266
rect 36343 125007 36993 125327
rect 6811 111610 18975 123778
rect 698512 101240 711002 113760
rect 6167 70054 19619 80934
rect 80222 6811 92390 18975
rect 136713 7143 144149 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19619
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18975
rect 624222 6811 636390 18975
use sky130_ef_io__corner_pad  mgmt_corner\[0\] $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1625505168
transform -1 0 40000 0 -1 40800
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_20um  FILLER_352 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1625505168
transform 0 -1 39593 1 0 40800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_148
timestamp 1625505168
transform -1 0 44000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_3 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1625505168
transform -1 0 59400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_2
timestamp 1625505168
transform -1 0 55400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_1
timestamp 1625505168
transform -1 0 51400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_149 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1625505168
transform -1 0 46000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_150 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1625505168
transform -1 0 47000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_152 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1625505168
transform -1 0 47400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_151
timestamp 1625505168
transform -1 0 47200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_6
timestamp 1625505168
transform -1 0 71400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_5
timestamp 1625505168
transform -1 0 67400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_4
timestamp 1625505168
transform -1 0 63400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_159
timestamp 1625505168
transform -1 0 75400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  mgmt_vssa_hvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1625505168
transform -1 0 93800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_160
timestamp 1625505168
transform -1 0 77400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_161
timestamp 1625505168
transform -1 0 78400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_163
timestamp 1625505168
transform -1 0 78800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_162
timestamp 1625505168
transform -1 0 78600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_165
timestamp 1625505168
transform -1 0 97800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_166
timestamp 1625505168
transform -1 0 99800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_167
timestamp 1625505168
transform -1 0 100800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_7
timestamp 1625505168
transform -1 0 105200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_169
timestamp 1625505168
transform -1 0 101200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_168
timestamp 1625505168
transform -1 0 101000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_8
timestamp 1625505168
transform -1 0 109200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_9
timestamp 1625505168
transform -1 0 113200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_10
timestamp 1625505168
transform -1 0 117200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_11
timestamp 1625505168
transform -1 0 121200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_12
timestamp 1625505168
transform -1 0 125200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_176
timestamp 1625505168
transform -1 0 129200 0 -1 39593
box 0 0 4000 39593
use sky130_fd_io__top_xres4v2  resetb_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1625505168
transform -1 0 147600 0 -1 40000
box -103 0 15124 40000
use sky130_ef_io__com_bus_slice_10um  FILLER_177
timestamp 1625505168
transform -1 0 131200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_178
timestamp 1625505168
transform -1 0 132200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_180
timestamp 1625505168
transform -1 0 132600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_179
timestamp 1625505168
transform -1 0 132400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_13
timestamp 1625505168
transform -1 0 159000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_183
timestamp 1625505168
transform -1 0 153600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_184
timestamp 1625505168
transform -1 0 154600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_186
timestamp 1625505168
transform -1 0 155000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_185
timestamp 1625505168
transform -1 0 154800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_182
timestamp 1625505168
transform -1 0 151600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_16
timestamp 1625505168
transform -1 0 171000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_15
timestamp 1625505168
transform -1 0 167000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_14
timestamp 1625505168
transform -1 0 163000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_18
timestamp 1625505168
transform -1 0 179000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_17
timestamp 1625505168
transform -1 0 175000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_194
timestamp 1625505168
transform -1 0 185000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_193
timestamp 1625505168
transform -1 0 183000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  clock_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1625505168
transform -1 0 202400 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_195
timestamp 1625505168
transform -1 0 186000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_197
timestamp 1625505168
transform -1 0 186400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_196
timestamp 1625505168
transform -1 0 186200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_19
timestamp 1625505168
transform -1 0 213800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_200
timestamp 1625505168
transform -1 0 208400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_201
timestamp 1625505168
transform -1 0 209400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_203
timestamp 1625505168
transform -1 0 209800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_202
timestamp 1625505168
transform -1 0 209600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_199
timestamp 1625505168
transform -1 0 206400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_23
timestamp 1625505168
transform -1 0 229800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_22
timestamp 1625505168
transform -1 0 225800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_21
timestamp 1625505168
transform -1 0 221800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_20
timestamp 1625505168
transform -1 0 217800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_24
timestamp 1625505168
transform -1 0 233800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__vssd_lvc_clamped_pad  mgmt_vssd_lvclmap_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1625505168
transform -1 0 256200 0 -1 39593
box 0 -2107 17239 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_211
timestamp 1625505168
transform -1 0 239800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_212
timestamp 1625505168
transform -1 0 240800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_214
timestamp 1625505168
transform -1 0 241200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_213
timestamp 1625505168
transform -1 0 241000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_210
timestamp 1625505168
transform -1 0 237800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_26
timestamp 1625505168
transform -1 0 271600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_25
timestamp 1625505168
transform -1 0 267600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_217
timestamp 1625505168
transform -1 0 262200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_218
timestamp 1625505168
transform -1 0 263200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_220
timestamp 1625505168
transform -1 0 263600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_219
timestamp 1625505168
transform -1 0 263400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_216
timestamp 1625505168
transform -1 0 260200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_30
timestamp 1625505168
transform -1 0 287600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_29
timestamp 1625505168
transform -1 0 283600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_28
timestamp 1625505168
transform -1 0 279600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_27
timestamp 1625505168
transform -1 0 275600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_csb_pad
timestamp 1625505168
transform -1 0 311000 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_228
timestamp 1625505168
transform -1 0 293600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_229
timestamp 1625505168
transform -1 0 294600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_231
timestamp 1625505168
transform -1 0 295000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_230
timestamp 1625505168
transform -1 0 294800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_227
timestamp 1625505168
transform -1 0 291600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_233
timestamp 1625505168
transform -1 0 315000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_234
timestamp 1625505168
transform -1 0 317000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_31
timestamp 1625505168
transform -1 0 322400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_235
timestamp 1625505168
transform -1 0 318000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_237
timestamp 1625505168
transform -1 0 318400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_236
timestamp 1625505168
transform -1 0 318200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_32
timestamp 1625505168
transform -1 0 326400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_33
timestamp 1625505168
transform -1 0 330400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_34
timestamp 1625505168
transform -1 0 334400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_35
timestamp 1625505168
transform -1 0 338400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_36
timestamp 1625505168
transform -1 0 342400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_clk_pad
timestamp 1625505168
transform -1 0 365800 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_245
timestamp 1625505168
transform -1 0 348400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_246
timestamp 1625505168
transform -1 0 349400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_248
timestamp 1625505168
transform -1 0 349800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_247
timestamp 1625505168
transform -1 0 349600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_244
timestamp 1625505168
transform -1 0 346400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_251
timestamp 1625505168
transform -1 0 371800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_250
timestamp 1625505168
transform -1 0 369800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_38
timestamp 1625505168
transform -1 0 381200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_37
timestamp 1625505168
transform -1 0 377200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_252
timestamp 1625505168
transform -1 0 372800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_254
timestamp 1625505168
transform -1 0 373200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_253
timestamp 1625505168
transform -1 0 373000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_42
timestamp 1625505168
transform -1 0 397200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_41
timestamp 1625505168
transform -1 0 393200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_40
timestamp 1625505168
transform -1 0 389200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_39
timestamp 1625505168
transform -1 0 385200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_io0_pad
timestamp 1625505168
transform -1 0 420600 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_262
timestamp 1625505168
transform -1 0 403200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_263
timestamp 1625505168
transform -1 0 404200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_265
timestamp 1625505168
transform -1 0 404600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_264
timestamp 1625505168
transform -1 0 404400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_261
timestamp 1625505168
transform -1 0 401200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_267
timestamp 1625505168
transform -1 0 424600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_45
timestamp 1625505168
transform -1 0 440000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_44
timestamp 1625505168
transform -1 0 436000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_43
timestamp 1625505168
transform -1 0 432000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_268
timestamp 1625505168
transform -1 0 426600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_269
timestamp 1625505168
transform -1 0 427600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_271
timestamp 1625505168
transform -1 0 428000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_270
timestamp 1625505168
transform -1 0 427800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_48
timestamp 1625505168
transform -1 0 452000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_47
timestamp 1625505168
transform -1 0 448000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_46
timestamp 1625505168
transform -1 0 444000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_278
timestamp 1625505168
transform -1 0 456000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_io1_pad
timestamp 1625505168
transform -1 0 475400 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_279
timestamp 1625505168
transform -1 0 458000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_280
timestamp 1625505168
transform -1 0 459000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_282
timestamp 1625505168
transform -1 0 459400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_281
timestamp 1625505168
transform -1 0 459200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_284
timestamp 1625505168
transform -1 0 479400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_285
timestamp 1625505168
transform -1 0 481400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_49
timestamp 1625505168
transform -1 0 486800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_286
timestamp 1625505168
transform -1 0 482400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_288
timestamp 1625505168
transform -1 0 482800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_287
timestamp 1625505168
transform -1 0 482600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_50
timestamp 1625505168
transform -1 0 490800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_51
timestamp 1625505168
transform -1 0 494800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_52
timestamp 1625505168
transform -1 0 498800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_53
timestamp 1625505168
transform -1 0 502800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_54
timestamp 1625505168
transform -1 0 506800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  gpio_pad
timestamp 1625505168
transform -1 0 530200 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_296
timestamp 1625505168
transform -1 0 512800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_297
timestamp 1625505168
transform -1 0 513800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_299
timestamp 1625505168
transform -1 0 514200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_298
timestamp 1625505168
transform -1 0 514000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_295
timestamp 1625505168
transform -1 0 510800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_55
timestamp 1625505168
transform -1 0 541600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_302
timestamp 1625505168
transform -1 0 536200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_303
timestamp 1625505168
transform -1 0 537200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_305
timestamp 1625505168
transform -1 0 537600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_304
timestamp 1625505168
transform -1 0 537400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_301
timestamp 1625505168
transform -1 0 534200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_57
timestamp 1625505168
transform -1 0 549600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_56
timestamp 1625505168
transform -1 0 545600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_60
timestamp 1625505168
transform -1 0 561600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_59
timestamp 1625505168
transform -1 0 557600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_58
timestamp 1625505168
transform -1 0 553600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_312
timestamp 1625505168
transform -1 0 565600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  mgmt_vssio_hvclamp_pad\[0\] $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1625505168
transform -1 0 584000 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_313
timestamp 1625505168
transform -1 0 567600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_314
timestamp 1625505168
transform -1 0 568600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_316
timestamp 1625505168
transform -1 0 569000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_315
timestamp 1625505168
transform -1 0 568800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_319
timestamp 1625505168
transform -1 0 590000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_320
timestamp 1625505168
transform -1 0 591000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_318
timestamp 1625505168
transform -1 0 588000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_64
timestamp 1625505168
transform -1 0 607400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_63
timestamp 1625505168
transform -1 0 603400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_62
timestamp 1625505168
transform -1 0 599400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_61
timestamp 1625505168
transform -1 0 595400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_322
timestamp 1625505168
transform -1 0 591400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_321
timestamp 1625505168
transform -1 0 591200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_66
timestamp 1625505168
transform -1 0 615400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_65
timestamp 1625505168
transform -1 0 611400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_330
timestamp 1625505168
transform -1 0 621400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_329
timestamp 1625505168
transform -1 0 619400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  mgmt_vdda_hvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1625505168
transform -1 0 637800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_331
timestamp 1625505168
transform -1 0 622400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_333
timestamp 1625505168
transform -1 0 622800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_332
timestamp 1625505168
transform -1 0 622600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_335
timestamp 1625505168
transform -1 0 641800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_336
timestamp 1625505168
transform -1 0 643800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_337
timestamp 1625505168
transform -1 0 644800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_338
timestamp 1625505168
transform -1 0 645000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_67
timestamp 1625505168
transform -1 0 649200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_339
timestamp 1625505168
transform -1 0 645200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_68
timestamp 1625505168
transform -1 0 653200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_69
timestamp 1625505168
transform -1 0 657200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_70
timestamp 1625505168
transform -1 0 661200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_71
timestamp 1625505168
transform -1 0 665200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_72
timestamp 1625505168
transform -1 0 669200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_346
timestamp 1625505168
transform -1 0 673200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_347
timestamp 1625505168
transform -1 0 675200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__corner_pad  mgmt_corner\[1\]
timestamp 1625505168
transform 0 1 676800 -1 0 40000
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_5um  FILLER_348
timestamp 1625505168
transform -1 0 676200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_349
timestamp 1625505168
transform -1 0 676400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_350
timestamp 1625505168
transform -1 0 676600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_351
timestamp 1625505168
transform -1 0 676800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_580
timestamp 1625505168
transform 0 1 678007 -1 0 44000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_356
timestamp 1625505168
transform 0 -1 39593 1 0 56800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_355
timestamp 1625505168
transform 0 -1 39593 1 0 52800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_354
timestamp 1625505168
transform 0 -1 39593 1 0 48800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_353
timestamp 1625505168
transform 0 -1 39593 1 0 44800
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_clamped_pad  mgmt_vccd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1625505168
transform 0 -1 39593 1 0 68000
box 0 -2107 17239 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_358
timestamp 1625505168
transform 0 -1 39593 1 0 64800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_359
timestamp 1625505168
transform 0 -1 39593 1 0 66800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_360
timestamp 1625505168
transform 0 -1 39593 1 0 67800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_357
timestamp 1625505168
transform 0 -1 39593 1 0 60800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_362
timestamp 1625505168
transform 0 -1 39593 1 0 83000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_581
timestamp 1625505168
transform 0 1 678007 -1 0 48000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_582
timestamp 1625505168
transform 0 1 678007 -1 0 52000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_583
timestamp 1625505168
transform 0 1 678007 -1 0 56000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_584
timestamp 1625505168
transform 0 1 678007 -1 0 60000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_585
timestamp 1625505168
transform 0 1 678007 -1 0 64000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_586
timestamp 1625505168
transform 0 1 678007 -1 0 68000
box 0 0 4000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_1 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1625505168
transform 0 1 678007 -1 0 70000
box 0 0 1000 39593
use sky130_ef_io__disconnect_vccd_slice_5um  disconnect_vccd_1 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1625505168
transform 0 1 678007 -1 0 71000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_587
timestamp 1625505168
transform 0 1 678007 -1 0 69000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_590
timestamp 1625505168
transform 0 1 678007 -1 0 75000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_591
timestamp 1625505168
transform 0 1 678007 -1 0 79000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_592
timestamp 1625505168
transform 0 1 678007 -1 0 83000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_593
timestamp 1625505168
transform 0 1 678007 -1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_366
timestamp 1625505168
transform 0 -1 39593 1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_365
timestamp 1625505168
transform 0 -1 39593 1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_364
timestamp 1625505168
transform 0 -1 39593 1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_363
timestamp 1625505168
transform 0 -1 39593 1 0 87000
box 0 0 4000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  mgmt_vddio_hvclamp_pad\[0\] $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1625505168
transform 0 -1 39593 1 0 110200
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_368
timestamp 1625505168
transform 0 -1 39593 1 0 107000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_369
timestamp 1625505168
transform 0 -1 39593 1 0 109000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_370
timestamp 1625505168
transform 0 -1 39593 1 0 110000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_367
timestamp 1625505168
transform 0 -1 39593 1 0 103000
box 0 0 4000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_2
timestamp 1625505168
transform 0 -1 39593 1 0 125200
box 0 0 1000 39593
use sky130_ef_io__disconnect_vccd_slice_5um  disconnect_vccd_2
timestamp 1625505168
transform 0 -1 39593 1 0 126200
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[0\]
timestamp 1625505168
transform 0 1 675407 -1 0 116000
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_597
timestamp 1625505168
transform 0 1 678007 -1 0 100000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_601
timestamp 1625505168
transform 0 1 678007 -1 0 128000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_600
timestamp 1625505168
transform 0 1 678007 -1 0 124000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_599
timestamp 1625505168
transform 0 1 678007 -1 0 120000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_596
timestamp 1625505168
transform 0 1 678007 -1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_595
timestamp 1625505168
transform 0 1 678007 -1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_594
timestamp 1625505168
transform 0 1 678007 -1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_374
timestamp 1625505168
transform 0 -1 39593 1 0 127200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_375
timestamp 1625505168
transform 0 -1 39593 1 0 131200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_376
timestamp 1625505168
transform 0 -1 39593 1 0 135200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_377
timestamp 1625505168
transform 0 -1 39593 1 0 139200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_378
timestamp 1625505168
transform 0 -1 39593 1 0 143200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_379
timestamp 1625505168
transform 0 -1 39593 1 0 147200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_380
timestamp 1625505168
transform 0 -1 39593 1 0 151200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_381
timestamp 1625505168
transform 0 -1 39593 1 0 155200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_382
timestamp 1625505168
transform 0 -1 39593 1 0 159200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_383
timestamp 1625505168
transform 0 -1 39593 1 0 163200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_384
timestamp 1625505168
transform 0 -1 39593 1 0 167200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[1\]
timestamp 1625505168
transform 0 1 675407 -1 0 161200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_606
timestamp 1625505168
transform 0 1 678007 -1 0 145000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_607
timestamp 1625505168
transform 0 1 678007 -1 0 145200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_610
timestamp 1625505168
transform 0 1 678007 -1 0 169200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_609
timestamp 1625505168
transform 0 1 678007 -1 0 165200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_605
timestamp 1625505168
transform 0 1 678007 -1 0 144000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_604
timestamp 1625505168
transform 0 1 678007 -1 0 140000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_603
timestamp 1625505168
transform 0 1 678007 -1 0 136000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_602
timestamp 1625505168
transform 0 1 678007 -1 0 132000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[12\]
timestamp 1625505168
transform 0 -1 42193 1 0 181600
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_387
timestamp 1625505168
transform 0 -1 39593 1 0 179200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_389
timestamp 1625505168
transform 0 -1 39593 1 0 181400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_388
timestamp 1625505168
transform 0 -1 39593 1 0 181200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_386
timestamp 1625505168
transform 0 -1 39593 1 0 175200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_385
timestamp 1625505168
transform 0 -1 39593 1 0 171200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_391
timestamp 1625505168
transform 0 -1 39593 1 0 197600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_394
timestamp 1625505168
transform 0 -1 39593 1 0 209600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_393
timestamp 1625505168
transform 0 -1 39593 1 0 205600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_392
timestamp 1625505168
transform 0 -1 39593 1 0 201600
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[2\]
timestamp 1625505168
transform 0 1 675407 -1 0 206200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_616
timestamp 1625505168
transform 0 1 678007 -1 0 190200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_619
timestamp 1625505168
transform 0 1 678007 -1 0 214200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_618
timestamp 1625505168
transform 0 1 678007 -1 0 210200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_615
timestamp 1625505168
transform 0 1 678007 -1 0 189200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_614
timestamp 1625505168
transform 0 1 678007 -1 0 185200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_613
timestamp 1625505168
transform 0 1 678007 -1 0 181200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_612
timestamp 1625505168
transform 0 1 678007 -1 0 177200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_611
timestamp 1625505168
transform 0 1 678007 -1 0 173200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[11\]
timestamp 1625505168
transform 0 -1 42193 1 0 224800
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_397
timestamp 1625505168
transform 0 -1 39593 1 0 221600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_398
timestamp 1625505168
transform 0 -1 39593 1 0 223600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_399
timestamp 1625505168
transform 0 -1 39593 1 0 224600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_396
timestamp 1625505168
transform 0 -1 39593 1 0 217600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_395
timestamp 1625505168
transform 0 -1 39593 1 0 213600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_401
timestamp 1625505168
transform 0 -1 39593 1 0 240800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_404
timestamp 1625505168
transform 0 -1 39593 1 0 252800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_403
timestamp 1625505168
transform 0 -1 39593 1 0 248800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_402
timestamp 1625505168
transform 0 -1 39593 1 0 244800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[3\]
timestamp 1625505168
transform 0 1 675407 -1 0 251400
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_625
timestamp 1625505168
transform 0 1 678007 -1 0 235200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_626
timestamp 1625505168
transform 0 1 678007 -1 0 235400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_628
timestamp 1625505168
transform 0 1 678007 -1 0 255400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_624
timestamp 1625505168
transform 0 1 678007 -1 0 234200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_623
timestamp 1625505168
transform 0 1 678007 -1 0 230200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_622
timestamp 1625505168
transform 0 1 678007 -1 0 226200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_621
timestamp 1625505168
transform 0 1 678007 -1 0 222200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_620
timestamp 1625505168
transform 0 1 678007 -1 0 218200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[10\]
timestamp 1625505168
transform 0 -1 42193 1 0 268000
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_407
timestamp 1625505168
transform 0 -1 39593 1 0 264800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_408
timestamp 1625505168
transform 0 -1 39593 1 0 266800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_409
timestamp 1625505168
transform 0 -1 39593 1 0 267800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_413
timestamp 1625505168
transform 0 -1 39593 1 0 292000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_412
timestamp 1625505168
transform 0 -1 39593 1 0 288000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_411
timestamp 1625505168
transform 0 -1 39593 1 0 284000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_406
timestamp 1625505168
transform 0 -1 39593 1 0 260800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_405
timestamp 1625505168
transform 0 -1 39593 1 0 256800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[4\]
timestamp 1625505168
transform 0 1 675407 -1 0 296400
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_635
timestamp 1625505168
transform 0 1 678007 -1 0 280400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_634
timestamp 1625505168
transform 0 1 678007 -1 0 279400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_633
timestamp 1625505168
transform 0 1 678007 -1 0 275400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_632
timestamp 1625505168
transform 0 1 678007 -1 0 271400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_631
timestamp 1625505168
transform 0 1 678007 -1 0 267400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_630
timestamp 1625505168
transform 0 1 678007 -1 0 263400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_629
timestamp 1625505168
transform 0 1 678007 -1 0 259400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[9\]
timestamp 1625505168
transform 0 -1 42193 1 0 311200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_417
timestamp 1625505168
transform 0 -1 39593 1 0 308000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_418
timestamp 1625505168
transform 0 -1 39593 1 0 310000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_419
timestamp 1625505168
transform 0 -1 39593 1 0 311000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_416
timestamp 1625505168
transform 0 -1 39593 1 0 304000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_415
timestamp 1625505168
transform 0 -1 39593 1 0 300000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_414
timestamp 1625505168
transform 0 -1 39593 1 0 296000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_421
timestamp 1625505168
transform 0 -1 39593 1 0 327200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_423
timestamp 1625505168
transform 0 -1 39593 1 0 335200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_422
timestamp 1625505168
transform 0 -1 39593 1 0 331200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[5\]
timestamp 1625505168
transform 0 1 675407 -1 0 341400
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_644
timestamp 1625505168
transform 0 1 678007 -1 0 325400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_643
timestamp 1625505168
transform 0 1 678007 -1 0 324400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_642
timestamp 1625505168
transform 0 1 678007 -1 0 320400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_641
timestamp 1625505168
transform 0 1 678007 -1 0 316400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_640
timestamp 1625505168
transform 0 1 678007 -1 0 312400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_639
timestamp 1625505168
transform 0 1 678007 -1 0 308400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_638
timestamp 1625505168
transform 0 1 678007 -1 0 304400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_637
timestamp 1625505168
transform 0 1 678007 -1 0 300400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_427
timestamp 1625505168
transform 0 -1 39593 1 0 351200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_428
timestamp 1625505168
transform 0 -1 39593 1 0 353200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_426
timestamp 1625505168
transform 0 -1 39593 1 0 347200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_425
timestamp 1625505168
transform 0 -1 39593 1 0 343200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_424
timestamp 1625505168
transform 0 -1 39593 1 0 339200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[8\]
timestamp 1625505168
transform 0 -1 42193 1 0 354400
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_1um  FILLER_429
timestamp 1625505168
transform 0 -1 39593 1 0 354200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_433
timestamp 1625505168
transform 0 -1 39593 1 0 378400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_432
timestamp 1625505168
transform 0 -1 39593 1 0 374400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_431
timestamp 1625505168
transform 0 -1 39593 1 0 370400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_646
timestamp 1625505168
transform 0 1 678007 -1 0 345400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_647
timestamp 1625505168
transform 0 1 678007 -1 0 349400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_648
timestamp 1625505168
transform 0 1 678007 -1 0 353400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_649
timestamp 1625505168
transform 0 1 678007 -1 0 357400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_653
timestamp 1625505168
transform 0 1 678007 -1 0 370400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_650
timestamp 1625505168
transform 0 1 678007 -1 0 361400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_651
timestamp 1625505168
transform 0 1 678007 -1 0 365400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_652
timestamp 1625505168
transform 0 1 678007 -1 0 369400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[6\]
timestamp 1625505168
transform 0 1 675407 -1 0 386600
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_1um  FILLER_654
timestamp 1625505168
transform 0 1 678007 -1 0 370600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_437
timestamp 1625505168
transform 0 -1 39593 1 0 394400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_436
timestamp 1625505168
transform 0 -1 39593 1 0 390400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_435
timestamp 1625505168
transform 0 -1 39593 1 0 386400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_434
timestamp 1625505168
transform 0 -1 39593 1 0 382400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[7\]
timestamp 1625505168
transform 0 -1 42193 1 0 397600
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_438
timestamp 1625505168
transform 0 -1 39593 1 0 396400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_439
timestamp 1625505168
transform 0 -1 39593 1 0 397400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_443
timestamp 1625505168
transform 0 -1 39593 1 0 421600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_442
timestamp 1625505168
transform 0 -1 39593 1 0 417600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_441
timestamp 1625505168
transform 0 -1 39593 1 0 413600
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user1_vssa_hvclamp_pad\[1\]
timestamp 1625505168
transform 0 1 678007 -1 0 430600
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_663
timestamp 1625505168
transform 0 1 678007 -1 0 415600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_658
timestamp 1625505168
transform 0 1 678007 -1 0 398600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_657
timestamp 1625505168
transform 0 1 678007 -1 0 394600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_656
timestamp 1625505168
transform 0 1 678007 -1 0 390600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_661
timestamp 1625505168
transform 0 1 678007 -1 0 410600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_660
timestamp 1625505168
transform 0 1 678007 -1 0 406600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_659
timestamp 1625505168
transform 0 1 678007 -1 0 402600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_662
timestamp 1625505168
transform 0 1 678007 -1 0 414600
box 0 0 4000 39593
use sky130_ef_io__vssd_lvc_clamped2_pad  user2_vssd_lvclmap_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1625505168
transform 0 -1 39593 1 0 440800
box -2195 -2184 17228 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_447
timestamp 1625505168
transform 0 -1 39593 1 0 437600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_448
timestamp 1625505168
transform 0 -1 39593 1 0 439600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_449
timestamp 1625505168
transform 0 -1 39593 1 0 440600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_446
timestamp 1625505168
transform 0 -1 39593 1 0 433600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_445
timestamp 1625505168
transform 0 -1 39593 1 0 429600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_444
timestamp 1625505168
transform 0 -1 39593 1 0 425600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_452
timestamp 1625505168
transform 0 -1 39593 1 0 459800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_451
timestamp 1625505168
transform 0 -1 39593 1 0 455800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_453
timestamp 1625505168
transform 0 -1 39593 1 0 463800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_665
timestamp 1625505168
transform 0 1 678007 -1 0 434600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_666
timestamp 1625505168
transform 0 1 678007 -1 0 438600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_667
timestamp 1625505168
transform 0 1 678007 -1 0 442600
box 0 0 4000 39593
use sky130_ef_io__vssd_lvc_clamped2_pad  user1_vssd_lvclmap_pad
timestamp 1625505168
transform 0 1 678007 -1 0 474800
box -2195 -2184 17228 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_672
timestamp 1625505168
transform 0 1 678007 -1 0 459600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_673
timestamp 1625505168
transform 0 1 678007 -1 0 459800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_668
timestamp 1625505168
transform 0 1 678007 -1 0 446600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_669
timestamp 1625505168
transform 0 1 678007 -1 0 450600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_670
timestamp 1625505168
transform 0 1 678007 -1 0 454600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_671
timestamp 1625505168
transform 0 1 678007 -1 0 458600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_456
timestamp 1625505168
transform 0 -1 39593 1 0 475800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_455
timestamp 1625505168
transform 0 -1 39593 1 0 471800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_454
timestamp 1625505168
transform 0 -1 39593 1 0 467800
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user2_vdda_hvclamp_pad
timestamp 1625505168
transform 0 -1 39593 1 0 483000
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_457
timestamp 1625505168
transform 0 -1 39593 1 0 479800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_458
timestamp 1625505168
transform 0 -1 39593 1 0 481800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_459
timestamp 1625505168
transform 0 -1 39593 1 0 482800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_463
timestamp 1625505168
transform 0 -1 39593 1 0 506000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_462
timestamp 1625505168
transform 0 -1 39593 1 0 502000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_461
timestamp 1625505168
transform 0 -1 39593 1 0 498000
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user1_vdda_hvclamp_pad\[1\]
timestamp 1625505168
transform 0 1 678007 -1 0 518800
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_682
timestamp 1625505168
transform 0 1 678007 -1 0 503800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_676
timestamp 1625505168
transform 0 1 678007 -1 0 482800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_675
timestamp 1625505168
transform 0 1 678007 -1 0 478800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_679
timestamp 1625505168
transform 0 1 678007 -1 0 494800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_678
timestamp 1625505168
transform 0 1 678007 -1 0 490800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_677
timestamp 1625505168
transform 0 1 678007 -1 0 486800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_681
timestamp 1625505168
transform 0 1 678007 -1 0 502800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_680
timestamp 1625505168
transform 0 1 678007 -1 0 498800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[6\]
timestamp 1625505168
transform 0 -1 42193 1 0 525200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_467
timestamp 1625505168
transform 0 -1 39593 1 0 522000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_468
timestamp 1625505168
transform 0 -1 39593 1 0 524000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_469
timestamp 1625505168
transform 0 -1 39593 1 0 525000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_466
timestamp 1625505168
transform 0 -1 39593 1 0 518000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_465
timestamp 1625505168
transform 0 -1 39593 1 0 514000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_464
timestamp 1625505168
transform 0 -1 39593 1 0 510000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_472
timestamp 1625505168
transform 0 -1 39593 1 0 545200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_471
timestamp 1625505168
transform 0 -1 39593 1 0 541200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[7\]
timestamp 1625505168
transform 0 1 675407 -1 0 563800
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_691
timestamp 1625505168
transform 0 1 678007 -1 0 547800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_690
timestamp 1625505168
transform 0 1 678007 -1 0 546800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_689
timestamp 1625505168
transform 0 1 678007 -1 0 542800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_688
timestamp 1625505168
transform 0 1 678007 -1 0 538800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_687
timestamp 1625505168
transform 0 1 678007 -1 0 534800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_686
timestamp 1625505168
transform 0 1 678007 -1 0 530800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_685
timestamp 1625505168
transform 0 1 678007 -1 0 526800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_684
timestamp 1625505168
transform 0 1 678007 -1 0 522800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_476
timestamp 1625505168
transform 0 -1 39593 1 0 561200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_475
timestamp 1625505168
transform 0 -1 39593 1 0 557200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_474
timestamp 1625505168
transform 0 -1 39593 1 0 553200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_473
timestamp 1625505168
transform 0 -1 39593 1 0 549200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[5\]
timestamp 1625505168
transform 0 -1 42193 1 0 568400
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_477
timestamp 1625505168
transform 0 -1 39593 1 0 565200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_478
timestamp 1625505168
transform 0 -1 39593 1 0 567200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_479
timestamp 1625505168
transform 0 -1 39593 1 0 568200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_482
timestamp 1625505168
transform 0 -1 39593 1 0 588400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_481
timestamp 1625505168
transform 0 -1 39593 1 0 584400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_699
timestamp 1625505168
transform 0 1 678007 -1 0 591800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_698
timestamp 1625505168
transform 0 1 678007 -1 0 587800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_697
timestamp 1625505168
transform 0 1 678007 -1 0 583800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_696
timestamp 1625505168
transform 0 1 678007 -1 0 579800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_695
timestamp 1625505168
transform 0 1 678007 -1 0 575800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_694
timestamp 1625505168
transform 0 1 678007 -1 0 571800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_693
timestamp 1625505168
transform 0 1 678007 -1 0 567800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_486
timestamp 1625505168
transform 0 -1 39593 1 0 604400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_485
timestamp 1625505168
transform 0 -1 39593 1 0 600400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_484
timestamp 1625505168
transform 0 -1 39593 1 0 596400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_483
timestamp 1625505168
transform 0 -1 39593 1 0 592400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[4\]
timestamp 1625505168
transform 0 -1 42193 1 0 611600
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_487
timestamp 1625505168
transform 0 -1 39593 1 0 608400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_488
timestamp 1625505168
transform 0 -1 39593 1 0 610400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_489
timestamp 1625505168
transform 0 -1 39593 1 0 611400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_492
timestamp 1625505168
transform 0 -1 39593 1 0 631600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_491
timestamp 1625505168
transform 0 -1 39593 1 0 627600
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[8\]
timestamp 1625505168
transform 0 1 675407 -1 0 609000
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_700
timestamp 1625505168
transform 0 1 678007 -1 0 592800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_701
timestamp 1625505168
transform 0 1 678007 -1 0 593000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_706
timestamp 1625505168
transform 0 1 678007 -1 0 625000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_705
timestamp 1625505168
transform 0 1 678007 -1 0 621000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_704
timestamp 1625505168
transform 0 1 678007 -1 0 617000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_703
timestamp 1625505168
transform 0 1 678007 -1 0 613000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_708
timestamp 1625505168
transform 0 1 678007 -1 0 633000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_707
timestamp 1625505168
transform 0 1 678007 -1 0 629000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_496
timestamp 1625505168
transform 0 -1 39593 1 0 647600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_495
timestamp 1625505168
transform 0 -1 39593 1 0 643600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_494
timestamp 1625505168
transform 0 -1 39593 1 0 639600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_493
timestamp 1625505168
transform 0 -1 39593 1 0 635600
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[3\]
timestamp 1625505168
transform 0 -1 42193 1 0 654800
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_497
timestamp 1625505168
transform 0 -1 39593 1 0 651600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_498
timestamp 1625505168
transform 0 -1 39593 1 0 653600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_499
timestamp 1625505168
transform 0 -1 39593 1 0 654600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_502
timestamp 1625505168
transform 0 -1 39593 1 0 674800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_501
timestamp 1625505168
transform 0 -1 39593 1 0 670800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[9\]
timestamp 1625505168
transform 0 1 675407 -1 0 654000
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_710
timestamp 1625505168
transform 0 1 678007 -1 0 638000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_717
timestamp 1625505168
transform 0 1 678007 -1 0 678000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_716
timestamp 1625505168
transform 0 1 678007 -1 0 674000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_715
timestamp 1625505168
transform 0 1 678007 -1 0 670000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_714
timestamp 1625505168
transform 0 1 678007 -1 0 666000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_713
timestamp 1625505168
transform 0 1 678007 -1 0 662000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_712
timestamp 1625505168
transform 0 1 678007 -1 0 658000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_709
timestamp 1625505168
transform 0 1 678007 -1 0 637000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[2\]
timestamp 1625505168
transform 0 -1 42193 1 0 698000
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_507
timestamp 1625505168
transform 0 -1 39593 1 0 694800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_508
timestamp 1625505168
transform 0 -1 39593 1 0 696800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_509
timestamp 1625505168
transform 0 -1 39593 1 0 697800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_506
timestamp 1625505168
transform 0 -1 39593 1 0 690800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_505
timestamp 1625505168
transform 0 -1 39593 1 0 686800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_504
timestamp 1625505168
transform 0 -1 39593 1 0 682800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_503
timestamp 1625505168
transform 0 -1 39593 1 0 678800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_511
timestamp 1625505168
transform 0 -1 39593 1 0 714000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[10\]
timestamp 1625505168
transform 0 1 675407 -1 0 699200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_719
timestamp 1625505168
transform 0 1 678007 -1 0 683000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_720
timestamp 1625505168
transform 0 1 678007 -1 0 683200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_726
timestamp 1625505168
transform 0 1 678007 -1 0 719200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_725
timestamp 1625505168
transform 0 1 678007 -1 0 715200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_724
timestamp 1625505168
transform 0 1 678007 -1 0 711200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_723
timestamp 1625505168
transform 0 1 678007 -1 0 707200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_722
timestamp 1625505168
transform 0 1 678007 -1 0 703200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_718
timestamp 1625505168
transform 0 1 678007 -1 0 682000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_515
timestamp 1625505168
transform 0 -1 39593 1 0 730000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_514
timestamp 1625505168
transform 0 -1 39593 1 0 726000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_513
timestamp 1625505168
transform 0 -1 39593 1 0 722000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_512
timestamp 1625505168
transform 0 -1 39593 1 0 718000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[1\]
timestamp 1625505168
transform 0 -1 42193 1 0 741200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_517
timestamp 1625505168
transform 0 -1 39593 1 0 738000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_518
timestamp 1625505168
transform 0 -1 39593 1 0 740000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_519
timestamp 1625505168
transform 0 -1 39593 1 0 741000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_516
timestamp 1625505168
transform 0 -1 39593 1 0 734000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_521
timestamp 1625505168
transform 0 -1 39593 1 0 757200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[11\]
timestamp 1625505168
transform 0 1 675407 -1 0 744200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_729
timestamp 1625505168
transform 0 1 678007 -1 0 728200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_728
timestamp 1625505168
transform 0 1 678007 -1 0 727200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_727
timestamp 1625505168
transform 0 1 678007 -1 0 723200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_732
timestamp 1625505168
transform 0 1 678007 -1 0 752200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_731
timestamp 1625505168
transform 0 1 678007 -1 0 748200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_734
timestamp 1625505168
transform 0 1 678007 -1 0 760200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_733
timestamp 1625505168
transform 0 1 678007 -1 0 756200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_525
timestamp 1625505168
transform 0 -1 39593 1 0 773200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_524
timestamp 1625505168
transform 0 -1 39593 1 0 769200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_523
timestamp 1625505168
transform 0 -1 39593 1 0 765200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_522
timestamp 1625505168
transform 0 -1 39593 1 0 761200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[0\]
timestamp 1625505168
transform 0 -1 42193 1 0 784400
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_527
timestamp 1625505168
transform 0 -1 39593 1 0 781200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_528
timestamp 1625505168
transform 0 -1 39593 1 0 783200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_529
timestamp 1625505168
transform 0 -1 39593 1 0 784200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_526
timestamp 1625505168
transform 0 -1 39593 1 0 777200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_531
timestamp 1625505168
transform 0 -1 39593 1 0 800400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[12\]
timestamp 1625505168
transform 0 1 675407 -1 0 789200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_738
timestamp 1625505168
transform 0 1 678007 -1 0 773200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_743
timestamp 1625505168
transform 0 1 678007 -1 0 805200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_742
timestamp 1625505168
transform 0 1 678007 -1 0 801200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_741
timestamp 1625505168
transform 0 1 678007 -1 0 797200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_740
timestamp 1625505168
transform 0 1 678007 -1 0 793200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_737
timestamp 1625505168
transform 0 1 678007 -1 0 772200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_736
timestamp 1625505168
transform 0 1 678007 -1 0 768200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_735
timestamp 1625505168
transform 0 1 678007 -1 0 764200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_535
timestamp 1625505168
transform 0 -1 39593 1 0 816400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_534
timestamp 1625505168
transform 0 -1 39593 1 0 812400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_533
timestamp 1625505168
transform 0 -1 39593 1 0 808400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_532
timestamp 1625505168
transform 0 -1 39593 1 0 804400
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user2_vssa_hvclamp_pad
timestamp 1625505168
transform 0 -1 39593 1 0 827600
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_537
timestamp 1625505168
transform 0 -1 39593 1 0 824400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_538
timestamp 1625505168
transform 0 -1 39593 1 0 826400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_539
timestamp 1625505168
transform 0 -1 39593 1 0 827400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_536
timestamp 1625505168
transform 0 -1 39593 1 0 820400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_541
timestamp 1625505168
transform 0 -1 39593 1 0 842600
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user1_vdda_hvclamp_pad\[0\]
timestamp 1625505168
transform 0 1 678007 -1 0 833400
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_747
timestamp 1625505168
transform 0 1 678007 -1 0 818200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_748
timestamp 1625505168
transform 0 1 678007 -1 0 818400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_752
timestamp 1625505168
transform 0 1 678007 -1 0 845400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_751
timestamp 1625505168
transform 0 1 678007 -1 0 841400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_750
timestamp 1625505168
transform 0 1 678007 -1 0 837400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_746
timestamp 1625505168
transform 0 1 678007 -1 0 817200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_745
timestamp 1625505168
transform 0 1 678007 -1 0 813200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_744
timestamp 1625505168
transform 0 1 678007 -1 0 809200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_545
timestamp 1625505168
transform 0 -1 39593 1 0 858600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_544
timestamp 1625505168
transform 0 -1 39593 1 0 854600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_543
timestamp 1625505168
transform 0 -1 39593 1 0 850600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_542
timestamp 1625505168
transform 0 -1 39593 1 0 846600
box 0 0 4000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  mgmt_vddio_hvclamp_pad\[1\]
timestamp 1625505168
transform 0 -1 39593 1 0 869800
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_547
timestamp 1625505168
transform 0 -1 39593 1 0 866600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_548
timestamp 1625505168
transform 0 -1 39593 1 0 868600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_549
timestamp 1625505168
transform 0 -1 39593 1 0 869600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_546
timestamp 1625505168
transform 0 -1 39593 1 0 862600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_551
timestamp 1625505168
transform 0 -1 39593 1 0 884800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[13\]
timestamp 1625505168
transform 0 1 675407 -1 0 878400
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_757
timestamp 1625505168
transform 0 1 678007 -1 0 862400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_760
timestamp 1625505168
transform 0 1 678007 -1 0 886400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_759
timestamp 1625505168
transform 0 1 678007 -1 0 882400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_756
timestamp 1625505168
transform 0 1 678007 -1 0 861400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_755
timestamp 1625505168
transform 0 1 678007 -1 0 857400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_754
timestamp 1625505168
transform 0 1 678007 -1 0 853400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_753
timestamp 1625505168
transform 0 1 678007 -1 0 849400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_556
timestamp 1625505168
transform 0 -1 39593 1 0 904800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_555
timestamp 1625505168
transform 0 -1 39593 1 0 900800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_554
timestamp 1625505168
transform 0 -1 39593 1 0 896800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_553
timestamp 1625505168
transform 0 -1 39593 1 0 892800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_552
timestamp 1625505168
transform 0 -1 39593 1 0 888800
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_clamped2_pad  user2_vccd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1625505168
transform 0 -1 39593 1 0 912000
box -2195 -2184 17228 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_557
timestamp 1625505168
transform 0 -1 39593 1 0 908800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_558
timestamp 1625505168
transform 0 -1 39593 1 0 910800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_559
timestamp 1625505168
transform 0 -1 39593 1 0 911800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_561
timestamp 1625505168
transform 0 -1 39593 1 0 927000
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_clamped2_pad  user1_vccd_lvclamp_pad
timestamp 1625505168
transform 0 1 678007 -1 0 922600
box -2195 -2184 17228 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_765
timestamp 1625505168
transform 0 1 678007 -1 0 906400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_764
timestamp 1625505168
transform 0 1 678007 -1 0 902400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_763
timestamp 1625505168
transform 0 1 678007 -1 0 898400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_762
timestamp 1625505168
transform 0 1 678007 -1 0 894400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_761
timestamp 1625505168
transform 0 1 678007 -1 0 890400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_766
timestamp 1625505168
transform 0 1 678007 -1 0 907400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_767
timestamp 1625505168
transform 0 1 678007 -1 0 907600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_769
timestamp 1625505168
transform 0 1 678007 -1 0 926600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_770
timestamp 1625505168
transform 0 1 678007 -1 0 930600
box 0 0 4000 39593
use sky130_ef_io__analog_pad  user2_analog_pad\[3\] $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1625505168
transform 0 -1 40000 1 0 955200
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_1um  FILLER_568
timestamp 1625505168
transform 0 -1 39593 1 0 955000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_565
timestamp 1625505168
transform 0 -1 39593 1 0 943000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_564
timestamp 1625505168
transform 0 -1 39593 1 0 939000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_563
timestamp 1625505168
transform 0 -1 39593 1 0 935000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_562
timestamp 1625505168
transform 0 -1 39593 1 0 931000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_567
timestamp 1625505168
transform 0 -1 39593 1 0 951000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_566
timestamp 1625505168
transform 0 -1 39593 1 0 947000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_570
timestamp 1625505168
transform 0 -1 39593 1 0 970200
box 0 0 4000 39593
use sky130_ef_io__analog_pad  user1_analog_pad\[3\]
timestamp 1625505168
transform 0 1 677600 -1 0 966600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_10um  FILLER_776
timestamp 1625505168
transform 0 1 678007 -1 0 968600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_777
timestamp 1625505168
transform 0 1 678007 -1 0 951600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_779
timestamp 1625505168
transform 0 1 678007 -1 0 972600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_775
timestamp 1625505168
transform 0 1 678007 -1 0 950600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_774
timestamp 1625505168
transform 0 1 678007 -1 0 946600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_773
timestamp 1625505168
transform 0 1 678007 -1 0 942600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_772
timestamp 1625505168
transform 0 1 678007 -1 0 938600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_771
timestamp 1625505168
transform 0 1 678007 -1 0 934600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_575
timestamp 1625505168
transform 0 -1 39593 1 0 990200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_574
timestamp 1625505168
transform 0 -1 39593 1 0 986200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_573
timestamp 1625505168
transform 0 -1 39593 1 0 982200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_572
timestamp 1625505168
transform 0 -1 39593 1 0 978200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_571
timestamp 1625505168
transform 0 -1 39593 1 0 974200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_576
timestamp 1625505168
transform 0 -1 39593 1 0 994200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_577
timestamp 1625505168
transform 0 -1 39593 1 0 996200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_579
timestamp 1625505168
transform 0 -1 39593 1 0 997400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_578
timestamp 1625505168
transform 0 -1 39593 1 0 997200
box 0 0 200 39593
use sky130_ef_io__corner_pad  user2_corner
timestamp 1625505168
transform 0 -1 40800 1 0 997600
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_20um  FILLER_5
timestamp 1625505168
transform 1 0 40800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_9
timestamp 1625505168
transform 1 0 56800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_8
timestamp 1625505168
transform 1 0 52800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_7
timestamp 1625505168
transform 1 0 48800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_6
timestamp 1625505168
transform 1 0 44800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_12
timestamp 1625505168
transform 1 0 68800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_11
timestamp 1625505168
transform 1 0 64800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_10
timestamp 1625505168
transform 1 0 60800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__analog_pad  user2_analog_pad\[2\]
timestamp 1625505168
transform 1 0 77200 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_1um  FILLER_15
timestamp 1625505168
transform 1 0 77000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_14
timestamp 1625505168
transform 1 0 76800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_13
timestamp 1625505168
transform 1 0 72800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_18
timestamp 1625505168
transform 1 0 96200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_17
timestamp 1625505168
transform 1 0 92200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_22
timestamp 1625505168
transform 1 0 112200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_21
timestamp 1625505168
transform 1 0 108200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_20
timestamp 1625505168
transform 1 0 104200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_19
timestamp 1625505168
transform 1 0 100200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_25
timestamp 1625505168
transform 1 0 124200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_24
timestamp 1625505168
transform 1 0 120200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_23
timestamp 1625505168
transform 1 0 116200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__analog_pad  user2_analog_pad\[1\]
timestamp 1625505168
transform 1 0 128600 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_1um  FILLER_27
timestamp 1625505168
transform 1 0 128400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_26
timestamp 1625505168
transform 1 0 128200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_32
timestamp 1625505168
transform 1 0 155600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_31
timestamp 1625505168
transform 1 0 151600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_30
timestamp 1625505168
transform 1 0 147600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_29
timestamp 1625505168
transform 1 0 143600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_35
timestamp 1625505168
transform 1 0 167600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_34
timestamp 1625505168
transform 1 0 163600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_33
timestamp 1625505168
transform 1 0 159600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__analog_pad  user2_analog_pad\[0\]
timestamp 1625505168
transform 1 0 180000 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_1um  FILLER_38
timestamp 1625505168
transform 1 0 179600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_39
timestamp 1625505168
transform 1 0 179800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_37
timestamp 1625505168
transform 1 0 175600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_36
timestamp 1625505168
transform 1 0 171600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_41
timestamp 1625505168
transform 1 0 195000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_44
timestamp 1625505168
transform 1 0 207000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_43
timestamp 1625505168
transform 1 0 203000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_42
timestamp 1625505168
transform 1 0 199000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__top_power_hvc  user2_analog_pad_with_clamp\[1\] $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1625505168
transform 1 0 221000 0 1 998007
box 0 -407 33800 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_47
timestamp 1625505168
transform 1 0 219000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_46
timestamp 1625505168
transform 1 0 215000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_45
timestamp 1625505168
transform 1 0 211000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_49
timestamp 1625505168
transform 1 0 254800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_50
timestamp 1625505168
transform 1 0 258800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_51
timestamp 1625505168
transform 1 0 262800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_52
timestamp 1625505168
transform 1 0 266800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_2
timestamp 1625505168
transform 1 0 272600 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_53
timestamp 1625505168
transform 1 0 270800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_54
timestamp 1625505168
transform 1 0 271800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_55
timestamp 1625505168
transform 1 0 272000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_56
timestamp 1625505168
transform 1 0 272200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_57
timestamp 1625505168
transform 1 0 272400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__top_power_hvc  user2_analog_pad_with_clamp\[0\]
timestamp 1625505168
transform 1 0 273600 0 1 998007
box 0 -407 33800 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_1
timestamp 1625505168
transform 1 0 308400 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_3
timestamp 1625505168
transform 1 0 307400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_60
timestamp 1625505168
transform 1 0 310400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_63
timestamp 1625505168
transform 1 0 322400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_62
timestamp 1625505168
transform 1 0 318400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_61
timestamp 1625505168
transform 1 0 314400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  mgmt_vssio_hvclamp_pad\[1\]
timestamp 1625505168
transform 1 0 333400 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_65
timestamp 1625505168
transform 1 0 330400 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_66
timestamp 1625505168
transform 1 0 332400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_64
timestamp 1625505168
transform 1 0 326400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_70
timestamp 1625505168
transform 1 0 356400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_69
timestamp 1625505168
transform 1 0 352400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_68
timestamp 1625505168
transform 1 0 348400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_0
timestamp 1625505168
transform 1 0 372400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__disconnect_vccd_slice_5um  disconnect_vccd_0
timestamp 1625505168
transform 1 0 373400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_0
timestamp 1625505168
transform 1 0 374400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_73
timestamp 1625505168
transform 1 0 368400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_72
timestamp 1625505168
transform 1 0 364400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_71
timestamp 1625505168
transform 1 0 360400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__top_power_hvc  user1_analog_pad_with_clamp
timestamp 1625505168
transform 1 0 375400 0 1 998007
box 0 -407 33800 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_0
timestamp 1625505168
transform 1 0 410200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_1
timestamp 1625505168
transform 1 0 409200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_78
timestamp 1625505168
transform 1 0 412200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_79
timestamp 1625505168
transform 1 0 416200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_80
timestamp 1625505168
transform 1 0 420200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_81
timestamp 1625505168
transform 1 0 424200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_82
timestamp 1625505168
transform 1 0 428200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_83
timestamp 1625505168
transform 1 0 432200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_84
timestamp 1625505168
transform 1 0 436200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_85
timestamp 1625505168
transform 1 0 440200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_86
timestamp 1625505168
transform 1 0 444200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_87
timestamp 1625505168
transform 1 0 448200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_88
timestamp 1625505168
transform 1 0 452200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_89
timestamp 1625505168
transform 1 0 456200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_90
timestamp 1625505168
transform 1 0 460200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__analog_pad  user1_analog_pad\[2\]
timestamp 1625505168
transform 1 0 473800 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_5um  FILLER_93
timestamp 1625505168
transform 1 0 472200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_96
timestamp 1625505168
transform 1 0 473600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_95
timestamp 1625505168
transform 1 0 473400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_94
timestamp 1625505168
transform 1 0 473200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_92
timestamp 1625505168
transform 1 0 468200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_91
timestamp 1625505168
transform 1 0 464200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_99
timestamp 1625505168
transform 1 0 492800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_98
timestamp 1625505168
transform 1 0 488800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_102
timestamp 1625505168
transform 1 0 504800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_101
timestamp 1625505168
transform 1 0 500800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_100
timestamp 1625505168
transform 1 0 496800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_106
timestamp 1625505168
transform 1 0 520800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_105
timestamp 1625505168
transform 1 0 516800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_104
timestamp 1625505168
transform 1 0 512800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_103
timestamp 1625505168
transform 1 0 508800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__analog_pad  user1_analog_pad\[1\]
timestamp 1625505168
transform 1 0 525200 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_1um  FILLER_108
timestamp 1625505168
transform 1 0 525000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_107
timestamp 1625505168
transform 1 0 524800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_112
timestamp 1625505168
transform 1 0 548200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_111
timestamp 1625505168
transform 1 0 544200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_110
timestamp 1625505168
transform 1 0 540200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_115
timestamp 1625505168
transform 1 0 560200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_114
timestamp 1625505168
transform 1 0 556200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_113
timestamp 1625505168
transform 1 0 552200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user1_vssa_hvclamp_pad\[0\]
timestamp 1625505168
transform 1 0 575600 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_118
timestamp 1625505168
transform 1 0 572200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_119
timestamp 1625505168
transform 1 0 574200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_121
timestamp 1625505168
transform 1 0 575400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_120
timestamp 1625505168
transform 1 0 575200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_117
timestamp 1625505168
transform 1 0 568200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_116
timestamp 1625505168
transform 1 0 564200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_123
timestamp 1625505168
transform 1 0 590600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_126
timestamp 1625505168
transform 1 0 602600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_125
timestamp 1625505168
transform 1 0 598600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_124
timestamp 1625505168
transform 1 0 594600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_130
timestamp 1625505168
transform 1 0 618600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_129
timestamp 1625505168
transform 1 0 614600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_128
timestamp 1625505168
transform 1 0 610600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_127
timestamp 1625505168
transform 1 0 606600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__analog_pad  user1_analog_pad\[0\]
timestamp 1625505168
transform 1 0 627000 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_1um  FILLER_133
timestamp 1625505168
transform 1 0 626800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_132
timestamp 1625505168
transform 1 0 626600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_131
timestamp 1625505168
transform 1 0 622600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_143
timestamp 1625505168
transform 1 0 674000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_142
timestamp 1625505168
transform 1 0 670000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_141
timestamp 1625505168
transform 1 0 666000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_140
timestamp 1625505168
transform 1 0 662000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_139
timestamp 1625505168
transform 1 0 658000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_138
timestamp 1625505168
transform 1 0 654000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_137
timestamp 1625505168
transform 1 0 650000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_136
timestamp 1625505168
transform 1 0 646000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_135
timestamp 1625505168
transform 1 0 642000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_784
timestamp 1625505168
transform 0 1 678007 -1 0 992600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_783
timestamp 1625505168
transform 0 1 678007 -1 0 988600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_782
timestamp 1625505168
transform 0 1 678007 -1 0 984600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_781
timestamp 1625505168
transform 0 1 678007 -1 0 980600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_780
timestamp 1625505168
transform 0 1 678007 -1 0 976600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_786
timestamp 1625505168
transform 0 1 678007 -1 0 996800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_785
timestamp 1625505168
transform 0 1 678007 -1 0 996600
box 0 0 4000 39593
use sky130_ef_io__corner_pad  user1_corner
timestamp 1625505168
transform 1 0 677600 0 1 996800
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_5um  FILLER_144
timestamp 1625505168
transform 1 0 676000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_147
timestamp 1625505168
transform 1 0 677400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_146
timestamp 1625505168
transform 1 0 677200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_145
timestamp 1625505168
transform 1 0 677000 0 1 998007
box 0 0 200 39593
<< labels >>
rlabel metal5 s 187640 6598 200180 19088 6 clock
port 0 nsew signal input
rlabel metal2 s 187327 41713 187383 42193 6 clock_core
port 1 nsew signal tristate
rlabel metal2 s 194043 41713 194099 42193 6 por
port 2 nsew signal input
rlabel metal5 s 351040 6598 363580 19088 6 flash_clk
port 3 nsew signal tristate
rlabel metal5 s 296240 6598 308780 19088 6 flash_csb
port 7 nsew signal tristate
rlabel metal5 s 405840 6598 418380 19088 6 flash_io0
port 11 nsew signal bidirectional
rlabel metal2 s 405527 41713 405583 42193 6 flash_io0_di_core
port 12 nsew signal tristate
rlabel metal2 s 416567 41713 416623 42193 6 flash_io0_do_core
port 13 nsew signal input
rlabel metal2 s 412243 41713 412299 42193 6 flash_io0_ieb_core
port 14 nsew signal input
rlabel metal2 s 419695 41713 419751 42193 6 flash_io0_oeb_core
port 15 nsew signal input
rlabel metal5 s 460640 6598 473180 19088 6 flash_io1
port 16 nsew signal bidirectional
rlabel metal2 s 460327 41713 460383 42193 6 flash_io1_di_core
port 17 nsew signal tristate
rlabel metal2 s 471367 41713 471423 42193 6 flash_io1_do_core
port 18 nsew signal input
rlabel metal2 s 467043 41713 467099 42193 6 flash_io1_ieb_core
port 19 nsew signal input
rlabel metal2 s 474495 41713 474551 42193 6 flash_io1_oeb_core
port 20 nsew signal input
rlabel metal5 s 515440 6598 527980 19088 6 gpio
port 21 nsew signal bidirectional
rlabel metal2 s 515127 41713 515183 42193 6 gpio_in_core
port 22 nsew signal tristate
rlabel metal2 s 521843 41713 521899 42193 6 gpio_inenb_core
port 23 nsew signal input
rlabel metal2 s 520647 41713 520703 42193 6 gpio_mode0_core
port 24 nsew signal input
rlabel metal2 s 524971 41713 525027 42193 6 gpio_mode1_core
port 25 nsew signal input
rlabel metal2 s 526167 41713 526223 42193 6 gpio_out_core
port 26 nsew signal input
rlabel metal2 s 529295 41713 529351 42193 6 gpio_outenb_core
port 27 nsew signal input
rlabel metal5 s 6167 70054 19619 80934 6 vccd_pad
port 28 nsew signal bidirectional
rlabel metal5 s 624222 6811 636390 18975 6 vdda_pad
port 29 nsew signal bidirectional
rlabel metal5 s 6811 111610 18975 123778 6 vddio_pad
port 30 nsew signal bidirectional
rlabel metal5 s 6811 871210 18975 883378 6 vddio_pad2
port 31 nsew signal bidirectional
rlabel metal5 s 80222 6811 92390 18975 6 vssa_pad
port 32 nsew signal bidirectional
rlabel metal5 s 243266 6167 254146 19619 6 vssd_pad
port 33 nsew signal bidirectional
rlabel metal5 s 570422 6811 582590 18975 6 vssio_pad
port 34 nsew signal bidirectional
rlabel metal5 s 334810 1018624 346978 1030788 6 vssio_pad2
port 35 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113780 6 mprj_io[0]
port 36 nsew signal bidirectional
rlabel metal2 s 675407 105803 675887 105859 6 mprj_io_analog_en[0]
port 37 nsew signal input
rlabel metal2 s 675407 107091 675887 107147 6 mprj_io_analog_pol[0]
port 38 nsew signal input
rlabel metal2 s 675407 110127 675887 110183 6 mprj_io_analog_sel[0]
port 39 nsew signal input
rlabel metal2 s 675407 106447 675887 106503 6 mprj_io_dm[0]
port 40 nsew signal input
rlabel metal2 s 675407 104607 675887 104663 6 mprj_io_dm[1]
port 41 nsew signal input
rlabel metal2 s 675407 110771 675887 110827 6 mprj_io_dm[2]
port 42 nsew signal input
rlabel metal2 s 675407 111415 675887 111471 6 mprj_io_holdover[0]
port 43 nsew signal input
rlabel metal2 s 675407 114451 675887 114507 6 mprj_io_ib_mode_sel[0]
port 44 nsew signal input
rlabel metal2 s 675407 107643 675887 107699 6 mprj_io_inp_dis[0]
port 45 nsew signal input
rlabel metal2 s 675407 115095 675887 115151 6 mprj_io_oeb[0]
port 46 nsew signal input
rlabel metal2 s 675407 111967 675887 112023 6 mprj_io_out[0]
port 47 nsew signal input
rlabel metal2 s 675407 102767 675887 102823 6 mprj_io_slow_sel[0]
port 48 nsew signal input
rlabel metal2 s 675407 113807 675887 113863 6 mprj_io_vtrip_sel[0]
port 49 nsew signal input
rlabel metal2 s 675407 100927 675887 100983 6 mprj_io_in[0]
port 50 nsew signal tristate
rlabel metal2 s 675407 115647 675887 115703 6 mprj_io_in_3v3[0]
port 51 nsew signal tristate
rlabel metal2 s 675407 686611 675887 686667 6 mprj_gpio_analog[3]
port 52 nsew signal bidirectional
rlabel metal2 s 675407 688451 675887 688507 6 mprj_gpio_noesd[3]
port 53 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696980 6 mprj_io[10]
port 54 nsew signal bidirectional
rlabel metal2 s 675407 689003 675887 689059 6 mprj_io_analog_en[10]
port 55 nsew signal input
rlabel metal2 s 675407 690291 675887 690347 6 mprj_io_analog_pol[10]
port 56 nsew signal input
rlabel metal2 s 675407 693327 675887 693383 6 mprj_io_analog_sel[10]
port 57 nsew signal input
rlabel metal2 s 675407 689647 675887 689703 6 mprj_io_dm[30]
port 58 nsew signal input
rlabel metal2 s 675407 687807 675887 687863 6 mprj_io_dm[31]
port 59 nsew signal input
rlabel metal2 s 675407 693971 675887 694027 6 mprj_io_dm[32]
port 60 nsew signal input
rlabel metal2 s 675407 694615 675887 694671 6 mprj_io_holdover[10]
port 61 nsew signal input
rlabel metal2 s 675407 697651 675887 697707 6 mprj_io_ib_mode_sel[10]
port 62 nsew signal input
rlabel metal2 s 675407 690843 675887 690899 6 mprj_io_inp_dis[10]
port 63 nsew signal input
rlabel metal2 s 675407 698295 675887 698351 6 mprj_io_oeb[10]
port 64 nsew signal input
rlabel metal2 s 675407 695167 675887 695223 6 mprj_io_out[10]
port 65 nsew signal input
rlabel metal2 s 675407 685967 675887 686023 6 mprj_io_slow_sel[10]
port 66 nsew signal input
rlabel metal2 s 675407 697007 675887 697063 6 mprj_io_vtrip_sel[10]
port 67 nsew signal input
rlabel metal2 s 675407 684127 675887 684183 6 mprj_io_in[10]
port 68 nsew signal tristate
rlabel metal2 s 675407 698847 675887 698903 6 mprj_io_in_3v3[10]
port 69 nsew signal tristate
rlabel metal2 s 675407 731611 675887 731667 6 mprj_gpio_analog[4]
port 70 nsew signal bidirectional
rlabel metal2 s 675407 733451 675887 733507 6 mprj_gpio_noesd[4]
port 71 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741980 6 mprj_io[11]
port 72 nsew signal bidirectional
rlabel metal2 s 675407 734003 675887 734059 6 mprj_io_analog_en[11]
port 73 nsew signal input
rlabel metal2 s 675407 735291 675887 735347 6 mprj_io_analog_pol[11]
port 74 nsew signal input
rlabel metal2 s 675407 738327 675887 738383 6 mprj_io_analog_sel[11]
port 75 nsew signal input
rlabel metal2 s 675407 734647 675887 734703 6 mprj_io_dm[33]
port 76 nsew signal input
rlabel metal2 s 675407 732807 675887 732863 6 mprj_io_dm[34]
port 77 nsew signal input
rlabel metal2 s 675407 738971 675887 739027 6 mprj_io_dm[35]
port 78 nsew signal input
rlabel metal2 s 675407 739615 675887 739671 6 mprj_io_holdover[11]
port 79 nsew signal input
rlabel metal2 s 675407 742651 675887 742707 6 mprj_io_ib_mode_sel[11]
port 80 nsew signal input
rlabel metal2 s 675407 735843 675887 735899 6 mprj_io_inp_dis[11]
port 81 nsew signal input
rlabel metal2 s 675407 743295 675887 743351 6 mprj_io_oeb[11]
port 82 nsew signal input
rlabel metal2 s 675407 740167 675887 740223 6 mprj_io_out[11]
port 83 nsew signal input
rlabel metal2 s 675407 730967 675887 731023 6 mprj_io_slow_sel[11]
port 84 nsew signal input
rlabel metal2 s 675407 742007 675887 742063 6 mprj_io_vtrip_sel[11]
port 85 nsew signal input
rlabel metal2 s 675407 729127 675887 729183 6 mprj_io_in[11]
port 86 nsew signal tristate
rlabel metal2 s 675407 743847 675887 743903 6 mprj_io_in_3v3[11]
port 87 nsew signal tristate
rlabel metal2 s 675407 776611 675887 776667 6 mprj_gpio_analog[5]
port 88 nsew signal bidirectional
rlabel metal2 s 675407 778451 675887 778507 6 mprj_gpio_noesd[5]
port 89 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786980 6 mprj_io[12]
port 90 nsew signal bidirectional
rlabel metal2 s 675407 779003 675887 779059 6 mprj_io_analog_en[12]
port 91 nsew signal input
rlabel metal2 s 675407 780291 675887 780347 6 mprj_io_analog_pol[12]
port 92 nsew signal input
rlabel metal2 s 675407 783327 675887 783383 6 mprj_io_analog_sel[12]
port 93 nsew signal input
rlabel metal2 s 675407 779647 675887 779703 6 mprj_io_dm[36]
port 94 nsew signal input
rlabel metal2 s 675407 777807 675887 777863 6 mprj_io_dm[37]
port 95 nsew signal input
rlabel metal2 s 675407 783971 675887 784027 6 mprj_io_dm[38]
port 96 nsew signal input
rlabel metal2 s 675407 784615 675887 784671 6 mprj_io_holdover[12]
port 97 nsew signal input
rlabel metal2 s 675407 787651 675887 787707 6 mprj_io_ib_mode_sel[12]
port 98 nsew signal input
rlabel metal2 s 675407 780843 675887 780899 6 mprj_io_inp_dis[12]
port 99 nsew signal input
rlabel metal2 s 675407 788295 675887 788351 6 mprj_io_oeb[12]
port 100 nsew signal input
rlabel metal2 s 675407 785167 675887 785223 6 mprj_io_out[12]
port 101 nsew signal input
rlabel metal2 s 675407 775967 675887 776023 6 mprj_io_slow_sel[12]
port 102 nsew signal input
rlabel metal2 s 675407 787007 675887 787063 6 mprj_io_vtrip_sel[12]
port 103 nsew signal input
rlabel metal2 s 675407 774127 675887 774183 6 mprj_io_in[12]
port 104 nsew signal tristate
rlabel metal2 s 675407 788847 675887 788903 6 mprj_io_in_3v3[12]
port 105 nsew signal tristate
rlabel metal2 s 675407 865811 675887 865867 6 mprj_gpio_analog[6]
port 106 nsew signal bidirectional
rlabel metal2 s 675407 867651 675887 867707 6 mprj_gpio_noesd[6]
port 107 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876180 6 mprj_io[13]
port 108 nsew signal bidirectional
rlabel metal2 s 675407 868203 675887 868259 6 mprj_io_analog_en[13]
port 109 nsew signal input
rlabel metal2 s 675407 869491 675887 869547 6 mprj_io_analog_pol[13]
port 110 nsew signal input
rlabel metal2 s 675407 872527 675887 872583 6 mprj_io_analog_sel[13]
port 111 nsew signal input
rlabel metal2 s 675407 868847 675887 868903 6 mprj_io_dm[39]
port 112 nsew signal input
rlabel metal2 s 675407 867007 675887 867063 6 mprj_io_dm[40]
port 113 nsew signal input
rlabel metal2 s 675407 873171 675887 873227 6 mprj_io_dm[41]
port 114 nsew signal input
rlabel metal2 s 675407 873815 675887 873871 6 mprj_io_holdover[13]
port 115 nsew signal input
rlabel metal2 s 675407 876851 675887 876907 6 mprj_io_ib_mode_sel[13]
port 116 nsew signal input
rlabel metal2 s 675407 870043 675887 870099 6 mprj_io_inp_dis[13]
port 117 nsew signal input
rlabel metal2 s 675407 877495 675887 877551 6 mprj_io_oeb[13]
port 118 nsew signal input
rlabel metal2 s 675407 874367 675887 874423 6 mprj_io_out[13]
port 119 nsew signal input
rlabel metal2 s 675407 865167 675887 865223 6 mprj_io_slow_sel[13]
port 120 nsew signal input
rlabel metal2 s 675407 876207 675887 876263 6 mprj_io_vtrip_sel[13]
port 121 nsew signal input
rlabel metal2 s 675407 863327 675887 863383 6 mprj_io_in[13]
port 122 nsew signal tristate
rlabel metal2 s 675407 878047 675887 878103 6 mprj_io_in_3v3[13]
port 123 nsew signal tristate
rlabel metal5 s 698512 146440 711002 158980 6 mprj_io[1]
port 124 nsew signal bidirectional
rlabel metal2 s 675407 151003 675887 151059 6 mprj_io_analog_en[1]
port 125 nsew signal input
rlabel metal2 s 675407 152291 675887 152347 6 mprj_io_analog_pol[1]
port 126 nsew signal input
rlabel metal2 s 675407 155327 675887 155383 6 mprj_io_analog_sel[1]
port 127 nsew signal input
rlabel metal2 s 675407 151647 675887 151703 6 mprj_io_dm[3]
port 128 nsew signal input
rlabel metal2 s 675407 149807 675887 149863 6 mprj_io_dm[4]
port 129 nsew signal input
rlabel metal2 s 675407 155971 675887 156027 6 mprj_io_dm[5]
port 130 nsew signal input
rlabel metal2 s 675407 156615 675887 156671 6 mprj_io_holdover[1]
port 131 nsew signal input
rlabel metal2 s 675407 159651 675887 159707 6 mprj_io_ib_mode_sel[1]
port 132 nsew signal input
rlabel metal2 s 675407 152843 675887 152899 6 mprj_io_inp_dis[1]
port 133 nsew signal input
rlabel metal2 s 675407 160295 675887 160351 6 mprj_io_oeb[1]
port 134 nsew signal input
rlabel metal2 s 675407 157167 675887 157223 6 mprj_io_out[1]
port 135 nsew signal input
rlabel metal2 s 675407 147967 675887 148023 6 mprj_io_slow_sel[1]
port 136 nsew signal input
rlabel metal2 s 675407 159007 675887 159063 6 mprj_io_vtrip_sel[1]
port 137 nsew signal input
rlabel metal2 s 675407 146127 675887 146183 6 mprj_io_in[1]
port 138 nsew signal tristate
rlabel metal2 s 675407 160847 675887 160903 6 mprj_io_in_3v3[1]
port 139 nsew signal tristate
rlabel metal5 s 698512 191440 711002 203980 6 mprj_io[2]
port 140 nsew signal bidirectional
rlabel metal2 s 675407 196003 675887 196059 6 mprj_io_analog_en[2]
port 141 nsew signal input
rlabel metal2 s 675407 197291 675887 197347 6 mprj_io_analog_pol[2]
port 142 nsew signal input
rlabel metal2 s 675407 200327 675887 200383 6 mprj_io_analog_sel[2]
port 143 nsew signal input
rlabel metal2 s 675407 196647 675887 196703 6 mprj_io_dm[6]
port 144 nsew signal input
rlabel metal2 s 675407 194807 675887 194863 6 mprj_io_dm[7]
port 145 nsew signal input
rlabel metal2 s 675407 200971 675887 201027 6 mprj_io_dm[8]
port 146 nsew signal input
rlabel metal2 s 675407 201615 675887 201671 6 mprj_io_holdover[2]
port 147 nsew signal input
rlabel metal2 s 675407 204651 675887 204707 6 mprj_io_ib_mode_sel[2]
port 148 nsew signal input
rlabel metal2 s 675407 197843 675887 197899 6 mprj_io_inp_dis[2]
port 149 nsew signal input
rlabel metal2 s 675407 205295 675887 205351 6 mprj_io_oeb[2]
port 150 nsew signal input
rlabel metal2 s 675407 202167 675887 202223 6 mprj_io_out[2]
port 151 nsew signal input
rlabel metal2 s 675407 192967 675887 193023 6 mprj_io_slow_sel[2]
port 152 nsew signal input
rlabel metal2 s 675407 204007 675887 204063 6 mprj_io_vtrip_sel[2]
port 153 nsew signal input
rlabel metal2 s 675407 191127 675887 191183 6 mprj_io_in[2]
port 154 nsew signal tristate
rlabel metal2 s 675407 205847 675887 205903 6 mprj_io_in_3v3[2]
port 155 nsew signal tristate
rlabel metal5 s 698512 236640 711002 249180 6 mprj_io[3]
port 156 nsew signal bidirectional
rlabel metal2 s 675407 241203 675887 241259 6 mprj_io_analog_en[3]
port 157 nsew signal input
rlabel metal2 s 675407 242491 675887 242547 6 mprj_io_analog_pol[3]
port 158 nsew signal input
rlabel metal2 s 675407 245527 675887 245583 6 mprj_io_analog_sel[3]
port 159 nsew signal input
rlabel metal2 s 675407 240007 675887 240063 6 mprj_io_dm[10]
port 160 nsew signal input
rlabel metal2 s 675407 246171 675887 246227 6 mprj_io_dm[11]
port 161 nsew signal input
rlabel metal2 s 675407 241847 675887 241903 6 mprj_io_dm[9]
port 162 nsew signal input
rlabel metal2 s 675407 246815 675887 246871 6 mprj_io_holdover[3]
port 163 nsew signal input
rlabel metal2 s 675407 249851 675887 249907 6 mprj_io_ib_mode_sel[3]
port 164 nsew signal input
rlabel metal2 s 675407 243043 675887 243099 6 mprj_io_inp_dis[3]
port 165 nsew signal input
rlabel metal2 s 675407 250495 675887 250551 6 mprj_io_oeb[3]
port 166 nsew signal input
rlabel metal2 s 675407 247367 675887 247423 6 mprj_io_out[3]
port 167 nsew signal input
rlabel metal2 s 675407 238167 675887 238223 6 mprj_io_slow_sel[3]
port 168 nsew signal input
rlabel metal2 s 675407 249207 675887 249263 6 mprj_io_vtrip_sel[3]
port 169 nsew signal input
rlabel metal2 s 675407 236327 675887 236383 6 mprj_io_in[3]
port 170 nsew signal tristate
rlabel metal2 s 675407 251047 675887 251103 6 mprj_io_in_3v3[3]
port 171 nsew signal tristate
rlabel metal5 s 698512 281640 711002 294180 6 mprj_io[4]
port 172 nsew signal bidirectional
rlabel metal2 s 675407 286203 675887 286259 6 mprj_io_analog_en[4]
port 173 nsew signal input
rlabel metal2 s 675407 287491 675887 287547 6 mprj_io_analog_pol[4]
port 174 nsew signal input
rlabel metal2 s 675407 290527 675887 290583 6 mprj_io_analog_sel[4]
port 175 nsew signal input
rlabel metal2 s 675407 286847 675887 286903 6 mprj_io_dm[12]
port 176 nsew signal input
rlabel metal2 s 675407 285007 675887 285063 6 mprj_io_dm[13]
port 177 nsew signal input
rlabel metal2 s 675407 291171 675887 291227 6 mprj_io_dm[14]
port 178 nsew signal input
rlabel metal2 s 675407 291815 675887 291871 6 mprj_io_holdover[4]
port 179 nsew signal input
rlabel metal2 s 675407 294851 675887 294907 6 mprj_io_ib_mode_sel[4]
port 180 nsew signal input
rlabel metal2 s 675407 288043 675887 288099 6 mprj_io_inp_dis[4]
port 181 nsew signal input
rlabel metal2 s 675407 295495 675887 295551 6 mprj_io_oeb[4]
port 182 nsew signal input
rlabel metal2 s 675407 292367 675887 292423 6 mprj_io_out[4]
port 183 nsew signal input
rlabel metal2 s 675407 283167 675887 283223 6 mprj_io_slow_sel[4]
port 184 nsew signal input
rlabel metal2 s 675407 294207 675887 294263 6 mprj_io_vtrip_sel[4]
port 185 nsew signal input
rlabel metal2 s 675407 281327 675887 281383 6 mprj_io_in[4]
port 186 nsew signal tristate
rlabel metal2 s 675407 296047 675887 296103 6 mprj_io_in_3v3[4]
port 187 nsew signal tristate
rlabel metal5 s 698512 326640 711002 339180 6 mprj_io[5]
port 188 nsew signal bidirectional
rlabel metal2 s 675407 331203 675887 331259 6 mprj_io_analog_en[5]
port 189 nsew signal input
rlabel metal2 s 675407 332491 675887 332547 6 mprj_io_analog_pol[5]
port 190 nsew signal input
rlabel metal2 s 675407 335527 675887 335583 6 mprj_io_analog_sel[5]
port 191 nsew signal input
rlabel metal2 s 675407 331847 675887 331903 6 mprj_io_dm[15]
port 192 nsew signal input
rlabel metal2 s 675407 330007 675887 330063 6 mprj_io_dm[16]
port 193 nsew signal input
rlabel metal2 s 675407 336171 675887 336227 6 mprj_io_dm[17]
port 194 nsew signal input
rlabel metal2 s 675407 336815 675887 336871 6 mprj_io_holdover[5]
port 195 nsew signal input
rlabel metal2 s 675407 339851 675887 339907 6 mprj_io_ib_mode_sel[5]
port 196 nsew signal input
rlabel metal2 s 675407 333043 675887 333099 6 mprj_io_inp_dis[5]
port 197 nsew signal input
rlabel metal2 s 675407 340495 675887 340551 6 mprj_io_oeb[5]
port 198 nsew signal input
rlabel metal2 s 675407 337367 675887 337423 6 mprj_io_out[5]
port 199 nsew signal input
rlabel metal2 s 675407 328167 675887 328223 6 mprj_io_slow_sel[5]
port 200 nsew signal input
rlabel metal2 s 675407 339207 675887 339263 6 mprj_io_vtrip_sel[5]
port 201 nsew signal input
rlabel metal2 s 675407 326327 675887 326383 6 mprj_io_in[5]
port 202 nsew signal tristate
rlabel metal2 s 675407 341047 675887 341103 6 mprj_io_in_3v3[5]
port 203 nsew signal tristate
rlabel metal5 s 698512 371840 711002 384380 6 mprj_io[6]
port 204 nsew signal bidirectional
rlabel metal2 s 675407 376403 675887 376459 6 mprj_io_analog_en[6]
port 205 nsew signal input
rlabel metal2 s 675407 377691 675887 377747 6 mprj_io_analog_pol[6]
port 206 nsew signal input
rlabel metal2 s 675407 380727 675887 380783 6 mprj_io_analog_sel[6]
port 207 nsew signal input
rlabel metal2 s 675407 377047 675887 377103 6 mprj_io_dm[18]
port 208 nsew signal input
rlabel metal2 s 675407 375207 675887 375263 6 mprj_io_dm[19]
port 209 nsew signal input
rlabel metal2 s 675407 381371 675887 381427 6 mprj_io_dm[20]
port 210 nsew signal input
rlabel metal2 s 675407 382015 675887 382071 6 mprj_io_holdover[6]
port 211 nsew signal input
rlabel metal2 s 675407 385051 675887 385107 6 mprj_io_ib_mode_sel[6]
port 212 nsew signal input
rlabel metal2 s 675407 378243 675887 378299 6 mprj_io_inp_dis[6]
port 213 nsew signal input
rlabel metal2 s 675407 385695 675887 385751 6 mprj_io_oeb[6]
port 214 nsew signal input
rlabel metal2 s 675407 382567 675887 382623 6 mprj_io_out[6]
port 215 nsew signal input
rlabel metal2 s 675407 373367 675887 373423 6 mprj_io_slow_sel[6]
port 216 nsew signal input
rlabel metal2 s 675407 384407 675887 384463 6 mprj_io_vtrip_sel[6]
port 217 nsew signal input
rlabel metal2 s 675407 371527 675887 371583 6 mprj_io_in[6]
port 218 nsew signal tristate
rlabel metal2 s 675407 386247 675887 386303 6 mprj_io_in_3v3[6]
port 219 nsew signal tristate
rlabel metal2 s 675407 551211 675887 551267 6 mprj_gpio_analog[0]
port 220 nsew signal bidirectional
rlabel metal2 s 675407 553051 675887 553107 6 mprj_gpio_noesd[0]
port 221 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561580 6 mprj_io[7]
port 222 nsew signal bidirectional
rlabel metal2 s 675407 553603 675887 553659 6 mprj_io_analog_en[7]
port 223 nsew signal input
rlabel metal2 s 675407 554891 675887 554947 6 mprj_io_analog_pol[7]
port 224 nsew signal input
rlabel metal2 s 675407 557927 675887 557983 6 mprj_io_analog_sel[7]
port 225 nsew signal input
rlabel metal2 s 675407 554247 675887 554303 6 mprj_io_dm[21]
port 226 nsew signal input
rlabel metal2 s 675407 552407 675887 552463 6 mprj_io_dm[22]
port 227 nsew signal input
rlabel metal2 s 675407 558571 675887 558627 6 mprj_io_dm[23]
port 228 nsew signal input
rlabel metal2 s 675407 559215 675887 559271 6 mprj_io_holdover[7]
port 229 nsew signal input
rlabel metal2 s 675407 562251 675887 562307 6 mprj_io_ib_mode_sel[7]
port 230 nsew signal input
rlabel metal2 s 675407 555443 675887 555499 6 mprj_io_inp_dis[7]
port 231 nsew signal input
rlabel metal2 s 675407 562895 675887 562951 6 mprj_io_oeb[7]
port 232 nsew signal input
rlabel metal2 s 675407 559767 675887 559823 6 mprj_io_out[7]
port 233 nsew signal input
rlabel metal2 s 675407 550567 675887 550623 6 mprj_io_slow_sel[7]
port 234 nsew signal input
rlabel metal2 s 675407 561607 675887 561663 6 mprj_io_vtrip_sel[7]
port 235 nsew signal input
rlabel metal2 s 675407 548727 675887 548783 6 mprj_io_in[7]
port 236 nsew signal tristate
rlabel metal2 s 675407 563447 675887 563503 6 mprj_io_in_3v3[7]
port 237 nsew signal tristate
rlabel metal2 s 675407 596411 675887 596467 6 mprj_gpio_analog[1]
port 238 nsew signal bidirectional
rlabel metal2 s 675407 598251 675887 598307 6 mprj_gpio_noesd[1]
port 239 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606780 6 mprj_io[8]
port 240 nsew signal bidirectional
rlabel metal2 s 675407 598803 675887 598859 6 mprj_io_analog_en[8]
port 241 nsew signal input
rlabel metal2 s 675407 600091 675887 600147 6 mprj_io_analog_pol[8]
port 242 nsew signal input
rlabel metal2 s 675407 603127 675887 603183 6 mprj_io_analog_sel[8]
port 243 nsew signal input
rlabel metal2 s 675407 599447 675887 599503 6 mprj_io_dm[24]
port 244 nsew signal input
rlabel metal2 s 675407 597607 675887 597663 6 mprj_io_dm[25]
port 245 nsew signal input
rlabel metal2 s 675407 603771 675887 603827 6 mprj_io_dm[26]
port 246 nsew signal input
rlabel metal2 s 675407 604415 675887 604471 6 mprj_io_holdover[8]
port 247 nsew signal input
rlabel metal2 s 675407 607451 675887 607507 6 mprj_io_ib_mode_sel[8]
port 248 nsew signal input
rlabel metal2 s 675407 600643 675887 600699 6 mprj_io_inp_dis[8]
port 249 nsew signal input
rlabel metal2 s 675407 608095 675887 608151 6 mprj_io_oeb[8]
port 250 nsew signal input
rlabel metal2 s 675407 604967 675887 605023 6 mprj_io_out[8]
port 251 nsew signal input
rlabel metal2 s 675407 595767 675887 595823 6 mprj_io_slow_sel[8]
port 252 nsew signal input
rlabel metal2 s 675407 606807 675887 606863 6 mprj_io_vtrip_sel[8]
port 253 nsew signal input
rlabel metal2 s 675407 593927 675887 593983 6 mprj_io_in[8]
port 254 nsew signal tristate
rlabel metal2 s 675407 608647 675887 608703 6 mprj_io_in_3v3[8]
port 255 nsew signal tristate
rlabel metal2 s 675407 641411 675887 641467 6 mprj_gpio_analog[2]
port 256 nsew signal bidirectional
rlabel metal2 s 675407 643251 675887 643307 6 mprj_gpio_noesd[2]
port 257 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651780 6 mprj_io[9]
port 258 nsew signal bidirectional
rlabel metal2 s 675407 643803 675887 643859 6 mprj_io_analog_en[9]
port 259 nsew signal input
rlabel metal2 s 675407 645091 675887 645147 6 mprj_io_analog_pol[9]
port 260 nsew signal input
rlabel metal2 s 675407 648127 675887 648183 6 mprj_io_analog_sel[9]
port 261 nsew signal input
rlabel metal2 s 675407 644447 675887 644503 6 mprj_io_dm[27]
port 262 nsew signal input
rlabel metal2 s 675407 642607 675887 642663 6 mprj_io_dm[28]
port 263 nsew signal input
rlabel metal2 s 675407 648771 675887 648827 6 mprj_io_dm[29]
port 264 nsew signal input
rlabel metal2 s 675407 649415 675887 649471 6 mprj_io_holdover[9]
port 265 nsew signal input
rlabel metal2 s 675407 652451 675887 652507 6 mprj_io_ib_mode_sel[9]
port 266 nsew signal input
rlabel metal2 s 675407 645643 675887 645699 6 mprj_io_inp_dis[9]
port 267 nsew signal input
rlabel metal2 s 675407 653095 675887 653151 6 mprj_io_oeb[9]
port 268 nsew signal input
rlabel metal2 s 675407 649967 675887 650023 6 mprj_io_out[9]
port 269 nsew signal input
rlabel metal2 s 675407 640767 675887 640823 6 mprj_io_slow_sel[9]
port 270 nsew signal input
rlabel metal2 s 675407 651807 675887 651863 6 mprj_io_vtrip_sel[9]
port 271 nsew signal input
rlabel metal2 s 675407 638927 675887 638983 6 mprj_io_in[9]
port 272 nsew signal tristate
rlabel metal2 s 675407 653647 675887 653703 6 mprj_io_in_3v3[9]
port 273 nsew signal tristate
rlabel metal2 s 41713 796933 42193 796989 6 mprj_gpio_analog[7]
port 274 nsew signal bidirectional
rlabel metal2 s 41713 795093 42193 795149 6 mprj_gpio_noesd[7]
port 275 nsew signal bidirectional
rlabel metal5 s 6598 786620 19088 799160 6 mprj_io[25]
port 276 nsew signal bidirectional
rlabel metal2 s 41713 794541 42193 794597 6 mprj_io_analog_en[14]
port 277 nsew signal input
rlabel metal2 s 41713 793253 42193 793309 6 mprj_io_analog_pol[14]
port 278 nsew signal input
rlabel metal2 s 41713 790217 42193 790273 6 mprj_io_analog_sel[14]
port 279 nsew signal input
rlabel metal2 s 41713 793897 42193 793953 6 mprj_io_dm[42]
port 280 nsew signal input
rlabel metal2 s 41713 795737 42193 795793 6 mprj_io_dm[43]
port 281 nsew signal input
rlabel metal2 s 41713 789573 42193 789629 6 mprj_io_dm[44]
port 282 nsew signal input
rlabel metal2 s 41713 788929 42193 788985 6 mprj_io_holdover[14]
port 283 nsew signal input
rlabel metal2 s 41713 785893 42193 785949 6 mprj_io_ib_mode_sel[14]
port 284 nsew signal input
rlabel metal2 s 41713 792701 42193 792757 6 mprj_io_inp_dis[14]
port 285 nsew signal input
rlabel metal2 s 41713 785249 42193 785305 6 mprj_io_oeb[14]
port 286 nsew signal input
rlabel metal2 s 41713 788377 42193 788433 6 mprj_io_out[14]
port 287 nsew signal input
rlabel metal2 s 41713 797577 42193 797633 6 mprj_io_slow_sel[14]
port 288 nsew signal input
rlabel metal2 s 41713 786537 42193 786593 6 mprj_io_vtrip_sel[14]
port 289 nsew signal input
rlabel metal2 s 41713 799417 42193 799473 6 mprj_io_in[14]
port 290 nsew signal tristate
rlabel metal2 s 41713 784697 42193 784753 6 mprj_io_in_3v3[14]
port 291 nsew signal tristate
rlabel metal2 s 41713 280533 42193 280589 6 mprj_gpio_analog[17]
port 292 nsew signal bidirectional
rlabel metal2 s 41713 278693 42193 278749 6 mprj_gpio_noesd[17]
port 293 nsew signal bidirectional
rlabel metal5 s 6598 270220 19088 282760 6 mprj_io[35]
port 294 nsew signal bidirectional
rlabel metal2 s 41713 278141 42193 278197 6 mprj_io_analog_en[24]
port 295 nsew signal input
rlabel metal2 s 41713 276853 42193 276909 6 mprj_io_analog_pol[24]
port 296 nsew signal input
rlabel metal2 s 41713 273817 42193 273873 6 mprj_io_analog_sel[24]
port 297 nsew signal input
rlabel metal2 s 41713 277497 42193 277553 6 mprj_io_dm[72]
port 298 nsew signal input
rlabel metal2 s 41713 279337 42193 279393 6 mprj_io_dm[73]
port 299 nsew signal input
rlabel metal2 s 41713 273173 42193 273229 6 mprj_io_dm[74]
port 300 nsew signal input
rlabel metal2 s 41713 272529 42193 272585 6 mprj_io_holdover[24]
port 301 nsew signal input
rlabel metal2 s 41713 269493 42193 269549 6 mprj_io_ib_mode_sel[24]
port 302 nsew signal input
rlabel metal2 s 41713 276301 42193 276357 6 mprj_io_inp_dis[24]
port 303 nsew signal input
rlabel metal2 s 41713 268849 42193 268905 6 mprj_io_oeb[24]
port 304 nsew signal input
rlabel metal2 s 41713 271977 42193 272033 6 mprj_io_out[24]
port 305 nsew signal input
rlabel metal2 s 41713 281177 42193 281233 6 mprj_io_slow_sel[24]
port 306 nsew signal input
rlabel metal2 s 41713 270137 42193 270193 6 mprj_io_vtrip_sel[24]
port 307 nsew signal input
rlabel metal2 s 41713 283017 42193 283073 6 mprj_io_in[24]
port 308 nsew signal tristate
rlabel metal2 s 41713 268297 42193 268353 6 mprj_io_in_3v3[24]
port 309 nsew signal tristate
rlabel metal5 s 6598 227020 19088 239560 6 mprj_io[36]
port 310 nsew signal bidirectional
rlabel metal2 s 41713 234941 42193 234997 6 mprj_io_analog_en[25]
port 311 nsew signal input
rlabel metal2 s 41713 233653 42193 233709 6 mprj_io_analog_pol[25]
port 312 nsew signal input
rlabel metal2 s 41713 230617 42193 230673 6 mprj_io_analog_sel[25]
port 313 nsew signal input
rlabel metal2 s 41713 234297 42193 234353 6 mprj_io_dm[75]
port 314 nsew signal input
rlabel metal2 s 41713 236137 42193 236193 6 mprj_io_dm[76]
port 315 nsew signal input
rlabel metal2 s 41713 229973 42193 230029 6 mprj_io_dm[77]
port 316 nsew signal input
rlabel metal2 s 41713 229329 42193 229385 6 mprj_io_holdover[25]
port 317 nsew signal input
rlabel metal2 s 41713 226293 42193 226349 6 mprj_io_ib_mode_sel[25]
port 318 nsew signal input
rlabel metal2 s 41713 233101 42193 233157 6 mprj_io_inp_dis[25]
port 319 nsew signal input
rlabel metal2 s 41713 225649 42193 225705 6 mprj_io_oeb[25]
port 320 nsew signal input
rlabel metal2 s 41713 228777 42193 228833 6 mprj_io_out[25]
port 321 nsew signal input
rlabel metal2 s 41713 237977 42193 238033 6 mprj_io_slow_sel[25]
port 322 nsew signal input
rlabel metal2 s 41713 226937 42193 226993 6 mprj_io_vtrip_sel[25]
port 323 nsew signal input
rlabel metal2 s 41713 239817 42193 239873 6 mprj_io_in[25]
port 324 nsew signal tristate
rlabel metal2 s 41713 225097 42193 225153 6 mprj_io_in_3v3[25]
port 325 nsew signal tristate
rlabel metal5 s 6598 183820 19088 196360 6 mprj_io[37]
port 326 nsew signal bidirectional
rlabel metal2 s 41713 191741 42193 191797 6 mprj_io_analog_en[26]
port 327 nsew signal input
rlabel metal2 s 41713 190453 42193 190509 6 mprj_io_analog_pol[26]
port 328 nsew signal input
rlabel metal2 s 41713 187417 42193 187473 6 mprj_io_analog_sel[26]
port 329 nsew signal input
rlabel metal2 s 41713 191097 42193 191153 6 mprj_io_dm[78]
port 330 nsew signal input
rlabel metal2 s 41713 192937 42193 192993 6 mprj_io_dm[79]
port 331 nsew signal input
rlabel metal2 s 41713 186773 42193 186829 6 mprj_io_dm[80]
port 332 nsew signal input
rlabel metal2 s 41713 186129 42193 186185 6 mprj_io_holdover[26]
port 333 nsew signal input
rlabel metal2 s 41713 183093 42193 183149 6 mprj_io_ib_mode_sel[26]
port 334 nsew signal input
rlabel metal2 s 41713 189901 42193 189957 6 mprj_io_inp_dis[26]
port 335 nsew signal input
rlabel metal2 s 41713 182449 42193 182505 6 mprj_io_oeb[26]
port 336 nsew signal input
rlabel metal2 s 41713 185577 42193 185633 6 mprj_io_out[26]
port 337 nsew signal input
rlabel metal2 s 41713 194777 42193 194833 6 mprj_io_slow_sel[26]
port 338 nsew signal input
rlabel metal2 s 41713 183737 42193 183793 6 mprj_io_vtrip_sel[26]
port 339 nsew signal input
rlabel metal2 s 41713 196617 42193 196673 6 mprj_io_in[26]
port 340 nsew signal tristate
rlabel metal2 s 41713 181897 42193 181953 6 mprj_io_in_3v3[26]
port 341 nsew signal tristate
rlabel metal2 s 41713 753733 42193 753789 6 mprj_gpio_analog[8]
port 342 nsew signal bidirectional
rlabel metal2 s 41713 751893 42193 751949 6 mprj_gpio_noesd[8]
port 343 nsew signal bidirectional
rlabel metal5 s 6598 743420 19088 755960 6 mprj_io[26]
port 344 nsew signal bidirectional
rlabel metal2 s 41713 751341 42193 751397 6 mprj_io_analog_en[15]
port 345 nsew signal input
rlabel metal2 s 41713 750053 42193 750109 6 mprj_io_analog_pol[15]
port 346 nsew signal input
rlabel metal2 s 41713 747017 42193 747073 6 mprj_io_analog_sel[15]
port 347 nsew signal input
rlabel metal2 s 41713 750697 42193 750753 6 mprj_io_dm[45]
port 348 nsew signal input
rlabel metal2 s 41713 752537 42193 752593 6 mprj_io_dm[46]
port 349 nsew signal input
rlabel metal2 s 41713 746373 42193 746429 6 mprj_io_dm[47]
port 350 nsew signal input
rlabel metal2 s 41713 745729 42193 745785 6 mprj_io_holdover[15]
port 351 nsew signal input
rlabel metal2 s 41713 742693 42193 742749 6 mprj_io_ib_mode_sel[15]
port 352 nsew signal input
rlabel metal2 s 41713 749501 42193 749557 6 mprj_io_inp_dis[15]
port 353 nsew signal input
rlabel metal2 s 41713 742049 42193 742105 6 mprj_io_oeb[15]
port 354 nsew signal input
rlabel metal2 s 41713 745177 42193 745233 6 mprj_io_out[15]
port 355 nsew signal input
rlabel metal2 s 41713 754377 42193 754433 6 mprj_io_slow_sel[15]
port 356 nsew signal input
rlabel metal2 s 41713 743337 42193 743393 6 mprj_io_vtrip_sel[15]
port 357 nsew signal input
rlabel metal2 s 41713 756217 42193 756273 6 mprj_io_in[15]
port 358 nsew signal tristate
rlabel metal2 s 41713 741497 42193 741553 6 mprj_io_in_3v3[15]
port 359 nsew signal tristate
rlabel metal2 s 41713 710533 42193 710589 6 mprj_gpio_analog[9]
port 360 nsew signal bidirectional
rlabel metal2 s 41713 708693 42193 708749 6 mprj_gpio_noesd[9]
port 361 nsew signal bidirectional
rlabel metal5 s 6598 700220 19088 712760 6 mprj_io[27]
port 362 nsew signal bidirectional
rlabel metal2 s 41713 708141 42193 708197 6 mprj_io_analog_en[16]
port 363 nsew signal input
rlabel metal2 s 41713 706853 42193 706909 6 mprj_io_analog_pol[16]
port 364 nsew signal input
rlabel metal2 s 41713 703817 42193 703873 6 mprj_io_analog_sel[16]
port 365 nsew signal input
rlabel metal2 s 41713 707497 42193 707553 6 mprj_io_dm[48]
port 366 nsew signal input
rlabel metal2 s 41713 709337 42193 709393 6 mprj_io_dm[49]
port 367 nsew signal input
rlabel metal2 s 41713 703173 42193 703229 6 mprj_io_dm[50]
port 368 nsew signal input
rlabel metal2 s 41713 702529 42193 702585 6 mprj_io_holdover[16]
port 369 nsew signal input
rlabel metal2 s 41713 699493 42193 699549 6 mprj_io_ib_mode_sel[16]
port 370 nsew signal input
rlabel metal2 s 41713 706301 42193 706357 6 mprj_io_inp_dis[16]
port 371 nsew signal input
rlabel metal2 s 41713 698849 42193 698905 6 mprj_io_oeb[16]
port 372 nsew signal input
rlabel metal2 s 41713 701977 42193 702033 6 mprj_io_out[16]
port 373 nsew signal input
rlabel metal2 s 41713 711177 42193 711233 6 mprj_io_slow_sel[16]
port 374 nsew signal input
rlabel metal2 s 41713 700137 42193 700193 6 mprj_io_vtrip_sel[16]
port 375 nsew signal input
rlabel metal2 s 41713 713017 42193 713073 6 mprj_io_in[16]
port 376 nsew signal tristate
rlabel metal2 s 41713 698297 42193 698353 6 mprj_io_in_3v3[16]
port 377 nsew signal tristate
rlabel metal2 s 41713 667333 42193 667389 6 mprj_gpio_analog[10]
port 378 nsew signal bidirectional
rlabel metal2 s 41713 665493 42193 665549 6 mprj_gpio_noesd[10]
port 379 nsew signal bidirectional
rlabel metal5 s 6598 657020 19088 669560 6 mprj_io[28]
port 380 nsew signal bidirectional
rlabel metal2 s 41713 664941 42193 664997 6 mprj_io_analog_en[17]
port 381 nsew signal input
rlabel metal2 s 41713 663653 42193 663709 6 mprj_io_analog_pol[17]
port 382 nsew signal input
rlabel metal2 s 41713 660617 42193 660673 6 mprj_io_analog_sel[17]
port 383 nsew signal input
rlabel metal2 s 41713 664297 42193 664353 6 mprj_io_dm[51]
port 384 nsew signal input
rlabel metal2 s 41713 666137 42193 666193 6 mprj_io_dm[52]
port 385 nsew signal input
rlabel metal2 s 41713 659973 42193 660029 6 mprj_io_dm[53]
port 386 nsew signal input
rlabel metal2 s 41713 659329 42193 659385 6 mprj_io_holdover[17]
port 387 nsew signal input
rlabel metal2 s 41713 656293 42193 656349 6 mprj_io_ib_mode_sel[17]
port 388 nsew signal input
rlabel metal2 s 41713 663101 42193 663157 6 mprj_io_inp_dis[17]
port 389 nsew signal input
rlabel metal2 s 41713 655649 42193 655705 6 mprj_io_oeb[17]
port 390 nsew signal input
rlabel metal2 s 41713 658777 42193 658833 6 mprj_io_out[17]
port 391 nsew signal input
rlabel metal2 s 41713 667977 42193 668033 6 mprj_io_slow_sel[17]
port 392 nsew signal input
rlabel metal2 s 41713 656937 42193 656993 6 mprj_io_vtrip_sel[17]
port 393 nsew signal input
rlabel metal2 s 41713 669817 42193 669873 6 mprj_io_in[17]
port 394 nsew signal tristate
rlabel metal2 s 41713 655097 42193 655153 6 mprj_io_in_3v3[17]
port 395 nsew signal tristate
rlabel metal2 s 41713 624133 42193 624189 6 mprj_gpio_analog[11]
port 396 nsew signal bidirectional
rlabel metal2 s 41713 622293 42193 622349 6 mprj_gpio_noesd[11]
port 397 nsew signal bidirectional
rlabel metal5 s 6598 613820 19088 626360 6 mprj_io[29]
port 398 nsew signal bidirectional
rlabel metal2 s 41713 621741 42193 621797 6 mprj_io_analog_en[18]
port 399 nsew signal input
rlabel metal2 s 41713 620453 42193 620509 6 mprj_io_analog_pol[18]
port 400 nsew signal input
rlabel metal2 s 41713 617417 42193 617473 6 mprj_io_analog_sel[18]
port 401 nsew signal input
rlabel metal2 s 41713 621097 42193 621153 6 mprj_io_dm[54]
port 402 nsew signal input
rlabel metal2 s 41713 622937 42193 622993 6 mprj_io_dm[55]
port 403 nsew signal input
rlabel metal2 s 41713 616773 42193 616829 6 mprj_io_dm[56]
port 404 nsew signal input
rlabel metal2 s 41713 616129 42193 616185 6 mprj_io_holdover[18]
port 405 nsew signal input
rlabel metal2 s 41713 613093 42193 613149 6 mprj_io_ib_mode_sel[18]
port 406 nsew signal input
rlabel metal2 s 41713 619901 42193 619957 6 mprj_io_inp_dis[18]
port 407 nsew signal input
rlabel metal2 s 41713 612449 42193 612505 6 mprj_io_oeb[18]
port 408 nsew signal input
rlabel metal2 s 41713 615577 42193 615633 6 mprj_io_out[18]
port 409 nsew signal input
rlabel metal2 s 41713 624777 42193 624833 6 mprj_io_slow_sel[18]
port 410 nsew signal input
rlabel metal2 s 41713 613737 42193 613793 6 mprj_io_vtrip_sel[18]
port 411 nsew signal input
rlabel metal2 s 41713 626617 42193 626673 6 mprj_io_in[18]
port 412 nsew signal tristate
rlabel metal2 s 41713 611897 42193 611953 6 mprj_io_in_3v3[18]
port 413 nsew signal tristate
rlabel metal2 s 41713 580933 42193 580989 6 mprj_gpio_analog[12]
port 414 nsew signal bidirectional
rlabel metal2 s 41713 579093 42193 579149 6 mprj_gpio_noesd[12]
port 415 nsew signal bidirectional
rlabel metal5 s 6598 570620 19088 583160 6 mprj_io[30]
port 416 nsew signal bidirectional
rlabel metal2 s 41713 578541 42193 578597 6 mprj_io_analog_en[19]
port 417 nsew signal input
rlabel metal2 s 41713 577253 42193 577309 6 mprj_io_analog_pol[19]
port 418 nsew signal input
rlabel metal2 s 41713 574217 42193 574273 6 mprj_io_analog_sel[19]
port 419 nsew signal input
rlabel metal2 s 41713 577897 42193 577953 6 mprj_io_dm[57]
port 420 nsew signal input
rlabel metal2 s 41713 579737 42193 579793 6 mprj_io_dm[58]
port 421 nsew signal input
rlabel metal2 s 41713 573573 42193 573629 6 mprj_io_dm[59]
port 422 nsew signal input
rlabel metal2 s 41713 572929 42193 572985 6 mprj_io_holdover[19]
port 423 nsew signal input
rlabel metal2 s 41713 569893 42193 569949 6 mprj_io_ib_mode_sel[19]
port 424 nsew signal input
rlabel metal2 s 41713 576701 42193 576757 6 mprj_io_inp_dis[19]
port 425 nsew signal input
rlabel metal2 s 41713 569249 42193 569305 6 mprj_io_oeb[19]
port 426 nsew signal input
rlabel metal2 s 41713 572377 42193 572433 6 mprj_io_out[19]
port 427 nsew signal input
rlabel metal2 s 41713 581577 42193 581633 6 mprj_io_slow_sel[19]
port 428 nsew signal input
rlabel metal2 s 41713 570537 42193 570593 6 mprj_io_vtrip_sel[19]
port 429 nsew signal input
rlabel metal2 s 41713 583417 42193 583473 6 mprj_io_in[19]
port 430 nsew signal tristate
rlabel metal2 s 41713 568697 42193 568753 6 mprj_io_in_3v3[19]
port 431 nsew signal tristate
rlabel metal2 s 41713 537733 42193 537789 6 mprj_gpio_analog[13]
port 432 nsew signal bidirectional
rlabel metal2 s 41713 535893 42193 535949 6 mprj_gpio_noesd[13]
port 433 nsew signal bidirectional
rlabel metal5 s 6598 527420 19088 539960 6 mprj_io[31]
port 434 nsew signal bidirectional
rlabel metal2 s 41713 535341 42193 535397 6 mprj_io_analog_en[20]
port 435 nsew signal input
rlabel metal2 s 41713 534053 42193 534109 6 mprj_io_analog_pol[20]
port 436 nsew signal input
rlabel metal2 s 41713 531017 42193 531073 6 mprj_io_analog_sel[20]
port 437 nsew signal input
rlabel metal2 s 41713 534697 42193 534753 6 mprj_io_dm[60]
port 438 nsew signal input
rlabel metal2 s 41713 536537 42193 536593 6 mprj_io_dm[61]
port 439 nsew signal input
rlabel metal2 s 41713 530373 42193 530429 6 mprj_io_dm[62]
port 440 nsew signal input
rlabel metal2 s 41713 529729 42193 529785 6 mprj_io_holdover[20]
port 441 nsew signal input
rlabel metal2 s 41713 526693 42193 526749 6 mprj_io_ib_mode_sel[20]
port 442 nsew signal input
rlabel metal2 s 41713 533501 42193 533557 6 mprj_io_inp_dis[20]
port 443 nsew signal input
rlabel metal2 s 41713 526049 42193 526105 6 mprj_io_oeb[20]
port 444 nsew signal input
rlabel metal2 s 41713 529177 42193 529233 6 mprj_io_out[20]
port 445 nsew signal input
rlabel metal2 s 41713 538377 42193 538433 6 mprj_io_slow_sel[20]
port 446 nsew signal input
rlabel metal2 s 41713 527337 42193 527393 6 mprj_io_vtrip_sel[20]
port 447 nsew signal input
rlabel metal2 s 41713 540217 42193 540273 6 mprj_io_in[20]
port 448 nsew signal tristate
rlabel metal2 s 41713 525497 42193 525553 6 mprj_io_in_3v3[20]
port 449 nsew signal tristate
rlabel metal2 s 41713 410133 42193 410189 6 mprj_gpio_analog[14]
port 450 nsew signal bidirectional
rlabel metal2 s 41713 408293 42193 408349 6 mprj_gpio_noesd[14]
port 451 nsew signal bidirectional
rlabel metal5 s 6598 399820 19088 412360 6 mprj_io[32]
port 452 nsew signal bidirectional
rlabel metal2 s 41713 407741 42193 407797 6 mprj_io_analog_en[21]
port 453 nsew signal input
rlabel metal2 s 41713 406453 42193 406509 6 mprj_io_analog_pol[21]
port 454 nsew signal input
rlabel metal2 s 41713 403417 42193 403473 6 mprj_io_analog_sel[21]
port 455 nsew signal input
rlabel metal2 s 41713 407097 42193 407153 6 mprj_io_dm[63]
port 456 nsew signal input
rlabel metal2 s 41713 408937 42193 408993 6 mprj_io_dm[64]
port 457 nsew signal input
rlabel metal2 s 41713 402773 42193 402829 6 mprj_io_dm[65]
port 458 nsew signal input
rlabel metal2 s 41713 402129 42193 402185 6 mprj_io_holdover[21]
port 459 nsew signal input
rlabel metal2 s 41713 399093 42193 399149 6 mprj_io_ib_mode_sel[21]
port 460 nsew signal input
rlabel metal2 s 41713 405901 42193 405957 6 mprj_io_inp_dis[21]
port 461 nsew signal input
rlabel metal2 s 41713 398449 42193 398505 6 mprj_io_oeb[21]
port 462 nsew signal input
rlabel metal2 s 41713 401577 42193 401633 6 mprj_io_out[21]
port 463 nsew signal input
rlabel metal2 s 41713 410777 42193 410833 6 mprj_io_slow_sel[21]
port 464 nsew signal input
rlabel metal2 s 41713 399737 42193 399793 6 mprj_io_vtrip_sel[21]
port 465 nsew signal input
rlabel metal2 s 41713 412617 42193 412673 6 mprj_io_in[21]
port 466 nsew signal tristate
rlabel metal2 s 41713 397897 42193 397953 6 mprj_io_in_3v3[21]
port 467 nsew signal tristate
rlabel metal2 s 41713 366933 42193 366989 6 mprj_gpio_analog[15]
port 468 nsew signal bidirectional
rlabel metal2 s 41713 365093 42193 365149 6 mprj_gpio_noesd[15]
port 469 nsew signal bidirectional
rlabel metal5 s 6598 356620 19088 369160 6 mprj_io[33]
port 470 nsew signal bidirectional
rlabel metal2 s 41713 364541 42193 364597 6 mprj_io_analog_en[22]
port 471 nsew signal input
rlabel metal2 s 41713 363253 42193 363309 6 mprj_io_analog_pol[22]
port 472 nsew signal input
rlabel metal2 s 41713 360217 42193 360273 6 mprj_io_analog_sel[22]
port 473 nsew signal input
rlabel metal2 s 41713 363897 42193 363953 6 mprj_io_dm[66]
port 474 nsew signal input
rlabel metal2 s 41713 365737 42193 365793 6 mprj_io_dm[67]
port 475 nsew signal input
rlabel metal2 s 41713 359573 42193 359629 6 mprj_io_dm[68]
port 476 nsew signal input
rlabel metal2 s 41713 358929 42193 358985 6 mprj_io_holdover[22]
port 477 nsew signal input
rlabel metal2 s 41713 355893 42193 355949 6 mprj_io_ib_mode_sel[22]
port 478 nsew signal input
rlabel metal2 s 41713 362701 42193 362757 6 mprj_io_inp_dis[22]
port 479 nsew signal input
rlabel metal2 s 41713 355249 42193 355305 6 mprj_io_oeb[22]
port 480 nsew signal input
rlabel metal2 s 41713 358377 42193 358433 6 mprj_io_out[22]
port 481 nsew signal input
rlabel metal2 s 41713 367577 42193 367633 6 mprj_io_slow_sel[22]
port 482 nsew signal input
rlabel metal2 s 41713 356537 42193 356593 6 mprj_io_vtrip_sel[22]
port 483 nsew signal input
rlabel metal2 s 41713 369417 42193 369473 6 mprj_io_in[22]
port 484 nsew signal tristate
rlabel metal2 s 41713 354697 42193 354753 6 mprj_io_in_3v3[22]
port 485 nsew signal tristate
rlabel metal2 s 41713 323733 42193 323789 6 mprj_gpio_analog[16]
port 486 nsew signal bidirectional
rlabel metal2 s 41713 321893 42193 321949 6 mprj_gpio_noesd[16]
port 487 nsew signal bidirectional
rlabel metal5 s 6598 313420 19088 325960 6 mprj_io[34]
port 488 nsew signal bidirectional
rlabel metal2 s 41713 321341 42193 321397 6 mprj_io_analog_en[23]
port 489 nsew signal input
rlabel metal2 s 41713 320053 42193 320109 6 mprj_io_analog_pol[23]
port 490 nsew signal input
rlabel metal2 s 41713 317017 42193 317073 6 mprj_io_analog_sel[23]
port 491 nsew signal input
rlabel metal2 s 41713 320697 42193 320753 6 mprj_io_dm[69]
port 492 nsew signal input
rlabel metal2 s 41713 322537 42193 322593 6 mprj_io_dm[70]
port 493 nsew signal input
rlabel metal2 s 41713 316373 42193 316429 6 mprj_io_dm[71]
port 494 nsew signal input
rlabel metal2 s 41713 315729 42193 315785 6 mprj_io_holdover[23]
port 495 nsew signal input
rlabel metal2 s 41713 312693 42193 312749 6 mprj_io_ib_mode_sel[23]
port 496 nsew signal input
rlabel metal2 s 41713 319501 42193 319557 6 mprj_io_inp_dis[23]
port 497 nsew signal input
rlabel metal2 s 41713 312049 42193 312105 6 mprj_io_oeb[23]
port 498 nsew signal input
rlabel metal2 s 41713 315177 42193 315233 6 mprj_io_out[23]
port 499 nsew signal input
rlabel metal2 s 41713 324377 42193 324433 6 mprj_io_slow_sel[23]
port 500 nsew signal input
rlabel metal2 s 41713 313337 42193 313393 6 mprj_io_vtrip_sel[23]
port 501 nsew signal input
rlabel metal2 s 41713 326217 42193 326273 6 mprj_io_in[23]
port 502 nsew signal tristate
rlabel metal2 s 41713 311497 42193 311553 6 mprj_io_in_3v3[23]
port 503 nsew signal tristate
rlabel metal2 s 145091 39706 145143 40000 6 porb_h
port 504 nsew signal input
rlabel metal5 s 136713 7143 144149 18309 6 resetb
port 505 nsew signal input
rlabel metal3 s 141667 38031 141813 39999 6 resetb_core_h
port 506 nsew signal tristate
rlabel metal4 s 132600 36323 132792 37013 6 vdda
port 507 nsew signal bidirectional
rlabel metal4 s 132600 28653 147600 28719 6 vssa
port 508 nsew signal bidirectional
rlabel metal4 s 132600 30762 132868 31674 6 vssd
port 509 nsew signal bidirectional
rlabel metal3 s 631944 997600 636944 1014070 6 mprj_analog[0]
port 510 nsew signal bidirectional
rlabel metal5 s 628410 1018624 640578 1030788 6 mprj_io[15]
port 511 nsew signal bidirectional
rlabel metal3 s 530144 997600 535144 1014070 6 mprj_analog[1]
port 512 nsew signal bidirectional
rlabel metal5 s 526610 1018624 538778 1030788 6 mprj_io[16]
port 513 nsew signal bidirectional
rlabel metal3 s 478744 997600 483744 1014070 6 mprj_analog[2]
port 514 nsew signal bidirectional
rlabel metal5 s 475210 1018624 487378 1030788 6 mprj_io[17]
port 515 nsew signal bidirectional
rlabel metal5 s 697980 909666 711432 920546 6 vccd1_pad
port 522 nsew signal bidirectional
rlabel metal5 s 698624 819822 710788 831990 6 vdda1_pad
port 523 nsew signal bidirectional
rlabel metal5 s 698624 505222 710788 517390 6 vdda1_pad2
port 524 nsew signal bidirectional
rlabel metal5 s 577010 1018624 589178 1030788 6 vssa1_pad
port 525 nsew signal bidirectional
rlabel metal5 s 698624 417022 710788 429190 6 vssa1_pad2
port 526 nsew signal bidirectional
rlabel metal4 s 679377 459800 680307 460054 6 vccd1
port 527 nsew signal bidirectional
rlabel metal4 s 680587 459800 681277 459992 6 vdda1
port 528 nsew signal bidirectional
rlabel metal4 s 688881 459800 688947 474800 6 vssa1
port 529 nsew signal bidirectional
rlabel metal3 s 678000 469900 685920 474700 6 vssd1
port 530 nsew signal bidirectional
rlabel metal5 s 697980 461866 711432 472746 6 vssd1_pad
port 531 nsew signal bidirectional
rlabel metal3 s 184944 997600 189944 1014070 6 mprj_analog[7]
port 532 nsew signal bidirectional
rlabel metal5 s 181410 1018624 193578 1030788 6 mprj_io[21]
port 533 nsew signal bidirectional
rlabel metal3 s 133544 997600 138544 1014070 6 mprj_analog[8]
port 534 nsew signal bidirectional
rlabel metal5 s 130010 1018624 142178 1030788 6 mprj_io[22]
port 535 nsew signal bidirectional
rlabel metal3 s 82144 997600 87144 1014070 6 mprj_analog[9]
port 536 nsew signal bidirectional
rlabel metal5 s 78610 1018624 90778 1030788 6 mprj_io[23]
port 537 nsew signal bidirectional
rlabel metal3 s 23530 960144 40000 965144 6 mprj_analog[10]
port 538 nsew signal bidirectional
rlabel metal5 s 6811 956610 18975 968778 6 mprj_io[24]
port 539 nsew signal bidirectional
rlabel metal3 s 240478 997600 254800 1000736 6 mprj_analog[6]
port 544 nsew signal bidirectional
rlabel metal2 s 240478 997600 245258 1002732 6 mprj_clamp_high[2]
port 545 nsew signal input
rlabel metal2 s 230499 997600 235279 998010 6 mprj_clamp_low[2]
port 546 nsew signal input
rlabel metal5 s 231810 1018624 243978 1030788 6 mprj_io[20]
port 547 nsew signal bidirectional
rlabel metal5 s 6167 914054 19619 924934 6 vccd2_pad
port 548 nsew signal bidirectional
rlabel metal5 s 6811 484410 18975 496578 6 vdda2_pad
port 549 nsew signal bidirectional
rlabel metal5 s 6811 829010 18975 841178 6 vssa2_pad
port 550 nsew signal bidirectional
rlabel metal4 s 38503 455546 39593 455800 6 vccd
port 551 nsew signal bidirectional
rlabel metal4 s 37293 455546 38223 455800 6 vccd2
port 552 nsew signal bidirectional
rlabel metal4 s 36323 455607 37013 455799 6 vdda2
port 553 nsew signal bidirectional
rlabel metal4 s 32933 455546 33623 455800 6 vddio
port 554 nsew signal bidirectional
rlabel metal4 s 28653 440800 28719 455800 6 vssa2
port 555 nsew signal bidirectional
rlabel metal3 s 31680 440900 39600 445700 6 vssd2
port 556 nsew signal bidirectional
rlabel metal5 s 6167 442854 19619 453734 6 vssd2_pad
port 557 nsew signal bidirectional
rlabel metal4 s 7 455645 4843 456093 6 vssio
port 558 nsew signal bidirectional
rlabel metal5 s 386210 1018624 398378 1030788 6 mprj_io[18]
port 521 nsew signal bidirectional
rlabel metal5 s 284410 1018624 296578 1030788 6 mprj_io[19]
port 543 nsew signal bidirectional
rlabel metal3 s 677600 956656 694070 961656 6 mprj_analog[3]
port 516 nsew signal bidirectional
rlabel metal5 s 698624 953022 710788 965190 6 mprj_io[14]
port 517 nsew signal bidirectional
rlabel metal3 s 293078 997600 307400 1000736 6 mprj_analog[5]
port 540 nsew signal bidirectional
rlabel metal2 s 293078 997600 297858 1002732 6 mprj_clamp_high[1]
port 541 nsew signal input
rlabel metal2 s 283099 997600 287879 998010 6 mprj_clamp_low[1]
port 542 nsew signal input
rlabel metal3 s 394878 997600 409200 1000736 6 mprj_analog[4]
port 518 nsew signal bidirectional
rlabel metal2 s 394878 997600 399658 1002732 6 mprj_clamp_high[0]
port 519 nsew signal input
rlabel metal2 s 384899 997600 389679 998010 6 mprj_clamp_low[0]
port 520 nsew signal input
rlabel metal2 306967 41713 307023 42193 0 flash_csb_core
port 559 nsew
rlabel metal2 357443 41713 357499 42193 0 flash_clk_ieb_core
port 560 nsew
rlabel metal2 364895 41713 364951 42193 0 flash_clk_oeb_core
port 561 nsew
rlabel metal2 361767 41713 361823 42193 0 flash_clk_core
port 562 nsew
rlabel metal2 310095 41713 310151 42193 0 flash_csb_oeb_core
port 563 nsew
rlabel metal2 302643 41713 302699 42193 0 flash_csb_ieb_core
port 564 nsew
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
