magic
tech sky130A
magscale 1 2
timestamp 1606493992
<< checkpaint >>
rect -1260 -1260 718860 1038860
<< pdiff >>
rect 77289 1034726 77323 1034752
rect 78523 1034726 78557 1034752
rect 128689 1034726 128723 1034752
rect 129923 1034726 129957 1034752
rect 180089 1034726 180123 1034752
rect 181323 1034726 181357 1034752
rect 231489 1034726 231523 1034752
rect 232723 1034726 232757 1034752
rect 283089 1034726 283123 1034752
rect 284323 1034726 284357 1034752
rect 384889 1034726 384923 1034752
rect 386123 1034726 386157 1034752
rect 473889 1034726 473923 1034752
rect 475123 1034726 475157 1034752
rect 525289 1034726 525323 1034752
rect 526523 1034726 526557 1034752
rect 627089 1034726 627123 1034752
rect 628323 1034726 628357 1034752
rect 82571 1032409 89682 1032431
rect 91517 1031619 91531 1032463
rect 133971 1032409 141082 1032431
rect 142917 1031619 142931 1032463
rect 185371 1032409 192482 1032431
rect 194317 1031619 194331 1032463
rect 236771 1032409 243882 1032431
rect 245717 1031619 245731 1032463
rect 288371 1032409 295482 1032431
rect 297317 1031619 297331 1032463
rect 390171 1032409 397282 1032431
rect 399117 1031619 399131 1032463
rect 479171 1032409 486282 1032431
rect 488117 1031619 488131 1032463
rect 530571 1032409 537682 1032431
rect 539517 1031619 539531 1032463
rect 632371 1032409 639482 1032431
rect 641317 1031619 641331 1032463
rect 91507 1031605 91531 1031619
rect 142907 1031605 142931 1031619
rect 194307 1031605 194331 1031619
rect 245707 1031605 245731 1031619
rect 297307 1031605 297331 1031619
rect 399107 1031605 399131 1031619
rect 488107 1031605 488131 1031619
rect 539507 1031605 539531 1031619
rect 641307 1031605 641331 1031619
rect 77501 1031579 89682 1031595
rect 89725 1031579 91531 1031605
rect 128901 1031579 141082 1031595
rect 141125 1031579 142931 1031605
rect 180301 1031579 192482 1031595
rect 192525 1031579 194331 1031605
rect 231701 1031579 243882 1031595
rect 243925 1031579 245731 1031605
rect 283301 1031579 295482 1031595
rect 295525 1031579 297331 1031605
rect 385101 1031579 397282 1031595
rect 397325 1031579 399131 1031605
rect 474101 1031579 486282 1031595
rect 486325 1031579 488131 1031605
rect 525501 1031579 537682 1031595
rect 537725 1031579 539531 1031605
rect 627301 1031579 639482 1031595
rect 639525 1031579 641331 1031605
rect 78136 1029211 78298 1030211
rect 90422 1029211 90463 1030211
rect 90984 1029211 91194 1030211
rect 129536 1029211 129698 1030211
rect 141822 1029211 141863 1030211
rect 142384 1029211 142594 1030211
rect 180936 1029211 181098 1030211
rect 193222 1029211 193263 1030211
rect 193784 1029211 193994 1030211
rect 232336 1029211 232498 1030211
rect 244622 1029211 244663 1030211
rect 245184 1029211 245394 1030211
rect 283936 1029211 284098 1030211
rect 296222 1029211 296263 1030211
rect 296784 1029211 296994 1030211
rect 385736 1029211 385898 1030211
rect 398022 1029211 398063 1030211
rect 398584 1029211 398794 1030211
rect 474736 1029211 474898 1030211
rect 487022 1029211 487063 1030211
rect 487584 1029211 487794 1030211
rect 526136 1029211 526298 1030211
rect 538422 1029211 538463 1030211
rect 538984 1029211 539194 1030211
rect 627936 1029211 628098 1030211
rect 640222 1029211 640263 1030211
rect 640784 1029211 640994 1030211
rect 78159 1027610 78299 1028610
rect 90422 1027610 90463 1028610
rect 90984 1027610 91194 1028610
rect 129559 1027610 129699 1028610
rect 141822 1027610 141863 1028610
rect 142384 1027610 142594 1028610
rect 180959 1027610 181099 1028610
rect 193222 1027610 193263 1028610
rect 193784 1027610 193994 1028610
rect 232359 1027610 232499 1028610
rect 244622 1027610 244663 1028610
rect 245184 1027610 245394 1028610
rect 283959 1027610 284099 1028610
rect 296222 1027610 296263 1028610
rect 296784 1027610 296994 1028610
rect 385759 1027610 385899 1028610
rect 398022 1027610 398063 1028610
rect 398584 1027610 398794 1028610
rect 474759 1027610 474899 1028610
rect 487022 1027610 487063 1028610
rect 487584 1027610 487794 1028610
rect 526159 1027610 526299 1028610
rect 538422 1027610 538463 1028610
rect 538984 1027610 539194 1028610
rect 627959 1027610 628099 1028610
rect 640222 1027610 640263 1028610
rect 640784 1027610 640994 1028610
rect 77035 1018110 77183 1022856
rect 77700 1020922 77726 1021922
rect 77771 1020922 77873 1021922
rect 90939 1020922 91094 1021922
rect 91264 1020922 91419 1021922
rect 77700 1019322 77726 1020322
rect 77771 1019322 77873 1020322
rect 90939 1019322 91094 1020322
rect 91264 1019322 91419 1020322
rect 128435 1018110 128583 1022856
rect 129100 1020922 129126 1021922
rect 129171 1020922 129273 1021922
rect 142339 1020922 142494 1021922
rect 142664 1020922 142819 1021922
rect 129100 1019322 129126 1020322
rect 129171 1019322 129273 1020322
rect 142339 1019322 142494 1020322
rect 142664 1019322 142819 1020322
rect 179835 1018110 179983 1022856
rect 180500 1020922 180526 1021922
rect 180571 1020922 180673 1021922
rect 193739 1020922 193894 1021922
rect 194064 1020922 194219 1021922
rect 180500 1019322 180526 1020322
rect 180571 1019322 180673 1020322
rect 193739 1019322 193894 1020322
rect 194064 1019322 194219 1020322
rect 231235 1018110 231383 1022856
rect 231900 1020922 231926 1021922
rect 231971 1020922 232073 1021922
rect 245139 1020922 245294 1021922
rect 245464 1020922 245619 1021922
rect 231900 1019322 231926 1020322
rect 231971 1019322 232073 1020322
rect 245139 1019322 245294 1020322
rect 245464 1019322 245619 1020322
rect 282835 1018110 282983 1022856
rect 283500 1020922 283526 1021922
rect 283571 1020922 283673 1021922
rect 296739 1020922 296894 1021922
rect 297064 1020922 297219 1021922
rect 283500 1019322 283526 1020322
rect 283571 1019322 283673 1020322
rect 296739 1019322 296894 1020322
rect 297064 1019322 297219 1020322
rect 384635 1018110 384783 1022856
rect 385300 1020922 385326 1021922
rect 385371 1020922 385473 1021922
rect 398539 1020922 398694 1021922
rect 398864 1020922 399019 1021922
rect 385300 1019322 385326 1020322
rect 385371 1019322 385473 1020322
rect 398539 1019322 398694 1020322
rect 398864 1019322 399019 1020322
rect 473635 1018110 473783 1022856
rect 474300 1020922 474326 1021922
rect 474371 1020922 474473 1021922
rect 487539 1020922 487694 1021922
rect 487864 1020922 488019 1021922
rect 474300 1019322 474326 1020322
rect 474371 1019322 474473 1020322
rect 487539 1019322 487694 1020322
rect 487864 1019322 488019 1020322
rect 525035 1018110 525183 1022856
rect 525700 1020922 525726 1021922
rect 525771 1020922 525873 1021922
rect 538939 1020922 539094 1021922
rect 539264 1020922 539419 1021922
rect 525700 1019322 525726 1020322
rect 525771 1019322 525873 1020322
rect 538939 1019322 539094 1020322
rect 539264 1019322 539419 1020322
rect 626835 1018110 626983 1022856
rect 627500 1020922 627526 1021922
rect 627571 1020922 627673 1021922
rect 640739 1020922 640894 1021922
rect 641064 1020922 641219 1021922
rect 627500 1019322 627526 1020322
rect 627571 1019322 627673 1020322
rect 640739 1019322 640894 1020322
rect 641064 1019322 641219 1020322
rect 77209 1018053 84133 1018084
rect 128609 1018053 135533 1018084
rect 180009 1018053 186933 1018084
rect 231409 1018053 238333 1018084
rect 283009 1018053 289933 1018084
rect 384809 1018053 391733 1018084
rect 473809 1018053 480733 1018084
rect 525209 1018053 532133 1018084
rect 627009 1018053 633933 1018084
rect 84137 1016817 85342 1016821
rect 135537 1016817 136742 1016821
rect 186937 1016817 188142 1016821
rect 238337 1016817 239542 1016821
rect 289937 1016817 291142 1016821
rect 391737 1016817 392942 1016821
rect 480737 1016817 481942 1016821
rect 532137 1016817 533342 1016821
rect 633937 1016817 635142 1016821
rect 77918 1016779 77974 1016791
rect 129318 1016779 129374 1016791
rect 180718 1016779 180774 1016791
rect 232118 1016779 232174 1016791
rect 283718 1016779 283774 1016791
rect 385518 1016779 385574 1016791
rect 474518 1016779 474574 1016791
rect 525918 1016779 525974 1016791
rect 627718 1016779 627774 1016791
rect 84763 1007758 85211 1007764
rect 87809 1007758 88283 1007764
rect 136163 1007758 136611 1007764
rect 139209 1007758 139683 1007764
rect 187563 1007758 188011 1007764
rect 190609 1007758 191083 1007764
rect 238963 1007758 239411 1007764
rect 242009 1007758 242483 1007764
rect 290563 1007758 291011 1007764
rect 293609 1007758 294083 1007764
rect 392363 1007758 392811 1007764
rect 395409 1007758 395883 1007764
rect 481363 1007758 481811 1007764
rect 484409 1007758 484883 1007764
rect 532763 1007758 533211 1007764
rect 535809 1007758 536283 1007764
rect 634563 1007758 635011 1007764
rect 637609 1007758 638083 1007764
rect 82935 1007645 88488 1007648
rect 134335 1007645 139888 1007648
rect 185735 1007645 191288 1007648
rect 237135 1007645 242688 1007648
rect 288735 1007645 294288 1007648
rect 390535 1007645 396088 1007648
rect 479535 1007645 485088 1007648
rect 530935 1007645 536488 1007648
rect 632735 1007645 638288 1007648
rect 83728 1007573 89477 1007585
rect 135128 1007573 140877 1007585
rect 186528 1007573 192277 1007585
rect 237928 1007573 243677 1007585
rect 289528 1007573 295277 1007585
rect 391328 1007573 397077 1007585
rect 480328 1007573 486077 1007585
rect 531728 1007573 537477 1007585
rect 633528 1007573 639277 1007585
rect 83728 1006882 83754 1007573
rect 135128 1006882 135154 1007573
rect 186528 1006882 186554 1007573
rect 237928 1006882 237954 1007573
rect 289528 1006882 289554 1007573
rect 391328 1006882 391354 1007573
rect 480328 1006882 480354 1007573
rect 531728 1006882 531754 1007573
rect 633528 1006882 633554 1007573
rect 83744 1006879 83754 1006882
rect 135144 1006879 135154 1006882
rect 186544 1006879 186554 1006882
rect 237944 1006879 237954 1006882
rect 289544 1006879 289554 1006882
rect 391344 1006879 391354 1006882
rect 480344 1006879 480354 1006882
rect 531744 1006879 531754 1006882
rect 633544 1006879 633554 1006882
rect 79916 1005803 79932 1006119
rect 81120 1005803 81138 1006119
rect 131316 1005803 131332 1006119
rect 132520 1005803 132538 1006119
rect 182716 1005803 182732 1006119
rect 183920 1005803 183938 1006119
rect 234116 1005803 234132 1006119
rect 235320 1005803 235338 1006119
rect 285716 1005803 285732 1006119
rect 286920 1005803 286938 1006119
rect 387516 1005803 387532 1006119
rect 388720 1005803 388738 1006119
rect 476516 1005803 476532 1006119
rect 477720 1005803 477738 1006119
rect 527916 1005803 527932 1006119
rect 529120 1005803 529138 1006119
rect 629716 1005803 629732 1006119
rect 630920 1005803 630938 1006119
rect 79916 1005777 79920 1005803
rect 131316 1005777 131320 1005803
rect 182716 1005777 182720 1005803
rect 234116 1005777 234120 1005803
rect 285716 1005777 285720 1005803
rect 387516 1005777 387520 1005803
rect 476516 1005777 476520 1005803
rect 527916 1005777 527920 1005803
rect 629716 1005777 629720 1005803
rect 79882 1005539 79920 1005777
rect 81140 1005539 81172 1005777
rect 131282 1005539 131320 1005777
rect 132540 1005539 132572 1005777
rect 182682 1005539 182720 1005777
rect 183940 1005539 183972 1005777
rect 234082 1005539 234120 1005777
rect 235340 1005539 235372 1005777
rect 285682 1005539 285720 1005777
rect 286940 1005539 286972 1005777
rect 387482 1005539 387520 1005777
rect 388740 1005539 388772 1005777
rect 476482 1005539 476520 1005777
rect 477740 1005539 477772 1005777
rect 527882 1005539 527920 1005777
rect 529140 1005539 529172 1005777
rect 629682 1005539 629720 1005777
rect 630940 1005539 630972 1005777
rect 80705 1001502 81195 1001529
rect 132105 1001502 132595 1001529
rect 183505 1001502 183995 1001529
rect 234905 1001502 235395 1001529
rect 286505 1001502 286995 1001529
rect 388305 1001502 388795 1001529
rect 477305 1001502 477795 1001529
rect 528705 1001502 529195 1001529
rect 630505 1001502 630995 1001529
rect 85213 998646 85239 998654
rect 88423 998646 88448 998654
rect 136613 998646 136639 998654
rect 139823 998646 139848 998654
rect 188013 998646 188039 998654
rect 191223 998646 191248 998654
rect 239413 998646 239439 998654
rect 242623 998646 242648 998654
rect 291013 998646 291039 998654
rect 294223 998646 294248 998654
rect 392813 998646 392839 998654
rect 396023 998646 396048 998654
rect 481813 998646 481839 998654
rect 485023 998646 485048 998654
rect 533213 998646 533239 998654
rect 536423 998646 536448 998654
rect 635013 998646 635039 998654
rect 638223 998646 638248 998654
rect 5137 969517 6021 969531
rect 5981 969507 6021 969517
rect 5995 967725 6021 969507
rect 15678 969264 16678 969419
rect 17278 969264 18278 969419
rect 7389 968984 8389 969194
rect 8990 968984 9990 969194
rect 15678 968939 16678 969094
rect 17278 968939 18278 969094
rect 7389 968422 8389 968463
rect 8990 968422 9990 968463
rect 5169 960571 5191 967682
rect 2848 956523 2874 956557
rect 6005 955501 6021 967682
rect 29836 965809 29842 966283
rect 20779 962137 20783 963342
rect 29836 962763 29842 963211
rect 7389 956136 8389 956298
rect 8990 956159 9990 956299
rect 15678 955771 16678 955873
rect 17278 955771 18278 955873
rect 15678 955700 16678 955726
rect 17278 955700 18278 955726
rect 2848 955289 2874 955323
rect 19516 955209 19547 962133
rect 29952 960935 29955 966488
rect 30015 961754 30027 967477
rect 698110 966617 702856 966765
rect 38946 966423 38954 966448
rect 696779 965826 696791 965882
rect 685539 963884 685777 963918
rect 685539 963880 686119 963884
rect 685803 963868 686119 963880
rect 38946 963213 38954 963239
rect 681502 962605 681529 963095
rect 685803 962662 686119 962680
rect 685539 962628 685777 962660
rect 30015 961744 30721 961754
rect 30015 961728 30718 961744
rect 686882 960056 687585 960072
rect 686879 960046 687585 960056
rect 31823 959140 32061 959172
rect 31481 959120 31797 959138
rect 36071 958705 36098 959195
rect 678646 958561 678654 958587
rect 31481 957920 31797 957932
rect 31481 957916 32061 957920
rect 31823 957882 32061 957916
rect 20809 955918 20821 955974
rect 678646 955352 678654 955377
rect 14744 955035 19490 955183
rect 687573 954323 687585 960046
rect 687645 955312 687648 960865
rect 698053 959667 698084 966591
rect 714726 966477 714752 966511
rect 699322 966074 700322 966100
rect 700922 966074 701922 966100
rect 699322 965927 700322 966029
rect 700922 965927 701922 966029
rect 707610 965501 708610 965641
rect 709211 965502 710211 965664
rect 687758 958589 687764 959037
rect 696817 958458 696821 959663
rect 687758 955517 687764 955991
rect 711579 954118 711595 966299
rect 714726 965243 714752 965277
rect 712409 954118 712431 961229
rect 707610 953337 708610 953378
rect 709211 953337 710211 953378
rect 699322 952706 700322 952861
rect 700922 952706 701922 952861
rect 707610 952606 708610 952816
rect 709211 952606 710211 952816
rect 699322 952381 700322 952536
rect 700922 952381 701922 952536
rect 711579 952293 711605 954075
rect 711579 952283 711619 952293
rect 711579 952269 712463 952283
rect 35930 919315 39318 919329
rect 678282 919187 681670 919245
rect 35930 915355 39318 915413
rect 678282 915271 681670 915285
rect 698110 877417 702856 877565
rect 696779 876626 696791 876682
rect 685539 874684 685777 874718
rect 685539 874680 686119 874684
rect 685803 874668 686119 874680
rect 681502 873405 681529 873895
rect 685803 873462 686119 873480
rect 685539 873428 685777 873460
rect 686882 870856 687585 870872
rect 686879 870846 687585 870856
rect 678646 869361 678654 869387
rect 678646 866152 678654 866177
rect 687573 865123 687585 870846
rect 687645 866112 687648 871665
rect 698053 870467 698084 877391
rect 714726 877277 714752 877311
rect 699322 876874 700322 876900
rect 700922 876874 701922 876900
rect 699322 876727 700322 876829
rect 700922 876727 701922 876829
rect 707610 876301 708610 876441
rect 709211 876302 710211 876464
rect 687758 869389 687764 869837
rect 696817 869258 696821 870463
rect 687758 866317 687764 866791
rect 711579 864918 711595 877099
rect 714726 876043 714752 876077
rect 712409 864918 712431 872029
rect 707610 864137 708610 864178
rect 709211 864137 710211 864178
rect 699322 863506 700322 863661
rect 700922 863506 701922 863661
rect 707610 863406 708610 863616
rect 709211 863406 710211 863616
rect 699322 863181 700322 863336
rect 700922 863181 701922 863336
rect 711579 863093 711605 864875
rect 711579 863083 711619 863093
rect 711579 863069 712463 863083
rect 5137 799717 6021 799731
rect 5981 799707 6021 799717
rect 5995 797925 6021 799707
rect 15678 799464 16678 799619
rect 17278 799464 18278 799619
rect 7389 799184 8389 799394
rect 8990 799184 9990 799394
rect 15678 799139 16678 799294
rect 17278 799139 18278 799294
rect 7389 798622 8389 798663
rect 8990 798622 9990 798663
rect 5169 790771 5191 797882
rect 2848 786723 2874 786757
rect 6005 785701 6021 797882
rect 29836 796009 29842 796483
rect 20779 792337 20783 793542
rect 29836 792963 29842 793411
rect 7389 786336 8389 786498
rect 8990 786359 9990 786499
rect 15678 785971 16678 786073
rect 17278 785971 18278 786073
rect 15678 785900 16678 785926
rect 17278 785900 18278 785926
rect 2848 785489 2874 785523
rect 19516 785409 19547 792333
rect 29952 791135 29955 796688
rect 30015 791954 30027 797677
rect 38946 796623 38954 796648
rect 38946 793413 38954 793439
rect 30015 791944 30721 791954
rect 30015 791928 30718 791944
rect 31823 789340 32061 789372
rect 31481 789320 31797 789338
rect 36071 788905 36098 789395
rect 698110 788217 702856 788365
rect 31481 788120 31797 788132
rect 31481 788116 32061 788120
rect 31823 788082 32061 788116
rect 696779 787426 696791 787482
rect 20809 786118 20821 786174
rect 685539 785484 685777 785518
rect 685539 785480 686119 785484
rect 685803 785468 686119 785480
rect 14744 785235 19490 785383
rect 681502 784205 681529 784695
rect 685803 784262 686119 784280
rect 685539 784228 685777 784260
rect 686882 781656 687585 781672
rect 686879 781646 687585 781656
rect 678646 780161 678654 780187
rect 678646 776952 678654 776977
rect 687573 775923 687585 781646
rect 687645 776912 687648 782465
rect 698053 781267 698084 788191
rect 714726 788077 714752 788111
rect 699322 787674 700322 787700
rect 700922 787674 701922 787700
rect 699322 787527 700322 787629
rect 700922 787527 701922 787629
rect 707610 787101 708610 787241
rect 709211 787102 710211 787264
rect 687758 780189 687764 780637
rect 696817 780058 696821 781263
rect 687758 777117 687764 777591
rect 711579 775718 711595 787899
rect 714726 786843 714752 786877
rect 712409 775718 712431 782829
rect 707610 774937 708610 774978
rect 709211 774937 710211 774978
rect 699322 774306 700322 774461
rect 700922 774306 701922 774461
rect 707610 774206 708610 774416
rect 709211 774206 710211 774416
rect 699322 773981 700322 774136
rect 700922 773981 701922 774136
rect 711579 773893 711605 775675
rect 711579 773883 711619 773893
rect 711579 773869 712463 773883
rect 5137 756517 6021 756531
rect 5981 756507 6021 756517
rect 5995 754725 6021 756507
rect 15678 756264 16678 756419
rect 17278 756264 18278 756419
rect 7389 755984 8389 756194
rect 8990 755984 9990 756194
rect 15678 755939 16678 756094
rect 17278 755939 18278 756094
rect 7389 755422 8389 755463
rect 8990 755422 9990 755463
rect 5169 747571 5191 754682
rect 2848 743523 2874 743557
rect 6005 742501 6021 754682
rect 29836 752809 29842 753283
rect 20779 749137 20783 750342
rect 29836 749763 29842 750211
rect 7389 743136 8389 743298
rect 8990 743159 9990 743299
rect 15678 742771 16678 742873
rect 17278 742771 18278 742873
rect 15678 742700 16678 742726
rect 17278 742700 18278 742726
rect 2848 742289 2874 742323
rect 19516 742209 19547 749133
rect 29952 747935 29955 753488
rect 30015 748754 30027 754477
rect 38946 753423 38954 753448
rect 38946 750213 38954 750239
rect 30015 748744 30721 748754
rect 30015 748728 30718 748744
rect 31823 746140 32061 746172
rect 31481 746120 31797 746138
rect 36071 745705 36098 746195
rect 31481 744920 31797 744932
rect 31481 744916 32061 744920
rect 31823 744882 32061 744916
rect 698110 743217 702856 743365
rect 20809 742918 20821 742974
rect 696779 742426 696791 742482
rect 14744 742035 19490 742183
rect 685539 740484 685777 740518
rect 685539 740480 686119 740484
rect 685803 740468 686119 740480
rect 681502 739205 681529 739695
rect 685803 739262 686119 739280
rect 685539 739228 685777 739260
rect 686882 736656 687585 736672
rect 686879 736646 687585 736656
rect 678646 735161 678654 735187
rect 678646 731952 678654 731977
rect 687573 730923 687585 736646
rect 687645 731912 687648 737465
rect 698053 736267 698084 743191
rect 714726 743077 714752 743111
rect 699322 742674 700322 742700
rect 700922 742674 701922 742700
rect 699322 742527 700322 742629
rect 700922 742527 701922 742629
rect 707610 742101 708610 742241
rect 709211 742102 710211 742264
rect 687758 735189 687764 735637
rect 696817 735058 696821 736263
rect 687758 732117 687764 732591
rect 711579 730718 711595 742899
rect 714726 741843 714752 741877
rect 712409 730718 712431 737829
rect 707610 729937 708610 729978
rect 709211 729937 710211 729978
rect 699322 729306 700322 729461
rect 700922 729306 701922 729461
rect 707610 729206 708610 729416
rect 709211 729206 710211 729416
rect 699322 728981 700322 729136
rect 700922 728981 701922 729136
rect 711579 728893 711605 730675
rect 711579 728883 711619 728893
rect 711579 728869 712463 728883
rect 5137 713317 6021 713331
rect 5981 713307 6021 713317
rect 5995 711525 6021 713307
rect 15678 713064 16678 713219
rect 17278 713064 18278 713219
rect 7389 712784 8389 712994
rect 8990 712784 9990 712994
rect 15678 712739 16678 712894
rect 17278 712739 18278 712894
rect 7389 712222 8389 712263
rect 8990 712222 9990 712263
rect 5169 704371 5191 711482
rect 2848 700323 2874 700357
rect 6005 699301 6021 711482
rect 29836 709609 29842 710083
rect 20779 705937 20783 707142
rect 29836 706563 29842 707011
rect 7389 699936 8389 700098
rect 8990 699959 9990 700099
rect 15678 699571 16678 699673
rect 17278 699571 18278 699673
rect 15678 699500 16678 699526
rect 17278 699500 18278 699526
rect 2848 699089 2874 699123
rect 19516 699009 19547 705933
rect 29952 704735 29955 710288
rect 30015 705554 30027 711277
rect 38946 710223 38954 710248
rect 38946 707013 38954 707039
rect 30015 705544 30721 705554
rect 30015 705528 30718 705544
rect 31823 702940 32061 702972
rect 31481 702920 31797 702938
rect 36071 702505 36098 702995
rect 31481 701720 31797 701732
rect 31481 701716 32061 701720
rect 31823 701682 32061 701716
rect 20809 699718 20821 699774
rect 14744 698835 19490 698983
rect 698110 698217 702856 698365
rect 696779 697426 696791 697482
rect 685539 695484 685777 695518
rect 685539 695480 686119 695484
rect 685803 695468 686119 695480
rect 681502 694205 681529 694695
rect 685803 694262 686119 694280
rect 685539 694228 685777 694260
rect 686882 691656 687585 691672
rect 686879 691646 687585 691656
rect 678646 690161 678654 690187
rect 678646 686952 678654 686977
rect 687573 685923 687585 691646
rect 687645 686912 687648 692465
rect 698053 691267 698084 698191
rect 714726 698077 714752 698111
rect 699322 697674 700322 697700
rect 700922 697674 701922 697700
rect 699322 697527 700322 697629
rect 700922 697527 701922 697629
rect 707610 697101 708610 697241
rect 709211 697102 710211 697264
rect 687758 690189 687764 690637
rect 696817 690058 696821 691263
rect 687758 687117 687764 687591
rect 711579 685718 711595 697899
rect 714726 696843 714752 696877
rect 712409 685718 712431 692829
rect 707610 684937 708610 684978
rect 709211 684937 710211 684978
rect 699322 684306 700322 684461
rect 700922 684306 701922 684461
rect 707610 684206 708610 684416
rect 709211 684206 710211 684416
rect 699322 683981 700322 684136
rect 700922 683981 701922 684136
rect 711579 683893 711605 685675
rect 711579 683883 711619 683893
rect 711579 683869 712463 683883
rect 5137 670117 6021 670131
rect 5981 670107 6021 670117
rect 5995 668325 6021 670107
rect 15678 669864 16678 670019
rect 17278 669864 18278 670019
rect 7389 669584 8389 669794
rect 8990 669584 9990 669794
rect 15678 669539 16678 669694
rect 17278 669539 18278 669694
rect 7389 669022 8389 669063
rect 8990 669022 9990 669063
rect 5169 661171 5191 668282
rect 2848 657123 2874 657157
rect 6005 656101 6021 668282
rect 29836 666409 29842 666883
rect 20779 662737 20783 663942
rect 29836 663363 29842 663811
rect 7389 656736 8389 656898
rect 8990 656759 9990 656899
rect 15678 656371 16678 656473
rect 17278 656371 18278 656473
rect 15678 656300 16678 656326
rect 17278 656300 18278 656326
rect 2848 655889 2874 655923
rect 19516 655809 19547 662733
rect 29952 661535 29955 667088
rect 30015 662354 30027 668077
rect 38946 667023 38954 667048
rect 38946 663813 38954 663839
rect 30015 662344 30721 662354
rect 30015 662328 30718 662344
rect 31823 659740 32061 659772
rect 31481 659720 31797 659738
rect 36071 659305 36098 659795
rect 31481 658520 31797 658532
rect 31481 658516 32061 658520
rect 31823 658482 32061 658516
rect 20809 656518 20821 656574
rect 14744 655635 19490 655783
rect 698110 653017 702856 653165
rect 696779 652226 696791 652282
rect 685539 650284 685777 650318
rect 685539 650280 686119 650284
rect 685803 650268 686119 650280
rect 681502 649005 681529 649495
rect 685803 649062 686119 649080
rect 685539 649028 685777 649060
rect 686882 646456 687585 646472
rect 686879 646446 687585 646456
rect 678646 644961 678654 644987
rect 678646 641752 678654 641777
rect 687573 640723 687585 646446
rect 687645 641712 687648 647265
rect 698053 646067 698084 652991
rect 714726 652877 714752 652911
rect 699322 652474 700322 652500
rect 700922 652474 701922 652500
rect 699322 652327 700322 652429
rect 700922 652327 701922 652429
rect 707610 651901 708610 652041
rect 709211 651902 710211 652064
rect 687758 644989 687764 645437
rect 696817 644858 696821 646063
rect 687758 641917 687764 642391
rect 711579 640518 711595 652699
rect 714726 651643 714752 651677
rect 712409 640518 712431 647629
rect 707610 639737 708610 639778
rect 709211 639737 710211 639778
rect 699322 639106 700322 639261
rect 700922 639106 701922 639261
rect 707610 639006 708610 639216
rect 709211 639006 710211 639216
rect 699322 638781 700322 638936
rect 700922 638781 701922 638936
rect 711579 638693 711605 640475
rect 711579 638683 711619 638693
rect 711579 638669 712463 638683
rect 5137 626917 6021 626931
rect 5981 626907 6021 626917
rect 5995 625125 6021 626907
rect 15678 626664 16678 626819
rect 17278 626664 18278 626819
rect 7389 626384 8389 626594
rect 8990 626384 9990 626594
rect 15678 626339 16678 626494
rect 17278 626339 18278 626494
rect 7389 625822 8389 625863
rect 8990 625822 9990 625863
rect 5169 617971 5191 625082
rect 2848 613923 2874 613957
rect 6005 612901 6021 625082
rect 29836 623209 29842 623683
rect 20779 619537 20783 620742
rect 29836 620163 29842 620611
rect 7389 613536 8389 613698
rect 8990 613559 9990 613699
rect 15678 613171 16678 613273
rect 17278 613171 18278 613273
rect 15678 613100 16678 613126
rect 17278 613100 18278 613126
rect 2848 612689 2874 612723
rect 19516 612609 19547 619533
rect 29952 618335 29955 623888
rect 30015 619154 30027 624877
rect 38946 623823 38954 623848
rect 38946 620613 38954 620639
rect 30015 619144 30721 619154
rect 30015 619128 30718 619144
rect 31823 616540 32061 616572
rect 31481 616520 31797 616538
rect 36071 616105 36098 616595
rect 31481 615320 31797 615332
rect 31481 615316 32061 615320
rect 31823 615282 32061 615316
rect 20809 613318 20821 613374
rect 14744 612435 19490 612583
rect 698110 608017 702856 608165
rect 696779 607226 696791 607282
rect 685539 605284 685777 605318
rect 685539 605280 686119 605284
rect 685803 605268 686119 605280
rect 681502 604005 681529 604495
rect 685803 604062 686119 604080
rect 685539 604028 685777 604060
rect 686882 601456 687585 601472
rect 686879 601446 687585 601456
rect 678646 599961 678654 599987
rect 678646 596752 678654 596777
rect 687573 595723 687585 601446
rect 687645 596712 687648 602265
rect 698053 601067 698084 607991
rect 714726 607877 714752 607911
rect 699322 607474 700322 607500
rect 700922 607474 701922 607500
rect 699322 607327 700322 607429
rect 700922 607327 701922 607429
rect 707610 606901 708610 607041
rect 709211 606902 710211 607064
rect 687758 599989 687764 600437
rect 696817 599858 696821 601063
rect 687758 596917 687764 597391
rect 711579 595518 711595 607699
rect 714726 606643 714752 606677
rect 712409 595518 712431 602629
rect 707610 594737 708610 594778
rect 709211 594737 710211 594778
rect 699322 594106 700322 594261
rect 700922 594106 701922 594261
rect 707610 594006 708610 594216
rect 709211 594006 710211 594216
rect 699322 593781 700322 593936
rect 700922 593781 701922 593936
rect 711579 593693 711605 595475
rect 711579 593683 711619 593693
rect 711579 593669 712463 593683
rect 5137 583717 6021 583731
rect 5981 583707 6021 583717
rect 5995 581925 6021 583707
rect 15678 583464 16678 583619
rect 17278 583464 18278 583619
rect 7389 583184 8389 583394
rect 8990 583184 9990 583394
rect 15678 583139 16678 583294
rect 17278 583139 18278 583294
rect 7389 582622 8389 582663
rect 8990 582622 9990 582663
rect 5169 574771 5191 581882
rect 2848 570723 2874 570757
rect 6005 569701 6021 581882
rect 29836 580009 29842 580483
rect 20779 576337 20783 577542
rect 29836 576963 29842 577411
rect 7389 570336 8389 570498
rect 8990 570359 9990 570499
rect 15678 569971 16678 570073
rect 17278 569971 18278 570073
rect 15678 569900 16678 569926
rect 17278 569900 18278 569926
rect 2848 569489 2874 569523
rect 19516 569409 19547 576333
rect 29952 575135 29955 580688
rect 30015 575954 30027 581677
rect 38946 580623 38954 580648
rect 38946 577413 38954 577439
rect 30015 575944 30721 575954
rect 30015 575928 30718 575944
rect 31823 573340 32061 573372
rect 31481 573320 31797 573338
rect 36071 572905 36098 573395
rect 31481 572120 31797 572132
rect 31481 572116 32061 572120
rect 31823 572082 32061 572116
rect 20809 570118 20821 570174
rect 14744 569235 19490 569383
rect 698110 562817 702856 562965
rect 696779 562026 696791 562082
rect 685539 560084 685777 560118
rect 685539 560080 686119 560084
rect 685803 560068 686119 560080
rect 681502 558805 681529 559295
rect 685803 558862 686119 558880
rect 685539 558828 685777 558860
rect 686882 556256 687585 556272
rect 686879 556246 687585 556256
rect 678646 554761 678654 554787
rect 678646 551552 678654 551577
rect 687573 550523 687585 556246
rect 687645 551512 687648 557065
rect 698053 555867 698084 562791
rect 714726 562677 714752 562711
rect 699322 562274 700322 562300
rect 700922 562274 701922 562300
rect 699322 562127 700322 562229
rect 700922 562127 701922 562229
rect 707610 561701 708610 561841
rect 709211 561702 710211 561864
rect 687758 554789 687764 555237
rect 696817 554658 696821 555863
rect 687758 551717 687764 552191
rect 711579 550318 711595 562499
rect 714726 561443 714752 561477
rect 712409 550318 712431 557429
rect 707610 549537 708610 549578
rect 709211 549537 710211 549578
rect 699322 548906 700322 549061
rect 700922 548906 701922 549061
rect 707610 548806 708610 549016
rect 709211 548806 710211 549016
rect 699322 548581 700322 548736
rect 700922 548581 701922 548736
rect 711579 548493 711605 550275
rect 711579 548483 711619 548493
rect 711579 548469 712463 548483
rect 5137 540517 6021 540531
rect 5981 540507 6021 540517
rect 5995 538725 6021 540507
rect 15678 540264 16678 540419
rect 17278 540264 18278 540419
rect 7389 539984 8389 540194
rect 8990 539984 9990 540194
rect 15678 539939 16678 540094
rect 17278 539939 18278 540094
rect 7389 539422 8389 539463
rect 8990 539422 9990 539463
rect 5169 531571 5191 538682
rect 2848 527523 2874 527557
rect 6005 526501 6021 538682
rect 29836 536809 29842 537283
rect 20779 533137 20783 534342
rect 29836 533763 29842 534211
rect 7389 527136 8389 527298
rect 8990 527159 9990 527299
rect 15678 526771 16678 526873
rect 17278 526771 18278 526873
rect 15678 526700 16678 526726
rect 17278 526700 18278 526726
rect 2848 526289 2874 526323
rect 19516 526209 19547 533133
rect 29952 531935 29955 537488
rect 30015 532754 30027 538477
rect 38946 537423 38954 537448
rect 38946 534213 38954 534239
rect 30015 532744 30721 532754
rect 30015 532728 30718 532744
rect 31823 530140 32061 530172
rect 31481 530120 31797 530138
rect 36071 529705 36098 530195
rect 31481 528920 31797 528932
rect 31481 528916 32061 528920
rect 31823 528882 32061 528916
rect 20809 526918 20821 526974
rect 14744 526035 19490 526183
rect 678282 471387 681670 471445
rect 678282 467471 681670 467485
rect 35930 448115 39318 448129
rect 35930 444155 39318 444213
rect 5137 412917 6021 412931
rect 5981 412907 6021 412917
rect 5995 411125 6021 412907
rect 15678 412664 16678 412819
rect 17278 412664 18278 412819
rect 7389 412384 8389 412594
rect 8990 412384 9990 412594
rect 15678 412339 16678 412494
rect 17278 412339 18278 412494
rect 7389 411822 8389 411863
rect 8990 411822 9990 411863
rect 5169 403971 5191 411082
rect 2848 399923 2874 399957
rect 6005 398901 6021 411082
rect 29836 409209 29842 409683
rect 20779 405537 20783 406742
rect 29836 406163 29842 406611
rect 7389 399536 8389 399698
rect 8990 399559 9990 399699
rect 15678 399171 16678 399273
rect 17278 399171 18278 399273
rect 15678 399100 16678 399126
rect 17278 399100 18278 399126
rect 2848 398689 2874 398723
rect 19516 398609 19547 405533
rect 29952 404335 29955 409888
rect 30015 405154 30027 410877
rect 38946 409823 38954 409848
rect 38946 406613 38954 406639
rect 30015 405144 30721 405154
rect 30015 405128 30718 405144
rect 31823 402540 32061 402572
rect 31481 402520 31797 402538
rect 36071 402105 36098 402595
rect 31481 401320 31797 401332
rect 31481 401316 32061 401320
rect 31823 401282 32061 401316
rect 20809 399318 20821 399374
rect 14744 398435 19490 398583
rect 698110 385617 702856 385765
rect 696779 384826 696791 384882
rect 685539 382884 685777 382918
rect 685539 382880 686119 382884
rect 685803 382868 686119 382880
rect 681502 381605 681529 382095
rect 685803 381662 686119 381680
rect 685539 381628 685777 381660
rect 686882 379056 687585 379072
rect 686879 379046 687585 379056
rect 678646 377561 678654 377587
rect 678646 374352 678654 374377
rect 687573 373323 687585 379046
rect 687645 374312 687648 379865
rect 698053 378667 698084 385591
rect 714726 385477 714752 385511
rect 699322 385074 700322 385100
rect 700922 385074 701922 385100
rect 699322 384927 700322 385029
rect 700922 384927 701922 385029
rect 707610 384501 708610 384641
rect 709211 384502 710211 384664
rect 687758 377589 687764 378037
rect 696817 377458 696821 378663
rect 687758 374517 687764 374991
rect 711579 373118 711595 385299
rect 714726 384243 714752 384277
rect 712409 373118 712431 380229
rect 707610 372337 708610 372378
rect 709211 372337 710211 372378
rect 699322 371706 700322 371861
rect 700922 371706 701922 371861
rect 707610 371606 708610 371816
rect 709211 371606 710211 371816
rect 699322 371381 700322 371536
rect 700922 371381 701922 371536
rect 711579 371293 711605 373075
rect 711579 371283 711619 371293
rect 711579 371269 712463 371283
rect 5137 369717 6021 369731
rect 5981 369707 6021 369717
rect 5995 367925 6021 369707
rect 15678 369464 16678 369619
rect 17278 369464 18278 369619
rect 7389 369184 8389 369394
rect 8990 369184 9990 369394
rect 15678 369139 16678 369294
rect 17278 369139 18278 369294
rect 7389 368622 8389 368663
rect 8990 368622 9990 368663
rect 5169 360771 5191 367882
rect 2848 356723 2874 356757
rect 6005 355701 6021 367882
rect 29836 366009 29842 366483
rect 20779 362337 20783 363542
rect 29836 362963 29842 363411
rect 7389 356336 8389 356498
rect 8990 356359 9990 356499
rect 15678 355971 16678 356073
rect 17278 355971 18278 356073
rect 15678 355900 16678 355926
rect 17278 355900 18278 355926
rect 2848 355489 2874 355523
rect 19516 355409 19547 362333
rect 29952 361135 29955 366688
rect 30015 361954 30027 367677
rect 38946 366623 38954 366648
rect 38946 363413 38954 363439
rect 30015 361944 30721 361954
rect 30015 361928 30718 361944
rect 31823 359340 32061 359372
rect 31481 359320 31797 359338
rect 36071 358905 36098 359395
rect 31481 358120 31797 358132
rect 31481 358116 32061 358120
rect 31823 358082 32061 358116
rect 20809 356118 20821 356174
rect 14744 355235 19490 355383
rect 698110 340417 702856 340565
rect 696779 339626 696791 339682
rect 685539 337684 685777 337718
rect 685539 337680 686119 337684
rect 685803 337668 686119 337680
rect 681502 336405 681529 336895
rect 685803 336462 686119 336480
rect 685539 336428 685777 336460
rect 686882 333856 687585 333872
rect 686879 333846 687585 333856
rect 678646 332361 678654 332387
rect 678646 329152 678654 329177
rect 687573 328123 687585 333846
rect 687645 329112 687648 334665
rect 698053 333467 698084 340391
rect 714726 340277 714752 340311
rect 699322 339874 700322 339900
rect 700922 339874 701922 339900
rect 699322 339727 700322 339829
rect 700922 339727 701922 339829
rect 707610 339301 708610 339441
rect 709211 339302 710211 339464
rect 687758 332389 687764 332837
rect 696817 332258 696821 333463
rect 687758 329317 687764 329791
rect 711579 327918 711595 340099
rect 714726 339043 714752 339077
rect 712409 327918 712431 335029
rect 707610 327137 708610 327178
rect 709211 327137 710211 327178
rect 5137 326517 6021 326531
rect 5981 326507 6021 326517
rect 5995 324725 6021 326507
rect 699322 326506 700322 326661
rect 700922 326506 701922 326661
rect 15678 326264 16678 326419
rect 17278 326264 18278 326419
rect 707610 326406 708610 326616
rect 709211 326406 710211 326616
rect 7389 325984 8389 326194
rect 8990 325984 9990 326194
rect 699322 326181 700322 326336
rect 700922 326181 701922 326336
rect 15678 325939 16678 326094
rect 17278 325939 18278 326094
rect 711579 326093 711605 327875
rect 711579 326083 711619 326093
rect 711579 326069 712463 326083
rect 7389 325422 8389 325463
rect 8990 325422 9990 325463
rect 5169 317571 5191 324682
rect 2848 313523 2874 313557
rect 6005 312501 6021 324682
rect 29836 322809 29842 323283
rect 20779 319137 20783 320342
rect 29836 319763 29842 320211
rect 7389 313136 8389 313298
rect 8990 313159 9990 313299
rect 15678 312771 16678 312873
rect 17278 312771 18278 312873
rect 15678 312700 16678 312726
rect 17278 312700 18278 312726
rect 2848 312289 2874 312323
rect 19516 312209 19547 319133
rect 29952 317935 29955 323488
rect 30015 318754 30027 324477
rect 38946 323423 38954 323448
rect 38946 320213 38954 320239
rect 30015 318744 30721 318754
rect 30015 318728 30718 318744
rect 31823 316140 32061 316172
rect 31481 316120 31797 316138
rect 36071 315705 36098 316195
rect 31481 314920 31797 314932
rect 31481 314916 32061 314920
rect 31823 314882 32061 314916
rect 20809 312918 20821 312974
rect 14744 312035 19490 312183
rect 698110 295417 702856 295565
rect 696779 294626 696791 294682
rect 685539 292684 685777 292718
rect 685539 292680 686119 292684
rect 685803 292668 686119 292680
rect 681502 291405 681529 291895
rect 685803 291462 686119 291480
rect 685539 291428 685777 291460
rect 686882 288856 687585 288872
rect 686879 288846 687585 288856
rect 678646 287361 678654 287387
rect 678646 284152 678654 284177
rect 5137 283317 6021 283331
rect 5981 283307 6021 283317
rect 5995 281525 6021 283307
rect 15678 283064 16678 283219
rect 17278 283064 18278 283219
rect 687573 283123 687585 288846
rect 687645 284112 687648 289665
rect 698053 288467 698084 295391
rect 714726 295277 714752 295311
rect 699322 294874 700322 294900
rect 700922 294874 701922 294900
rect 699322 294727 700322 294829
rect 700922 294727 701922 294829
rect 707610 294301 708610 294441
rect 709211 294302 710211 294464
rect 687758 287389 687764 287837
rect 696817 287258 696821 288463
rect 687758 284317 687764 284791
rect 7389 282784 8389 282994
rect 8990 282784 9990 282994
rect 711579 282918 711595 295099
rect 714726 294043 714752 294077
rect 712409 282918 712431 290029
rect 15678 282739 16678 282894
rect 17278 282739 18278 282894
rect 7389 282222 8389 282263
rect 8990 282222 9990 282263
rect 707610 282137 708610 282178
rect 709211 282137 710211 282178
rect 699322 281506 700322 281661
rect 700922 281506 701922 281661
rect 5169 274371 5191 281482
rect 2848 270323 2874 270357
rect 6005 269301 6021 281482
rect 707610 281406 708610 281616
rect 709211 281406 710211 281616
rect 29836 279609 29842 280083
rect 20779 275937 20783 277142
rect 29836 276563 29842 277011
rect 7389 269936 8389 270098
rect 8990 269959 9990 270099
rect 15678 269571 16678 269673
rect 17278 269571 18278 269673
rect 15678 269500 16678 269526
rect 17278 269500 18278 269526
rect 2848 269089 2874 269123
rect 19516 269009 19547 275933
rect 29952 274735 29955 280288
rect 30015 275554 30027 281277
rect 699322 281181 700322 281336
rect 700922 281181 701922 281336
rect 711579 281093 711605 282875
rect 711579 281083 711619 281093
rect 711579 281069 712463 281083
rect 38946 280223 38954 280248
rect 38946 277013 38954 277039
rect 30015 275544 30721 275554
rect 30015 275528 30718 275544
rect 31823 272940 32061 272972
rect 31481 272920 31797 272938
rect 36071 272505 36098 272995
rect 31481 271720 31797 271732
rect 31481 271716 32061 271720
rect 31823 271682 32061 271716
rect 20809 269718 20821 269774
rect 14744 268835 19490 268983
rect 698110 250417 702856 250565
rect 696779 249626 696791 249682
rect 685539 247684 685777 247718
rect 685539 247680 686119 247684
rect 685803 247668 686119 247680
rect 681502 246405 681529 246895
rect 685803 246462 686119 246480
rect 685539 246428 685777 246460
rect 686882 243856 687585 243872
rect 686879 243846 687585 243856
rect 678646 242361 678654 242387
rect 5137 240117 6021 240131
rect 5981 240107 6021 240117
rect 5995 238325 6021 240107
rect 15678 239864 16678 240019
rect 17278 239864 18278 240019
rect 7389 239584 8389 239794
rect 8990 239584 9990 239794
rect 15678 239539 16678 239694
rect 17278 239539 18278 239694
rect 678646 239152 678654 239177
rect 7389 239022 8389 239063
rect 8990 239022 9990 239063
rect 5169 231171 5191 238282
rect 2848 227123 2874 227157
rect 6005 226101 6021 238282
rect 687573 238123 687585 243846
rect 687645 239112 687648 244665
rect 698053 243467 698084 250391
rect 714726 250277 714752 250311
rect 699322 249874 700322 249900
rect 700922 249874 701922 249900
rect 699322 249727 700322 249829
rect 700922 249727 701922 249829
rect 707610 249301 708610 249441
rect 709211 249302 710211 249464
rect 687758 242389 687764 242837
rect 696817 242258 696821 243463
rect 687758 239317 687764 239791
rect 29836 236409 29842 236883
rect 20779 232737 20783 233942
rect 29836 233363 29842 233811
rect 7389 226736 8389 226898
rect 8990 226759 9990 226899
rect 15678 226371 16678 226473
rect 17278 226371 18278 226473
rect 15678 226300 16678 226326
rect 17278 226300 18278 226326
rect 2848 225889 2874 225923
rect 19516 225809 19547 232733
rect 29952 231535 29955 237088
rect 30015 232354 30027 238077
rect 711579 237918 711595 250099
rect 714726 249043 714752 249077
rect 712409 237918 712431 245029
rect 707610 237137 708610 237178
rect 709211 237137 710211 237178
rect 38946 237023 38954 237048
rect 699322 236506 700322 236661
rect 700922 236506 701922 236661
rect 707610 236406 708610 236616
rect 709211 236406 710211 236616
rect 699322 236181 700322 236336
rect 700922 236181 701922 236336
rect 711579 236093 711605 237875
rect 711579 236083 711619 236093
rect 711579 236069 712463 236083
rect 38946 233813 38954 233839
rect 30015 232344 30721 232354
rect 30015 232328 30718 232344
rect 31823 229740 32061 229772
rect 31481 229720 31797 229738
rect 36071 229305 36098 229795
rect 31481 228520 31797 228532
rect 31481 228516 32061 228520
rect 31823 228482 32061 228516
rect 20809 226518 20821 226574
rect 14744 225635 19490 225783
rect 698110 205217 702856 205365
rect 696779 204426 696791 204482
rect 685539 202484 685777 202518
rect 685539 202480 686119 202484
rect 685803 202468 686119 202480
rect 681502 201205 681529 201695
rect 685803 201262 686119 201280
rect 685539 201228 685777 201260
rect 686882 198656 687585 198672
rect 686879 198646 687585 198656
rect 678646 197161 678654 197187
rect 5137 196917 6021 196931
rect 5981 196907 6021 196917
rect 5995 195125 6021 196907
rect 15678 196664 16678 196819
rect 17278 196664 18278 196819
rect 7389 196384 8389 196594
rect 8990 196384 9990 196594
rect 15678 196339 16678 196494
rect 17278 196339 18278 196494
rect 7389 195822 8389 195863
rect 8990 195822 9990 195863
rect 5169 187971 5191 195082
rect 2848 183923 2874 183957
rect 6005 182901 6021 195082
rect 29836 193209 29842 193683
rect 20779 189537 20783 190742
rect 29836 190163 29842 190611
rect 7389 183536 8389 183698
rect 8990 183559 9990 183699
rect 15678 183171 16678 183273
rect 17278 183171 18278 183273
rect 15678 183100 16678 183126
rect 17278 183100 18278 183126
rect 2848 182689 2874 182723
rect 19516 182609 19547 189533
rect 29952 188335 29955 193888
rect 30015 189154 30027 194877
rect 678646 193952 678654 193977
rect 38946 193823 38954 193848
rect 687573 192923 687585 198646
rect 687645 193912 687648 199465
rect 698053 198267 698084 205191
rect 714726 205077 714752 205111
rect 699322 204674 700322 204700
rect 700922 204674 701922 204700
rect 699322 204527 700322 204629
rect 700922 204527 701922 204629
rect 707610 204101 708610 204241
rect 709211 204102 710211 204264
rect 687758 197189 687764 197637
rect 696817 197058 696821 198263
rect 687758 194117 687764 194591
rect 711579 192718 711595 204899
rect 714726 203843 714752 203877
rect 712409 192718 712431 199829
rect 707610 191937 708610 191978
rect 709211 191937 710211 191978
rect 699322 191306 700322 191461
rect 700922 191306 701922 191461
rect 707610 191206 708610 191416
rect 709211 191206 710211 191416
rect 699322 190981 700322 191136
rect 700922 190981 701922 191136
rect 711579 190893 711605 192675
rect 711579 190883 711619 190893
rect 711579 190869 712463 190883
rect 38946 190613 38954 190639
rect 30015 189144 30721 189154
rect 30015 189128 30718 189144
rect 31823 186540 32061 186572
rect 31481 186520 31797 186538
rect 36071 186105 36098 186595
rect 31481 185320 31797 185332
rect 31481 185316 32061 185320
rect 31823 185282 32061 185316
rect 20809 183318 20821 183374
rect 14744 182435 19490 182583
rect 698110 160217 702856 160365
rect 696779 159426 696791 159482
rect 685539 157484 685777 157518
rect 685539 157480 686119 157484
rect 685803 157468 686119 157480
rect 681502 156205 681529 156695
rect 685803 156262 686119 156280
rect 685539 156228 685777 156260
rect 686882 153656 687585 153672
rect 686879 153646 687585 153656
rect 678646 152161 678654 152187
rect 678646 148952 678654 148977
rect 687573 147923 687585 153646
rect 687645 148912 687648 154465
rect 698053 153267 698084 160191
rect 714726 160077 714752 160111
rect 699322 159674 700322 159700
rect 700922 159674 701922 159700
rect 699322 159527 700322 159629
rect 700922 159527 701922 159629
rect 707610 159101 708610 159241
rect 709211 159102 710211 159264
rect 687758 152189 687764 152637
rect 696817 152058 696821 153263
rect 687758 149117 687764 149591
rect 711579 147718 711595 159899
rect 714726 158843 714752 158877
rect 712409 147718 712431 154829
rect 707610 146937 708610 146978
rect 709211 146937 710211 146978
rect 699322 146306 700322 146461
rect 700922 146306 701922 146461
rect 707610 146206 708610 146416
rect 709211 146206 710211 146416
rect 699322 145981 700322 146136
rect 700922 145981 701922 146136
rect 711579 145893 711605 147675
rect 711579 145883 711619 145893
rect 711579 145869 712463 145883
rect 698110 115017 702856 115165
rect 696779 114226 696791 114282
rect 685539 112284 685777 112318
rect 685539 112280 686119 112284
rect 685803 112268 686119 112280
rect 681502 111005 681529 111495
rect 685803 111062 686119 111080
rect 685539 111028 685777 111060
rect 686882 108456 687585 108472
rect 686879 108446 687585 108456
rect 678646 106961 678654 106987
rect 678646 103752 678654 103777
rect 687573 102723 687585 108446
rect 687645 103712 687648 109265
rect 698053 108067 698084 114991
rect 714726 114877 714752 114911
rect 699322 114474 700322 114500
rect 700922 114474 701922 114500
rect 699322 114327 700322 114429
rect 700922 114327 701922 114429
rect 707610 113901 708610 114041
rect 709211 113902 710211 114064
rect 687758 106989 687764 107437
rect 696817 106858 696821 108063
rect 687758 103917 687764 104391
rect 711579 102518 711595 114699
rect 714726 113643 714752 113677
rect 712409 102518 712431 109629
rect 707610 101737 708610 101778
rect 709211 101737 710211 101778
rect 699322 101106 700322 101261
rect 700922 101106 701922 101261
rect 707610 101006 708610 101216
rect 709211 101006 710211 101216
rect 699322 100781 700322 100936
rect 700922 100781 701922 100936
rect 711579 100693 711605 102475
rect 711579 100683 711619 100693
rect 711579 100669 712463 100683
rect 35930 75315 39318 75329
rect 35930 71355 39318 71413
rect 190152 38946 190177 38954
rect 193361 38946 193387 38954
rect 146187 38280 146453 38291
rect 144718 36866 144738 37390
rect 197405 36071 197895 36098
rect 248871 35930 248885 39318
rect 252787 35930 252845 39318
rect 298752 38946 298777 38954
rect 301961 38946 301987 38954
rect 353552 38946 353577 38954
rect 356761 38946 356787 38954
rect 408352 38946 408377 38954
rect 411561 38946 411587 38954
rect 463152 38946 463177 38954
rect 466361 38946 466387 38954
rect 517952 38946 517977 38954
rect 521161 38946 521187 38954
rect 306005 36071 306495 36098
rect 360805 36071 361295 36098
rect 415605 36071 416095 36098
rect 470405 36071 470895 36098
rect 525205 36071 525695 36098
rect 143407 35902 143463 35923
rect 143407 35793 143429 35902
rect 197428 31823 197460 32061
rect 198680 31823 198718 32061
rect 306028 31823 306060 32061
rect 307280 31823 307318 32061
rect 360828 31823 360860 32061
rect 362080 31823 362118 32061
rect 415628 31823 415660 32061
rect 416880 31823 416918 32061
rect 470428 31823 470460 32061
rect 471680 31823 471718 32061
rect 525228 31823 525260 32061
rect 526480 31823 526518 32061
rect 198680 31797 198684 31823
rect 307280 31797 307284 31823
rect 362080 31797 362084 31823
rect 416880 31797 416884 31823
rect 471680 31797 471684 31823
rect 526480 31797 526484 31823
rect 197462 31481 197480 31797
rect 198668 31481 198684 31797
rect 306062 31481 306080 31797
rect 307268 31481 307284 31797
rect 360862 31481 360880 31797
rect 362068 31481 362084 31797
rect 415662 31481 415680 31797
rect 416868 31481 416884 31797
rect 470462 31481 470480 31797
rect 471668 31481 471684 31797
rect 525262 31481 525280 31797
rect 526468 31481 526484 31797
rect 194846 30718 194856 30721
rect 303446 30718 303456 30721
rect 358246 30718 358256 30721
rect 413046 30718 413056 30721
rect 467846 30718 467856 30721
rect 522646 30718 522656 30721
rect 194846 30027 194872 30718
rect 303446 30027 303472 30718
rect 358246 30027 358272 30718
rect 413046 30027 413072 30718
rect 467846 30027 467872 30718
rect 522646 30027 522672 30718
rect 189123 30015 194872 30027
rect 297723 30015 303472 30027
rect 352523 30015 358272 30027
rect 407323 30015 413072 30027
rect 462123 30015 467872 30027
rect 516923 30015 522672 30027
rect 190112 29952 195665 29955
rect 298712 29952 304265 29955
rect 353512 29952 359065 29955
rect 408312 29952 413865 29955
rect 463112 29952 468665 29955
rect 517912 29952 523465 29955
rect 190317 29836 190791 29842
rect 193389 29836 193837 29842
rect 298917 29836 299391 29842
rect 301989 29836 302437 29842
rect 353717 29836 354191 29842
rect 356789 29836 357237 29842
rect 408517 29836 408991 29842
rect 411589 29836 412037 29842
rect 463317 29836 463791 29842
rect 466389 29836 466837 29842
rect 518117 29836 518591 29842
rect 521189 29836 521637 29842
rect 200626 20809 200682 20821
rect 309226 20809 309282 20821
rect 364026 20809 364082 20821
rect 418826 20809 418882 20821
rect 473626 20809 473682 20821
rect 528426 20809 528482 20821
rect 193258 20779 194463 20783
rect 301858 20779 303063 20783
rect 356658 20779 357863 20783
rect 411458 20779 412663 20783
rect 466258 20779 467463 20783
rect 521058 20779 522263 20783
rect 147509 19547 147573 19618
rect 194467 19516 201391 19547
rect 303067 19516 309991 19547
rect 357867 19516 364791 19547
rect 412667 19516 419591 19547
rect 467467 19516 474391 19547
rect 522267 19516 529191 19547
rect 133241 17478 133396 18478
rect 133566 17478 133721 18478
rect 146787 17478 146889 18478
rect 146934 17478 146960 18478
rect 187181 17278 187336 18278
rect 187506 17278 187661 18278
rect 200727 17278 200829 18278
rect 200874 17278 200900 18278
rect 133241 15878 133396 16878
rect 133566 15878 133721 16878
rect 146787 15878 146889 16878
rect 146934 15878 146960 16878
rect 187181 15678 187336 16678
rect 187506 15678 187661 16678
rect 200727 15678 200829 16678
rect 200874 15678 200900 16678
rect 201417 14744 201565 19490
rect 295781 17278 295936 18278
rect 296106 17278 296261 18278
rect 309327 17278 309429 18278
rect 309474 17278 309500 18278
rect 295781 15678 295936 16678
rect 296106 15678 296261 16678
rect 309327 15678 309429 16678
rect 309474 15678 309500 16678
rect 310017 14744 310165 19490
rect 350581 17278 350736 18278
rect 350906 17278 351061 18278
rect 364127 17278 364229 18278
rect 364274 17278 364300 18278
rect 350581 15678 350736 16678
rect 350906 15678 351061 16678
rect 364127 15678 364229 16678
rect 364274 15678 364300 16678
rect 364817 14744 364965 19490
rect 405381 17278 405536 18278
rect 405706 17278 405861 18278
rect 418927 17278 419029 18278
rect 419074 17278 419100 18278
rect 405381 15678 405536 16678
rect 405706 15678 405861 16678
rect 418927 15678 419029 16678
rect 419074 15678 419100 16678
rect 419617 14744 419765 19490
rect 460181 17278 460336 18278
rect 460506 17278 460661 18278
rect 473727 17278 473829 18278
rect 473874 17278 473900 18278
rect 460181 15678 460336 16678
rect 460506 15678 460661 16678
rect 473727 15678 473829 16678
rect 473874 15678 473900 16678
rect 474417 14744 474565 19490
rect 514981 17278 515136 18278
rect 515306 17278 515461 18278
rect 528527 17278 528629 18278
rect 528674 17278 528700 18278
rect 514981 15678 515136 16678
rect 515306 15678 515461 16678
rect 528527 15678 528629 16678
rect 528674 15678 528700 16678
rect 529217 14744 529365 19490
rect 133606 8990 133816 9990
rect 134337 8990 134378 9990
rect 146501 8990 146641 9990
rect 187406 8990 187616 9990
rect 188137 8990 188178 9990
rect 200301 8990 200441 9990
rect 296006 8990 296216 9990
rect 296737 8990 296778 9990
rect 308901 8990 309041 9990
rect 350806 8990 351016 9990
rect 351537 8990 351578 9990
rect 363701 8990 363841 9990
rect 405606 8990 405816 9990
rect 406337 8990 406378 9990
rect 418501 8990 418641 9990
rect 460406 8990 460616 9990
rect 461137 8990 461178 9990
rect 473301 8990 473441 9990
rect 515206 8990 515416 9990
rect 515937 8990 515978 9990
rect 528101 8990 528241 9990
rect 133606 7389 133816 8389
rect 134337 7389 134378 8389
rect 146502 7389 146664 8389
rect 187406 7389 187616 8389
rect 188137 7389 188178 8389
rect 200302 7389 200464 8389
rect 296006 7389 296216 8389
rect 296737 7389 296778 8389
rect 308902 7389 309064 8389
rect 350806 7389 351016 8389
rect 351537 7389 351578 8389
rect 363702 7389 363864 8389
rect 405606 7389 405816 8389
rect 406337 7389 406378 8389
rect 418502 7389 418664 8389
rect 460406 7389 460616 8389
rect 461137 7389 461178 8389
rect 473302 7389 473464 8389
rect 515206 7389 515416 8389
rect 515937 7389 515978 8389
rect 528102 7389 528264 8389
rect 187069 5995 188875 6021
rect 188918 6005 201099 6021
rect 295669 5995 297475 6021
rect 297518 6005 309699 6021
rect 350469 5995 352275 6021
rect 352318 6005 364499 6021
rect 405269 5995 407075 6021
rect 407118 6005 419299 6021
rect 460069 5995 461875 6021
rect 461918 6005 474099 6021
rect 514869 5995 516675 6021
rect 516718 6005 528899 6021
rect 187069 5981 187093 5995
rect 295669 5981 295693 5995
rect 350469 5981 350493 5995
rect 405269 5981 405293 5995
rect 460069 5981 460093 5995
rect 514869 5981 514893 5995
rect 187069 5137 187083 5981
rect 188918 5169 196029 5191
rect 295669 5137 295683 5981
rect 297518 5169 304629 5191
rect 350469 5137 350483 5981
rect 352318 5169 359429 5191
rect 405269 5137 405283 5981
rect 407118 5169 414229 5191
rect 460069 5137 460083 5981
rect 461918 5169 469029 5191
rect 514869 5137 514883 5981
rect 516718 5169 523829 5191
rect 200043 2848 200077 2874
rect 201277 2848 201311 2874
rect 308643 2848 308677 2874
rect 309877 2848 309911 2874
rect 363443 2848 363477 2874
rect 364677 2848 364711 2874
rect 418243 2848 418277 2874
rect 419477 2848 419511 2874
rect 473043 2848 473077 2874
rect 474277 2848 474311 2874
rect 527843 2848 527877 2874
rect 529077 2848 529111 2874
<< metal1 >>
rect 84010 995596 84016 995648
rect 84068 995636 84074 995648
rect 91738 995636 91744 995648
rect 84068 995608 91744 995636
rect 84068 995596 84074 995608
rect 91738 995596 91744 995608
rect 91796 995596 91802 995648
rect 238202 995596 238208 995648
rect 238260 995636 238266 995648
rect 245930 995636 245936 995648
rect 238260 995608 245936 995636
rect 238260 995596 238266 995608
rect 245930 995596 245936 995608
rect 245988 995596 245994 995648
rect 531958 995596 531964 995648
rect 532016 995636 532022 995648
rect 539686 995636 539692 995648
rect 532016 995608 539692 995636
rect 532016 995596 532022 995608
rect 539686 995596 539692 995608
rect 539744 995596 539750 995648
rect 135346 995460 135352 995512
rect 135404 995500 135410 995512
rect 143166 995500 143172 995512
rect 135404 995472 143172 995500
rect 135404 995460 135410 995472
rect 143166 995460 143172 995472
rect 143224 995460 143230 995512
rect 633802 995460 633808 995512
rect 633860 995500 633866 995512
rect 641530 995500 641536 995512
rect 633860 995472 641536 995500
rect 633860 995460 633866 995472
rect 641530 995460 641536 995472
rect 641588 995460 641594 995512
rect 289630 995256 289636 995308
rect 289688 995296 289694 995308
rect 297634 995296 297640 995308
rect 289688 995268 297640 995296
rect 289688 995256 289694 995268
rect 297634 995256 297640 995268
rect 297692 995256 297698 995308
rect 391474 995256 391480 995308
rect 391532 995296 391538 995308
rect 399478 995296 399484 995308
rect 391532 995268 399484 995296
rect 391532 995256 391538 995268
rect 399478 995256 399484 995268
rect 399536 995256 399542 995308
rect 480438 995256 480444 995308
rect 480496 995296 480502 995308
rect 488442 995296 488448 995308
rect 480496 995268 488448 995296
rect 480496 995256 480502 995268
rect 488442 995256 488448 995268
rect 488500 995256 488506 995308
rect 82630 992060 82636 992112
rect 82688 992100 82694 992112
rect 89990 992100 89996 992112
rect 82688 992072 89996 992100
rect 82688 992060 82694 992072
rect 89990 992060 89996 992072
rect 90048 992060 90054 992112
rect 79502 990768 79508 990820
rect 79560 990808 79566 990820
rect 130930 990808 130936 990820
rect 79560 990780 130936 990808
rect 79560 990768 79566 990780
rect 130930 990768 130936 990780
rect 130988 990808 130994 990820
rect 131114 990808 131120 990820
rect 130988 990780 131120 990808
rect 130988 990768 130994 990780
rect 131114 990768 131120 990780
rect 131172 990768 131178 990820
rect 186682 990768 186688 990820
rect 186740 990808 186746 990820
rect 194686 990808 194692 990820
rect 186740 990780 194692 990808
rect 186740 990768 186746 990780
rect 194686 990768 194692 990780
rect 194744 990768 194750 990820
rect 194778 990768 194784 990820
rect 194836 990808 194842 990820
rect 233050 990808 233056 990820
rect 194836 990780 233056 990808
rect 194836 990768 194842 990780
rect 233050 990768 233056 990780
rect 233108 990808 233114 990820
rect 284662 990808 284668 990820
rect 233108 990780 284668 990808
rect 233108 990768 233114 990780
rect 284662 990768 284668 990780
rect 284720 990808 284726 990820
rect 386506 990808 386512 990820
rect 284720 990780 386512 990808
rect 284720 990768 284726 990780
rect 386506 990768 386512 990780
rect 386564 990768 386570 990820
rect 486602 990768 486608 990820
rect 486660 990808 486666 990820
rect 538030 990808 538036 990820
rect 486660 990780 538036 990808
rect 486660 990768 486666 990780
rect 538030 990768 538036 990780
rect 538088 990808 538094 990820
rect 639782 990808 639788 990820
rect 538088 990780 639788 990808
rect 538088 990768 538094 990780
rect 639782 990768 639788 990780
rect 639840 990768 639846 990820
rect 78858 990700 78864 990752
rect 78916 990740 78922 990752
rect 130286 990740 130292 990752
rect 78916 990712 130292 990740
rect 78916 990700 78922 990712
rect 130286 990700 130292 990712
rect 130344 990700 130350 990752
rect 182358 990700 182364 990752
rect 182416 990740 182422 990752
rect 200022 990740 200028 990752
rect 182416 990712 200028 990740
rect 182416 990700 182422 990712
rect 200022 990700 200028 990712
rect 200080 990700 200086 990752
rect 244182 990700 244188 990752
rect 244240 990740 244246 990752
rect 295794 990740 295800 990752
rect 244240 990712 295800 990740
rect 244240 990700 244246 990712
rect 295794 990700 295800 990712
rect 295852 990740 295858 990752
rect 397454 990740 397460 990752
rect 295852 990712 397460 990740
rect 295852 990700 295858 990712
rect 397454 990700 397460 990712
rect 397512 990700 397518 990752
rect 474734 990700 474740 990752
rect 474792 990740 474798 990752
rect 475470 990740 475476 990752
rect 474792 990712 475476 990740
rect 474792 990700 474798 990712
rect 475470 990700 475476 990712
rect 475528 990740 475534 990752
rect 526898 990740 526904 990752
rect 475528 990712 526904 990740
rect 475528 990700 475534 990712
rect 526898 990700 526904 990712
rect 526956 990740 526962 990752
rect 626534 990740 626540 990752
rect 526956 990712 626540 990740
rect 526956 990700 526962 990712
rect 626534 990700 626540 990712
rect 626592 990700 626598 990752
rect 89990 990632 89996 990684
rect 90048 990672 90054 990684
rect 141418 990672 141424 990684
rect 90048 990644 141424 990672
rect 90048 990632 90054 990644
rect 141418 990632 141424 990644
rect 141476 990672 141482 990684
rect 192846 990672 192852 990684
rect 141476 990644 192852 990672
rect 141476 990632 141482 990644
rect 192846 990632 192852 990644
rect 192904 990632 192910 990684
rect 233602 990632 233608 990684
rect 233660 990672 233666 990684
rect 245562 990672 245568 990684
rect 233660 990644 245568 990672
rect 233660 990632 233666 990644
rect 245562 990632 245568 990644
rect 245620 990632 245626 990684
rect 285306 990672 285312 990684
rect 275940 990644 285312 990672
rect 79502 990604 79508 990616
rect 45756 990576 79508 990604
rect 42242 990360 42248 990412
rect 42300 990400 42306 990412
rect 45756 990400 45784 990576
rect 79502 990564 79508 990576
rect 79560 990564 79566 990616
rect 130286 990564 130292 990616
rect 130344 990604 130350 990616
rect 181714 990604 181720 990616
rect 130344 990576 181720 990604
rect 130344 990564 130350 990576
rect 181714 990564 181720 990576
rect 181772 990564 181778 990616
rect 275940 990604 275968 990644
rect 285306 990632 285312 990644
rect 285364 990632 285370 990684
rect 387150 990672 387156 990684
rect 372540 990644 387156 990672
rect 314470 990604 314476 990616
rect 256712 990576 275968 990604
rect 295352 990576 314476 990604
rect 182358 990536 182364 990548
rect 179340 990508 182364 990536
rect 131114 990428 131120 990480
rect 131172 990468 131178 990480
rect 132494 990468 132500 990480
rect 131172 990440 132500 990468
rect 131172 990428 131178 990440
rect 132494 990428 132500 990440
rect 132552 990428 132558 990480
rect 160002 990468 160008 990480
rect 151832 990440 160008 990468
rect 151832 990400 151860 990440
rect 160002 990428 160008 990440
rect 160060 990428 160066 990480
rect 179340 990468 179368 990508
rect 182358 990496 182364 990508
rect 182416 990496 182422 990548
rect 192846 990496 192852 990548
rect 192904 990536 192910 990548
rect 244182 990536 244188 990548
rect 192904 990508 244188 990536
rect 192904 990496 192910 990508
rect 244182 990496 244188 990508
rect 244240 990496 244246 990548
rect 245562 990496 245568 990548
rect 245620 990536 245626 990548
rect 256712 990536 256740 990576
rect 245620 990508 256740 990536
rect 245620 990496 245626 990508
rect 285306 990496 285312 990548
rect 285364 990536 285370 990548
rect 295352 990536 295380 990576
rect 314470 990564 314476 990576
rect 314528 990564 314534 990616
rect 314746 990564 314752 990616
rect 314804 990604 314810 990616
rect 372540 990604 372568 990644
rect 387150 990632 387156 990644
rect 387208 990672 387214 990684
rect 476114 990672 476120 990684
rect 387208 990644 476120 990672
rect 387208 990632 387214 990644
rect 476114 990632 476120 990644
rect 476172 990672 476178 990684
rect 527542 990672 527548 990684
rect 476172 990644 527548 990672
rect 476172 990632 476178 990644
rect 527542 990632 527548 990644
rect 527600 990672 527606 990684
rect 629294 990672 629300 990684
rect 527600 990644 629300 990672
rect 527600 990632 527606 990644
rect 629294 990632 629300 990644
rect 629352 990672 629358 990684
rect 630950 990672 630956 990684
rect 629352 990644 630956 990672
rect 629352 990632 629358 990644
rect 630950 990632 630956 990644
rect 631008 990632 631014 990684
rect 314804 990576 328500 990604
rect 314804 990564 314810 990576
rect 328472 990548 328500 990576
rect 353312 990576 372568 990604
rect 285364 990508 295380 990536
rect 285364 990496 285370 990508
rect 328454 990496 328460 990548
rect 328512 990496 328518 990548
rect 347682 990496 347688 990548
rect 347740 990536 347746 990548
rect 353312 990536 353340 990576
rect 386506 990564 386512 990616
rect 386564 990604 386570 990616
rect 474734 990604 474740 990616
rect 386564 990576 474740 990604
rect 386564 990564 386570 990576
rect 474734 990564 474740 990576
rect 474792 990564 474798 990616
rect 347740 990508 353340 990536
rect 347740 990496 347746 990508
rect 397454 990496 397460 990548
rect 397512 990536 397518 990548
rect 486602 990536 486608 990548
rect 397512 990508 486608 990536
rect 397512 990496 397518 990508
rect 486602 990496 486608 990508
rect 486660 990496 486666 990548
rect 171060 990440 179368 990468
rect 42300 990372 45784 990400
rect 151740 990372 151860 990400
rect 42300 990360 42306 990372
rect 42702 990292 42708 990344
rect 42760 990332 42766 990344
rect 63402 990332 63408 990344
rect 42760 990304 63408 990332
rect 42760 990292 42766 990304
rect 63402 990292 63408 990304
rect 63460 990292 63466 990344
rect 140774 990292 140780 990344
rect 140832 990332 140838 990344
rect 151740 990332 151768 990372
rect 160094 990360 160100 990412
rect 160152 990400 160158 990412
rect 171060 990400 171088 990440
rect 181714 990428 181720 990480
rect 181772 990468 181778 990480
rect 194778 990468 194784 990480
rect 181772 990440 194784 990468
rect 181772 990428 181778 990440
rect 194778 990428 194784 990440
rect 194836 990428 194842 990480
rect 160152 990372 171088 990400
rect 160152 990360 160158 990372
rect 140832 990304 151768 990332
rect 140832 990292 140838 990304
rect 200022 990292 200028 990344
rect 200080 990332 200086 990344
rect 233602 990332 233608 990344
rect 200080 990304 233608 990332
rect 200080 990292 200086 990304
rect 233602 990292 233608 990304
rect 233660 990292 233666 990344
rect 275830 990292 275836 990344
rect 275888 990332 275894 990344
rect 289722 990332 289728 990344
rect 275888 990304 289728 990332
rect 275888 990292 275894 990304
rect 289722 990292 289728 990304
rect 289780 990292 289786 990344
rect 328362 990292 328368 990344
rect 328420 990332 328426 990344
rect 328420 990304 328500 990332
rect 328420 990292 328426 990304
rect 328472 990276 328500 990304
rect 42426 990224 42432 990276
rect 42484 990264 42490 990276
rect 42484 990236 45876 990264
rect 42484 990224 42490 990236
rect 45848 990196 45876 990236
rect 45922 990224 45928 990276
rect 45980 990264 45986 990276
rect 77294 990264 77300 990276
rect 45980 990236 77300 990264
rect 45980 990224 45986 990236
rect 77294 990224 77300 990236
rect 77352 990224 77358 990276
rect 121362 990264 121368 990276
rect 102060 990236 121368 990264
rect 78858 990196 78864 990208
rect 45848 990168 78864 990196
rect 78858 990156 78864 990168
rect 78916 990156 78922 990208
rect 82906 990156 82912 990208
rect 82964 990196 82970 990208
rect 102060 990196 102088 990236
rect 121362 990224 121368 990236
rect 121420 990224 121426 990276
rect 121454 990224 121460 990276
rect 121512 990264 121518 990276
rect 121512 990236 125548 990264
rect 121512 990224 121518 990236
rect 82964 990168 102088 990196
rect 125520 990196 125548 990236
rect 328454 990224 328460 990276
rect 328512 990224 328518 990276
rect 125520 990168 140728 990196
rect 82964 990156 82970 990168
rect 63402 990088 63408 990140
rect 63460 990128 63466 990140
rect 82630 990128 82636 990140
rect 63460 990100 82636 990128
rect 63460 990088 63466 990100
rect 82630 990088 82636 990100
rect 82688 990088 82694 990140
rect 140700 990128 140728 990168
rect 198734 990156 198740 990208
rect 198792 990196 198798 990208
rect 198792 990168 218008 990196
rect 198792 990156 198798 990168
rect 160002 990128 160008 990140
rect 140700 990100 160008 990128
rect 160002 990088 160008 990100
rect 160060 990088 160066 990140
rect 160094 990088 160100 990140
rect 160152 990128 160158 990140
rect 160152 990100 161428 990128
rect 160152 990088 160158 990100
rect 161400 990060 161428 990100
rect 179230 990088 179236 990140
rect 179288 990088 179294 990140
rect 179506 990088 179512 990140
rect 179564 990128 179570 990140
rect 198642 990128 198648 990140
rect 179564 990100 198648 990128
rect 179564 990088 179570 990100
rect 198642 990088 198648 990100
rect 198700 990088 198706 990140
rect 217980 990128 218008 990168
rect 231854 990156 231860 990208
rect 231912 990196 231918 990208
rect 256602 990196 256608 990208
rect 231912 990168 256608 990196
rect 231912 990156 231918 990168
rect 256602 990156 256608 990168
rect 256660 990156 256666 990208
rect 256786 990156 256792 990208
rect 256844 990196 256850 990208
rect 256844 990168 270448 990196
rect 256844 990156 256850 990168
rect 231762 990128 231768 990140
rect 217980 990100 231768 990128
rect 231762 990088 231768 990100
rect 231820 990088 231826 990140
rect 270420 990128 270448 990168
rect 295260 990168 314608 990196
rect 275830 990128 275836 990140
rect 270420 990100 275836 990128
rect 275830 990088 275836 990100
rect 275888 990088 275894 990140
rect 289722 990088 289728 990140
rect 289780 990128 289786 990140
rect 295260 990128 295288 990168
rect 289780 990100 295288 990128
rect 314580 990128 314608 990168
rect 639782 990156 639788 990208
rect 639840 990196 639846 990208
rect 673546 990196 673552 990208
rect 639840 990168 673552 990196
rect 639840 990156 639846 990168
rect 673546 990156 673552 990168
rect 673604 990156 673610 990208
rect 328178 990128 328184 990140
rect 314580 990100 328184 990128
rect 289780 990088 289786 990100
rect 328178 990088 328184 990100
rect 328236 990088 328242 990140
rect 626534 990088 626540 990140
rect 626592 990088 626598 990140
rect 628650 990088 628656 990140
rect 628708 990088 628714 990140
rect 630950 990088 630956 990140
rect 631008 990128 631014 990140
rect 673638 990128 673644 990140
rect 631008 990100 673644 990128
rect 631008 990088 631014 990100
rect 673638 990088 673644 990100
rect 673696 990088 673702 990140
rect 179248 990060 179276 990088
rect 161400 990032 179276 990060
rect 626552 990060 626580 990088
rect 628668 990060 628696 990088
rect 673454 990060 673460 990072
rect 626552 990032 673460 990060
rect 673454 990020 673460 990032
rect 673512 990020 673518 990072
rect 41782 969348 41788 969400
rect 41840 969388 41846 969400
rect 42334 969388 42340 969400
rect 41840 969360 42340 969388
rect 41840 969348 41846 969360
rect 42334 969348 42340 969360
rect 42392 969348 42398 969400
rect 41782 968464 41788 968516
rect 41840 968504 41846 968516
rect 42702 968504 42708 968516
rect 41840 968476 42708 968504
rect 41840 968464 41846 968476
rect 42702 968464 42708 968476
rect 42760 968464 42766 968516
rect 673454 965268 673460 965320
rect 673512 965308 673518 965320
rect 675386 965308 675392 965320
rect 673512 965280 675392 965308
rect 673512 965268 673518 965280
rect 675386 965268 675392 965280
rect 675444 965268 675450 965320
rect 673638 964724 673644 964776
rect 673696 964764 673702 964776
rect 675386 964764 675392 964776
rect 673696 964736 675392 964764
rect 673696 964724 673702 964736
rect 675386 964724 675392 964736
rect 675444 964724 675450 964776
rect 41782 962412 41788 962464
rect 41840 962452 41846 962464
rect 42334 962452 42340 962464
rect 41840 962424 42340 962452
rect 41840 962412 41846 962424
rect 42334 962412 42340 962424
rect 42392 962412 42398 962464
rect 41782 956428 41788 956480
rect 41840 956468 41846 956480
rect 42426 956468 42432 956480
rect 41840 956440 42432 956468
rect 41840 956428 41846 956440
rect 42426 956428 42432 956440
rect 42484 956428 42490 956480
rect 673546 953300 673552 953352
rect 673604 953340 673610 953352
rect 675386 953340 675392 953352
rect 673604 953312 675392 953340
rect 673604 953300 673610 953312
rect 675386 953300 675392 953312
rect 675444 953300 675450 953352
rect 42426 950784 42432 950836
rect 42484 950824 42490 950836
rect 42702 950824 42708 950836
rect 42484 950796 42708 950824
rect 42484 950784 42490 950796
rect 42702 950784 42708 950796
rect 42760 950784 42766 950836
rect 42426 946636 42432 946688
rect 42484 946676 42490 946688
rect 42610 946676 42616 946688
rect 42484 946648 42616 946676
rect 42484 946636 42490 946648
rect 42610 946636 42616 946648
rect 42668 946636 42674 946688
rect 44266 930112 44272 930164
rect 44324 930152 44330 930164
rect 45462 930152 45468 930164
rect 44324 930124 45468 930152
rect 44324 930112 44330 930124
rect 45462 930112 45468 930124
rect 45520 930112 45526 930164
rect 39666 922904 39672 922956
rect 39724 922944 39730 922956
rect 44266 922944 44272 922956
rect 39724 922916 44272 922944
rect 39724 922904 39730 922916
rect 44266 922904 44272 922916
rect 44324 922904 44330 922956
rect 39850 921748 39856 921800
rect 39908 921788 39914 921800
rect 42242 921788 42248 921800
rect 39908 921760 42248 921788
rect 39908 921748 39914 921760
rect 42242 921748 42248 921760
rect 42300 921748 42306 921800
rect 39850 916240 39856 916292
rect 39908 916280 39914 916292
rect 41414 916280 41420 916292
rect 39908 916252 41420 916280
rect 39908 916240 39914 916252
rect 41414 916240 41420 916252
rect 41472 916240 41478 916292
rect 42702 913588 42708 913640
rect 42760 913588 42766 913640
rect 42720 913492 42748 913588
rect 42794 913492 42800 913504
rect 42720 913464 42800 913492
rect 42794 913452 42800 913464
rect 42852 913452 42858 913504
rect 673638 910732 673644 910784
rect 673696 910772 673702 910784
rect 677778 910772 677784 910784
rect 673696 910744 677784 910772
rect 673696 910732 673702 910744
rect 677778 910732 677784 910744
rect 677836 910732 677842 910784
rect 42426 885912 42432 885964
rect 42484 885952 42490 885964
rect 42610 885952 42616 885964
rect 42484 885924 42616 885952
rect 42484 885912 42490 885924
rect 42610 885912 42616 885924
rect 42668 885912 42674 885964
rect 673454 876120 673460 876172
rect 673512 876160 673518 876172
rect 675386 876160 675392 876172
rect 673512 876132 675392 876160
rect 673512 876120 673518 876132
rect 675386 876120 675392 876132
rect 675444 876120 675450 876172
rect 41414 875576 41420 875628
rect 41472 875616 41478 875628
rect 42242 875616 42248 875628
rect 41472 875588 42248 875616
rect 41472 875576 41478 875588
rect 42242 875576 42248 875588
rect 42300 875576 42306 875628
rect 673638 875508 673644 875560
rect 673696 875548 673702 875560
rect 675386 875548 675392 875560
rect 673696 875520 675392 875548
rect 673696 875508 673702 875520
rect 675386 875508 675392 875520
rect 675444 875508 675450 875560
rect 675202 870136 675208 870188
rect 675260 870176 675266 870188
rect 675386 870176 675392 870188
rect 675260 870148 675392 870176
rect 675260 870136 675266 870148
rect 675386 870136 675392 870148
rect 675444 870136 675450 870188
rect 673546 864968 673552 865020
rect 673604 865008 673610 865020
rect 675386 865008 675392 865020
rect 673604 864980 675392 865008
rect 673604 864968 673610 864980
rect 675386 864968 675392 864980
rect 675444 864968 675450 865020
rect 674650 862792 674656 862844
rect 674708 862832 674714 862844
rect 675294 862832 675300 862844
rect 674708 862804 675300 862832
rect 674708 862792 674714 862804
rect 675294 862792 675300 862804
rect 675352 862792 675358 862844
rect 673914 850552 673920 850604
rect 673972 850592 673978 850604
rect 674650 850592 674656 850604
rect 673972 850564 674656 850592
rect 673972 850552 673978 850564
rect 674650 850552 674656 850564
rect 674708 850552 674714 850604
rect 42610 850008 42616 850060
rect 42668 850048 42674 850060
rect 42702 850048 42708 850060
rect 42668 850020 42708 850048
rect 42668 850008 42674 850020
rect 42702 850008 42708 850020
rect 42760 850008 42766 850060
rect 42610 830764 42616 830816
rect 42668 830804 42674 830816
rect 42794 830804 42800 830816
rect 42668 830776 42800 830804
rect 42668 830764 42674 830776
rect 42794 830764 42800 830776
rect 42852 830764 42858 830816
rect 673730 830764 673736 830816
rect 673788 830804 673794 830816
rect 674006 830804 674012 830816
rect 673788 830776 674012 830804
rect 673788 830764 673794 830776
rect 674006 830764 674012 830776
rect 674064 830764 674070 830816
rect 673822 816960 673828 817012
rect 673880 817000 673886 817012
rect 674006 817000 674012 817012
rect 673880 816972 674012 817000
rect 673880 816960 673886 816972
rect 674006 816960 674012 816972
rect 674064 816960 674070 817012
rect 672810 811384 672816 811436
rect 672868 811424 672874 811436
rect 673086 811424 673092 811436
rect 672868 811396 673092 811424
rect 672868 811384 672874 811396
rect 673086 811384 673092 811396
rect 673144 811384 673150 811436
rect 42518 807440 42524 807492
rect 42576 807440 42582 807492
rect 42536 807288 42564 807440
rect 42518 807236 42524 807288
rect 42576 807236 42582 807288
rect 42242 806352 42248 806404
rect 42300 806392 42306 806404
rect 42610 806392 42616 806404
rect 42300 806364 42616 806392
rect 42300 806352 42306 806364
rect 42610 806352 42616 806364
rect 42668 806352 42674 806404
rect 42334 804244 42340 804296
rect 42392 804284 42398 804296
rect 42794 804284 42800 804296
rect 42392 804256 42800 804284
rect 42392 804244 42398 804256
rect 42794 804244 42800 804256
rect 42852 804244 42858 804296
rect 41782 798124 41788 798176
rect 41840 798164 41846 798176
rect 42334 798164 42340 798176
rect 41840 798136 42340 798164
rect 41840 798124 41846 798136
rect 42334 798124 42340 798136
rect 42392 798124 42398 798176
rect 674006 797580 674012 797632
rect 674064 797620 674070 797632
rect 675294 797620 675300 797632
rect 674064 797592 675300 797620
rect 674064 797580 674070 797592
rect 675294 797580 675300 797592
rect 675352 797580 675358 797632
rect 41782 787856 41788 787908
rect 41840 787896 41846 787908
rect 42242 787896 42248 787908
rect 41840 787868 42248 787896
rect 41840 787856 41846 787868
rect 42242 787856 42248 787868
rect 42300 787896 42306 787908
rect 42610 787896 42616 787908
rect 42300 787868 42616 787896
rect 42300 787856 42306 787868
rect 42610 787856 42616 787868
rect 42668 787856 42674 787908
rect 41782 787584 41788 787636
rect 41840 787624 41846 787636
rect 42518 787624 42524 787636
rect 41840 787596 42524 787624
rect 41840 787584 41846 787596
rect 42518 787584 42524 787596
rect 42576 787584 42582 787636
rect 673454 785272 673460 785324
rect 673512 785312 673518 785324
rect 675386 785312 675392 785324
rect 673512 785284 675392 785312
rect 673512 785272 673518 785284
rect 675386 785272 675392 785284
rect 675444 785272 675450 785324
rect 672994 778336 673000 778388
rect 673052 778336 673058 778388
rect 673012 778308 673040 778336
rect 673178 778308 673184 778320
rect 673012 778280 673184 778308
rect 673178 778268 673184 778280
rect 673236 778268 673242 778320
rect 673546 774868 673552 774920
rect 673604 774908 673610 774920
rect 675386 774908 675392 774920
rect 673604 774880 675392 774908
rect 673604 774868 673610 774880
rect 675386 774868 675392 774880
rect 675444 774868 675450 774920
rect 673086 772760 673092 772812
rect 673144 772800 673150 772812
rect 673178 772800 673184 772812
rect 673144 772772 673184 772800
rect 673144 772760 673150 772772
rect 673178 772760 673184 772772
rect 673236 772760 673242 772812
rect 41782 754468 41788 754520
rect 41840 754508 41846 754520
rect 42426 754508 42432 754520
rect 41840 754480 42432 754508
rect 41840 754468 41846 754480
rect 42426 754468 42432 754480
rect 42484 754468 42490 754520
rect 41782 744404 41788 744456
rect 41840 744444 41846 744456
rect 42426 744444 42432 744456
rect 41840 744416 42432 744444
rect 41840 744404 41846 744416
rect 42426 744404 42432 744416
rect 42484 744444 42490 744456
rect 42610 744444 42616 744456
rect 42484 744416 42616 744444
rect 42484 744404 42490 744416
rect 42610 744404 42616 744416
rect 42668 744404 42674 744456
rect 673822 741888 673828 741940
rect 673880 741928 673886 741940
rect 675386 741928 675392 741940
rect 673880 741900 675392 741928
rect 673880 741888 673886 741900
rect 675386 741888 675392 741900
rect 675444 741888 675450 741940
rect 673454 741344 673460 741396
rect 673512 741384 673518 741396
rect 675386 741384 675392 741396
rect 673512 741356 675392 741384
rect 673512 741344 673518 741356
rect 675386 741344 675392 741356
rect 675444 741344 675450 741396
rect 673178 739752 673184 739764
rect 673104 739724 673184 739752
rect 673104 739560 673132 739724
rect 673178 739712 673184 739724
rect 673236 739712 673242 739764
rect 673086 739508 673092 739560
rect 673144 739508 673150 739560
rect 673454 736584 673460 736636
rect 673512 736624 673518 736636
rect 675294 736624 675300 736636
rect 673512 736596 675300 736624
rect 673512 736584 673518 736596
rect 675294 736584 675300 736596
rect 675352 736584 675358 736636
rect 42242 730804 42248 730856
rect 42300 730844 42306 730856
rect 42610 730844 42616 730856
rect 42300 730816 42616 730844
rect 42300 730804 42306 730816
rect 42610 730804 42616 730816
rect 42668 730804 42674 730856
rect 673546 730124 673552 730176
rect 673604 730164 673610 730176
rect 673914 730164 673920 730176
rect 673604 730136 673920 730164
rect 673604 730124 673610 730136
rect 673914 730124 673920 730136
rect 673972 730164 673978 730176
rect 675386 730164 675392 730176
rect 673972 730136 675392 730164
rect 673972 730124 673978 730136
rect 675386 730124 675392 730136
rect 675444 730124 675450 730176
rect 673730 720332 673736 720384
rect 673788 720372 673794 720384
rect 673914 720372 673920 720384
rect 673788 720344 673920 720372
rect 673788 720332 673794 720344
rect 673914 720332 673920 720344
rect 673972 720332 673978 720384
rect 672810 712036 672816 712088
rect 672868 712076 672874 712088
rect 672994 712076 673000 712088
rect 672868 712048 673000 712076
rect 672868 712036 672874 712048
rect 672994 712036 673000 712048
rect 673052 712036 673058 712088
rect 41782 711288 41788 711340
rect 41840 711288 41846 711340
rect 41800 711260 41828 711288
rect 42702 711260 42708 711272
rect 41800 711232 42708 711260
rect 42702 711220 42708 711232
rect 42760 711220 42766 711272
rect 673454 710676 673460 710728
rect 673512 710716 673518 710728
rect 675294 710716 675300 710728
rect 673512 710688 675300 710716
rect 673512 710676 673518 710688
rect 675294 710676 675300 710688
rect 675352 710676 675358 710728
rect 42334 708704 42340 708756
rect 42392 708744 42398 708756
rect 42610 708744 42616 708756
rect 42392 708716 42616 708744
rect 42392 708704 42398 708716
rect 42610 708704 42616 708716
rect 42668 708704 42674 708756
rect 673822 701128 673828 701140
rect 673656 701100 673828 701128
rect 673656 701072 673684 701100
rect 673822 701088 673828 701100
rect 673880 701088 673886 701140
rect 673638 701020 673644 701072
rect 673696 701020 673702 701072
rect 41782 700952 41788 701004
rect 41840 700992 41846 701004
rect 42334 700992 42340 701004
rect 41840 700964 42340 700992
rect 41840 700952 41846 700964
rect 42334 700952 42340 700964
rect 42392 700992 42398 701004
rect 42518 700992 42524 701004
rect 42392 700964 42524 700992
rect 42392 700952 42398 700964
rect 42518 700952 42524 700964
rect 42576 700952 42582 701004
rect 673638 695920 673644 695972
rect 673696 695960 673702 695972
rect 673822 695960 673828 695972
rect 673696 695932 673828 695960
rect 673696 695920 673702 695932
rect 673822 695920 673828 695932
rect 673880 695960 673886 695972
rect 675386 695960 675392 695972
rect 673880 695932 675392 695960
rect 673880 695920 673886 695932
rect 675386 695920 675392 695932
rect 675444 695920 675450 695972
rect 42702 695444 42708 695496
rect 42760 695484 42766 695496
rect 42978 695484 42984 695496
rect 42760 695456 42984 695484
rect 42760 695444 42766 695456
rect 42978 695444 42984 695456
rect 43036 695444 43042 695496
rect 672810 692792 672816 692844
rect 672868 692832 672874 692844
rect 673178 692832 673184 692844
rect 672868 692804 673184 692832
rect 672868 692792 672874 692804
rect 673178 692792 673184 692804
rect 673236 692792 673242 692844
rect 673454 681708 673460 681760
rect 673512 681748 673518 681760
rect 675202 681748 675208 681760
rect 673512 681720 675208 681748
rect 673512 681708 673518 681720
rect 675202 681708 675208 681720
rect 675260 681708 675266 681760
rect 42794 676200 42800 676252
rect 42852 676240 42858 676252
rect 42978 676240 42984 676252
rect 42852 676212 42984 676240
rect 42852 676200 42858 676212
rect 42978 676200 42984 676212
rect 43036 676200 43042 676252
rect 672994 676132 673000 676184
rect 673052 676172 673058 676184
rect 673086 676172 673092 676184
rect 673052 676144 673092 676172
rect 673052 676132 673058 676144
rect 673086 676132 673092 676144
rect 673144 676132 673150 676184
rect 673638 676132 673644 676184
rect 673696 676172 673702 676184
rect 673914 676172 673920 676184
rect 673696 676144 673920 676172
rect 673696 676132 673702 676144
rect 673914 676132 673920 676144
rect 673972 676132 673978 676184
rect 42334 672256 42340 672308
rect 42392 672296 42398 672308
rect 42518 672296 42524 672308
rect 42392 672268 42524 672296
rect 42392 672256 42398 672268
rect 42518 672256 42524 672268
rect 42576 672256 42582 672308
rect 41782 669060 41788 669112
rect 41840 669100 41846 669112
rect 42426 669100 42432 669112
rect 41840 669072 42432 669100
rect 41840 669060 41846 669072
rect 42426 669060 42432 669072
rect 42484 669100 42490 669112
rect 42794 669100 42800 669112
rect 42484 669072 42800 669100
rect 42484 669060 42490 669072
rect 42794 669060 42800 669072
rect 42852 669060 42858 669112
rect 41782 657636 41788 657688
rect 41840 657676 41846 657688
rect 42334 657676 42340 657688
rect 41840 657648 42340 657676
rect 41840 657636 41846 657648
rect 42334 657636 42340 657648
rect 42392 657676 42398 657688
rect 42610 657676 42616 657688
rect 42392 657648 42616 657676
rect 42392 657636 42398 657648
rect 42610 657636 42616 657648
rect 42668 657636 42674 657688
rect 42242 657092 42248 657144
rect 42300 657132 42306 657144
rect 42702 657132 42708 657144
rect 42300 657104 42708 657132
rect 42300 657092 42306 657104
rect 42702 657092 42708 657104
rect 42760 657092 42766 657144
rect 673086 656888 673092 656940
rect 673144 656928 673150 656940
rect 673178 656928 673184 656940
rect 673144 656900 673184 656928
rect 673144 656888 673150 656900
rect 673178 656888 673184 656900
rect 673236 656888 673242 656940
rect 673546 656888 673552 656940
rect 673604 656928 673610 656940
rect 673914 656928 673920 656940
rect 673604 656900 673920 656928
rect 673604 656888 673610 656900
rect 673914 656888 673920 656900
rect 673972 656888 673978 656940
rect 673454 651720 673460 651772
rect 673512 651760 673518 651772
rect 673822 651760 673828 651772
rect 673512 651732 673828 651760
rect 673512 651720 673518 651732
rect 673822 651720 673828 651732
rect 673880 651760 673886 651772
rect 675386 651760 675392 651772
rect 673880 651732 675392 651760
rect 673880 651720 673886 651732
rect 675386 651720 675392 651732
rect 675444 651720 675450 651772
rect 673546 651108 673552 651160
rect 673604 651148 673610 651160
rect 673822 651148 673828 651160
rect 673604 651120 673828 651148
rect 673604 651108 673610 651120
rect 673822 651108 673828 651120
rect 673880 651148 673886 651160
rect 675386 651148 675392 651160
rect 673880 651120 675392 651148
rect 673880 651108 673886 651120
rect 675386 651108 675392 651120
rect 675444 651108 675450 651160
rect 673546 639684 673552 639736
rect 673604 639724 673610 639736
rect 673730 639724 673736 639736
rect 673604 639696 673736 639724
rect 673604 639684 673610 639696
rect 673730 639684 673736 639696
rect 673788 639724 673794 639736
rect 675386 639724 675392 639736
rect 673788 639696 675392 639724
rect 673788 639684 673794 639696
rect 675386 639684 675392 639696
rect 675444 639684 675450 639736
rect 672810 637508 672816 637560
rect 672868 637548 672874 637560
rect 673086 637548 673092 637560
rect 672868 637520 673092 637548
rect 672868 637508 672874 637520
rect 673086 637508 673092 637520
rect 673144 637508 673150 637560
rect 673730 637508 673736 637560
rect 673788 637548 673794 637560
rect 674006 637548 674012 637560
rect 673788 637520 674012 637548
rect 673788 637508 673794 637520
rect 674006 637508 674012 637520
rect 674064 637508 674070 637560
rect 41782 625880 41788 625932
rect 41840 625920 41846 625932
rect 42518 625920 42524 625932
rect 41840 625892 42524 625920
rect 41840 625880 41846 625892
rect 42518 625880 42524 625892
rect 42576 625880 42582 625932
rect 42242 618468 42248 618520
rect 42300 618508 42306 618520
rect 42794 618508 42800 618520
rect 42300 618480 42800 618508
rect 42300 618468 42306 618480
rect 42794 618468 42800 618480
rect 42852 618468 42858 618520
rect 672810 618264 672816 618316
rect 672868 618304 672874 618316
rect 672994 618304 673000 618316
rect 672868 618276 673000 618304
rect 672868 618264 672874 618276
rect 672994 618264 673000 618276
rect 673052 618264 673058 618316
rect 673730 618264 673736 618316
rect 673788 618304 673794 618316
rect 673914 618304 673920 618316
rect 673788 618276 673920 618304
rect 673788 618264 673794 618276
rect 673914 618264 673920 618276
rect 673972 618264 673978 618316
rect 41782 614116 41788 614168
rect 41840 614156 41846 614168
rect 42334 614156 42340 614168
rect 41840 614128 42340 614156
rect 41840 614116 41846 614128
rect 42334 614116 42340 614128
rect 42392 614116 42398 614168
rect 673454 606704 673460 606756
rect 673512 606744 673518 606756
rect 673822 606744 673828 606756
rect 673512 606716 673828 606744
rect 673512 606704 673518 606716
rect 673822 606704 673828 606716
rect 673880 606744 673886 606756
rect 675386 606744 675392 606756
rect 673880 606716 675392 606744
rect 673880 606704 673886 606716
rect 675386 606704 675392 606716
rect 675444 606704 675450 606756
rect 672810 605820 672816 605872
rect 672868 605860 672874 605872
rect 672994 605860 673000 605872
rect 672868 605832 673000 605860
rect 672868 605820 672874 605832
rect 672994 605820 673000 605832
rect 673052 605820 673058 605872
rect 673914 605616 673920 605668
rect 673972 605656 673978 605668
rect 675294 605656 675300 605668
rect 673972 605628 675300 605656
rect 673972 605616 673978 605628
rect 675294 605616 675300 605628
rect 675352 605616 675358 605668
rect 673638 604460 673644 604512
rect 673696 604500 673702 604512
rect 673914 604500 673920 604512
rect 673696 604472 673920 604500
rect 673696 604460 673702 604472
rect 673914 604460 673920 604472
rect 673972 604460 673978 604512
rect 42610 604392 42616 604444
rect 42668 604392 42674 604444
rect 42628 604364 42656 604392
rect 42702 604364 42708 604376
rect 42628 604336 42708 604364
rect 42702 604324 42708 604336
rect 42760 604324 42766 604376
rect 672810 596164 672816 596216
rect 672868 596204 672874 596216
rect 672994 596204 673000 596216
rect 672868 596176 673000 596204
rect 672868 596164 672874 596176
rect 672994 596164 673000 596176
rect 673052 596164 673058 596216
rect 672810 596028 672816 596080
rect 672868 596068 672874 596080
rect 672994 596068 673000 596080
rect 672868 596040 673000 596068
rect 672868 596028 672874 596040
rect 672994 596028 673000 596040
rect 673052 596028 673058 596080
rect 673546 594872 673552 594924
rect 673604 594912 673610 594924
rect 675386 594912 675392 594924
rect 673604 594884 675392 594912
rect 673604 594872 673610 594884
rect 675386 594872 675392 594884
rect 675444 594872 675450 594924
rect 672810 585080 672816 585132
rect 672868 585120 672874 585132
rect 672994 585120 673000 585132
rect 672868 585092 673000 585120
rect 672868 585080 672874 585092
rect 672994 585080 673000 585092
rect 673052 585080 673058 585132
rect 41782 581680 41788 581732
rect 41840 581720 41846 581732
rect 42702 581720 42708 581732
rect 41840 581692 42708 581720
rect 41840 581680 41846 581692
rect 42702 581680 42708 581692
rect 42760 581680 42766 581732
rect 41782 571616 41788 571668
rect 41840 571656 41846 571668
rect 42518 571656 42524 571668
rect 41840 571628 42524 571656
rect 41840 571616 41846 571628
rect 42518 571616 42524 571628
rect 42576 571616 42582 571668
rect 673822 561484 673828 561536
rect 673880 561524 673886 561536
rect 675386 561524 675392 561536
rect 673880 561496 675392 561524
rect 673880 561484 673886 561496
rect 675386 561484 675392 561496
rect 675444 561484 675450 561536
rect 673454 559920 673460 559972
rect 673512 559960 673518 559972
rect 673638 559960 673644 559972
rect 673512 559932 673644 559960
rect 673512 559920 673518 559932
rect 673638 559920 673644 559932
rect 673696 559960 673702 559972
rect 675386 559960 675392 559972
rect 673696 559932 675392 559960
rect 673696 559920 673702 559932
rect 675386 559920 675392 559932
rect 675444 559920 675450 559972
rect 673546 550468 673552 550520
rect 673604 550508 673610 550520
rect 675386 550508 675392 550520
rect 673604 550480 675392 550508
rect 673604 550468 673610 550480
rect 675386 550468 675392 550480
rect 675444 550468 675450 550520
rect 42426 546456 42432 546508
rect 42484 546496 42490 546508
rect 42610 546496 42616 546508
rect 42484 546468 42616 546496
rect 42484 546456 42490 546468
rect 42610 546456 42616 546468
rect 42668 546456 42674 546508
rect 41782 538500 41788 538552
rect 41840 538540 41846 538552
rect 42426 538540 42432 538552
rect 41840 538512 42432 538540
rect 41840 538500 41846 538512
rect 42426 538500 42432 538512
rect 42484 538500 42490 538552
rect 672902 538228 672908 538280
rect 672960 538268 672966 538280
rect 673086 538268 673092 538280
rect 672960 538240 673092 538268
rect 672960 538228 672966 538240
rect 673086 538228 673092 538240
rect 673144 538228 673150 538280
rect 41782 527756 41788 527808
rect 41840 527796 41846 527808
rect 42518 527796 42524 527808
rect 41840 527768 42524 527796
rect 41840 527756 41846 527768
rect 42518 527756 42524 527768
rect 42576 527756 42582 527808
rect 672902 527008 672908 527060
rect 672960 527048 672966 527060
rect 673178 527048 673184 527060
rect 672960 527020 673184 527048
rect 672960 527008 672966 527020
rect 673178 527008 673184 527020
rect 673236 527008 673242 527060
rect 672994 499536 673000 499588
rect 673052 499576 673058 499588
rect 673270 499576 673276 499588
rect 673052 499548 673276 499576
rect 673052 499536 673058 499548
rect 673270 499536 673276 499548
rect 673328 499536 673334 499588
rect 672994 482944 673000 482996
rect 673052 482984 673058 482996
rect 673270 482984 673276 482996
rect 673052 482956 673276 482984
rect 673052 482944 673058 482956
rect 673270 482944 673276 482956
rect 673328 482944 673334 482996
rect 673454 463632 673460 463684
rect 673512 463672 673518 463684
rect 677686 463672 677692 463684
rect 673512 463644 677692 463672
rect 673512 463632 673518 463644
rect 677686 463632 677692 463644
rect 677744 463632 677750 463684
rect 39390 458192 39396 458244
rect 39448 458232 39454 458244
rect 44266 458232 44272 458244
rect 39448 458204 44272 458232
rect 39448 458192 39454 458204
rect 44266 458192 44272 458204
rect 44324 458192 44330 458244
rect 39850 448264 39856 448316
rect 39908 448304 39914 448316
rect 42242 448304 42248 448316
rect 39908 448276 42248 448304
rect 39908 448264 39914 448276
rect 42242 448264 42248 448276
rect 42300 448264 42306 448316
rect 676214 440172 676220 440224
rect 676272 440212 676278 440224
rect 677686 440212 677692 440224
rect 676272 440184 677692 440212
rect 676272 440172 676278 440184
rect 677686 440172 677692 440184
rect 677744 440172 677750 440224
rect 42242 413380 42248 413432
rect 42300 413420 42306 413432
rect 42610 413420 42616 413432
rect 42300 413392 42616 413420
rect 42300 413380 42306 413392
rect 42610 413380 42616 413392
rect 42668 413380 42674 413432
rect 672810 412496 672816 412548
rect 672868 412536 672874 412548
rect 676214 412536 676220 412548
rect 672868 412508 676220 412536
rect 672868 412496 672874 412508
rect 676214 412496 676220 412508
rect 676272 412496 676278 412548
rect 41782 410932 41788 410984
rect 41840 410972 41846 410984
rect 42426 410972 42432 410984
rect 41840 410944 42432 410972
rect 41840 410932 41846 410944
rect 42426 410932 42432 410944
rect 42484 410932 42490 410984
rect 42242 405356 42248 405408
rect 42300 405396 42306 405408
rect 42518 405396 42524 405408
rect 42300 405368 42524 405396
rect 42300 405356 42306 405368
rect 42518 405356 42524 405368
rect 42576 405356 42582 405408
rect 41782 400800 41788 400852
rect 41840 400840 41846 400852
rect 42610 400840 42616 400852
rect 41840 400812 42616 400840
rect 41840 400800 41846 400812
rect 42610 400800 42616 400812
rect 42668 400800 42674 400852
rect 42242 400120 42248 400172
rect 42300 400160 42306 400172
rect 42518 400160 42524 400172
rect 42300 400132 42524 400160
rect 42300 400120 42306 400132
rect 42518 400120 42524 400132
rect 42576 400120 42582 400172
rect 672718 386316 672724 386368
rect 672776 386356 672782 386368
rect 672902 386356 672908 386368
rect 672776 386328 672908 386356
rect 672776 386316 672782 386328
rect 672902 386316 672908 386328
rect 672960 386316 672966 386368
rect 673546 384004 673552 384056
rect 673604 384044 673610 384056
rect 675386 384044 675392 384056
rect 673604 384016 675392 384044
rect 673604 384004 673610 384016
rect 675386 384004 675392 384016
rect 675444 384004 675450 384056
rect 673454 382576 673460 382628
rect 673512 382616 673518 382628
rect 673638 382616 673644 382628
rect 673512 382588 673644 382616
rect 673512 382576 673518 382588
rect 673638 382576 673644 382588
rect 673696 382616 673702 382628
rect 675294 382616 675300 382628
rect 673696 382588 675300 382616
rect 673696 382576 673702 382588
rect 675294 382576 675300 382588
rect 675352 382576 675358 382628
rect 673914 372308 673920 372360
rect 673972 372348 673978 372360
rect 675386 372348 675392 372360
rect 673972 372320 675392 372348
rect 673972 372308 673978 372320
rect 675386 372308 675392 372320
rect 675444 372308 675450 372360
rect 41782 368636 41788 368688
rect 41840 368676 41846 368688
rect 42426 368676 42432 368688
rect 41840 368648 42432 368676
rect 41840 368636 41846 368648
rect 42426 368636 42432 368648
rect 42484 368636 42490 368688
rect 42242 357620 42248 357672
rect 42300 357660 42306 357672
rect 42610 357660 42616 357672
rect 42300 357632 42616 357660
rect 42300 357620 42306 357632
rect 42610 357620 42616 357632
rect 42668 357620 42674 357672
rect 41782 356668 41788 356720
rect 41840 356708 41846 356720
rect 42518 356708 42524 356720
rect 41840 356680 42524 356708
rect 41840 356668 41846 356680
rect 42518 356668 42524 356680
rect 42576 356668 42582 356720
rect 672718 353336 672724 353388
rect 672776 353336 672782 353388
rect 672736 353252 672764 353336
rect 672718 353200 672724 353252
rect 672776 353200 672782 353252
rect 672718 347692 672724 347744
rect 672776 347732 672782 347744
rect 672902 347732 672908 347744
rect 672776 347704 672908 347732
rect 672776 347692 672782 347704
rect 672902 347692 672908 347704
rect 672960 347692 672966 347744
rect 42242 342184 42248 342236
rect 42300 342224 42306 342236
rect 42610 342224 42616 342236
rect 42300 342196 42616 342224
rect 42300 342184 42306 342196
rect 42610 342184 42616 342196
rect 42668 342184 42674 342236
rect 673454 338512 673460 338564
rect 673512 338552 673518 338564
rect 673638 338552 673644 338564
rect 673512 338524 673644 338552
rect 673512 338512 673518 338524
rect 673638 338512 673644 338524
rect 673696 338552 673702 338564
rect 675386 338552 675392 338564
rect 673696 338524 675392 338552
rect 673696 338512 673702 338524
rect 675386 338512 675392 338524
rect 675444 338512 675450 338564
rect 672534 328448 672540 328500
rect 672592 328488 672598 328500
rect 672902 328488 672908 328500
rect 672592 328460 672908 328488
rect 672592 328448 672598 328460
rect 672902 328448 672908 328460
rect 672960 328448 672966 328500
rect 42610 328380 42616 328432
rect 42668 328420 42674 328432
rect 42886 328420 42892 328432
rect 42668 328392 42892 328420
rect 42668 328380 42674 328392
rect 42886 328380 42892 328392
rect 42944 328380 42950 328432
rect 673822 327088 673828 327140
rect 673880 327128 673886 327140
rect 675386 327128 675392 327140
rect 673880 327100 675392 327128
rect 673880 327088 673886 327100
rect 675386 327088 675392 327100
rect 675444 327088 675450 327140
rect 41782 324504 41788 324556
rect 41840 324544 41846 324556
rect 42426 324544 42432 324556
rect 41840 324516 42432 324544
rect 41840 324504 41846 324516
rect 42426 324504 42432 324516
rect 42484 324544 42490 324556
rect 42702 324544 42708 324556
rect 42484 324516 42708 324544
rect 42484 324504 42490 324516
rect 42702 324504 42708 324516
rect 42760 324504 42766 324556
rect 672534 316004 672540 316056
rect 672592 316044 672598 316056
rect 672718 316044 672724 316056
rect 672592 316016 672724 316044
rect 672592 316004 672598 316016
rect 672718 316004 672724 316016
rect 672776 316004 672782 316056
rect 42886 315120 42892 315172
rect 42944 315120 42950 315172
rect 41782 315052 41788 315104
rect 41840 315092 41846 315104
rect 42904 315092 42932 315120
rect 41840 315064 42932 315092
rect 41840 315052 41846 315064
rect 41782 314440 41788 314492
rect 41840 314480 41846 314492
rect 42334 314480 42340 314492
rect 41840 314452 42340 314480
rect 41840 314440 41846 314452
rect 42334 314440 42340 314452
rect 42392 314480 42398 314492
rect 42518 314480 42524 314492
rect 42392 314452 42524 314480
rect 42392 314440 42398 314452
rect 42518 314440 42524 314452
rect 42576 314440 42582 314492
rect 42426 313556 42432 313608
rect 42484 313596 42490 313608
rect 42702 313596 42708 313608
rect 42484 313568 42708 313596
rect 42484 313556 42490 313568
rect 42702 313556 42708 313568
rect 42760 313556 42766 313608
rect 42702 309068 42708 309120
rect 42760 309108 42766 309120
rect 42886 309108 42892 309120
rect 42760 309080 42892 309108
rect 42760 309068 42766 309080
rect 42886 309068 42892 309080
rect 42944 309068 42950 309120
rect 672442 306348 672448 306400
rect 672500 306388 672506 306400
rect 672718 306388 672724 306400
rect 672500 306360 672724 306388
rect 672500 306348 672506 306360
rect 672718 306348 672724 306360
rect 672776 306348 672782 306400
rect 673546 293564 673552 293616
rect 673604 293604 673610 293616
rect 675386 293604 675392 293616
rect 673604 293576 675392 293604
rect 673604 293564 673610 293576
rect 675386 293564 675392 293576
rect 675444 293564 675450 293616
rect 42702 289824 42708 289876
rect 42760 289864 42766 289876
rect 42978 289864 42984 289876
rect 42760 289836 42984 289864
rect 42760 289824 42766 289836
rect 42978 289824 42984 289836
rect 43036 289824 43042 289876
rect 673638 283024 673644 283076
rect 673696 283064 673702 283076
rect 675386 283064 675392 283076
rect 673696 283036 675392 283064
rect 673696 283024 673702 283036
rect 675386 283024 675392 283036
rect 675444 283024 675450 283076
rect 41782 282276 41788 282328
rect 41840 282316 41846 282328
rect 42426 282316 42432 282328
rect 41840 282288 42432 282316
rect 41840 282276 41846 282288
rect 42426 282276 42432 282288
rect 42484 282276 42490 282328
rect 42610 277176 42616 277228
rect 42668 277216 42674 277228
rect 42978 277216 42984 277228
rect 42668 277188 42984 277216
rect 42668 277176 42674 277188
rect 42978 277176 42984 277188
rect 43036 277176 43042 277228
rect 672626 276060 672632 276072
rect 672552 276032 672632 276060
rect 672552 276004 672580 276032
rect 672626 276020 672632 276032
rect 672684 276020 672690 276072
rect 672534 275952 672540 276004
rect 672592 275952 672598 276004
rect 41782 271464 41788 271516
rect 41840 271504 41846 271516
rect 42610 271504 42616 271516
rect 41840 271476 42616 271504
rect 41840 271464 41846 271476
rect 42610 271464 42616 271476
rect 42668 271464 42674 271516
rect 42610 270512 42616 270564
rect 42668 270552 42674 270564
rect 42702 270552 42708 270564
rect 42668 270524 42708 270552
rect 42668 270512 42674 270524
rect 42702 270512 42708 270524
rect 42760 270512 42766 270564
rect 672534 260788 672540 260840
rect 672592 260828 672598 260840
rect 672902 260828 672908 260840
rect 672592 260800 672908 260828
rect 672592 260788 672598 260800
rect 672902 260788 672908 260800
rect 672960 260788 672966 260840
rect 673638 256640 673644 256692
rect 673696 256680 673702 256692
rect 674006 256680 674012 256692
rect 673696 256652 674012 256680
rect 673696 256640 673702 256652
rect 674006 256640 674012 256652
rect 674064 256640 674070 256692
rect 672718 251200 672724 251252
rect 672776 251240 672782 251252
rect 672902 251240 672908 251252
rect 672776 251212 672908 251240
rect 672776 251200 672782 251212
rect 672902 251200 672908 251212
rect 672960 251200 672966 251252
rect 672534 251064 672540 251116
rect 672592 251104 672598 251116
rect 672718 251104 672724 251116
rect 672592 251076 672724 251104
rect 672592 251064 672598 251076
rect 672718 251064 672724 251076
rect 672776 251064 672782 251116
rect 673546 248140 673552 248192
rect 673604 248180 673610 248192
rect 675386 248180 675392 248192
rect 673604 248152 675392 248180
rect 673604 248140 673610 248152
rect 675386 248140 675392 248152
rect 675444 248140 675450 248192
rect 673454 247460 673460 247512
rect 673512 247500 673518 247512
rect 673730 247500 673736 247512
rect 673512 247472 673736 247500
rect 673512 247460 673518 247472
rect 673730 247460 673736 247472
rect 673788 247500 673794 247512
rect 675386 247500 675392 247512
rect 673788 247472 675392 247500
rect 673788 247460 673794 247472
rect 675386 247460 675392 247472
rect 675444 247460 675450 247512
rect 42150 245624 42156 245676
rect 42208 245664 42214 245676
rect 42334 245664 42340 245676
rect 42208 245636 42340 245664
rect 42208 245624 42214 245636
rect 42334 245624 42340 245636
rect 42392 245624 42398 245676
rect 42150 240592 42156 240644
rect 42208 240632 42214 240644
rect 42702 240632 42708 240644
rect 42208 240604 42708 240632
rect 42208 240592 42214 240604
rect 42702 240592 42708 240604
rect 42760 240592 42766 240644
rect 41782 238076 41788 238128
rect 41840 238116 41846 238128
rect 42426 238116 42432 238128
rect 41840 238088 42432 238116
rect 41840 238076 41846 238088
rect 42426 238076 42432 238088
rect 42484 238116 42490 238128
rect 42610 238116 42616 238128
rect 42484 238088 42616 238116
rect 42484 238076 42490 238088
rect 42610 238076 42616 238088
rect 42668 238076 42674 238128
rect 674006 237736 674012 237788
rect 674064 237776 674070 237788
rect 675386 237776 675392 237788
rect 674064 237748 675392 237776
rect 674064 237736 674070 237748
rect 675386 237736 675392 237748
rect 675444 237736 675450 237788
rect 673822 231820 673828 231872
rect 673880 231860 673886 231872
rect 674006 231860 674012 231872
rect 673880 231832 674012 231860
rect 673880 231820 673886 231832
rect 674006 231820 674012 231832
rect 674064 231820 674070 231872
rect 41782 228624 41788 228676
rect 41840 228664 41846 228676
rect 42426 228664 42432 228676
rect 41840 228636 42432 228664
rect 41840 228624 41846 228636
rect 42426 228624 42432 228636
rect 42484 228664 42490 228676
rect 42886 228664 42892 228676
rect 42484 228636 42892 228664
rect 42484 228624 42490 228636
rect 42886 228624 42892 228636
rect 42944 228624 42950 228676
rect 41782 228012 41788 228064
rect 41840 228052 41846 228064
rect 42242 228052 42248 228064
rect 41840 228024 42248 228052
rect 41840 228012 41846 228024
rect 42242 228012 42248 228024
rect 42300 228052 42306 228064
rect 42702 228052 42708 228064
rect 42300 228024 42708 228052
rect 42300 228012 42306 228024
rect 42702 228012 42708 228024
rect 42760 228012 42766 228064
rect 673546 206728 673552 206780
rect 673604 206768 673610 206780
rect 675294 206768 675300 206780
rect 673604 206740 675300 206768
rect 673604 206728 673610 206740
rect 675294 206728 675300 206740
rect 675352 206728 675358 206780
rect 673730 202920 673736 202972
rect 673788 202960 673794 202972
rect 673914 202960 673920 202972
rect 673788 202932 673920 202960
rect 673788 202920 673794 202932
rect 673914 202920 673920 202932
rect 673972 202960 673978 202972
rect 675386 202960 675392 202972
rect 673972 202932 675392 202960
rect 673972 202920 673978 202932
rect 675386 202920 675392 202932
rect 675444 202920 675450 202972
rect 42426 198636 42432 198688
rect 42484 198676 42490 198688
rect 42794 198676 42800 198688
rect 42484 198648 42800 198676
rect 42484 198636 42490 198648
rect 42794 198636 42800 198648
rect 42852 198636 42858 198688
rect 42242 197344 42248 197396
rect 42300 197384 42306 197396
rect 42518 197384 42524 197396
rect 42300 197356 42524 197384
rect 42300 197344 42306 197356
rect 42518 197344 42524 197356
rect 42576 197344 42582 197396
rect 41782 195848 41788 195900
rect 41840 195888 41846 195900
rect 42610 195888 42616 195900
rect 41840 195860 42616 195888
rect 41840 195848 41846 195860
rect 42610 195848 42616 195860
rect 42668 195888 42674 195900
rect 44634 195888 44640 195900
rect 42668 195860 44640 195888
rect 42668 195848 42674 195860
rect 44634 195848 44640 195860
rect 44692 195848 44698 195900
rect 673638 193196 673644 193248
rect 673696 193236 673702 193248
rect 674006 193236 674012 193248
rect 673696 193208 674012 193236
rect 673696 193196 673702 193208
rect 674006 193196 674012 193208
rect 674064 193196 674070 193248
rect 673638 191904 673644 191956
rect 673696 191944 673702 191956
rect 675386 191944 675392 191956
rect 673696 191916 675392 191944
rect 673696 191904 673702 191916
rect 675386 191904 675392 191916
rect 675444 191904 675450 191956
rect 42334 188300 42340 188352
rect 42392 188340 42398 188352
rect 42794 188340 42800 188352
rect 42392 188312 42800 188340
rect 42392 188300 42398 188312
rect 42794 188300 42800 188312
rect 42852 188300 42858 188352
rect 41782 184832 41788 184884
rect 41840 184872 41846 184884
rect 42242 184872 42248 184884
rect 41840 184844 42248 184872
rect 41840 184832 41846 184844
rect 42242 184832 42248 184844
rect 42300 184872 42306 184884
rect 42518 184872 42524 184884
rect 42300 184844 42524 184872
rect 42300 184832 42306 184844
rect 42518 184832 42524 184844
rect 42576 184832 42582 184884
rect 44542 173952 44548 174004
rect 44600 173992 44606 174004
rect 44726 173992 44732 174004
rect 44600 173964 44732 173992
rect 44600 173952 44606 173964
rect 44726 173952 44732 173964
rect 44784 173952 44790 174004
rect 42334 173884 42340 173936
rect 42392 173924 42398 173936
rect 42886 173924 42892 173936
rect 42392 173896 42892 173924
rect 42392 173884 42398 173896
rect 42886 173884 42892 173896
rect 42944 173884 42950 173936
rect 672718 173884 672724 173936
rect 672776 173924 672782 173936
rect 672902 173924 672908 173936
rect 672776 173896 672908 173924
rect 672776 173884 672782 173896
rect 672902 173884 672908 173896
rect 672960 173884 672966 173936
rect 44450 171028 44456 171080
rect 44508 171068 44514 171080
rect 44726 171068 44732 171080
rect 44508 171040 44732 171068
rect 44508 171028 44514 171040
rect 44726 171028 44732 171040
rect 44784 171028 44790 171080
rect 42518 160080 42524 160132
rect 42576 160120 42582 160132
rect 42886 160120 42892 160132
rect 42576 160092 42892 160120
rect 42576 160080 42582 160092
rect 42886 160080 42892 160092
rect 42944 160080 42950 160132
rect 673454 158312 673460 158364
rect 673512 158352 673518 158364
rect 675386 158352 675392 158364
rect 673512 158324 675392 158352
rect 673512 158312 673518 158324
rect 675386 158312 675392 158324
rect 675444 158312 675450 158364
rect 673546 157292 673552 157344
rect 673604 157332 673610 157344
rect 673914 157332 673920 157344
rect 673604 157304 673920 157332
rect 673604 157292 673610 157304
rect 673914 157292 673920 157304
rect 673972 157332 673978 157344
rect 675386 157332 675392 157344
rect 673972 157304 675392 157332
rect 673972 157292 673978 157304
rect 675386 157292 675392 157304
rect 675444 157292 675450 157344
rect 672534 156544 672540 156596
rect 672592 156584 672598 156596
rect 672718 156584 672724 156596
rect 672592 156556 672724 156584
rect 672592 156544 672598 156556
rect 672718 156544 672724 156556
rect 672776 156544 672782 156596
rect 44450 151784 44456 151836
rect 44508 151824 44514 151836
rect 44634 151824 44640 151836
rect 44508 151796 44640 151824
rect 44508 151784 44514 151796
rect 44634 151784 44640 151796
rect 44692 151784 44698 151836
rect 673638 147840 673644 147892
rect 673696 147880 673702 147892
rect 674006 147880 674012 147892
rect 673696 147852 674012 147880
rect 673696 147840 673702 147852
rect 674006 147840 674012 147852
rect 674064 147880 674070 147892
rect 675386 147880 675392 147892
rect 674064 147852 675392 147880
rect 674064 147840 674070 147852
rect 675386 147840 675392 147852
rect 675444 147840 675450 147892
rect 42334 140768 42340 140820
rect 42392 140808 42398 140820
rect 42518 140808 42524 140820
rect 42392 140780 42524 140808
rect 42392 140768 42398 140780
rect 42518 140768 42524 140780
rect 42576 140768 42582 140820
rect 44634 140768 44640 140820
rect 44692 140768 44698 140820
rect 44652 140672 44680 140768
rect 44726 140672 44732 140684
rect 44652 140644 44732 140672
rect 44726 140632 44732 140644
rect 44784 140632 44790 140684
rect 42150 131044 42156 131096
rect 42208 131084 42214 131096
rect 42334 131084 42340 131096
rect 42208 131056 42340 131084
rect 42208 131044 42214 131056
rect 42334 131044 42340 131056
rect 42392 131044 42398 131096
rect 44726 121564 44732 121576
rect 44652 121536 44732 121564
rect 44652 121440 44680 121536
rect 44726 121524 44732 121536
rect 44784 121524 44790 121576
rect 44634 121388 44640 121440
rect 44692 121388 44698 121440
rect 672718 115880 672724 115932
rect 672776 115920 672782 115932
rect 672810 115920 672816 115932
rect 672776 115892 672816 115920
rect 672776 115880 672782 115892
rect 672810 115880 672816 115892
rect 672868 115880 672874 115932
rect 673454 112752 673460 112804
rect 673512 112792 673518 112804
rect 675386 112792 675392 112804
rect 673512 112764 675392 112792
rect 673512 112752 673518 112764
rect 675386 112752 675392 112764
rect 675444 112752 675450 112804
rect 673546 112072 673552 112124
rect 673604 112112 673610 112124
rect 675386 112112 675392 112124
rect 673604 112084 675392 112112
rect 673604 112072 673610 112084
rect 675386 112072 675392 112084
rect 675444 112072 675450 112124
rect 672810 102184 672816 102196
rect 672736 102156 672816 102184
rect 672736 102128 672764 102156
rect 672810 102144 672816 102156
rect 672868 102144 672874 102196
rect 673638 102144 673644 102196
rect 673696 102184 673702 102196
rect 673822 102184 673828 102196
rect 673696 102156 673828 102184
rect 673696 102144 673702 102156
rect 673822 102144 673828 102156
rect 673880 102144 673886 102196
rect 672718 102076 672724 102128
rect 672776 102076 672782 102128
rect 673638 102008 673644 102060
rect 673696 102048 673702 102060
rect 675386 102048 675392 102060
rect 673696 102020 675392 102048
rect 673696 102008 673702 102020
rect 675386 102008 675392 102020
rect 675444 102008 675450 102060
rect 44266 96568 44272 96620
rect 44324 96608 44330 96620
rect 44542 96608 44548 96620
rect 44324 96580 44548 96608
rect 44324 96568 44330 96580
rect 44542 96568 44548 96580
rect 44600 96568 44606 96620
rect 672810 82900 672816 82952
rect 672868 82900 672874 82952
rect 672828 82748 672856 82900
rect 672810 82696 672816 82748
rect 672868 82696 672874 82748
rect 44266 77256 44272 77308
rect 44324 77296 44330 77308
rect 44358 77296 44364 77308
rect 44324 77268 44364 77296
rect 44324 77256 44330 77268
rect 44358 77256 44364 77268
rect 44416 77256 44422 77308
rect 39666 75216 39672 75268
rect 39724 75216 39730 75268
rect 39684 74996 39712 75216
rect 39666 74944 39672 74996
rect 39724 74944 39730 74996
rect 39574 67940 39580 67992
rect 39632 67980 39638 67992
rect 41414 67980 41420 67992
rect 39632 67952 41420 67980
rect 39632 67940 39638 67952
rect 41414 67940 41420 67952
rect 41472 67940 41478 67992
rect 41414 64608 41420 64660
rect 41472 64648 41478 64660
rect 42702 64648 42708 64660
rect 41472 64620 42708 64648
rect 41472 64608 41478 64620
rect 42702 64608 42708 64620
rect 42760 64608 42766 64660
rect 39666 52368 39672 52420
rect 39724 52408 39730 52420
rect 39850 52408 39856 52420
rect 39724 52380 39856 52408
rect 39724 52368 39730 52380
rect 39850 52368 39856 52380
rect 39908 52368 39914 52420
rect 45462 47880 45468 47932
rect 45520 47920 45526 47932
rect 195974 47920 195980 47932
rect 45520 47892 195980 47920
rect 45520 47880 45526 47892
rect 195974 47880 195980 47892
rect 196032 47880 196038 47932
rect 516318 47880 516324 47932
rect 516376 47920 516382 47932
rect 673638 47920 673644 47932
rect 516376 47892 673644 47920
rect 516376 47880 516382 47892
rect 673638 47880 673644 47892
rect 673696 47880 673702 47932
rect 39850 47812 39856 47864
rect 39908 47852 39914 47864
rect 189166 47852 189172 47864
rect 39908 47824 189172 47852
rect 39908 47812 39914 47824
rect 189166 47812 189172 47824
rect 189224 47812 189230 47864
rect 414198 47852 414204 47864
rect 411180 47824 414204 47852
rect 45554 47744 45560 47796
rect 45612 47784 45618 47796
rect 149054 47784 149060 47796
rect 45612 47756 149060 47784
rect 45612 47744 45618 47756
rect 149054 47744 149060 47756
rect 149112 47784 149118 47796
rect 150894 47784 150900 47796
rect 149112 47756 150900 47784
rect 149112 47744 149118 47756
rect 150894 47744 150900 47756
rect 150952 47744 150958 47796
rect 39758 47676 39764 47728
rect 39816 47716 39822 47728
rect 86402 47716 86408 47728
rect 39816 47688 86408 47716
rect 39816 47676 39822 47688
rect 86402 47676 86408 47688
rect 86460 47676 86466 47728
rect 411180 47716 411208 47824
rect 414198 47812 414204 47824
rect 414256 47852 414262 47864
rect 425054 47852 425060 47864
rect 414256 47824 425060 47852
rect 414256 47812 414262 47824
rect 425054 47812 425060 47824
rect 425112 47812 425118 47864
rect 430758 47812 430764 47864
rect 430816 47852 430822 47864
rect 430816 47824 444328 47852
rect 430816 47812 430822 47824
rect 444300 47784 444328 47824
rect 529842 47812 529848 47864
rect 529900 47852 529906 47864
rect 673454 47852 673460 47864
rect 529900 47824 673460 47852
rect 529900 47812 529906 47824
rect 673454 47812 673460 47824
rect 673512 47812 673518 47864
rect 444300 47756 449848 47784
rect 391952 47688 411208 47716
rect 449820 47716 449848 47756
rect 528646 47744 528652 47796
rect 528704 47784 528710 47796
rect 672810 47784 672816 47796
rect 528704 47756 672816 47784
rect 528704 47744 528710 47756
rect 672810 47744 672816 47756
rect 672868 47744 672874 47796
rect 466454 47716 466460 47728
rect 449820 47688 466460 47716
rect 192846 47472 192852 47524
rect 192904 47512 192910 47524
rect 201494 47512 201500 47524
rect 192904 47484 201500 47512
rect 192904 47472 192910 47484
rect 201494 47472 201500 47484
rect 201552 47472 201558 47524
rect 358814 47472 358820 47524
rect 358872 47512 358878 47524
rect 359366 47512 359372 47524
rect 358872 47484 359372 47512
rect 358872 47472 358878 47484
rect 359366 47472 359372 47484
rect 359424 47512 359430 47524
rect 391952 47512 391980 47688
rect 466454 47676 466460 47688
rect 466512 47676 466518 47728
rect 480162 47540 480168 47592
rect 480220 47580 480226 47592
rect 483014 47580 483020 47592
rect 480220 47552 483020 47580
rect 480220 47540 480226 47552
rect 483014 47540 483020 47552
rect 483072 47540 483078 47592
rect 422294 47512 422300 47524
rect 359424 47484 391980 47512
rect 411640 47484 422300 47512
rect 359424 47472 359430 47484
rect 328454 47444 328460 47456
rect 315776 47416 328460 47444
rect 248322 47336 248328 47388
rect 248380 47376 248386 47388
rect 248380 47348 276152 47376
rect 248380 47336 248386 47348
rect 276124 47308 276152 47348
rect 307570 47308 307576 47320
rect 206848 47280 276060 47308
rect 276124 47280 307576 47308
rect 199654 47200 199660 47252
rect 199712 47240 199718 47252
rect 206848 47240 206876 47280
rect 199712 47212 206876 47240
rect 199712 47200 199718 47212
rect 206922 47200 206928 47252
rect 206980 47240 206986 47252
rect 240134 47240 240140 47252
rect 206980 47212 240140 47240
rect 206980 47200 206986 47212
rect 240134 47200 240140 47212
rect 240192 47200 240198 47252
rect 150894 47132 150900 47184
rect 150952 47172 150958 47184
rect 192846 47172 192852 47184
rect 150952 47144 192852 47172
rect 150952 47132 150958 47144
rect 192846 47132 192852 47144
rect 192904 47132 192910 47184
rect 200850 47132 200856 47184
rect 200908 47172 200914 47184
rect 242894 47172 242900 47184
rect 200908 47144 242900 47172
rect 200908 47132 200914 47144
rect 242894 47132 242900 47144
rect 242952 47132 242958 47184
rect 276032 47172 276060 47280
rect 307570 47268 307576 47280
rect 307628 47308 307634 47320
rect 315776 47308 315804 47416
rect 328454 47404 328460 47416
rect 328512 47404 328518 47456
rect 411254 47404 411260 47456
rect 411312 47444 411318 47456
rect 411640 47444 411668 47484
rect 422294 47472 422300 47484
rect 422352 47472 422358 47524
rect 441522 47472 441528 47524
rect 441580 47512 441586 47524
rect 460934 47512 460940 47524
rect 441580 47484 460940 47512
rect 441580 47472 441586 47484
rect 460934 47472 460940 47484
rect 460992 47472 460998 47524
rect 411312 47416 411668 47444
rect 424980 47416 430620 47444
rect 411312 47404 411318 47416
rect 342254 47336 342260 47388
rect 342312 47376 342318 47388
rect 358722 47376 358728 47388
rect 342312 47348 358728 47376
rect 342312 47336 342318 47348
rect 358722 47336 358728 47348
rect 358780 47376 358786 47388
rect 361482 47376 361488 47388
rect 358780 47348 361488 47376
rect 358780 47336 358786 47348
rect 361482 47336 361488 47348
rect 361540 47336 361546 47388
rect 417234 47336 417240 47388
rect 417292 47376 417298 47388
rect 424980 47376 425008 47416
rect 417292 47348 425008 47376
rect 430592 47376 430620 47416
rect 488626 47404 488632 47456
rect 488684 47444 488690 47456
rect 516318 47444 516324 47456
rect 488684 47416 516324 47444
rect 488684 47404 488690 47416
rect 516318 47404 516324 47416
rect 516376 47404 516382 47456
rect 430592 47348 449848 47376
rect 417292 47336 417298 47348
rect 307628 47280 315804 47308
rect 307628 47268 307634 47280
rect 334066 47268 334072 47320
rect 334124 47308 334130 47320
rect 362402 47308 362408 47320
rect 334124 47280 362408 47308
rect 334124 47268 334130 47280
rect 362402 47268 362408 47280
rect 362460 47308 362466 47320
rect 391934 47308 391940 47320
rect 362460 47280 391940 47308
rect 362460 47268 362466 47280
rect 391934 47268 391940 47280
rect 391992 47268 391998 47320
rect 422294 47268 422300 47320
rect 422352 47308 422358 47320
rect 441522 47308 441528 47320
rect 422352 47280 441528 47308
rect 422352 47268 422358 47280
rect 441522 47268 441528 47280
rect 441580 47268 441586 47320
rect 449820 47308 449848 47348
rect 474642 47336 474648 47388
rect 474700 47376 474706 47388
rect 524414 47376 524420 47388
rect 474700 47348 524420 47376
rect 474700 47336 474706 47348
rect 524414 47336 524420 47348
rect 524472 47336 524478 47388
rect 453482 47308 453488 47320
rect 449820 47280 453488 47308
rect 453482 47268 453488 47280
rect 453540 47268 453546 47320
rect 309410 47200 309416 47252
rect 309468 47240 309474 47252
rect 352558 47240 352564 47252
rect 309468 47212 352564 47240
rect 309468 47200 309474 47212
rect 352558 47200 352564 47212
rect 352616 47200 352622 47252
rect 364242 47200 364248 47252
rect 364300 47240 364306 47252
rect 407390 47240 407396 47252
rect 364300 47212 407396 47240
rect 364300 47200 364306 47212
rect 407390 47200 407396 47212
rect 407448 47200 407454 47252
rect 419074 47200 419080 47252
rect 419132 47240 419138 47252
rect 462130 47240 462136 47252
rect 419132 47212 462136 47240
rect 419132 47200 419138 47212
rect 462130 47200 462136 47212
rect 462188 47200 462194 47252
rect 466454 47200 466460 47252
rect 466512 47240 466518 47252
rect 468938 47240 468944 47252
rect 466512 47212 468944 47240
rect 466512 47200 466518 47212
rect 468938 47200 468944 47212
rect 468996 47240 469002 47252
rect 469214 47240 469220 47252
rect 468996 47212 469220 47240
rect 468996 47200 469002 47212
rect 469214 47200 469220 47212
rect 469272 47200 469278 47252
rect 473814 47200 473820 47252
rect 473872 47240 473878 47252
rect 516962 47240 516968 47252
rect 473872 47212 516968 47240
rect 473872 47200 473878 47212
rect 516962 47200 516968 47212
rect 517020 47200 517026 47252
rect 527450 47240 527456 47252
rect 517440 47212 527456 47240
rect 289814 47172 289820 47184
rect 276032 47144 289820 47172
rect 289814 47132 289820 47144
rect 289872 47132 289878 47184
rect 305914 47132 305920 47184
rect 305972 47172 305978 47184
rect 351914 47172 351920 47184
rect 305972 47144 351920 47172
rect 305972 47132 305978 47144
rect 351914 47132 351920 47144
rect 351972 47132 351978 47184
rect 360562 47132 360568 47184
rect 360620 47172 360626 47184
rect 406746 47172 406752 47184
rect 360620 47144 406752 47172
rect 360620 47132 360626 47144
rect 406746 47132 406752 47144
rect 406804 47172 406810 47184
rect 411162 47172 411168 47184
rect 406804 47144 411168 47172
rect 406804 47132 406810 47144
rect 411162 47132 411168 47144
rect 411220 47132 411226 47184
rect 417878 47132 417884 47184
rect 417936 47172 417942 47184
rect 468294 47172 468300 47184
rect 417936 47144 468300 47172
rect 417936 47132 417942 47144
rect 468294 47132 468300 47144
rect 468352 47172 468358 47184
rect 517440 47172 517468 47212
rect 527450 47200 527456 47212
rect 527508 47240 527514 47252
rect 529842 47240 529848 47252
rect 527508 47212 529848 47240
rect 527508 47200 527514 47212
rect 529842 47200 529848 47212
rect 529900 47200 529906 47252
rect 468352 47144 517468 47172
rect 468352 47132 468358 47144
rect 524414 47132 524420 47184
rect 524472 47172 524478 47184
rect 526806 47172 526812 47184
rect 524472 47144 526812 47172
rect 524472 47132 524478 47144
rect 526806 47132 526812 47144
rect 526864 47172 526870 47184
rect 634814 47172 634820 47184
rect 526864 47144 634820 47172
rect 526864 47132 526870 47144
rect 634814 47132 634820 47144
rect 634872 47132 634878 47184
rect 186682 47064 186688 47116
rect 186740 47104 186746 47116
rect 194686 47104 194692 47116
rect 186740 47076 194692 47104
rect 186740 47064 186746 47076
rect 194686 47064 194692 47076
rect 194744 47064 194750 47116
rect 199010 47064 199016 47116
rect 199068 47104 199074 47116
rect 247310 47104 247316 47116
rect 199068 47076 247316 47104
rect 199068 47064 199074 47076
rect 247310 47064 247316 47076
rect 247368 47104 247374 47116
rect 248322 47104 248328 47116
rect 247368 47076 248328 47104
rect 247368 47064 247374 47076
rect 248322 47064 248328 47076
rect 248380 47064 248386 47116
rect 309042 47064 309048 47116
rect 309100 47104 309106 47116
rect 342254 47104 342260 47116
rect 309100 47076 342260 47104
rect 309100 47064 309106 47076
rect 342254 47064 342260 47076
rect 342312 47064 342318 47116
rect 361482 47064 361488 47116
rect 361540 47104 361546 47116
rect 363046 47104 363052 47116
rect 361540 47076 363052 47104
rect 361540 47064 361546 47076
rect 363046 47064 363052 47076
rect 363104 47104 363110 47116
rect 411070 47104 411076 47116
rect 363104 47076 411076 47104
rect 363104 47064 363110 47076
rect 411070 47064 411076 47076
rect 411128 47064 411134 47116
rect 523770 47104 523776 47116
rect 507780 47076 523776 47104
rect 195974 46996 195980 47048
rect 196032 47036 196038 47048
rect 304534 47036 304540 47048
rect 196032 47008 304540 47036
rect 196032 46996 196038 47008
rect 304534 46996 304540 47008
rect 304592 47036 304598 47048
rect 358814 47036 358820 47048
rect 304592 47008 358820 47036
rect 304592 46996 304598 47008
rect 358814 46996 358820 47008
rect 358872 46996 358878 47048
rect 391934 46996 391940 47048
rect 391992 47036 391998 47048
rect 410978 47036 410984 47048
rect 391992 47008 410984 47036
rect 391992 46996 391998 47008
rect 410978 46996 410984 47008
rect 411036 46996 411042 47048
rect 469214 46996 469220 47048
rect 469272 47036 469278 47048
rect 507780 47036 507808 47076
rect 523770 47064 523776 47076
rect 523828 47064 523834 47116
rect 569126 47104 569132 47116
rect 546420 47076 569132 47104
rect 546420 47036 546448 47076
rect 569126 47064 569132 47076
rect 569184 47064 569190 47116
rect 469272 47008 478000 47036
rect 469272 46996 469278 47008
rect 86402 46928 86408 46980
rect 86460 46968 86466 46980
rect 199010 46968 199016 46980
rect 86460 46940 199016 46968
rect 86460 46928 86466 46940
rect 199010 46928 199016 46940
rect 199068 46928 199074 46980
rect 201494 46928 201500 46980
rect 201552 46968 201558 46980
rect 206922 46968 206928 46980
rect 201552 46940 206928 46968
rect 201552 46928 201558 46940
rect 206922 46928 206928 46940
rect 206980 46928 206986 46980
rect 453482 46928 453488 46980
rect 453540 46968 453546 46980
rect 471974 46968 471980 46980
rect 453540 46940 471980 46968
rect 453540 46928 453546 46940
rect 471974 46928 471980 46940
rect 472032 46968 472038 46980
rect 474642 46968 474648 46980
rect 472032 46940 474648 46968
rect 472032 46928 472038 46940
rect 474642 46928 474648 46940
rect 474700 46928 474706 46980
rect 477972 46968 478000 47008
rect 488552 47008 507808 47036
rect 527192 47008 546448 47036
rect 488552 46968 488580 47008
rect 477972 46940 488580 46968
rect 514478 46928 514484 46980
rect 514536 46968 514542 46980
rect 522482 46968 522488 46980
rect 514536 46940 522488 46968
rect 514536 46928 514542 46940
rect 522482 46928 522488 46940
rect 522540 46928 522546 46980
rect 523770 46928 523776 46980
rect 523828 46968 523834 46980
rect 527192 46968 527220 47008
rect 523828 46940 527220 46968
rect 523828 46928 523834 46940
rect 42242 45636 42248 45688
rect 42300 45676 42306 45688
rect 143534 45676 143540 45688
rect 42300 45648 143540 45676
rect 42300 45636 42306 45648
rect 143534 45636 143540 45648
rect 143592 45636 143598 45688
rect 42702 45568 42708 45620
rect 42760 45608 42766 45620
rect 140958 45608 140964 45620
rect 42760 45580 140964 45608
rect 42760 45568 42766 45580
rect 140958 45568 140964 45580
rect 141016 45568 141022 45620
rect 242894 45500 242900 45552
rect 242952 45540 242958 45552
rect 297726 45540 297732 45552
rect 242952 45512 297732 45540
rect 242952 45500 242958 45512
rect 297726 45500 297732 45512
rect 297784 45500 297790 45552
rect 579154 45500 579160 45552
rect 579212 45540 579218 45552
rect 673546 45540 673552 45552
rect 579212 45512 673552 45540
rect 579212 45500 579218 45512
rect 673546 45500 673552 45512
rect 673604 45500 673610 45552
rect 410978 45364 410984 45416
rect 411036 45404 411042 45416
rect 417234 45404 417240 45416
rect 411036 45376 417240 45404
rect 411036 45364 411042 45376
rect 417234 45364 417240 45376
rect 417292 45364 417298 45416
rect 411070 44412 411076 44464
rect 411128 44452 411134 44464
rect 413554 44452 413560 44464
rect 411128 44424 413560 44452
rect 411128 44412 411134 44424
rect 413554 44412 413560 44424
rect 413612 44412 413618 44464
rect 143534 44208 143540 44260
rect 143592 44248 143598 44260
rect 145098 44248 145104 44260
rect 143592 44220 145104 44248
rect 143592 44208 143598 44220
rect 145098 44208 145104 44220
rect 145156 44248 145162 44260
rect 195330 44248 195336 44260
rect 145156 44220 195336 44248
rect 145156 44208 145162 44220
rect 195330 44208 195336 44220
rect 195388 44208 195394 44260
rect 140958 44140 140964 44192
rect 141016 44180 141022 44192
rect 254026 44180 254032 44192
rect 141016 44152 254032 44180
rect 141016 44140 141022 44152
rect 254026 44140 254032 44152
rect 254084 44180 254090 44192
rect 569218 44180 569224 44192
rect 254084 44152 569224 44180
rect 254084 44140 254090 44152
rect 569218 44140 569224 44152
rect 569276 44140 569282 44192
rect 303890 42236 303896 42288
rect 303948 42276 303954 42288
rect 308214 42276 308220 42288
rect 303948 42248 308220 42276
rect 303948 42236 303954 42248
rect 308214 42236 308220 42248
rect 308272 42236 308278 42288
rect 413554 42236 413560 42288
rect 413612 42276 413618 42288
rect 417878 42276 417884 42288
rect 413612 42248 417884 42276
rect 413612 42236 413618 42248
rect 417878 42236 417884 42248
rect 417936 42236 417942 42288
rect 302234 41964 302240 42016
rect 302292 42004 302298 42016
rect 304994 42004 305000 42016
rect 302292 41976 305000 42004
rect 302292 41964 302298 41976
rect 304994 41964 305000 41976
rect 305052 41964 305058 42016
rect 411530 42004 411536 42016
rect 410260 41976 411536 42004
rect 410260 41948 410288 41976
rect 411530 41964 411536 41976
rect 411588 42004 411594 42016
rect 414566 42004 414572 42016
rect 411588 41976 414572 42004
rect 411588 41964 411594 41976
rect 414566 41964 414572 41976
rect 414624 42004 414630 42016
rect 415854 42004 415860 42016
rect 414624 41976 415860 42004
rect 414624 41964 414630 41976
rect 415854 41964 415860 41976
rect 415912 42004 415918 42016
rect 418246 42004 418252 42016
rect 415912 41976 418252 42004
rect 415912 41964 415918 41976
rect 418246 41964 418252 41976
rect 418304 41964 418310 42016
rect 466362 42004 466368 42016
rect 465092 41976 466368 42004
rect 465092 41948 465120 41976
rect 466362 41964 466368 41976
rect 466420 42004 466426 42016
rect 469398 42004 469404 42016
rect 466420 41976 469404 42004
rect 466420 41964 466426 41976
rect 469398 41964 469404 41976
rect 469456 42004 469462 42016
rect 470686 42004 470692 42016
rect 469456 41976 470692 42004
rect 469456 41964 469462 41976
rect 470686 41964 470692 41976
rect 470744 42004 470750 42016
rect 473078 42004 473084 42016
rect 470744 41976 473084 42004
rect 470744 41964 470750 41976
rect 473078 41964 473084 41976
rect 473136 41964 473142 42016
rect 352650 41896 352656 41948
rect 352708 41936 352714 41948
rect 355502 41936 355508 41948
rect 352708 41908 355508 41936
rect 352708 41896 352714 41908
rect 355502 41896 355508 41908
rect 355560 41896 355566 41948
rect 356974 41896 356980 41948
rect 357032 41936 357038 41948
rect 359826 41936 359832 41948
rect 357032 41908 359832 41936
rect 357032 41896 357038 41908
rect 359826 41896 359832 41908
rect 359884 41936 359890 41948
rect 361114 41936 361120 41948
rect 359884 41908 361120 41936
rect 359884 41896 359890 41908
rect 361114 41896 361120 41908
rect 361172 41896 361178 41948
rect 407482 41896 407488 41948
rect 407540 41936 407546 41948
rect 410242 41936 410248 41948
rect 407540 41908 410248 41936
rect 407540 41896 407546 41908
rect 410242 41896 410248 41908
rect 410300 41896 410306 41948
rect 411162 41896 411168 41948
rect 411220 41936 411226 41948
rect 411220 41908 415624 41936
rect 411220 41896 411226 41908
rect 189258 41828 189264 41880
rect 189316 41868 189322 41880
rect 191098 41868 191104 41880
rect 189316 41840 191104 41868
rect 189316 41828 189322 41840
rect 191098 41828 191104 41840
rect 191156 41868 191162 41880
rect 192294 41868 192300 41880
rect 191156 41840 192300 41868
rect 191156 41828 191162 41840
rect 192294 41828 192300 41840
rect 192352 41868 192358 41880
rect 192352 41840 193628 41868
rect 192352 41828 192358 41840
rect 193600 41812 193628 41840
rect 195422 41828 195428 41880
rect 195480 41868 195486 41880
rect 199562 41868 199568 41880
rect 195480 41840 199568 41868
rect 195480 41828 195486 41840
rect 199562 41828 199568 41840
rect 199620 41828 199626 41880
rect 297910 41828 297916 41880
rect 297968 41868 297974 41880
rect 300670 41868 300676 41880
rect 297968 41840 300676 41868
rect 297968 41828 297974 41840
rect 300670 41828 300676 41840
rect 300728 41828 300734 41880
rect 352006 41828 352012 41880
rect 352064 41868 352070 41880
rect 354306 41868 354312 41880
rect 352064 41840 354312 41868
rect 352064 41828 352070 41840
rect 354306 41828 354312 41840
rect 354364 41868 354370 41880
rect 360470 41868 360476 41880
rect 354364 41840 360476 41868
rect 354364 41828 354370 41840
rect 360470 41828 360476 41840
rect 360528 41828 360534 41880
rect 188614 41760 188620 41812
rect 188672 41800 188678 41812
rect 192754 41800 192760 41812
rect 188672 41772 192760 41800
rect 188672 41760 188678 41772
rect 192754 41760 192760 41772
rect 192812 41760 192818 41812
rect 193582 41760 193588 41812
rect 193640 41800 193646 41812
rect 196434 41800 196440 41812
rect 193640 41772 196440 41800
rect 193640 41760 193646 41772
rect 196434 41760 196440 41772
rect 196492 41760 196498 41812
rect 198458 41760 198464 41812
rect 198516 41800 198522 41812
rect 200114 41800 200120 41812
rect 198516 41772 200120 41800
rect 198516 41760 198522 41772
rect 200114 41760 200120 41772
rect 200172 41760 200178 41812
rect 295426 41760 295432 41812
rect 295484 41800 295490 41812
rect 303154 41800 303160 41812
rect 295484 41772 303160 41800
rect 295484 41760 295490 41772
rect 303154 41760 303160 41772
rect 303212 41760 303218 41812
rect 305270 41760 305276 41812
rect 305328 41800 305334 41812
rect 306558 41800 306564 41812
rect 305328 41772 306564 41800
rect 305328 41760 305334 41772
rect 306558 41760 306564 41772
rect 306616 41800 306622 41812
rect 308674 41800 308680 41812
rect 306616 41772 308680 41800
rect 306616 41760 306622 41772
rect 308674 41760 308680 41772
rect 308732 41760 308738 41812
rect 350166 41760 350172 41812
rect 350224 41800 350230 41812
rect 357986 41800 357992 41812
rect 350224 41772 357992 41800
rect 350224 41760 350230 41772
rect 357986 41760 357992 41772
rect 358044 41760 358050 41812
rect 361132 41800 361160 41896
rect 409322 41828 409328 41880
rect 409380 41868 409386 41880
rect 412358 41868 412364 41880
rect 409380 41840 412364 41868
rect 409380 41828 409386 41840
rect 412358 41828 412364 41840
rect 412416 41868 412422 41880
rect 415486 41868 415492 41880
rect 412416 41840 415492 41868
rect 412416 41828 412422 41840
rect 415486 41828 415492 41840
rect 415544 41828 415550 41880
rect 415596 41868 415624 41908
rect 462314 41896 462320 41948
rect 462372 41936 462378 41948
rect 465074 41936 465080 41948
rect 462372 41908 465080 41936
rect 462372 41896 462378 41908
rect 465074 41896 465080 41908
rect 465132 41896 465138 41948
rect 465994 41896 466000 41948
rect 466052 41936 466058 41948
rect 474366 41936 474372 41948
rect 466052 41908 474372 41936
rect 466052 41896 466058 41908
rect 474366 41896 474372 41908
rect 474424 41896 474430 41948
rect 523218 41896 523224 41948
rect 523276 41936 523282 41948
rect 527358 41936 527364 41948
rect 523276 41908 527364 41936
rect 523276 41896 523282 41908
rect 527358 41896 527364 41908
rect 527416 41896 527422 41948
rect 419534 41868 419540 41880
rect 415596 41840 419540 41868
rect 419534 41828 419540 41840
rect 419592 41828 419598 41880
rect 464154 41828 464160 41880
rect 464212 41868 464218 41880
rect 466914 41868 466920 41880
rect 464212 41840 466920 41868
rect 464212 41828 464218 41840
rect 466914 41828 466920 41840
rect 466972 41868 466978 41880
rect 466972 41840 468432 41868
rect 466972 41828 466978 41840
rect 363506 41800 363512 41812
rect 361132 41772 363512 41800
rect 363506 41760 363512 41772
rect 363564 41760 363570 41812
rect 404998 41760 405004 41812
rect 405056 41800 405062 41812
rect 412726 41800 412732 41812
rect 405056 41772 412732 41800
rect 405056 41760 405062 41772
rect 412726 41760 412732 41772
rect 412784 41760 412790 41812
rect 459830 41760 459836 41812
rect 459888 41800 459894 41812
rect 467558 41800 467564 41812
rect 459888 41772 467564 41800
rect 459888 41760 459894 41772
rect 467558 41760 467564 41772
rect 467616 41760 467622 41812
rect 468404 41800 468432 41840
rect 468478 41828 468484 41880
rect 468536 41868 468542 41880
rect 472526 41868 472532 41880
rect 468536 41840 472532 41868
rect 468536 41828 468542 41840
rect 472526 41828 472532 41840
rect 472584 41828 472590 41880
rect 518894 41828 518900 41880
rect 518952 41868 518958 41880
rect 524874 41868 524880 41880
rect 518952 41840 524880 41868
rect 518952 41828 518958 41840
rect 524874 41828 524880 41840
rect 524932 41828 524938 41880
rect 470042 41800 470048 41812
rect 468404 41772 470048 41800
rect 470042 41760 470048 41772
rect 470100 41760 470106 41812
rect 517054 41760 517060 41812
rect 517112 41800 517118 41812
rect 520090 41800 520096 41812
rect 517112 41772 520096 41800
rect 517112 41760 517118 41772
rect 520090 41760 520096 41772
rect 520148 41800 520154 41812
rect 521378 41800 521384 41812
rect 520148 41772 521384 41800
rect 520148 41760 520154 41772
rect 521378 41760 521384 41772
rect 521436 41800 521442 41812
rect 524414 41800 524420 41812
rect 521436 41772 524420 41800
rect 521436 41760 521442 41772
rect 524414 41760 524420 41772
rect 524472 41800 524478 41812
rect 525702 41800 525708 41812
rect 524472 41772 525708 41800
rect 524472 41760 524478 41772
rect 525702 41760 525708 41772
rect 525760 41800 525766 41812
rect 527910 41800 527916 41812
rect 525760 41772 527916 41800
rect 525760 41760 525766 41772
rect 527910 41760 527916 41772
rect 527968 41760 527974 41812
rect 253934 41556 253940 41608
rect 253992 41596 253998 41608
rect 253992 41568 256740 41596
rect 253992 41556 253998 41568
rect 256712 41528 256740 41568
rect 256712 41500 275968 41528
rect 275940 41460 275968 41500
rect 290182 41460 290188 41472
rect 275940 41432 290188 41460
rect 290182 41420 290188 41432
rect 290240 41420 290246 41472
rect 133092 40196 133098 40248
rect 133150 40236 133156 40248
rect 143810 40236 143816 40248
rect 133150 40208 143816 40236
rect 133150 40196 133156 40208
rect 143810 40196 143816 40208
rect 143868 40196 143874 40248
rect 140990 40060 140996 40112
rect 141048 40100 141054 40112
rect 143066 40100 143072 40112
rect 141048 40072 143072 40100
rect 141048 40060 141054 40072
rect 142586 39950 142614 40072
rect 143066 40060 143072 40072
rect 143124 40100 143130 40112
rect 143350 40100 143356 40112
rect 143124 40072 143356 40100
rect 143124 40060 143130 40072
rect 143350 40060 143356 40072
rect 143408 40100 143414 40112
rect 143408 40072 144684 40100
rect 143408 40060 143414 40072
rect 144656 39984 144684 40072
rect 252094 39652 252100 39704
rect 252152 39692 252158 39704
rect 254026 39692 254032 39704
rect 252152 39664 254032 39692
rect 252152 39652 252158 39664
rect 254026 39652 254032 39664
rect 254084 39652 254090 39704
<< via1 >>
rect 84016 995596 84068 995648
rect 91744 995596 91796 995648
rect 238208 995596 238260 995648
rect 245936 995596 245988 995648
rect 531964 995596 532016 995648
rect 539692 995596 539744 995648
rect 135352 995460 135404 995512
rect 143172 995460 143224 995512
rect 633808 995460 633860 995512
rect 641536 995460 641588 995512
rect 289636 995256 289688 995308
rect 297640 995256 297692 995308
rect 391480 995256 391532 995308
rect 399484 995256 399536 995308
rect 480444 995256 480496 995308
rect 488448 995256 488500 995308
rect 82636 992060 82688 992112
rect 89996 992060 90048 992112
rect 79508 990768 79560 990820
rect 130936 990768 130988 990820
rect 131120 990768 131172 990820
rect 186688 990768 186740 990820
rect 194692 990768 194744 990820
rect 194784 990768 194836 990820
rect 233056 990768 233108 990820
rect 284668 990768 284720 990820
rect 386512 990768 386564 990820
rect 486608 990768 486660 990820
rect 538036 990768 538088 990820
rect 639788 990768 639840 990820
rect 78864 990700 78916 990752
rect 130292 990700 130344 990752
rect 182364 990700 182416 990752
rect 200028 990700 200080 990752
rect 244188 990700 244240 990752
rect 295800 990700 295852 990752
rect 397460 990700 397512 990752
rect 474740 990700 474792 990752
rect 475476 990700 475528 990752
rect 526904 990700 526956 990752
rect 626540 990700 626592 990752
rect 89996 990632 90048 990684
rect 141424 990632 141476 990684
rect 192852 990632 192904 990684
rect 233608 990632 233660 990684
rect 245568 990632 245620 990684
rect 42248 990360 42300 990412
rect 79508 990564 79560 990616
rect 130292 990564 130344 990616
rect 181720 990564 181772 990616
rect 285312 990632 285364 990684
rect 131120 990428 131172 990480
rect 132500 990428 132552 990480
rect 160008 990428 160060 990480
rect 182364 990496 182416 990548
rect 192852 990496 192904 990548
rect 244188 990496 244240 990548
rect 245568 990496 245620 990548
rect 285312 990496 285364 990548
rect 314476 990564 314528 990616
rect 314752 990564 314804 990616
rect 387156 990632 387208 990684
rect 476120 990632 476172 990684
rect 527548 990632 527600 990684
rect 629300 990632 629352 990684
rect 630956 990632 631008 990684
rect 328460 990496 328512 990548
rect 347688 990496 347740 990548
rect 386512 990564 386564 990616
rect 474740 990564 474792 990616
rect 397460 990496 397512 990548
rect 486608 990496 486660 990548
rect 42708 990292 42760 990344
rect 63408 990292 63460 990344
rect 140780 990292 140832 990344
rect 160100 990360 160152 990412
rect 181720 990428 181772 990480
rect 194784 990428 194836 990480
rect 200028 990292 200080 990344
rect 233608 990292 233660 990344
rect 275836 990292 275888 990344
rect 289728 990292 289780 990344
rect 328368 990292 328420 990344
rect 42432 990224 42484 990276
rect 45928 990224 45980 990276
rect 77300 990224 77352 990276
rect 78864 990156 78916 990208
rect 82912 990156 82964 990208
rect 121368 990224 121420 990276
rect 121460 990224 121512 990276
rect 328460 990224 328512 990276
rect 63408 990088 63460 990140
rect 82636 990088 82688 990140
rect 198740 990156 198792 990208
rect 160008 990088 160060 990140
rect 160100 990088 160152 990140
rect 179236 990088 179288 990140
rect 179512 990088 179564 990140
rect 198648 990088 198700 990140
rect 231860 990156 231912 990208
rect 256608 990156 256660 990208
rect 256792 990156 256844 990208
rect 231768 990088 231820 990140
rect 275836 990088 275888 990140
rect 289728 990088 289780 990140
rect 639788 990156 639840 990208
rect 673552 990156 673604 990208
rect 328184 990088 328236 990140
rect 626540 990088 626592 990140
rect 628656 990088 628708 990140
rect 630956 990088 631008 990140
rect 673644 990088 673696 990140
rect 673460 990020 673512 990072
rect 41788 969348 41840 969400
rect 42340 969348 42392 969400
rect 41788 968464 41840 968516
rect 42708 968464 42760 968516
rect 673460 965268 673512 965320
rect 675392 965268 675444 965320
rect 673644 964724 673696 964776
rect 675392 964724 675444 964776
rect 41788 962412 41840 962464
rect 42340 962412 42392 962464
rect 41788 956428 41840 956480
rect 42432 956428 42484 956480
rect 673552 953300 673604 953352
rect 675392 953300 675444 953352
rect 42432 950784 42484 950836
rect 42708 950784 42760 950836
rect 42432 946636 42484 946688
rect 42616 946636 42668 946688
rect 44272 930112 44324 930164
rect 45468 930112 45520 930164
rect 39672 922904 39724 922956
rect 44272 922904 44324 922956
rect 39856 921748 39908 921800
rect 42248 921748 42300 921800
rect 39856 916240 39908 916292
rect 41420 916240 41472 916292
rect 42708 913588 42760 913640
rect 42800 913452 42852 913504
rect 673644 910732 673696 910784
rect 677784 910732 677836 910784
rect 42432 885912 42484 885964
rect 42616 885912 42668 885964
rect 673460 876120 673512 876172
rect 675392 876120 675444 876172
rect 41420 875576 41472 875628
rect 42248 875576 42300 875628
rect 673644 875508 673696 875560
rect 675392 875508 675444 875560
rect 675208 870136 675260 870188
rect 675392 870136 675444 870188
rect 673552 864968 673604 865020
rect 675392 864968 675444 865020
rect 674656 862792 674708 862844
rect 675300 862792 675352 862844
rect 673920 850552 673972 850604
rect 674656 850552 674708 850604
rect 42616 850008 42668 850060
rect 42708 850008 42760 850060
rect 42616 830764 42668 830816
rect 42800 830764 42852 830816
rect 673736 830764 673788 830816
rect 674012 830764 674064 830816
rect 673828 816960 673880 817012
rect 674012 816960 674064 817012
rect 672816 811384 672868 811436
rect 673092 811384 673144 811436
rect 42524 807440 42576 807492
rect 42524 807236 42576 807288
rect 42248 806352 42300 806404
rect 42616 806352 42668 806404
rect 42340 804244 42392 804296
rect 42800 804244 42852 804296
rect 41788 798124 41840 798176
rect 42340 798124 42392 798176
rect 674012 797580 674064 797632
rect 675300 797580 675352 797632
rect 41788 787856 41840 787908
rect 42248 787856 42300 787908
rect 42616 787856 42668 787908
rect 41788 787584 41840 787636
rect 42524 787584 42576 787636
rect 673460 785272 673512 785324
rect 675392 785272 675444 785324
rect 673000 778336 673052 778388
rect 673184 778268 673236 778320
rect 673552 774868 673604 774920
rect 675392 774868 675444 774920
rect 673092 772760 673144 772812
rect 673184 772760 673236 772812
rect 41788 754468 41840 754520
rect 42432 754468 42484 754520
rect 41788 744404 41840 744456
rect 42432 744404 42484 744456
rect 42616 744404 42668 744456
rect 673828 741888 673880 741940
rect 675392 741888 675444 741940
rect 673460 741344 673512 741396
rect 675392 741344 675444 741396
rect 673184 739712 673236 739764
rect 673092 739508 673144 739560
rect 673460 736584 673512 736636
rect 675300 736584 675352 736636
rect 42248 730804 42300 730856
rect 42616 730804 42668 730856
rect 673552 730124 673604 730176
rect 673920 730124 673972 730176
rect 675392 730124 675444 730176
rect 673736 720332 673788 720384
rect 673920 720332 673972 720384
rect 672816 712036 672868 712088
rect 673000 712036 673052 712088
rect 41788 711288 41840 711340
rect 42708 711220 42760 711272
rect 673460 710676 673512 710728
rect 675300 710676 675352 710728
rect 42340 708704 42392 708756
rect 42616 708704 42668 708756
rect 673828 701088 673880 701140
rect 673644 701020 673696 701072
rect 41788 700952 41840 701004
rect 42340 700952 42392 701004
rect 42524 700952 42576 701004
rect 673644 695920 673696 695972
rect 673828 695920 673880 695972
rect 675392 695920 675444 695972
rect 42708 695444 42760 695496
rect 42984 695444 43036 695496
rect 672816 692792 672868 692844
rect 673184 692792 673236 692844
rect 673460 681708 673512 681760
rect 675208 681708 675260 681760
rect 42800 676200 42852 676252
rect 42984 676200 43036 676252
rect 673000 676132 673052 676184
rect 673092 676132 673144 676184
rect 673644 676132 673696 676184
rect 673920 676132 673972 676184
rect 42340 672256 42392 672308
rect 42524 672256 42576 672308
rect 41788 669060 41840 669112
rect 42432 669060 42484 669112
rect 42800 669060 42852 669112
rect 41788 657636 41840 657688
rect 42340 657636 42392 657688
rect 42616 657636 42668 657688
rect 42248 657092 42300 657144
rect 42708 657092 42760 657144
rect 673092 656888 673144 656940
rect 673184 656888 673236 656940
rect 673552 656888 673604 656940
rect 673920 656888 673972 656940
rect 673460 651720 673512 651772
rect 673828 651720 673880 651772
rect 675392 651720 675444 651772
rect 673552 651108 673604 651160
rect 673828 651108 673880 651160
rect 675392 651108 675444 651160
rect 673552 639684 673604 639736
rect 673736 639684 673788 639736
rect 675392 639684 675444 639736
rect 672816 637508 672868 637560
rect 673092 637508 673144 637560
rect 673736 637508 673788 637560
rect 674012 637508 674064 637560
rect 41788 625880 41840 625932
rect 42524 625880 42576 625932
rect 42248 618468 42300 618520
rect 42800 618468 42852 618520
rect 672816 618264 672868 618316
rect 673000 618264 673052 618316
rect 673736 618264 673788 618316
rect 673920 618264 673972 618316
rect 41788 614116 41840 614168
rect 42340 614116 42392 614168
rect 673460 606704 673512 606756
rect 673828 606704 673880 606756
rect 675392 606704 675444 606756
rect 672816 605820 672868 605872
rect 673000 605820 673052 605872
rect 673920 605616 673972 605668
rect 675300 605616 675352 605668
rect 673644 604460 673696 604512
rect 673920 604460 673972 604512
rect 42616 604392 42668 604444
rect 42708 604324 42760 604376
rect 672816 596164 672868 596216
rect 673000 596164 673052 596216
rect 672816 596028 672868 596080
rect 673000 596028 673052 596080
rect 673552 594872 673604 594924
rect 675392 594872 675444 594924
rect 672816 585080 672868 585132
rect 673000 585080 673052 585132
rect 41788 581680 41840 581732
rect 42708 581680 42760 581732
rect 41788 571616 41840 571668
rect 42524 571616 42576 571668
rect 673828 561484 673880 561536
rect 675392 561484 675444 561536
rect 673460 559920 673512 559972
rect 673644 559920 673696 559972
rect 675392 559920 675444 559972
rect 673552 550468 673604 550520
rect 675392 550468 675444 550520
rect 42432 546456 42484 546508
rect 42616 546456 42668 546508
rect 41788 538500 41840 538552
rect 42432 538500 42484 538552
rect 672908 538228 672960 538280
rect 673092 538228 673144 538280
rect 41788 527756 41840 527808
rect 42524 527756 42576 527808
rect 672908 527008 672960 527060
rect 673184 527008 673236 527060
rect 673000 499536 673052 499588
rect 673276 499536 673328 499588
rect 673000 482944 673052 482996
rect 673276 482944 673328 482996
rect 673460 463632 673512 463684
rect 677692 463632 677744 463684
rect 39396 458192 39448 458244
rect 44272 458192 44324 458244
rect 39856 448264 39908 448316
rect 42248 448264 42300 448316
rect 676220 440172 676272 440224
rect 677692 440172 677744 440224
rect 42248 413380 42300 413432
rect 42616 413380 42668 413432
rect 672816 412496 672868 412548
rect 676220 412496 676272 412548
rect 41788 410932 41840 410984
rect 42432 410932 42484 410984
rect 42248 405356 42300 405408
rect 42524 405356 42576 405408
rect 41788 400800 41840 400852
rect 42616 400800 42668 400852
rect 42248 400120 42300 400172
rect 42524 400120 42576 400172
rect 672724 386316 672776 386368
rect 672908 386316 672960 386368
rect 673552 384004 673604 384056
rect 675392 384004 675444 384056
rect 673460 382576 673512 382628
rect 673644 382576 673696 382628
rect 675300 382576 675352 382628
rect 673920 372308 673972 372360
rect 675392 372308 675444 372360
rect 41788 368636 41840 368688
rect 42432 368636 42484 368688
rect 42248 357620 42300 357672
rect 42616 357620 42668 357672
rect 41788 356668 41840 356720
rect 42524 356668 42576 356720
rect 672724 353336 672776 353388
rect 672724 353200 672776 353252
rect 672724 347692 672776 347744
rect 672908 347692 672960 347744
rect 42248 342184 42300 342236
rect 42616 342184 42668 342236
rect 673460 338512 673512 338564
rect 673644 338512 673696 338564
rect 675392 338512 675444 338564
rect 672540 328448 672592 328500
rect 672908 328448 672960 328500
rect 42616 328380 42668 328432
rect 42892 328380 42944 328432
rect 673828 327088 673880 327140
rect 675392 327088 675444 327140
rect 41788 324504 41840 324556
rect 42432 324504 42484 324556
rect 42708 324504 42760 324556
rect 672540 316004 672592 316056
rect 672724 316004 672776 316056
rect 42892 315120 42944 315172
rect 41788 315052 41840 315104
rect 41788 314440 41840 314492
rect 42340 314440 42392 314492
rect 42524 314440 42576 314492
rect 42432 313556 42484 313608
rect 42708 313556 42760 313608
rect 42708 309068 42760 309120
rect 42892 309068 42944 309120
rect 672448 306348 672500 306400
rect 672724 306348 672776 306400
rect 673552 293564 673604 293616
rect 675392 293564 675444 293616
rect 42708 289824 42760 289876
rect 42984 289824 43036 289876
rect 673644 283024 673696 283076
rect 675392 283024 675444 283076
rect 41788 282276 41840 282328
rect 42432 282276 42484 282328
rect 42616 277176 42668 277228
rect 42984 277176 43036 277228
rect 672632 276020 672684 276072
rect 672540 275952 672592 276004
rect 41788 271464 41840 271516
rect 42616 271464 42668 271516
rect 42616 270512 42668 270564
rect 42708 270512 42760 270564
rect 672540 260788 672592 260840
rect 672908 260788 672960 260840
rect 673644 256640 673696 256692
rect 674012 256640 674064 256692
rect 672724 251200 672776 251252
rect 672908 251200 672960 251252
rect 672540 251064 672592 251116
rect 672724 251064 672776 251116
rect 673552 248140 673604 248192
rect 675392 248140 675444 248192
rect 673460 247460 673512 247512
rect 673736 247460 673788 247512
rect 675392 247460 675444 247512
rect 42156 245624 42208 245676
rect 42340 245624 42392 245676
rect 42156 240592 42208 240644
rect 42708 240592 42760 240644
rect 41788 238076 41840 238128
rect 42432 238076 42484 238128
rect 42616 238076 42668 238128
rect 674012 237736 674064 237788
rect 675392 237736 675444 237788
rect 673828 231820 673880 231872
rect 674012 231820 674064 231872
rect 41788 228624 41840 228676
rect 42432 228624 42484 228676
rect 42892 228624 42944 228676
rect 41788 228012 41840 228064
rect 42248 228012 42300 228064
rect 42708 228012 42760 228064
rect 673552 206728 673604 206780
rect 675300 206728 675352 206780
rect 673736 202920 673788 202972
rect 673920 202920 673972 202972
rect 675392 202920 675444 202972
rect 42432 198636 42484 198688
rect 42800 198636 42852 198688
rect 42248 197344 42300 197396
rect 42524 197344 42576 197396
rect 41788 195848 41840 195900
rect 42616 195848 42668 195900
rect 44640 195848 44692 195900
rect 673644 193196 673696 193248
rect 674012 193196 674064 193248
rect 673644 191904 673696 191956
rect 675392 191904 675444 191956
rect 42340 188300 42392 188352
rect 42800 188300 42852 188352
rect 41788 184832 41840 184884
rect 42248 184832 42300 184884
rect 42524 184832 42576 184884
rect 44548 173952 44600 174004
rect 44732 173952 44784 174004
rect 42340 173884 42392 173936
rect 42892 173884 42944 173936
rect 672724 173884 672776 173936
rect 672908 173884 672960 173936
rect 44456 171028 44508 171080
rect 44732 171028 44784 171080
rect 42524 160080 42576 160132
rect 42892 160080 42944 160132
rect 673460 158312 673512 158364
rect 675392 158312 675444 158364
rect 673552 157292 673604 157344
rect 673920 157292 673972 157344
rect 675392 157292 675444 157344
rect 672540 156544 672592 156596
rect 672724 156544 672776 156596
rect 44456 151784 44508 151836
rect 44640 151784 44692 151836
rect 673644 147840 673696 147892
rect 674012 147840 674064 147892
rect 675392 147840 675444 147892
rect 42340 140768 42392 140820
rect 42524 140768 42576 140820
rect 44640 140768 44692 140820
rect 44732 140632 44784 140684
rect 42156 131044 42208 131096
rect 42340 131044 42392 131096
rect 44732 121524 44784 121576
rect 44640 121388 44692 121440
rect 672724 115880 672776 115932
rect 672816 115880 672868 115932
rect 673460 112752 673512 112804
rect 675392 112752 675444 112804
rect 673552 112072 673604 112124
rect 675392 112072 675444 112124
rect 672816 102144 672868 102196
rect 673644 102144 673696 102196
rect 673828 102144 673880 102196
rect 672724 102076 672776 102128
rect 673644 102008 673696 102060
rect 675392 102008 675444 102060
rect 44272 96568 44324 96620
rect 44548 96568 44600 96620
rect 672816 82900 672868 82952
rect 672816 82696 672868 82748
rect 44272 77256 44324 77308
rect 44364 77256 44416 77308
rect 39672 75216 39724 75268
rect 39672 74944 39724 74996
rect 39580 67940 39632 67992
rect 41420 67940 41472 67992
rect 41420 64608 41472 64660
rect 42708 64608 42760 64660
rect 39672 52368 39724 52420
rect 39856 52368 39908 52420
rect 45468 47880 45520 47932
rect 195980 47880 196032 47932
rect 516324 47880 516376 47932
rect 673644 47880 673696 47932
rect 39856 47812 39908 47864
rect 189172 47812 189224 47864
rect 45560 47744 45612 47796
rect 149060 47744 149112 47796
rect 150900 47744 150952 47796
rect 39764 47676 39816 47728
rect 86408 47676 86460 47728
rect 414204 47812 414256 47864
rect 425060 47812 425112 47864
rect 430764 47812 430816 47864
rect 529848 47812 529900 47864
rect 673460 47812 673512 47864
rect 528652 47744 528704 47796
rect 672816 47744 672868 47796
rect 192852 47472 192904 47524
rect 201500 47472 201552 47524
rect 358820 47472 358872 47524
rect 359372 47472 359424 47524
rect 466460 47676 466512 47728
rect 480168 47540 480220 47592
rect 483020 47540 483072 47592
rect 248328 47336 248380 47388
rect 199660 47200 199712 47252
rect 206928 47200 206980 47252
rect 240140 47200 240192 47252
rect 150900 47132 150952 47184
rect 192852 47132 192904 47184
rect 200856 47132 200908 47184
rect 242900 47132 242952 47184
rect 307576 47268 307628 47320
rect 328460 47404 328512 47456
rect 411260 47404 411312 47456
rect 422300 47472 422352 47524
rect 441528 47472 441580 47524
rect 460940 47472 460992 47524
rect 342260 47336 342312 47388
rect 358728 47336 358780 47388
rect 361488 47336 361540 47388
rect 417240 47336 417292 47388
rect 488632 47404 488684 47456
rect 516324 47404 516376 47456
rect 334072 47268 334124 47320
rect 362408 47268 362460 47320
rect 391940 47268 391992 47320
rect 422300 47268 422352 47320
rect 441528 47268 441580 47320
rect 474648 47336 474700 47388
rect 524420 47336 524472 47388
rect 453488 47268 453540 47320
rect 309416 47200 309468 47252
rect 352564 47200 352616 47252
rect 364248 47200 364300 47252
rect 407396 47200 407448 47252
rect 419080 47200 419132 47252
rect 462136 47200 462188 47252
rect 466460 47200 466512 47252
rect 468944 47200 468996 47252
rect 469220 47200 469272 47252
rect 473820 47200 473872 47252
rect 516968 47200 517020 47252
rect 289820 47132 289872 47184
rect 305920 47132 305972 47184
rect 351920 47132 351972 47184
rect 360568 47132 360620 47184
rect 406752 47132 406804 47184
rect 411168 47132 411220 47184
rect 417884 47132 417936 47184
rect 468300 47132 468352 47184
rect 527456 47200 527508 47252
rect 529848 47200 529900 47252
rect 524420 47132 524472 47184
rect 526812 47132 526864 47184
rect 634820 47132 634872 47184
rect 186688 47064 186740 47116
rect 194692 47064 194744 47116
rect 199016 47064 199068 47116
rect 247316 47064 247368 47116
rect 248328 47064 248380 47116
rect 309048 47064 309100 47116
rect 342260 47064 342312 47116
rect 361488 47064 361540 47116
rect 363052 47064 363104 47116
rect 411076 47064 411128 47116
rect 195980 46996 196032 47048
rect 304540 46996 304592 47048
rect 358820 46996 358872 47048
rect 391940 46996 391992 47048
rect 410984 46996 411036 47048
rect 469220 46996 469272 47048
rect 523776 47064 523828 47116
rect 569132 47064 569184 47116
rect 86408 46928 86460 46980
rect 199016 46928 199068 46980
rect 201500 46928 201552 46980
rect 206928 46928 206980 46980
rect 453488 46928 453540 46980
rect 471980 46928 472032 46980
rect 474648 46928 474700 46980
rect 514484 46928 514536 46980
rect 522488 46928 522540 46980
rect 523776 46928 523828 46980
rect 42248 45636 42300 45688
rect 143540 45636 143592 45688
rect 42708 45568 42760 45620
rect 140964 45568 141016 45620
rect 242900 45500 242952 45552
rect 297732 45500 297784 45552
rect 579160 45500 579212 45552
rect 673552 45500 673604 45552
rect 410984 45364 411036 45416
rect 417240 45364 417292 45416
rect 411076 44412 411128 44464
rect 413560 44412 413612 44464
rect 143540 44208 143592 44260
rect 145104 44208 145156 44260
rect 195336 44208 195388 44260
rect 140964 44140 141016 44192
rect 254032 44140 254084 44192
rect 569224 44140 569276 44192
rect 303896 42236 303948 42288
rect 308220 42236 308272 42288
rect 413560 42236 413612 42288
rect 417884 42236 417936 42288
rect 302240 41964 302292 42016
rect 305000 41964 305052 42016
rect 411536 41964 411588 42016
rect 414572 41964 414624 42016
rect 415860 41964 415912 42016
rect 418252 41964 418304 42016
rect 466368 41964 466420 42016
rect 469404 41964 469456 42016
rect 470692 41964 470744 42016
rect 473084 41964 473136 42016
rect 352656 41896 352708 41948
rect 355508 41896 355560 41948
rect 356980 41896 357032 41948
rect 359832 41896 359884 41948
rect 361120 41896 361172 41948
rect 407488 41896 407540 41948
rect 410248 41896 410300 41948
rect 411168 41896 411220 41948
rect 189264 41828 189316 41880
rect 191104 41828 191156 41880
rect 192300 41828 192352 41880
rect 195428 41828 195480 41880
rect 199568 41828 199620 41880
rect 297916 41828 297968 41880
rect 300676 41828 300728 41880
rect 352012 41828 352064 41880
rect 354312 41828 354364 41880
rect 360476 41828 360528 41880
rect 188620 41760 188672 41812
rect 192760 41760 192812 41812
rect 193588 41760 193640 41812
rect 196440 41760 196492 41812
rect 198464 41760 198516 41812
rect 200120 41760 200172 41812
rect 295432 41760 295484 41812
rect 303160 41760 303212 41812
rect 305276 41760 305328 41812
rect 306564 41760 306616 41812
rect 308680 41760 308732 41812
rect 350172 41760 350224 41812
rect 357992 41760 358044 41812
rect 409328 41828 409380 41880
rect 412364 41828 412416 41880
rect 415492 41828 415544 41880
rect 462320 41896 462372 41948
rect 465080 41896 465132 41948
rect 466000 41896 466052 41948
rect 474372 41896 474424 41948
rect 523224 41896 523276 41948
rect 527364 41896 527416 41948
rect 419540 41828 419592 41880
rect 464160 41828 464212 41880
rect 466920 41828 466972 41880
rect 363512 41760 363564 41812
rect 405004 41760 405056 41812
rect 412732 41760 412784 41812
rect 459836 41760 459888 41812
rect 467564 41760 467616 41812
rect 468484 41828 468536 41880
rect 472532 41828 472584 41880
rect 518900 41828 518952 41880
rect 524880 41828 524932 41880
rect 470048 41760 470100 41812
rect 517060 41760 517112 41812
rect 520096 41760 520148 41812
rect 521384 41760 521436 41812
rect 524420 41760 524472 41812
rect 525708 41760 525760 41812
rect 527916 41760 527968 41812
rect 253940 41556 253992 41608
rect 290188 41420 290240 41472
rect 133098 40196 133150 40248
rect 143816 40196 143868 40248
rect 140996 40060 141048 40112
rect 143072 40060 143124 40112
rect 143356 40060 143408 40112
rect 252100 39652 252152 39704
rect 254032 39652 254084 39704
<< metal2 >>
rect 328550 997384 328606 997393
rect 328550 997319 328606 997328
rect 77049 995407 77105 995887
rect 77693 995407 77749 995887
rect 78337 995407 78393 995887
rect 78876 990758 78904 995452
rect 79520 990826 79548 995452
rect 80177 995407 80233 995887
rect 80729 995407 80785 995887
rect 81373 995407 81429 995887
rect 82017 995407 82073 995887
rect 82569 995407 82625 995887
rect 83213 995407 83269 995887
rect 84016 995648 84068 995654
rect 84016 995590 84068 995596
rect 84028 995466 84056 995590
rect 83858 995438 84056 995466
rect 84501 995407 84557 995887
rect 85053 995407 85109 995887
rect 85697 995407 85753 995887
rect 86341 995407 86397 995887
rect 87537 995407 87593 995887
rect 88733 995407 88789 995887
rect 89377 995407 89433 995887
rect 90008 992118 90036 995452
rect 91217 995407 91273 995887
rect 91744 995648 91796 995654
rect 91744 995590 91796 995596
rect 91756 995466 91784 995590
rect 91756 995438 91862 995466
rect 128449 995407 128505 995887
rect 129093 995407 129149 995887
rect 129737 995407 129793 995887
rect 82636 992112 82688 992118
rect 82636 992054 82688 992060
rect 89996 992112 90048 992118
rect 89996 992054 90048 992060
rect 79508 990820 79560 990826
rect 79508 990762 79560 990768
rect 78864 990752 78916 990758
rect 78864 990694 78916 990700
rect 42248 990412 42300 990418
rect 42248 990354 42300 990360
rect 41722 969870 41828 969898
rect 41800 969406 41828 969870
rect 41788 969400 41840 969406
rect 41788 969342 41840 969348
rect 41713 969217 42193 969273
rect 41788 968516 41840 968522
rect 41788 968458 41840 968464
rect 41800 968063 41828 968458
rect 41722 968035 41828 968063
rect 41713 967377 42193 967433
rect 41713 966733 42193 966789
rect 41713 965537 42193 965593
rect 41713 964341 42193 964397
rect 41713 963697 42193 963753
rect 41713 963053 42193 963109
rect 41713 962501 42193 962557
rect 41788 962464 41840 962470
rect 41788 962406 41840 962412
rect 41800 961874 41828 962406
rect 41722 961846 41828 961874
rect 41713 961213 42193 961269
rect 41713 960569 42193 960625
rect 41713 960017 42193 960073
rect 41713 959373 42193 959429
rect 41713 958729 42193 958785
rect 41713 958177 42193 958233
rect 41722 957547 41828 957575
rect 41800 957386 41828 957547
rect 42260 957386 42288 990354
rect 42708 990344 42760 990350
rect 42708 990286 42760 990292
rect 63408 990344 63460 990350
rect 63408 990286 63460 990292
rect 77298 990312 77354 990321
rect 42432 990276 42484 990282
rect 42432 990218 42484 990224
rect 42340 969400 42392 969406
rect 42340 969342 42392 969348
rect 42352 962470 42380 969342
rect 42340 962464 42392 962470
rect 42340 962406 42392 962412
rect 41800 957358 42288 957386
rect 41722 956903 41828 956931
rect 41800 956486 41828 956903
rect 41788 956480 41840 956486
rect 41788 956422 41840 956428
rect 41713 956337 42193 956393
rect 41713 955693 42193 955749
rect 41713 955049 42193 955105
rect 39330 922962 39712 922978
rect 39330 922956 39724 922962
rect 39330 922950 39672 922956
rect 39672 922898 39724 922904
rect 39670 922312 39726 922321
rect 39670 922247 39726 922256
rect 39684 920281 39712 922247
rect 42260 921806 42288 957358
rect 42444 956486 42472 990218
rect 42720 968522 42748 990286
rect 45928 990276 45980 990282
rect 45928 990218 45980 990224
rect 45466 990176 45522 990185
rect 45466 990111 45522 990120
rect 42708 968516 42760 968522
rect 42708 968458 42760 968464
rect 42432 956480 42484 956486
rect 42432 956422 42484 956428
rect 42444 950994 42472 956422
rect 42444 950966 42564 950994
rect 42432 950836 42484 950842
rect 42432 950778 42484 950784
rect 42444 946694 42472 950778
rect 42432 946688 42484 946694
rect 42432 946630 42484 946636
rect 39856 921800 39908 921806
rect 39856 921742 39908 921748
rect 42248 921800 42300 921806
rect 42248 921742 42300 921748
rect 39670 920272 39726 920281
rect 39670 920207 39726 920216
rect 39868 919034 39896 921742
rect 39567 919006 39896 919034
rect 39868 916298 39896 919006
rect 39856 916292 39908 916298
rect 39856 916234 39908 916240
rect 41420 916292 41472 916298
rect 41420 916234 41472 916240
rect 39330 912206 39712 912234
rect 39684 908177 39712 912206
rect 39670 908168 39726 908177
rect 39670 908103 39726 908112
rect 40130 877568 40186 877577
rect 40130 877503 40186 877512
rect 40144 870097 40172 877503
rect 41432 875634 41460 916234
rect 42432 885964 42484 885970
rect 42432 885906 42484 885912
rect 41420 875628 41472 875634
rect 41420 875570 41472 875576
rect 42248 875628 42300 875634
rect 42248 875570 42300 875576
rect 41432 875129 41460 875570
rect 41418 875120 41474 875129
rect 41418 875055 41474 875064
rect 40130 870088 40186 870097
rect 40130 870023 40186 870032
rect 40498 830784 40554 830793
rect 40498 830719 40554 830728
rect 39606 827750 39712 827778
rect 39684 827529 39712 827750
rect 39670 827520 39726 827529
rect 39670 827455 39726 827464
rect 40512 811617 40540 830719
rect 40498 811608 40554 811617
rect 40498 811543 40554 811552
rect 42260 806410 42288 875570
rect 42444 866697 42472 885906
rect 42430 866688 42486 866697
rect 42430 866623 42486 866632
rect 42536 807498 42564 950966
rect 42720 950842 42748 968458
rect 42708 950836 42760 950842
rect 42708 950778 42760 950784
rect 42616 946688 42668 946694
rect 42616 946630 42668 946636
rect 42628 927466 42656 946630
rect 45480 930170 45508 990111
rect 44272 930164 44324 930170
rect 44272 930106 44324 930112
rect 45468 930164 45520 930170
rect 45468 930106 45520 930112
rect 42628 927438 42748 927466
rect 42720 913646 42748 927438
rect 44284 922962 44312 930106
rect 44272 922956 44324 922962
rect 44272 922898 44324 922904
rect 42708 913640 42760 913646
rect 42708 913582 42760 913588
rect 42800 913504 42852 913510
rect 42800 913446 42852 913452
rect 42812 894418 42840 913446
rect 42812 894390 42932 894418
rect 42904 886009 42932 894390
rect 42614 886000 42670 886009
rect 42614 885935 42616 885944
rect 42668 885935 42670 885944
rect 42890 886000 42946 886009
rect 42890 885935 42946 885944
rect 42616 885906 42668 885912
rect 44178 870088 44234 870097
rect 44178 870023 44234 870032
rect 42706 866688 42762 866697
rect 42706 866623 42762 866632
rect 42720 850066 42748 866623
rect 42616 850060 42668 850066
rect 42616 850002 42668 850008
rect 42708 850060 42760 850066
rect 42708 850002 42760 850008
rect 42628 830822 42656 850002
rect 42616 830816 42668 830822
rect 42616 830758 42668 830764
rect 42800 830816 42852 830822
rect 42800 830758 42852 830764
rect 42524 807492 42576 807498
rect 42524 807434 42576 807440
rect 42524 807288 42576 807294
rect 42524 807230 42576 807236
rect 42248 806404 42300 806410
rect 42248 806346 42300 806352
rect 42340 804296 42392 804302
rect 42340 804238 42392 804244
rect 41722 800075 41828 800103
rect 41800 799898 41828 800075
rect 41800 799870 42288 799898
rect 41713 799417 42193 799473
rect 41722 798238 41828 798266
rect 41800 798182 41828 798238
rect 41788 798176 41840 798182
rect 41788 798118 41840 798124
rect 41713 797577 42193 797633
rect 41713 796933 42193 796989
rect 41713 795737 42193 795793
rect 41713 794541 42193 794597
rect 41713 793897 42193 793953
rect 41713 793253 42193 793309
rect 41713 792701 42193 792757
rect 42260 792282 42288 799870
rect 42352 798182 42380 804238
rect 42340 798176 42392 798182
rect 42340 798118 42392 798124
rect 41800 792254 42288 792282
rect 41800 792099 41828 792254
rect 41722 792071 41828 792099
rect 41713 791413 42193 791469
rect 41713 790769 42193 790825
rect 41713 790217 42193 790273
rect 41713 789573 42193 789629
rect 41713 788929 42193 788985
rect 41713 788377 42193 788433
rect 41788 787908 41840 787914
rect 41788 787850 41840 787856
rect 42248 787908 42300 787914
rect 42248 787850 42300 787856
rect 41800 787794 41828 787850
rect 41722 787766 41828 787794
rect 41788 787636 41840 787642
rect 41788 787578 41840 787584
rect 41800 787114 41828 787578
rect 41722 787086 41828 787114
rect 41713 786537 42193 786593
rect 41713 785893 42193 785949
rect 41713 785249 42193 785305
rect 39854 778560 39910 778569
rect 39854 778495 39910 778504
rect 39868 772857 39896 778495
rect 39854 772848 39910 772857
rect 39854 772783 39910 772792
rect 42260 757058 42288 787850
rect 42352 757194 42380 798118
rect 42536 787658 42564 807230
rect 42616 806404 42668 806410
rect 42616 806346 42668 806352
rect 42628 787914 42656 806346
rect 42812 804302 42840 830758
rect 42800 804296 42852 804302
rect 42800 804238 42852 804244
rect 42616 787908 42668 787914
rect 42616 787850 42668 787856
rect 42536 787642 42656 787658
rect 42524 787636 42656 787642
rect 42576 787630 42656 787636
rect 42524 787578 42576 787584
rect 42352 757166 42472 757194
rect 42260 757030 42380 757058
rect 41722 756894 42288 756922
rect 41713 756217 42193 756273
rect 41722 755035 41828 755063
rect 41800 754526 41828 755035
rect 41788 754520 41840 754526
rect 41788 754462 41840 754468
rect 41713 754377 42193 754433
rect 41713 753733 42193 753789
rect 41713 752537 42193 752593
rect 41713 751341 42193 751397
rect 41713 750697 42193 750753
rect 41713 750053 42193 750109
rect 41713 749501 42193 749557
rect 42260 749034 42288 756894
rect 41800 749006 42288 749034
rect 41800 748898 41828 749006
rect 41722 748870 41828 748898
rect 41713 748213 42193 748269
rect 41713 747569 42193 747625
rect 41713 747017 42193 747073
rect 41713 746373 42193 746429
rect 41713 745729 42193 745785
rect 41713 745177 42193 745233
rect 42352 744575 42380 757030
rect 42444 754526 42472 757166
rect 42432 754520 42484 754526
rect 42484 754468 42564 754474
rect 42432 754462 42564 754468
rect 42444 754446 42564 754462
rect 41722 744547 42380 744575
rect 41788 744456 41840 744462
rect 41788 744398 41840 744404
rect 41800 743931 41828 744398
rect 41722 743903 41828 743931
rect 41713 743337 42193 743393
rect 41713 742693 42193 742749
rect 41713 742049 42193 742105
rect 42260 730862 42288 744547
rect 42432 744456 42484 744462
rect 42432 744398 42484 744404
rect 42248 730856 42300 730862
rect 42248 730798 42300 730804
rect 41722 713675 42288 713703
rect 41713 713017 42193 713073
rect 41722 711835 41828 711863
rect 41800 711346 41828 711835
rect 41788 711340 41840 711346
rect 41788 711282 41840 711288
rect 41713 711177 42193 711233
rect 41713 710533 42193 710589
rect 41713 709337 42193 709393
rect 41713 708141 42193 708197
rect 41713 707497 42193 707553
rect 41713 706853 42193 706909
rect 41713 706301 42193 706357
rect 42260 705786 42288 713675
rect 42340 708756 42392 708762
rect 42340 708698 42392 708704
rect 41800 705758 42288 705786
rect 41800 705699 41828 705758
rect 41722 705671 41828 705699
rect 41713 705013 42193 705069
rect 41713 704369 42193 704425
rect 41713 703817 42193 703873
rect 41713 703173 42193 703229
rect 41713 702529 42193 702585
rect 41713 701977 42193 702033
rect 41722 701347 41828 701375
rect 41800 701010 41828 701347
rect 42352 701010 42380 708698
rect 41788 701004 41840 701010
rect 41788 700946 41840 700952
rect 42340 701004 42392 701010
rect 42340 700946 42392 700952
rect 42444 700754 42472 744398
rect 42536 731082 42564 754446
rect 42628 744462 42656 787630
rect 42616 744456 42668 744462
rect 42616 744398 42668 744404
rect 42536 731054 42840 731082
rect 42616 730856 42668 730862
rect 42616 730798 42668 730804
rect 42628 708762 42656 730798
rect 42708 711272 42760 711278
rect 42812 711226 42840 731054
rect 42760 711220 42840 711226
rect 42708 711214 42840 711220
rect 42720 711198 42840 711214
rect 42616 708756 42668 708762
rect 42616 708698 42668 708704
rect 42524 701004 42576 701010
rect 42524 700946 42576 700952
rect 41722 700726 42472 700754
rect 41713 700137 42193 700193
rect 41713 699493 42193 699549
rect 41713 698849 42193 698905
rect 42340 672308 42392 672314
rect 42340 672250 42392 672256
rect 41722 670475 42288 670503
rect 41713 669817 42193 669873
rect 41788 669112 41840 669118
rect 41788 669054 41840 669060
rect 41800 668658 41828 669054
rect 41722 668630 41828 668658
rect 41713 667977 42193 668033
rect 41713 667333 42193 667389
rect 41713 666137 42193 666193
rect 41713 664941 42193 664997
rect 41713 664297 42193 664353
rect 41713 663653 42193 663709
rect 41713 663101 42193 663157
rect 42260 662538 42288 670475
rect 41708 662510 42288 662538
rect 41708 662485 41736 662510
rect 41713 661813 42193 661869
rect 41713 661169 42193 661225
rect 41713 660617 42193 660673
rect 41713 659973 42193 660029
rect 41713 659329 42193 659385
rect 41713 658777 42193 658833
rect 41722 658158 41828 658186
rect 41800 657694 41828 658158
rect 42352 657694 42380 672250
rect 42444 672058 42472 700726
rect 42536 672314 42564 700946
rect 42720 695502 42748 711198
rect 42708 695496 42760 695502
rect 42708 695438 42760 695444
rect 42984 695496 43036 695502
rect 42984 695438 43036 695444
rect 42996 676258 43024 695438
rect 42800 676252 42852 676258
rect 42800 676194 42852 676200
rect 42984 676252 43036 676258
rect 42984 676194 43036 676200
rect 42524 672308 42576 672314
rect 42524 672250 42576 672256
rect 42444 672030 42564 672058
rect 42432 669112 42484 669118
rect 42432 669054 42484 669060
rect 42536 669066 42564 672030
rect 42812 669118 42840 676194
rect 42800 669112 42852 669118
rect 41788 657688 41840 657694
rect 41788 657630 41840 657636
rect 42340 657688 42392 657694
rect 42340 657630 42392 657636
rect 41722 657478 41920 657506
rect 41892 657098 41920 657478
rect 42260 657150 42288 657181
rect 42248 657144 42300 657150
rect 41892 657092 42248 657098
rect 41892 657086 42300 657092
rect 41892 657070 42288 657086
rect 41713 656937 42193 656993
rect 41713 656293 42193 656349
rect 41713 655649 42193 655705
rect 42260 633434 42288 657070
rect 42444 652746 42472 669054
rect 42536 669038 42748 669066
rect 42800 669054 42852 669060
rect 42616 657688 42668 657694
rect 42616 657630 42668 657636
rect 42628 656962 42656 657630
rect 42720 657150 42748 669038
rect 42708 657144 42760 657150
rect 42708 657086 42760 657092
rect 42628 656934 42748 656962
rect 42352 652718 42472 652746
rect 42352 633570 42380 652718
rect 42720 643090 42748 656934
rect 42720 643062 42840 643090
rect 42352 633542 42564 633570
rect 42260 633406 42380 633434
rect 41722 627286 42288 627314
rect 41713 626617 42193 626673
rect 41788 625932 41840 625938
rect 41788 625874 41840 625880
rect 41800 625463 41828 625874
rect 41722 625435 41828 625463
rect 41713 624777 42193 624833
rect 41713 624133 42193 624189
rect 41713 622937 42193 622993
rect 41713 621741 42193 621797
rect 41713 621097 42193 621153
rect 41713 620453 42193 620509
rect 41713 619901 42193 619957
rect 42260 619426 42288 627286
rect 41800 619398 42288 619426
rect 41800 619290 41828 619398
rect 41722 619262 41828 619290
rect 41713 618613 42193 618669
rect 42248 618520 42300 618526
rect 42248 618462 42300 618468
rect 41713 617969 42193 618025
rect 41713 617417 42193 617473
rect 41713 616773 42193 616829
rect 41713 616129 42193 616185
rect 41713 615577 42193 615633
rect 41708 614938 41736 614961
rect 42260 614938 42288 618462
rect 41708 614910 42288 614938
rect 41722 614303 41828 614331
rect 41800 614174 41828 614303
rect 41788 614168 41840 614174
rect 41788 614110 41840 614116
rect 41713 613737 42193 613793
rect 41713 613093 42193 613149
rect 41713 612449 42193 612505
rect 42260 584202 42288 614910
rect 42352 614174 42380 633406
rect 42536 625938 42564 633542
rect 42524 625932 42576 625938
rect 42524 625874 42576 625880
rect 42536 625818 42564 625874
rect 42536 625790 42656 625818
rect 42340 614168 42392 614174
rect 42340 614110 42392 614116
rect 42352 584338 42380 614110
rect 42628 604450 42656 625790
rect 42812 618526 42840 643062
rect 42800 618520 42852 618526
rect 42800 618462 42852 618468
rect 42616 604444 42668 604450
rect 42616 604386 42668 604392
rect 42708 604376 42760 604382
rect 42708 604318 42760 604324
rect 42352 584310 42564 584338
rect 42260 584174 42380 584202
rect 41722 584075 42288 584103
rect 41713 583417 42193 583473
rect 41722 582235 41828 582263
rect 41800 581738 41828 582235
rect 41788 581732 41840 581738
rect 41788 581674 41840 581680
rect 41713 581577 42193 581633
rect 41713 580933 42193 580989
rect 41713 579737 42193 579793
rect 41713 578541 42193 578597
rect 41713 577897 42193 577953
rect 41713 577253 42193 577309
rect 41713 576701 42193 576757
rect 42260 576178 42288 584075
rect 41892 576150 42288 576178
rect 41892 576099 41920 576150
rect 41722 576071 41920 576099
rect 41713 575413 42193 575469
rect 41713 574769 42193 574825
rect 41713 574217 42193 574273
rect 41713 573573 42193 573629
rect 41713 572929 42193 572985
rect 41713 572377 42193 572433
rect 42352 571775 42380 584174
rect 41722 571747 42380 571775
rect 41788 571668 41840 571674
rect 41788 571610 41840 571616
rect 41800 571146 41828 571610
rect 41722 571118 41828 571146
rect 41713 570537 42193 570593
rect 41713 569893 42193 569949
rect 41713 569249 42193 569305
rect 40222 550624 40278 550633
rect 40222 550559 40278 550568
rect 40236 546417 40264 550559
rect 40222 546408 40278 546417
rect 40222 546343 40278 546352
rect 42260 541090 42288 571747
rect 42536 571674 42564 584310
rect 42720 581738 42748 604318
rect 42708 581732 42760 581738
rect 42708 581674 42760 581680
rect 42524 571668 42576 571674
rect 42524 571610 42576 571616
rect 42432 546508 42484 546514
rect 42432 546450 42484 546456
rect 42260 541062 42380 541090
rect 41722 540875 42288 540903
rect 41713 540217 42193 540273
rect 41722 539022 41828 539050
rect 41800 538558 41828 539022
rect 41788 538552 41840 538558
rect 41788 538494 41840 538500
rect 41713 538377 42193 538433
rect 41713 537733 42193 537789
rect 41713 536537 42193 536593
rect 41713 535341 42193 535397
rect 41713 534697 42193 534753
rect 41713 534053 42193 534109
rect 41713 533501 42193 533557
rect 42260 532930 42288 540875
rect 41708 532902 42288 532930
rect 41708 532885 41736 532902
rect 41713 532213 42193 532269
rect 41713 531569 42193 531625
rect 41713 531017 42193 531073
rect 41713 530373 42193 530429
rect 41713 529729 42193 529785
rect 41713 529177 42193 529233
rect 42352 528850 42380 541062
rect 42444 538558 42472 546450
rect 42432 538552 42484 538558
rect 42432 538494 42484 538500
rect 41800 528822 42380 528850
rect 41800 528578 41828 528822
rect 41722 528550 41828 528578
rect 41722 527903 41828 527931
rect 41800 527814 41828 527903
rect 41788 527808 41840 527814
rect 41788 527750 41840 527756
rect 41713 527337 42193 527393
rect 41713 526693 42193 526749
rect 41713 526049 42193 526105
rect 39606 493190 39804 493218
rect 39776 492969 39804 493190
rect 39762 492960 39818 492969
rect 39762 492895 39818 492904
rect 39396 458244 39448 458250
rect 39396 458186 39448 458192
rect 39408 451874 39436 458186
rect 39946 455424 40002 455433
rect 39946 455359 40002 455368
rect 39670 451888 39726 451897
rect 39330 451846 39670 451874
rect 39670 451823 39726 451832
rect 39856 448316 39908 448322
rect 39856 448258 39908 448264
rect 39868 447794 39896 448258
rect 39567 447766 39896 447794
rect 39670 441008 39726 441017
rect 39330 440966 39670 440994
rect 39960 440994 39988 455359
rect 42260 448322 42288 528822
rect 42248 448316 42300 448322
rect 42248 448258 42300 448264
rect 39726 440966 39988 440994
rect 39670 440943 39726 440952
rect 42260 413438 42288 448258
rect 42248 413432 42300 413438
rect 42248 413374 42300 413380
rect 41722 413275 42288 413303
rect 41713 412617 42193 412673
rect 41722 411454 41828 411482
rect 41800 410990 41828 411454
rect 41788 410984 41840 410990
rect 41788 410926 41840 410932
rect 41713 410777 42193 410833
rect 41713 410133 42193 410189
rect 41713 408937 42193 408993
rect 41713 407741 42193 407797
rect 41713 407097 42193 407153
rect 41713 406453 42193 406509
rect 41713 405901 42193 405957
rect 42260 405498 42288 413275
rect 42444 410990 42472 538494
rect 42536 527814 42564 571610
rect 42720 546666 42748 581674
rect 42628 546638 42748 546666
rect 42628 546514 42656 546638
rect 42616 546508 42668 546514
rect 42616 546450 42668 546456
rect 42524 527808 42576 527814
rect 42524 527750 42576 527756
rect 42432 410984 42484 410990
rect 42432 410926 42484 410932
rect 41892 405470 42288 405498
rect 41892 405299 41920 405470
rect 42248 405408 42300 405414
rect 42248 405350 42300 405356
rect 41722 405271 41920 405299
rect 41713 404613 42193 404669
rect 41713 403969 42193 404025
rect 41713 403417 42193 403473
rect 41713 402773 42193 402829
rect 41713 402129 42193 402185
rect 41713 401577 42193 401633
rect 41722 400947 41828 400975
rect 41800 400858 41828 400947
rect 41788 400852 41840 400858
rect 41788 400794 41840 400800
rect 42260 400330 42288 405350
rect 41722 400302 42288 400330
rect 42260 400178 42288 400302
rect 42248 400172 42300 400178
rect 42248 400114 42300 400120
rect 41713 399737 42193 399793
rect 41713 399093 42193 399149
rect 41713 398449 42193 398505
rect 41722 370075 42288 370103
rect 41713 369417 42193 369473
rect 41788 368688 41840 368694
rect 41788 368630 41840 368636
rect 41800 368263 41828 368630
rect 41722 368235 41828 368263
rect 41713 367577 42193 367633
rect 41713 366933 42193 366989
rect 41713 365737 42193 365793
rect 41713 364541 42193 364597
rect 41713 363897 42193 363953
rect 41713 363253 42193 363309
rect 41713 362701 42193 362757
rect 42260 362250 42288 370075
rect 42444 368694 42472 410926
rect 42536 405414 42564 527750
rect 42616 413432 42668 413438
rect 42616 413374 42668 413380
rect 42524 405408 42576 405414
rect 42524 405350 42576 405356
rect 42628 400858 42656 413374
rect 42616 400852 42668 400858
rect 42616 400794 42668 400800
rect 42524 400172 42576 400178
rect 42524 400114 42576 400120
rect 42432 368688 42484 368694
rect 42432 368630 42484 368636
rect 41800 362222 42288 362250
rect 41800 362114 41828 362222
rect 41722 362086 41828 362114
rect 41713 361413 42193 361469
rect 41713 360769 42193 360825
rect 41713 360217 42193 360273
rect 41713 359573 42193 359629
rect 41713 358929 42193 358985
rect 41713 358377 42193 358433
rect 41722 357734 41920 357762
rect 41892 357626 41920 357734
rect 42260 357678 42288 357709
rect 42248 357672 42300 357678
rect 41892 357620 42248 357626
rect 41892 357614 42300 357620
rect 41892 357598 42288 357614
rect 41722 357103 41828 357131
rect 41800 356726 41828 357103
rect 41788 356720 41840 356726
rect 41788 356662 41840 356668
rect 41713 356537 42193 356593
rect 41713 355893 42193 355949
rect 41713 355249 42193 355305
rect 42260 342242 42288 357598
rect 42248 342236 42300 342242
rect 42248 342178 42300 342184
rect 41722 326862 42288 326890
rect 41713 326217 42193 326273
rect 41722 325035 41828 325063
rect 41800 324562 41828 325035
rect 41788 324556 41840 324562
rect 41788 324498 41840 324504
rect 41713 324377 42193 324433
rect 41713 323733 42193 323789
rect 41713 322537 42193 322593
rect 41713 321341 42193 321397
rect 41713 320697 42193 320753
rect 41713 320053 42193 320109
rect 41713 319501 42193 319557
rect 42260 318899 42288 326862
rect 42444 324562 42472 368630
rect 42536 356726 42564 400114
rect 42628 357678 42656 400794
rect 42616 357672 42668 357678
rect 42616 357614 42668 357620
rect 42524 356720 42576 356726
rect 42524 356662 42576 356668
rect 42432 324556 42484 324562
rect 42432 324498 42484 324504
rect 41953 318871 42288 318899
rect 41713 318213 42193 318269
rect 41713 317569 42193 317625
rect 41713 317017 42193 317073
rect 41713 316373 42193 316429
rect 41713 315729 42193 315785
rect 41713 315177 42193 315233
rect 41788 315104 41840 315110
rect 41788 315046 41840 315052
rect 41800 314575 41828 315046
rect 41722 314547 41828 314575
rect 42536 314498 42564 356662
rect 42616 342236 42668 342242
rect 42616 342178 42668 342184
rect 42628 328438 42656 342178
rect 42616 328432 42668 328438
rect 42616 328374 42668 328380
rect 42892 328432 42944 328438
rect 42892 328374 42944 328380
rect 42708 324556 42760 324562
rect 42708 324498 42760 324504
rect 41788 314492 41840 314498
rect 41788 314434 41840 314440
rect 42340 314492 42392 314498
rect 42340 314434 42392 314440
rect 42524 314492 42576 314498
rect 42524 314434 42576 314440
rect 41800 313931 41828 314434
rect 41722 313903 41828 313931
rect 41713 313337 42193 313393
rect 41713 312693 42193 312749
rect 41713 312049 42193 312105
rect 41722 283675 41828 283703
rect 41800 283506 41828 283675
rect 41800 283478 42288 283506
rect 41713 283017 42193 283073
rect 41788 282328 41840 282334
rect 41788 282270 41840 282276
rect 41800 281874 41828 282270
rect 41722 281846 41828 281874
rect 41713 281177 42193 281233
rect 41713 280533 42193 280589
rect 41713 279337 42193 279393
rect 41713 278141 42193 278197
rect 41713 277497 42193 277553
rect 41713 276853 42193 276909
rect 41713 276301 42193 276357
rect 42260 275722 42288 283478
rect 41694 275713 41750 275722
rect 41694 275648 41750 275657
rect 42246 275713 42302 275722
rect 42246 275648 42302 275657
rect 41713 275013 42193 275069
rect 41713 274369 42193 274425
rect 41713 273817 42193 273873
rect 41713 273173 42193 273229
rect 41713 272529 42193 272585
rect 41713 271977 42193 272033
rect 41788 271516 41840 271522
rect 41788 271458 41840 271464
rect 41800 271402 41828 271458
rect 41722 271374 41828 271402
rect 42352 270722 42380 314434
rect 42720 313614 42748 324498
rect 42904 315194 42932 328374
rect 42904 315178 43024 315194
rect 42892 315172 43024 315178
rect 42944 315166 43024 315172
rect 42892 315114 42944 315120
rect 42432 313608 42484 313614
rect 42432 313550 42484 313556
rect 42708 313608 42760 313614
rect 42708 313550 42760 313556
rect 42444 282334 42472 313550
rect 42996 309210 43024 315166
rect 42904 309182 43024 309210
rect 42904 309126 42932 309182
rect 42708 309120 42760 309126
rect 42708 309062 42760 309068
rect 42892 309120 42944 309126
rect 42892 309062 42944 309068
rect 42720 289882 42748 309062
rect 42708 289876 42760 289882
rect 42708 289818 42760 289824
rect 42984 289876 43036 289882
rect 42984 289818 43036 289824
rect 42432 282328 42484 282334
rect 42432 282270 42484 282276
rect 41722 270694 42380 270722
rect 41713 270137 42193 270193
rect 41713 269493 42193 269549
rect 41713 268849 42193 268905
rect 42352 245682 42380 270694
rect 42156 245676 42208 245682
rect 42156 245618 42208 245624
rect 42340 245676 42392 245682
rect 42340 245618 42392 245624
rect 42168 240650 42196 245618
rect 42156 240644 42208 240650
rect 42156 240586 42208 240592
rect 41722 240502 42288 240530
rect 41713 239817 42193 239873
rect 41722 238635 41828 238663
rect 41800 238134 41828 238635
rect 41788 238128 41840 238134
rect 41788 238070 41840 238076
rect 41713 237977 42193 238033
rect 41713 237333 42193 237389
rect 41713 236137 42193 236193
rect 41713 234941 42193 234997
rect 41713 234297 42193 234353
rect 41713 233653 42193 233709
rect 41713 233101 42193 233157
rect 42260 232642 42288 240502
rect 42444 238134 42472 282270
rect 42996 277234 43024 289818
rect 42616 277228 42668 277234
rect 42616 277170 42668 277176
rect 42984 277228 43036 277234
rect 42984 277170 43036 277176
rect 42628 271522 42656 277170
rect 42616 271516 42668 271522
rect 42616 271458 42668 271464
rect 42628 270570 42656 271458
rect 42616 270564 42668 270570
rect 42616 270506 42668 270512
rect 42708 270564 42760 270570
rect 42708 270506 42760 270512
rect 42720 256714 42748 270506
rect 42536 256686 42748 256714
rect 42536 245562 42564 256686
rect 42536 245534 42932 245562
rect 42708 240644 42760 240650
rect 42708 240586 42760 240592
rect 42432 238128 42484 238134
rect 42432 238070 42484 238076
rect 42616 238128 42668 238134
rect 42616 238070 42668 238076
rect 41892 232614 42288 232642
rect 41892 232506 41920 232614
rect 41722 232478 41920 232506
rect 41713 231813 42193 231869
rect 41713 231169 42193 231225
rect 41713 230617 42193 230673
rect 41713 229973 42193 230029
rect 41713 229329 42193 229385
rect 41713 228777 42193 228833
rect 41788 228676 41840 228682
rect 41788 228618 41840 228624
rect 42432 228676 42484 228682
rect 42432 228618 42484 228624
rect 41800 228154 41828 228618
rect 41722 228126 41828 228154
rect 41788 228064 41840 228070
rect 41788 228006 41840 228012
rect 42248 228064 42300 228070
rect 42248 228006 42300 228012
rect 41800 227531 41828 228006
rect 41722 227503 41828 227531
rect 41713 226937 42193 226993
rect 41713 226293 42193 226349
rect 41713 225649 42193 225705
rect 42260 197402 42288 228006
rect 42444 198694 42472 228618
rect 42432 198688 42484 198694
rect 42432 198630 42484 198636
rect 42248 197396 42300 197402
rect 42248 197338 42300 197344
rect 42524 197396 42576 197402
rect 42524 197338 42576 197344
rect 41722 197254 42288 197282
rect 41713 196617 42193 196673
rect 41788 195900 41840 195906
rect 41788 195842 41840 195848
rect 41800 195463 41828 195842
rect 41722 195435 41828 195463
rect 41713 194777 42193 194833
rect 41713 194133 42193 194189
rect 41713 192937 42193 192993
rect 41713 191741 42193 191797
rect 41713 191097 42193 191153
rect 41713 190453 42193 190509
rect 41713 189901 42193 189957
rect 42260 189394 42288 197254
rect 41800 189366 42288 189394
rect 41800 189299 41828 189366
rect 41722 189271 41828 189299
rect 41713 188613 42193 188669
rect 42340 188352 42392 188358
rect 42340 188294 42392 188300
rect 41713 187969 42193 188025
rect 41713 187417 42193 187473
rect 41713 186773 42193 186829
rect 41713 186129 42193 186185
rect 41713 185577 42193 185633
rect 42352 184998 42380 188294
rect 41694 184989 41750 184998
rect 41694 184924 41750 184933
rect 42338 184989 42394 184998
rect 42338 184924 42394 184933
rect 41788 184884 41840 184890
rect 41788 184826 41840 184832
rect 42248 184884 42300 184890
rect 42248 184826 42300 184832
rect 41800 184331 41828 184826
rect 41722 184303 41828 184331
rect 41713 183737 42193 183793
rect 41713 183093 42193 183149
rect 41713 182449 42193 182505
rect 42156 131096 42208 131102
rect 42156 131038 42208 131044
rect 39606 120278 39804 120306
rect 39776 120193 39804 120278
rect 39762 120184 39818 120193
rect 39762 120119 39818 120128
rect 42168 115977 42196 131038
rect 41418 115968 41474 115977
rect 41418 115903 41474 115912
rect 42154 115968 42210 115977
rect 42154 115903 42210 115912
rect 39394 84280 39450 84289
rect 39394 84215 39450 84224
rect 39408 79098 39436 84215
rect 39316 79070 39528 79098
rect 39316 78948 39344 79070
rect 39500 78962 39528 79070
rect 39500 78934 39712 78962
rect 39684 75274 39712 78934
rect 39672 75268 39724 75274
rect 39672 75210 39724 75216
rect 39592 75126 39804 75154
rect 39592 75018 39620 75126
rect 39567 74990 39620 75018
rect 39672 74996 39724 75002
rect 39672 74938 39724 74944
rect 39330 68190 39620 68218
rect 39592 67998 39620 68190
rect 39580 67992 39632 67998
rect 39580 67934 39632 67940
rect 39684 52426 39712 74938
rect 39672 52420 39724 52426
rect 39672 52362 39724 52368
rect 39776 47734 39804 75126
rect 41432 67998 41460 115903
rect 41420 67992 41472 67998
rect 41420 67934 41472 67940
rect 41432 64666 41460 67934
rect 41420 64660 41472 64666
rect 41420 64602 41472 64608
rect 39856 52420 39908 52426
rect 39856 52362 39908 52368
rect 39868 47870 39896 52362
rect 39856 47864 39908 47870
rect 39856 47806 39908 47812
rect 39764 47728 39816 47734
rect 39764 47670 39816 47676
rect 42260 45694 42288 184826
rect 42352 173942 42380 184924
rect 42536 184890 42564 197338
rect 42628 195906 42656 238070
rect 42720 228070 42748 240586
rect 42904 228682 42932 245534
rect 42892 228676 42944 228682
rect 42892 228618 42944 228624
rect 42708 228064 42760 228070
rect 42708 228006 42760 228012
rect 42800 198688 42852 198694
rect 42800 198630 42852 198636
rect 42616 195900 42668 195906
rect 42616 195842 42668 195848
rect 42812 188358 42840 198630
rect 42800 188352 42852 188358
rect 42800 188294 42852 188300
rect 42524 184884 42576 184890
rect 42524 184826 42576 184832
rect 42340 173936 42392 173942
rect 42340 173878 42392 173884
rect 42892 173936 42944 173942
rect 42892 173878 42944 173884
rect 42904 160138 42932 173878
rect 42524 160132 42576 160138
rect 42524 160074 42576 160080
rect 42892 160132 42944 160138
rect 42892 160074 42944 160080
rect 42536 140826 42564 160074
rect 42340 140820 42392 140826
rect 42340 140762 42392 140768
rect 42524 140820 42576 140826
rect 42524 140762 42576 140768
rect 42352 131102 42380 140762
rect 42340 131096 42392 131102
rect 42340 131038 42392 131044
rect 44192 120193 44220 870023
rect 44284 458250 44312 922898
rect 44362 917280 44418 917289
rect 44362 917215 44418 917224
rect 44272 458244 44324 458250
rect 44272 458186 44324 458192
rect 44376 448633 44404 917215
rect 45834 877568 45890 877577
rect 45940 877554 45968 990218
rect 63420 990146 63448 990286
rect 77298 990247 77300 990256
rect 77352 990247 77354 990256
rect 77300 990218 77352 990224
rect 78876 990214 78904 990694
rect 79520 990622 79548 990762
rect 79508 990616 79560 990622
rect 79508 990558 79560 990564
rect 78864 990208 78916 990214
rect 78864 990150 78916 990156
rect 82648 990146 82676 992054
rect 90008 990690 90036 992054
rect 130304 990758 130332 995452
rect 130948 990826 130976 995452
rect 131577 995407 131633 995887
rect 132129 995407 132185 995887
rect 132773 995407 132829 995887
rect 133417 995407 133473 995887
rect 133969 995407 134025 995887
rect 134613 995407 134669 995887
rect 135352 995512 135404 995518
rect 135286 995460 135352 995466
rect 135286 995454 135404 995460
rect 135286 995438 135392 995454
rect 135901 995407 135957 995887
rect 136453 995407 136509 995887
rect 137097 995407 137153 995887
rect 137741 995407 137797 995887
rect 138937 995407 138993 995887
rect 140133 995407 140189 995887
rect 140777 995407 140833 995887
rect 130936 990820 130988 990826
rect 130936 990762 130988 990768
rect 131120 990820 131172 990826
rect 131120 990762 131172 990768
rect 130292 990752 130344 990758
rect 130292 990694 130344 990700
rect 89996 990684 90048 990690
rect 89996 990626 90048 990632
rect 130304 990622 130332 990694
rect 130292 990616 130344 990622
rect 130292 990558 130344 990564
rect 131132 990486 131160 990762
rect 141436 990690 141464 995452
rect 142617 995407 142673 995887
rect 143172 995512 143224 995518
rect 143224 995460 143290 995466
rect 143172 995454 143290 995460
rect 143184 995438 143290 995454
rect 179849 995407 179905 995887
rect 180493 995407 180549 995887
rect 181137 995407 181193 995887
rect 181717 995438 181760 995466
rect 182361 995438 182404 995466
rect 141424 990684 141476 990690
rect 141424 990626 141476 990632
rect 181732 990622 181760 995438
rect 182376 990758 182404 995438
rect 182977 995407 183033 995887
rect 183529 995407 183585 995887
rect 184173 995407 184229 995887
rect 184817 995407 184873 995887
rect 185369 995407 185425 995887
rect 186013 995407 186069 995887
rect 186685 995438 186728 995466
rect 186700 990826 186728 995438
rect 187301 995407 187357 995887
rect 187853 995407 187909 995887
rect 188497 995407 188553 995887
rect 189141 995407 189197 995887
rect 190337 995407 190393 995887
rect 191533 995407 191589 995887
rect 192177 995407 192233 995887
rect 192849 995438 192892 995466
rect 186688 990820 186740 990826
rect 186688 990762 186740 990768
rect 182364 990752 182416 990758
rect 182364 990694 182416 990700
rect 181720 990616 181772 990622
rect 181720 990558 181772 990564
rect 181732 990486 181760 990558
rect 182376 990554 182404 990694
rect 192864 990690 192892 995438
rect 194017 995407 194073 995887
rect 194689 995438 194732 995466
rect 194704 990826 194732 995438
rect 231249 995407 231305 995887
rect 231893 995407 231949 995887
rect 232537 995407 232593 995887
rect 233068 995438 233117 995466
rect 233620 995438 233761 995466
rect 233068 990826 233096 995438
rect 194692 990820 194744 990826
rect 194692 990762 194744 990768
rect 194784 990820 194836 990826
rect 194784 990762 194836 990768
rect 233056 990820 233108 990826
rect 233056 990762 233108 990768
rect 192852 990684 192904 990690
rect 192852 990626 192904 990632
rect 192864 990554 192892 990626
rect 182364 990548 182416 990554
rect 182364 990490 182416 990496
rect 192852 990548 192904 990554
rect 192852 990490 192904 990496
rect 194796 990486 194824 990762
rect 200028 990752 200080 990758
rect 200028 990694 200080 990700
rect 131120 990480 131172 990486
rect 132500 990480 132552 990486
rect 131120 990422 131172 990428
rect 132498 990448 132500 990457
rect 160008 990480 160060 990486
rect 132552 990448 132554 990457
rect 132498 990383 132554 990392
rect 140778 990448 140834 990457
rect 181720 990480 181772 990486
rect 160060 990428 160140 990434
rect 160008 990422 160140 990428
rect 181720 990422 181772 990428
rect 194784 990480 194836 990486
rect 194784 990422 194836 990428
rect 160020 990418 160140 990422
rect 160020 990412 160152 990418
rect 160020 990406 160100 990412
rect 140778 990383 140834 990392
rect 140792 990350 140820 990383
rect 160100 990354 160152 990360
rect 200040 990350 200068 990694
rect 233620 990690 233648 995438
rect 234377 995407 234433 995887
rect 234929 995407 234985 995887
rect 235573 995407 235629 995887
rect 236217 995407 236273 995887
rect 236769 995407 236825 995887
rect 237413 995407 237469 995887
rect 238208 995648 238260 995654
rect 238208 995590 238260 995596
rect 238220 995466 238248 995590
rect 238085 995438 238248 995466
rect 238701 995407 238757 995887
rect 239253 995407 239309 995887
rect 239897 995407 239953 995887
rect 240541 995407 240597 995887
rect 241737 995407 241793 995887
rect 242933 995407 242989 995887
rect 243577 995407 243633 995887
rect 244200 995438 244249 995466
rect 244200 990758 244228 995438
rect 245417 995407 245473 995887
rect 245936 995648 245988 995654
rect 245936 995590 245988 995596
rect 245948 995466 245976 995590
rect 245948 995438 246089 995466
rect 282849 995407 282905 995887
rect 283493 995407 283549 995887
rect 284137 995407 284193 995887
rect 284680 990826 284708 995452
rect 284668 990820 284720 990826
rect 284668 990762 284720 990768
rect 244188 990752 244240 990758
rect 244188 990694 244240 990700
rect 233608 990684 233660 990690
rect 233608 990626 233660 990632
rect 233620 990350 233648 990626
rect 244200 990554 244228 990694
rect 285324 990690 285352 995452
rect 285977 995407 286033 995887
rect 286529 995407 286585 995887
rect 287173 995407 287229 995887
rect 287817 995407 287873 995887
rect 288369 995407 288425 995887
rect 289013 995407 289069 995887
rect 289648 995314 289676 995452
rect 290301 995407 290357 995887
rect 290853 995407 290909 995887
rect 291497 995407 291553 995887
rect 292141 995407 292197 995887
rect 293337 995407 293393 995887
rect 294533 995407 294589 995887
rect 295177 995407 295233 995887
rect 289636 995308 289688 995314
rect 289636 995250 289688 995256
rect 295812 990758 295840 995452
rect 297017 995407 297073 995887
rect 297652 995314 297680 995452
rect 297640 995308 297692 995314
rect 297640 995250 297692 995256
rect 295800 990752 295852 990758
rect 295800 990694 295852 990700
rect 245568 990684 245620 990690
rect 245568 990626 245620 990632
rect 285312 990684 285364 990690
rect 285312 990626 285364 990632
rect 245580 990554 245608 990626
rect 285324 990554 285352 990626
rect 314476 990616 314528 990622
rect 314752 990616 314804 990622
rect 314528 990564 314752 990570
rect 314476 990558 314804 990564
rect 244188 990548 244240 990554
rect 244188 990490 244240 990496
rect 245568 990548 245620 990554
rect 245568 990490 245620 990496
rect 285312 990548 285364 990554
rect 314488 990542 314792 990558
rect 328460 990548 328512 990554
rect 285312 990490 285364 990496
rect 328564 990536 328592 997319
rect 347686 997112 347742 997121
rect 347686 997047 347742 997056
rect 347700 990554 347728 997047
rect 585704 996441 585732 997628
rect 672630 996568 672686 996577
rect 672630 996503 672686 996512
rect 585690 996432 585746 996441
rect 585690 996367 585746 996376
rect 672446 996432 672502 996441
rect 672446 996367 672502 996376
rect 384649 995407 384705 995887
rect 385293 995407 385349 995887
rect 385937 995407 385993 995887
rect 386524 990826 386552 995452
rect 386512 990820 386564 990826
rect 386512 990762 386564 990768
rect 386524 990622 386552 990762
rect 387168 990690 387196 995452
rect 387777 995407 387833 995887
rect 388329 995407 388385 995887
rect 388973 995407 389029 995887
rect 389617 995407 389673 995887
rect 390169 995407 390225 995887
rect 390813 995407 390869 995887
rect 391492 995314 391520 995452
rect 392101 995407 392157 995887
rect 392653 995407 392709 995887
rect 393297 995407 393353 995887
rect 393941 995407 393997 995887
rect 395137 995407 395193 995887
rect 396333 995407 396389 995887
rect 396977 995407 397033 995887
rect 397472 995438 397670 995466
rect 391480 995308 391532 995314
rect 391480 995250 391532 995256
rect 397472 990758 397500 995438
rect 398817 995407 398873 995887
rect 399496 995314 399524 995452
rect 473649 995407 473705 995887
rect 474293 995407 474349 995887
rect 474937 995407 474993 995887
rect 399484 995308 399536 995314
rect 399484 995250 399536 995256
rect 475488 990758 475516 995452
rect 397460 990752 397512 990758
rect 397460 990694 397512 990700
rect 474740 990752 474792 990758
rect 474740 990694 474792 990700
rect 475476 990752 475528 990758
rect 475476 990694 475528 990700
rect 387156 990684 387208 990690
rect 387156 990626 387208 990632
rect 386512 990616 386564 990622
rect 386512 990558 386564 990564
rect 397472 990554 397500 990694
rect 474752 990622 474780 990694
rect 476132 990690 476160 995452
rect 476777 995407 476833 995887
rect 477329 995407 477385 995887
rect 477973 995407 478029 995887
rect 478617 995407 478673 995887
rect 479169 995407 479225 995887
rect 479813 995407 479869 995887
rect 480456 995314 480484 995452
rect 481101 995407 481157 995887
rect 481653 995407 481709 995887
rect 482297 995407 482353 995887
rect 482941 995407 482997 995887
rect 484137 995407 484193 995887
rect 485333 995407 485389 995887
rect 485977 995407 486033 995887
rect 480444 995308 480496 995314
rect 480444 995250 480496 995256
rect 486620 990826 486648 995452
rect 487817 995407 487873 995887
rect 488460 995314 488488 995452
rect 525049 995407 525105 995887
rect 525693 995407 525749 995887
rect 526337 995407 526393 995887
rect 488448 995308 488500 995314
rect 488448 995250 488500 995256
rect 486608 990820 486660 990826
rect 486608 990762 486660 990768
rect 476120 990684 476172 990690
rect 476120 990626 476172 990632
rect 474740 990616 474792 990622
rect 474740 990558 474792 990564
rect 486620 990554 486648 990762
rect 526916 990758 526944 995452
rect 526904 990752 526956 990758
rect 526904 990694 526956 990700
rect 527560 990690 527588 995452
rect 528177 995407 528233 995887
rect 528729 995407 528785 995887
rect 529373 995407 529429 995887
rect 530017 995407 530073 995887
rect 530569 995407 530625 995887
rect 531213 995407 531269 995887
rect 531964 995648 532016 995654
rect 531964 995590 532016 995596
rect 531976 995466 532004 995590
rect 531898 995438 532004 995466
rect 532501 995407 532557 995887
rect 533053 995407 533109 995887
rect 533697 995407 533753 995887
rect 534341 995407 534397 995887
rect 535537 995407 535593 995887
rect 536733 995407 536789 995887
rect 537377 995407 537433 995887
rect 538048 990826 538076 995452
rect 539217 995407 539273 995887
rect 539692 995648 539744 995654
rect 539692 995590 539744 995596
rect 539704 995466 539732 995590
rect 539704 995438 539902 995466
rect 626849 995407 626905 995887
rect 627493 995407 627549 995887
rect 628137 995407 628193 995887
rect 628668 995438 628717 995466
rect 629312 995438 629361 995466
rect 538036 990820 538088 990826
rect 538036 990762 538088 990768
rect 626540 990752 626592 990758
rect 626540 990694 626592 990700
rect 527548 990684 527600 990690
rect 527548 990626 527600 990632
rect 328512 990508 328592 990536
rect 347688 990548 347740 990554
rect 328460 990490 328512 990496
rect 347688 990490 347740 990496
rect 397460 990548 397512 990554
rect 397460 990490 397512 990496
rect 486608 990548 486660 990554
rect 486608 990490 486660 990496
rect 328196 990406 328408 990434
rect 140780 990344 140832 990350
rect 82910 990312 82966 990321
rect 121380 990282 121500 990298
rect 140780 990286 140832 990292
rect 200028 990344 200080 990350
rect 200028 990286 200080 990292
rect 233608 990344 233660 990350
rect 233608 990286 233660 990292
rect 275836 990344 275888 990350
rect 275836 990286 275888 990292
rect 289728 990344 289780 990350
rect 289728 990286 289780 990292
rect 82910 990247 82966 990256
rect 121368 990276 121512 990282
rect 82924 990214 82952 990247
rect 121420 990270 121460 990276
rect 121368 990218 121420 990224
rect 121460 990218 121512 990224
rect 82912 990208 82964 990214
rect 198740 990208 198792 990214
rect 82912 990150 82964 990156
rect 160020 990146 160140 990162
rect 179248 990146 179552 990162
rect 198660 990156 198740 990162
rect 231860 990208 231912 990214
rect 198660 990150 198792 990156
rect 231780 990156 231860 990162
rect 231780 990150 231912 990156
rect 256608 990208 256660 990214
rect 256792 990208 256844 990214
rect 256660 990156 256792 990162
rect 256608 990150 256844 990156
rect 198660 990146 198780 990150
rect 231780 990146 231900 990150
rect 63408 990140 63460 990146
rect 63408 990082 63460 990088
rect 82636 990140 82688 990146
rect 82636 990082 82688 990088
rect 160008 990140 160152 990146
rect 160060 990134 160100 990140
rect 160008 990082 160060 990088
rect 160100 990082 160152 990088
rect 179236 990140 179564 990146
rect 179288 990134 179512 990140
rect 179236 990082 179288 990088
rect 179512 990082 179564 990088
rect 198648 990140 198780 990146
rect 198700 990134 198780 990140
rect 231768 990140 231900 990146
rect 198648 990082 198700 990088
rect 231820 990134 231900 990140
rect 256620 990134 256832 990150
rect 275848 990146 275876 990286
rect 289740 990146 289768 990286
rect 328196 990146 328224 990406
rect 328380 990350 328408 990406
rect 328368 990344 328420 990350
rect 328368 990286 328420 990292
rect 328458 990312 328514 990321
rect 328458 990247 328460 990256
rect 328512 990247 328514 990256
rect 328460 990218 328512 990224
rect 626552 990146 626580 990694
rect 628668 990146 628696 995438
rect 629312 990690 629340 995438
rect 629977 995407 630033 995887
rect 630529 995407 630585 995887
rect 631173 995407 631229 995887
rect 631817 995407 631873 995887
rect 632369 995407 632425 995887
rect 633013 995407 633069 995887
rect 633808 995512 633860 995518
rect 633685 995460 633808 995466
rect 633685 995454 633860 995460
rect 633685 995438 633848 995454
rect 634301 995407 634357 995887
rect 634853 995407 634909 995887
rect 635497 995407 635553 995887
rect 636141 995407 636197 995887
rect 637337 995407 637393 995887
rect 638533 995407 638589 995887
rect 639177 995407 639233 995887
rect 639800 995438 639849 995466
rect 639800 990826 639828 995438
rect 641017 995407 641073 995887
rect 641536 995512 641588 995518
rect 641588 995460 641689 995466
rect 641536 995454 641689 995460
rect 641548 995438 641689 995454
rect 639788 990820 639840 990826
rect 639788 990762 639840 990768
rect 629300 990684 629352 990690
rect 629300 990626 629352 990632
rect 630956 990684 631008 990690
rect 630956 990626 631008 990632
rect 630968 990146 630996 990626
rect 639800 990214 639828 990762
rect 639788 990208 639840 990214
rect 639788 990150 639840 990156
rect 275836 990140 275888 990146
rect 231768 990082 231820 990088
rect 275836 990082 275888 990088
rect 289728 990140 289780 990146
rect 289728 990082 289780 990088
rect 328184 990140 328236 990146
rect 328184 990082 328236 990088
rect 626540 990140 626592 990146
rect 626540 990082 626592 990088
rect 628656 990140 628708 990146
rect 628656 990082 628708 990088
rect 630956 990140 631008 990146
rect 630956 990082 631008 990088
rect 45890 877526 45968 877554
rect 45834 877503 45890 877512
rect 44638 835272 44694 835281
rect 44638 835207 44694 835216
rect 44454 828064 44510 828073
rect 44454 827999 44510 828008
rect 44468 488617 44496 827999
rect 44652 493241 44680 835207
rect 672460 828730 672488 996367
rect 672538 828744 672594 828753
rect 672460 828702 672538 828730
rect 672460 823698 672488 828702
rect 672538 828679 672594 828688
rect 672644 826169 672672 996503
rect 673552 990208 673604 990214
rect 673552 990150 673604 990156
rect 673460 990072 673512 990078
rect 673460 990014 673512 990020
rect 673472 965326 673500 990014
rect 673460 965320 673512 965326
rect 673460 965262 673512 965268
rect 673366 908168 673422 908177
rect 673366 908103 673422 908112
rect 672630 826160 672686 826169
rect 672630 826095 672686 826104
rect 673274 826160 673330 826169
rect 673274 826095 673330 826104
rect 672538 823712 672594 823721
rect 672460 823670 672538 823698
rect 672538 823647 672594 823656
rect 673182 823712 673238 823721
rect 673182 823647 673238 823656
rect 673196 816898 673224 823647
rect 673104 816870 673224 816898
rect 673104 811442 673132 816870
rect 672816 811436 672868 811442
rect 672816 811378 672868 811384
rect 673092 811436 673144 811442
rect 673092 811378 673144 811384
rect 672828 792169 672856 811378
rect 672814 792160 672870 792169
rect 672814 792095 672870 792104
rect 672998 792160 673054 792169
rect 672998 792095 673054 792104
rect 673012 778394 673040 792095
rect 673000 778388 673052 778394
rect 673000 778330 673052 778336
rect 673184 778320 673236 778326
rect 673184 778262 673236 778268
rect 673196 772834 673224 778262
rect 673104 772818 673224 772834
rect 673092 772812 673236 772818
rect 673144 772806 673184 772812
rect 673092 772754 673144 772760
rect 673184 772754 673236 772760
rect 673104 772723 673132 772754
rect 673196 739770 673224 772754
rect 673184 739764 673236 739770
rect 673184 739706 673236 739712
rect 673092 739560 673144 739566
rect 673092 739502 673144 739508
rect 673104 721449 673132 739502
rect 673090 721440 673146 721449
rect 673090 721375 673146 721384
rect 672998 714912 673054 714921
rect 672998 714847 673054 714856
rect 673012 712094 673040 714847
rect 672816 712088 672868 712094
rect 672816 712030 672868 712036
rect 673000 712088 673052 712094
rect 673000 712030 673052 712036
rect 672828 692850 672856 712030
rect 672816 692844 672868 692850
rect 672816 692786 672868 692792
rect 673184 692844 673236 692850
rect 673184 692786 673236 692792
rect 673196 681714 673224 692786
rect 673012 681686 673224 681714
rect 673012 676190 673040 681686
rect 673000 676184 673052 676190
rect 673000 676126 673052 676132
rect 673092 676184 673144 676190
rect 673092 676126 673144 676132
rect 673104 656946 673132 676126
rect 673092 656940 673144 656946
rect 673092 656882 673144 656888
rect 673184 656940 673236 656946
rect 673184 656882 673236 656888
rect 673196 643090 673224 656882
rect 673104 643062 673224 643090
rect 673104 637566 673132 643062
rect 672816 637560 672868 637566
rect 672816 637502 672868 637508
rect 673092 637560 673144 637566
rect 673092 637502 673144 637508
rect 672828 618322 672856 637502
rect 672816 618316 672868 618322
rect 672816 618258 672868 618264
rect 673000 618316 673052 618322
rect 673000 618258 673052 618264
rect 673012 605878 673040 618258
rect 672816 605872 672868 605878
rect 672816 605814 672868 605820
rect 673000 605872 673052 605878
rect 673000 605814 673052 605820
rect 672828 596222 672856 605814
rect 672816 596216 672868 596222
rect 672816 596158 672868 596164
rect 673000 596216 673052 596222
rect 673000 596158 673052 596164
rect 673012 596086 673040 596158
rect 672816 596080 672868 596086
rect 672816 596022 672868 596028
rect 673000 596080 673052 596086
rect 673000 596022 673052 596028
rect 672828 585138 672856 596022
rect 672816 585132 672868 585138
rect 672816 585074 672868 585080
rect 673000 585132 673052 585138
rect 673000 585074 673052 585080
rect 673012 576858 673040 585074
rect 673012 576830 673132 576858
rect 673104 538286 673132 576830
rect 672908 538280 672960 538286
rect 672908 538222 672960 538228
rect 673092 538280 673144 538286
rect 673092 538222 673144 538228
rect 672920 527066 672948 538222
rect 672908 527060 672960 527066
rect 672908 527002 672960 527008
rect 673184 527060 673236 527066
rect 673184 527002 673236 527008
rect 673196 514185 673224 527002
rect 672998 514176 673054 514185
rect 672998 514111 673054 514120
rect 673182 514176 673238 514185
rect 673182 514111 673238 514120
rect 673012 509153 673040 514111
rect 673288 511465 673316 826095
rect 673090 511456 673146 511465
rect 673090 511391 673146 511400
rect 673274 511456 673330 511465
rect 673274 511391 673330 511400
rect 672998 509144 673054 509153
rect 672998 509079 673054 509088
rect 673012 499594 673040 509079
rect 673000 499588 673052 499594
rect 673000 499530 673052 499536
rect 44638 493232 44694 493241
rect 44638 493167 44694 493176
rect 44454 488608 44510 488617
rect 44454 488543 44510 488552
rect 673000 482996 673052 483002
rect 673000 482938 673052 482944
rect 673012 463729 673040 482938
rect 672998 463720 673054 463729
rect 672998 463655 673054 463664
rect 44362 448624 44418 448633
rect 44362 448559 44418 448568
rect 673104 427961 673132 511391
rect 673276 499588 673328 499594
rect 673276 499530 673328 499536
rect 673288 483002 673316 499530
rect 673276 482996 673328 483002
rect 673276 482938 673328 482944
rect 673380 467537 673408 908103
rect 673472 876178 673500 965262
rect 673564 953358 673592 990150
rect 673644 990140 673696 990146
rect 673644 990082 673696 990088
rect 673656 964782 673684 990082
rect 675407 966695 675887 966751
rect 675407 966051 675887 966107
rect 675407 965407 675887 965463
rect 675392 965320 675444 965326
rect 675392 965262 675444 965268
rect 675404 964883 675432 965262
rect 673644 964776 673696 964782
rect 673644 964718 673696 964724
rect 675392 964776 675444 964782
rect 675392 964718 675444 964724
rect 673552 953352 673604 953358
rect 673552 953294 673604 953300
rect 673460 876172 673512 876178
rect 673460 876114 673512 876120
rect 673564 865026 673592 953294
rect 673656 910790 673684 964718
rect 675404 964239 675432 964718
rect 675407 963567 675887 963623
rect 675407 963015 675887 963071
rect 675407 962371 675887 962427
rect 675407 961727 675887 961783
rect 675407 961175 675887 961231
rect 675407 960531 675887 960587
rect 675312 959901 675418 959929
rect 675312 951810 675340 959901
rect 675407 959243 675887 959299
rect 675407 958691 675887 958747
rect 675407 958047 675887 958103
rect 675407 957403 675887 957459
rect 675407 956207 675887 956263
rect 675407 955011 675887 955067
rect 675407 954367 675887 954423
rect 675404 953358 675432 953751
rect 675392 953352 675444 953358
rect 675392 953294 675444 953300
rect 675407 952527 675887 952583
rect 675404 951810 675432 951932
rect 675312 951782 675432 951810
rect 677874 918640 677930 918649
rect 677930 918598 678086 918626
rect 677874 918575 677930 918584
rect 677598 915376 677654 915385
rect 677598 915311 677654 915320
rect 677612 912801 677640 915311
rect 677796 913974 678046 914002
rect 677598 912792 677654 912801
rect 677598 912727 677654 912736
rect 677796 910790 677824 913974
rect 678018 913716 678046 913974
rect 677874 912792 677930 912801
rect 677874 912727 677930 912736
rect 673644 910784 673696 910790
rect 673644 910726 673696 910732
rect 677784 910784 677836 910790
rect 677784 910726 677836 910732
rect 673656 875566 673684 910726
rect 677888 908177 677916 912727
rect 677874 908168 677930 908177
rect 677874 908103 677930 908112
rect 677782 907760 677838 907769
rect 677838 907718 678086 907746
rect 677782 907695 677838 907704
rect 675407 877495 675887 877551
rect 675407 876851 675887 876907
rect 675407 876207 675887 876263
rect 675392 876172 675444 876178
rect 675392 876114 675444 876120
rect 675404 875697 675432 876114
rect 675312 875683 675432 875697
rect 675312 875669 675418 875683
rect 673644 875560 673696 875566
rect 673644 875502 673696 875508
rect 675208 870188 675260 870194
rect 675208 870130 675260 870136
rect 673552 865020 673604 865026
rect 673552 864962 673604 864968
rect 673460 785324 673512 785330
rect 673460 785266 673512 785272
rect 673472 741402 673500 785266
rect 673564 774926 673592 864962
rect 674656 862844 674708 862850
rect 674656 862786 674708 862792
rect 674668 850610 674696 862786
rect 675220 862730 675248 870130
rect 675312 862850 675340 875669
rect 675392 875560 675444 875566
rect 675392 875502 675444 875508
rect 675404 875039 675432 875502
rect 675407 874367 675887 874423
rect 675407 873815 675887 873871
rect 675407 873171 675887 873227
rect 675407 872527 675887 872583
rect 675407 871975 675887 872031
rect 675407 871331 675887 871387
rect 675404 870194 675432 870740
rect 675392 870188 675444 870194
rect 675392 870130 675444 870136
rect 675407 870043 675887 870099
rect 675407 869491 675887 869547
rect 675407 868847 675887 868903
rect 675407 868203 675887 868259
rect 675407 867007 675887 867063
rect 675407 865811 675887 865867
rect 675407 865167 675887 865223
rect 675392 865020 675444 865026
rect 675392 864962 675444 864968
rect 675404 864551 675432 864962
rect 675407 863327 675887 863383
rect 675300 862844 675352 862850
rect 675300 862786 675352 862792
rect 675220 862702 675418 862730
rect 673920 850604 673972 850610
rect 673920 850546 673972 850552
rect 674656 850604 674708 850610
rect 674656 850546 674708 850552
rect 673932 850105 673960 850546
rect 673734 850096 673790 850105
rect 673734 850031 673790 850040
rect 673918 850096 673974 850105
rect 673918 850031 673974 850040
rect 673748 830822 673776 850031
rect 673736 830816 673788 830822
rect 673736 830758 673788 830764
rect 674012 830816 674064 830822
rect 674012 830758 674064 830764
rect 674024 817018 674052 830758
rect 673828 817012 673880 817018
rect 673828 816954 673880 816960
rect 674012 817012 674064 817018
rect 674012 816954 674064 816960
rect 673840 797722 673868 816954
rect 673840 797694 674052 797722
rect 674024 797638 674052 797694
rect 674012 797632 674064 797638
rect 674012 797574 674064 797580
rect 675300 797632 675352 797638
rect 675300 797574 675352 797580
rect 675312 786497 675340 797574
rect 675407 788295 675887 788351
rect 675407 787651 675887 787707
rect 675407 787007 675887 787063
rect 675220 786469 675418 786497
rect 673552 774920 673604 774926
rect 673552 774862 673604 774868
rect 673460 741396 673512 741402
rect 673460 741338 673512 741344
rect 673460 736636 673512 736642
rect 673460 736578 673512 736584
rect 673472 710734 673500 736578
rect 673564 730182 673592 774862
rect 675220 772857 675248 786469
rect 675404 785330 675432 785839
rect 675392 785324 675444 785330
rect 675392 785266 675444 785272
rect 675407 785167 675887 785223
rect 675407 784615 675887 784671
rect 675407 783971 675887 784027
rect 675407 783327 675887 783383
rect 675407 782775 675887 782831
rect 675407 782131 675887 782187
rect 675312 781510 675418 781538
rect 675312 773514 675340 781510
rect 675407 780843 675887 780899
rect 675407 780291 675887 780347
rect 675407 779647 675887 779703
rect 675407 779003 675887 779059
rect 675407 777807 675887 777863
rect 675407 776611 675887 776667
rect 675407 775967 675887 776023
rect 675404 774926 675432 775351
rect 675392 774920 675444 774926
rect 675392 774862 675444 774868
rect 675407 774127 675887 774183
rect 675312 773486 675418 773514
rect 673826 772848 673882 772857
rect 673826 772783 673882 772792
rect 675206 772848 675262 772857
rect 675206 772783 675262 772792
rect 673840 741946 673868 772783
rect 675407 743295 675887 743351
rect 675407 742651 675887 742707
rect 675407 742007 675887 742063
rect 673828 741940 673880 741946
rect 673828 741882 673880 741888
rect 675392 741940 675444 741946
rect 675392 741882 675444 741888
rect 673552 730176 673604 730182
rect 673552 730118 673604 730124
rect 673736 720384 673788 720390
rect 673736 720326 673788 720332
rect 673460 710728 673512 710734
rect 673460 710670 673512 710676
rect 673644 701072 673696 701078
rect 673644 701014 673696 701020
rect 673656 695978 673684 701014
rect 673644 695972 673696 695978
rect 673644 695914 673696 695920
rect 673748 685409 673776 720326
rect 673840 701146 673868 741882
rect 675404 741483 675432 741882
rect 675392 741396 675444 741402
rect 675392 741338 675444 741344
rect 675404 740874 675432 741338
rect 675312 740860 675432 740874
rect 675312 740846 675418 740860
rect 675312 736642 675340 740846
rect 675407 740167 675887 740223
rect 675407 739615 675887 739671
rect 675407 738971 675887 739027
rect 675407 738327 675887 738383
rect 675407 737775 675887 737831
rect 675407 737131 675887 737187
rect 675300 736636 675352 736642
rect 675300 736578 675352 736584
rect 675312 736494 675418 736522
rect 673920 730176 673972 730182
rect 673920 730118 673972 730124
rect 673932 720390 673960 730118
rect 675312 729042 675340 736494
rect 675407 735843 675887 735899
rect 675407 735291 675887 735347
rect 675407 734647 675887 734703
rect 675407 734003 675887 734059
rect 675407 732807 675887 732863
rect 675407 731611 675887 731667
rect 675407 730967 675887 731023
rect 675404 730182 675432 730351
rect 675392 730176 675444 730182
rect 675392 730118 675444 730124
rect 675407 729127 675887 729183
rect 675312 729014 675432 729042
rect 675404 728484 675432 729014
rect 673920 720384 673972 720390
rect 673920 720326 673972 720332
rect 675300 710728 675352 710734
rect 675300 710670 675352 710676
rect 673828 701140 673880 701146
rect 673828 701082 673880 701088
rect 673828 695972 673880 695978
rect 673828 695914 673880 695920
rect 673734 685400 673790 685409
rect 673734 685335 673790 685344
rect 673460 681760 673512 681766
rect 673512 681708 673684 681714
rect 673460 681702 673684 681708
rect 673472 681686 673684 681702
rect 673656 676190 673684 681686
rect 673644 676184 673696 676190
rect 673644 676126 673696 676132
rect 673552 656940 673604 656946
rect 673552 656882 673604 656888
rect 673460 651772 673512 651778
rect 673460 651714 673512 651720
rect 673472 606762 673500 651714
rect 673564 651166 673592 656882
rect 673552 651160 673604 651166
rect 673552 651102 673604 651108
rect 673748 639742 673776 685335
rect 673840 651778 673868 695914
rect 675312 695858 675340 710670
rect 675407 698295 675887 698351
rect 675407 697651 675887 697707
rect 675407 697007 675887 697063
rect 675404 695978 675432 696483
rect 675392 695972 675444 695978
rect 675392 695914 675444 695920
rect 675312 695844 675418 695858
rect 675312 695830 675432 695844
rect 675404 695314 675432 695830
rect 675220 695286 675432 695314
rect 675220 681766 675248 695286
rect 675407 695167 675887 695223
rect 675407 694615 675887 694671
rect 675407 693971 675887 694027
rect 675407 693327 675887 693383
rect 675407 692775 675887 692831
rect 675407 692131 675887 692187
rect 675312 691614 675432 691642
rect 675312 683525 675340 691614
rect 675404 691492 675432 691614
rect 675407 690843 675887 690899
rect 675407 690291 675887 690347
rect 675407 689647 675887 689703
rect 675407 689003 675887 689059
rect 675407 687807 675887 687863
rect 675407 686611 675887 686667
rect 675407 685967 675887 686023
rect 675390 685400 675446 685409
rect 675390 685335 675446 685344
rect 675407 684127 675887 684183
rect 675312 683497 675418 683525
rect 675208 681760 675260 681766
rect 675208 681702 675260 681708
rect 673920 676184 673972 676190
rect 673920 676126 673972 676132
rect 673932 656946 673960 676126
rect 673920 656940 673972 656946
rect 673920 656882 673972 656888
rect 675407 653095 675887 653151
rect 675407 652451 675887 652507
rect 675407 651807 675887 651863
rect 673828 651772 673880 651778
rect 673828 651714 673880 651720
rect 675392 651772 675444 651778
rect 675392 651714 675444 651720
rect 675404 651283 675432 651714
rect 673828 651160 673880 651166
rect 673828 651102 673880 651108
rect 675392 651160 675444 651166
rect 675392 651102 675444 651108
rect 673840 643090 673868 651102
rect 675404 650639 675432 651102
rect 675407 649967 675887 650023
rect 675407 649415 675887 649471
rect 675407 648771 675887 648827
rect 675407 648127 675887 648183
rect 675407 647575 675887 647631
rect 675407 646931 675887 646987
rect 675404 645810 675432 646340
rect 675312 645782 675432 645810
rect 673840 643062 674052 643090
rect 673552 639736 673604 639742
rect 673552 639678 673604 639684
rect 673736 639736 673788 639742
rect 673736 639678 673788 639684
rect 673460 606756 673512 606762
rect 673460 606698 673512 606704
rect 673564 594930 673592 639678
rect 674024 637566 674052 643062
rect 675312 638330 675340 645782
rect 675407 645643 675887 645699
rect 675407 645091 675887 645147
rect 675407 644447 675887 644503
rect 675407 643803 675887 643859
rect 675407 642607 675887 642663
rect 675407 641411 675887 641467
rect 675407 640767 675887 640823
rect 675404 639742 675432 640151
rect 675392 639736 675444 639742
rect 675392 639678 675444 639684
rect 675407 638927 675887 638983
rect 675312 638302 675418 638330
rect 673736 637560 673788 637566
rect 673736 637502 673788 637508
rect 674012 637560 674064 637566
rect 674012 637502 674064 637508
rect 673748 618322 673776 637502
rect 673736 618316 673788 618322
rect 673736 618258 673788 618264
rect 673920 618316 673972 618322
rect 673920 618258 673972 618264
rect 673828 606756 673880 606762
rect 673828 606698 673880 606704
rect 673644 604512 673696 604518
rect 673644 604454 673696 604460
rect 673552 594924 673604 594930
rect 673552 594866 673604 594872
rect 673460 559972 673512 559978
rect 673460 559914 673512 559920
rect 673366 467528 673422 467537
rect 673366 467463 673422 467472
rect 673274 463720 673330 463729
rect 673472 463690 673500 559914
rect 673564 550526 673592 594866
rect 673656 559978 673684 604454
rect 673840 561542 673868 606698
rect 673932 605674 673960 618258
rect 675407 608095 675887 608151
rect 675407 607451 675887 607507
rect 675407 606807 675887 606863
rect 675392 606756 675444 606762
rect 675392 606698 675444 606704
rect 675404 606283 675432 606698
rect 673920 605668 673972 605674
rect 673920 605610 673972 605616
rect 675300 605668 675352 605674
rect 675352 605625 675418 605653
rect 675300 605610 675352 605616
rect 673932 604518 673960 605610
rect 675407 604967 675887 605023
rect 673920 604512 673972 604518
rect 673920 604454 673972 604460
rect 675407 604415 675887 604471
rect 675407 603771 675887 603827
rect 675407 603127 675887 603183
rect 675407 602575 675887 602631
rect 675407 601931 675887 601987
rect 675312 601310 675418 601338
rect 675312 593314 675340 601310
rect 675407 600643 675887 600699
rect 675407 600091 675887 600147
rect 675407 599447 675887 599503
rect 675407 598803 675887 598859
rect 675407 597607 675887 597663
rect 675407 596411 675887 596467
rect 675407 595767 675887 595823
rect 675404 594930 675432 595151
rect 675392 594924 675444 594930
rect 675392 594866 675444 594872
rect 675407 593927 675887 593983
rect 675312 593286 675418 593314
rect 675407 562895 675887 562951
rect 675407 562251 675887 562307
rect 675407 561607 675887 561663
rect 673828 561536 673880 561542
rect 673828 561478 673880 561484
rect 675392 561536 675444 561542
rect 675392 561478 675444 561484
rect 675404 561068 675432 561478
rect 675404 559978 675432 560439
rect 673644 559972 673696 559978
rect 673644 559914 673696 559920
rect 675392 559972 675444 559978
rect 675392 559914 675444 559920
rect 675407 559767 675887 559823
rect 675407 559215 675887 559271
rect 675407 558571 675887 558627
rect 675407 557927 675887 557983
rect 675407 557375 675887 557431
rect 675407 556731 675887 556787
rect 675312 556101 675418 556129
rect 673552 550520 673604 550526
rect 673552 550462 673604 550468
rect 675312 548125 675340 556101
rect 675407 555443 675887 555499
rect 675407 554891 675887 554947
rect 675407 554247 675887 554303
rect 675407 553603 675887 553659
rect 675407 552407 675887 552463
rect 675407 551211 675887 551267
rect 675407 550567 675887 550623
rect 675392 550520 675444 550526
rect 675392 550462 675444 550468
rect 675404 549951 675432 550462
rect 675407 548727 675887 548783
rect 675312 548097 675418 548125
rect 678058 480176 678114 480185
rect 678058 480111 678114 480120
rect 678072 470778 678100 480111
rect 677888 470764 678100 470778
rect 677888 470750 678086 470764
rect 677888 469985 677916 470750
rect 677874 469976 677930 469985
rect 677874 469911 677930 469920
rect 677704 465990 678032 466018
rect 677704 463690 677732 465990
rect 673274 463655 673330 463664
rect 673460 463684 673512 463690
rect 673288 449970 673316 463655
rect 673460 463626 673512 463632
rect 677692 463684 677744 463690
rect 677692 463626 677744 463632
rect 673288 449942 673408 449970
rect 673090 427952 673146 427961
rect 673090 427887 673146 427896
rect 673380 420889 673408 449942
rect 673366 420880 673422 420889
rect 673366 420815 673422 420824
rect 672816 412548 672868 412554
rect 672816 412490 672868 412496
rect 672828 411210 672856 412490
rect 672736 411182 672856 411210
rect 672736 392057 672764 411182
rect 672722 392048 672778 392057
rect 672722 391983 672778 391992
rect 672722 386472 672778 386481
rect 672722 386407 672778 386416
rect 672736 386374 672764 386407
rect 672724 386368 672776 386374
rect 672724 386310 672776 386316
rect 672908 386368 672960 386374
rect 672908 386310 672960 386316
rect 672920 372450 672948 386310
rect 673472 382634 673500 463626
rect 677704 459870 678086 459898
rect 677704 440230 677732 459870
rect 676220 440224 676272 440230
rect 676220 440166 676272 440172
rect 677692 440224 677744 440230
rect 677692 440166 677744 440172
rect 676232 412554 676260 440166
rect 677414 427952 677470 427961
rect 677414 427887 677470 427896
rect 677428 425762 677456 427887
rect 677598 425776 677654 425785
rect 677428 425734 677598 425762
rect 677598 425711 677654 425720
rect 676220 412548 676272 412554
rect 676220 412490 676272 412496
rect 675407 385695 675887 385751
rect 675407 385051 675887 385107
rect 675407 384407 675887 384463
rect 673552 384056 673604 384062
rect 673552 383998 673604 384004
rect 675392 384056 675444 384062
rect 675392 383998 675444 384004
rect 673460 382628 673512 382634
rect 673460 382570 673512 382576
rect 672736 372422 672948 372450
rect 672736 353394 672764 372422
rect 672724 353388 672776 353394
rect 672724 353330 672776 353336
rect 672724 353252 672776 353258
rect 672724 353194 672776 353200
rect 672736 347750 672764 353194
rect 672724 347744 672776 347750
rect 672724 347686 672776 347692
rect 672908 347744 672960 347750
rect 672908 347686 672960 347692
rect 672920 328506 672948 347686
rect 673564 338745 673592 383998
rect 675404 383860 675432 383998
rect 675312 383225 675418 383253
rect 675312 382634 675340 383225
rect 673644 382628 673696 382634
rect 673644 382570 673696 382576
rect 675300 382628 675352 382634
rect 675300 382570 675352 382576
rect 673550 338736 673606 338745
rect 673550 338671 673606 338680
rect 673460 338564 673512 338570
rect 673460 338506 673512 338512
rect 672540 328500 672592 328506
rect 672540 328442 672592 328448
rect 672908 328500 672960 328506
rect 672908 328442 672960 328448
rect 672552 316062 672580 328442
rect 672540 316056 672592 316062
rect 672540 315998 672592 316004
rect 672724 316056 672776 316062
rect 672724 315998 672776 316004
rect 672736 306406 672764 315998
rect 672448 306400 672500 306406
rect 672448 306342 672500 306348
rect 672724 306400 672776 306406
rect 672724 306342 672776 306348
rect 672460 295474 672488 306342
rect 672538 295488 672594 295497
rect 672460 295446 672538 295474
rect 672538 295423 672594 295432
rect 672630 295216 672686 295225
rect 672630 295151 672686 295160
rect 672644 276078 672672 295151
rect 673472 293049 673500 338506
rect 673564 293622 673592 338671
rect 673656 338570 673684 382570
rect 675407 382567 675887 382623
rect 675407 382015 675887 382071
rect 675407 381371 675887 381427
rect 675407 380727 675887 380783
rect 675407 380175 675887 380231
rect 675407 379531 675887 379587
rect 675312 378901 675418 378929
rect 673920 372360 673972 372366
rect 673920 372302 673972 372308
rect 673644 338564 673696 338570
rect 673644 338506 673696 338512
rect 673932 334098 673960 372302
rect 675312 370925 675340 378901
rect 675407 378243 675887 378299
rect 675407 377691 675887 377747
rect 675407 377047 675887 377103
rect 675407 376403 675887 376459
rect 675407 375207 675887 375263
rect 675407 373367 675887 373423
rect 675404 372366 675432 372751
rect 675392 372360 675444 372366
rect 675392 372302 675444 372308
rect 675407 371527 675887 371583
rect 675312 370897 675418 370925
rect 675407 340495 675887 340551
rect 675407 339851 675887 339907
rect 675407 339207 675887 339263
rect 675390 338736 675446 338745
rect 675390 338671 675446 338680
rect 675392 338564 675444 338570
rect 675392 338506 675444 338512
rect 675404 338028 675432 338506
rect 675407 337367 675887 337423
rect 675407 336815 675887 336871
rect 675407 336171 675887 336227
rect 675407 335527 675887 335583
rect 675407 334975 675887 335031
rect 675407 334331 675887 334387
rect 673840 334070 673960 334098
rect 673840 327146 673868 334070
rect 675312 333701 675418 333729
rect 673828 327140 673880 327146
rect 673828 327082 673880 327088
rect 673840 314650 673868 327082
rect 675312 325725 675340 333701
rect 675407 333043 675887 333099
rect 675407 332491 675887 332547
rect 675407 331847 675887 331903
rect 675407 331203 675887 331259
rect 675407 330007 675887 330063
rect 675407 328167 675887 328223
rect 675404 327146 675432 327556
rect 675392 327140 675444 327146
rect 675392 327082 675444 327088
rect 675407 326327 675887 326383
rect 675312 325697 675418 325725
rect 673748 314622 673868 314650
rect 673748 295338 673776 314622
rect 675407 295495 675887 295551
rect 673656 295310 673776 295338
rect 673552 293616 673604 293622
rect 673552 293558 673604 293564
rect 673458 293040 673514 293049
rect 673458 292975 673514 292984
rect 672632 276072 672684 276078
rect 672632 276014 672684 276020
rect 672540 276004 672592 276010
rect 672540 275946 672592 275952
rect 672552 260846 672580 275946
rect 672540 260840 672592 260846
rect 672540 260782 672592 260788
rect 672908 260840 672960 260846
rect 672908 260782 672960 260788
rect 672920 251258 672948 260782
rect 672724 251252 672776 251258
rect 672724 251194 672776 251200
rect 672908 251252 672960 251258
rect 672908 251194 672960 251200
rect 672736 251122 672764 251194
rect 672540 251116 672592 251122
rect 672540 251058 672592 251064
rect 672724 251116 672776 251122
rect 672724 251058 672776 251064
rect 672552 218090 672580 251058
rect 673472 247518 673500 292975
rect 673564 248198 673592 293558
rect 673656 283082 673684 295310
rect 675407 294851 675887 294907
rect 675407 294207 675887 294263
rect 675404 293622 675432 293692
rect 675392 293616 675444 293622
rect 675392 293558 675444 293564
rect 675390 293040 675446 293049
rect 675390 292975 675446 292984
rect 675407 292367 675887 292423
rect 675407 291815 675887 291871
rect 675407 291171 675887 291227
rect 675407 290527 675887 290583
rect 675407 289975 675887 290031
rect 675407 289331 675887 289387
rect 675312 288701 675418 288729
rect 673644 283076 673696 283082
rect 673644 283018 673696 283024
rect 673656 256698 673684 283018
rect 675312 280725 675340 288701
rect 675407 288043 675887 288099
rect 675407 287491 675887 287547
rect 675407 286847 675887 286903
rect 675407 286203 675887 286259
rect 675407 285007 675887 285063
rect 675407 283167 675887 283223
rect 675392 283076 675444 283082
rect 675392 283018 675444 283024
rect 675404 282540 675432 283018
rect 675407 281327 675887 281383
rect 675312 280697 675418 280725
rect 673644 256692 673696 256698
rect 673644 256634 673696 256640
rect 674012 256692 674064 256698
rect 674012 256634 674064 256640
rect 673552 248192 673604 248198
rect 673552 248134 673604 248140
rect 673460 247512 673512 247518
rect 673460 247454 673512 247460
rect 672552 218062 672672 218090
rect 672644 198778 672672 218062
rect 673564 206786 673592 248134
rect 673736 247512 673788 247518
rect 673736 247454 673788 247460
rect 673552 206780 673604 206786
rect 673552 206722 673604 206728
rect 673564 198778 673592 206722
rect 673748 202978 673776 247454
rect 674024 237794 674052 256634
rect 675407 250495 675887 250551
rect 675407 249851 675887 249907
rect 675407 249207 675887 249263
rect 675404 248198 675432 248676
rect 675392 248192 675444 248198
rect 675392 248134 675444 248140
rect 675404 247518 675432 248039
rect 675392 247512 675444 247518
rect 675392 247454 675444 247460
rect 675407 247367 675887 247423
rect 675407 246815 675887 246871
rect 675407 246171 675887 246227
rect 675407 245527 675887 245583
rect 675407 244975 675887 245031
rect 675407 244331 675887 244387
rect 675312 243701 675418 243729
rect 674012 237788 674064 237794
rect 674012 237730 674064 237736
rect 674024 231878 674052 237730
rect 675312 235725 675340 243701
rect 675407 243043 675887 243099
rect 675407 242491 675887 242547
rect 675407 241847 675887 241903
rect 675407 241203 675887 241259
rect 675407 240007 675887 240063
rect 675407 238167 675887 238223
rect 675392 237788 675444 237794
rect 675392 237730 675444 237736
rect 675404 237524 675432 237730
rect 675407 236327 675887 236383
rect 675312 235697 675418 235725
rect 673828 231872 673880 231878
rect 673828 231814 673880 231820
rect 674012 231872 674064 231878
rect 674012 231814 674064 231820
rect 673840 212537 673868 231814
rect 673826 212528 673882 212537
rect 673826 212463 673882 212472
rect 674010 212528 674066 212537
rect 674010 212463 674066 212472
rect 673736 202972 673788 202978
rect 673736 202914 673788 202920
rect 673920 202972 673972 202978
rect 673920 202914 673972 202920
rect 672552 198750 672672 198778
rect 673472 198750 673592 198778
rect 44640 195900 44692 195906
rect 44640 195842 44692 195848
rect 44652 183546 44680 195842
rect 672552 193225 672580 198750
rect 672538 193216 672594 193225
rect 672538 193151 672594 193160
rect 672906 193216 672962 193225
rect 672906 193151 672962 193160
rect 44560 183518 44680 183546
rect 44560 174010 44588 183518
rect 44548 174004 44600 174010
rect 44548 173946 44600 173952
rect 44732 174004 44784 174010
rect 44732 173946 44784 173952
rect 44744 171086 44772 173946
rect 672920 173942 672948 193151
rect 672724 173936 672776 173942
rect 672724 173878 672776 173884
rect 672908 173936 672960 173942
rect 672908 173878 672960 173884
rect 44456 171080 44508 171086
rect 44456 171022 44508 171028
rect 44732 171080 44784 171086
rect 44732 171022 44784 171028
rect 44468 151842 44496 171022
rect 672736 156602 672764 173878
rect 673472 158370 673500 198750
rect 673644 193248 673696 193254
rect 673644 193190 673696 193196
rect 673656 191962 673684 193190
rect 673644 191956 673696 191962
rect 673644 191898 673696 191904
rect 673460 158364 673512 158370
rect 673460 158306 673512 158312
rect 672540 156596 672592 156602
rect 672540 156538 672592 156544
rect 672724 156596 672776 156602
rect 672724 156538 672776 156544
rect 44456 151836 44508 151842
rect 44456 151778 44508 151784
rect 44640 151836 44692 151842
rect 44640 151778 44692 151784
rect 44652 140826 44680 151778
rect 44640 140820 44692 140826
rect 44640 140762 44692 140768
rect 672552 140706 672580 156538
rect 44732 140684 44784 140690
rect 672552 140678 672672 140706
rect 44732 140626 44784 140632
rect 44744 121582 44772 140626
rect 44732 121576 44784 121582
rect 44732 121518 44784 121524
rect 44640 121440 44692 121446
rect 44640 121382 44692 121388
rect 672644 121394 672672 140678
rect 44178 120184 44234 120193
rect 44178 120119 44234 120128
rect 44192 110537 44220 120119
rect 44178 110528 44234 110537
rect 44178 110463 44234 110472
rect 44652 102082 44680 121382
rect 672644 121366 672764 121394
rect 672736 115938 672764 121366
rect 672724 115932 672776 115938
rect 672724 115874 672776 115880
rect 672816 115932 672868 115938
rect 672816 115874 672868 115880
rect 45466 110528 45522 110537
rect 45466 110463 45522 110472
rect 44560 102054 44680 102082
rect 44560 96626 44588 102054
rect 44272 96620 44324 96626
rect 44272 96562 44324 96568
rect 44548 96620 44600 96626
rect 44548 96562 44600 96568
rect 44284 77314 44312 96562
rect 44272 77308 44324 77314
rect 44272 77250 44324 77256
rect 44364 77308 44416 77314
rect 44364 77250 44416 77256
rect 44270 75848 44326 75857
rect 44376 75834 44404 77250
rect 44326 75806 44404 75834
rect 44270 75783 44326 75792
rect 44284 73273 44312 75783
rect 44270 73264 44326 73273
rect 44270 73199 44326 73208
rect 44284 68241 44312 73199
rect 44270 68232 44326 68241
rect 44270 68167 44326 68176
rect 42708 64660 42760 64666
rect 42708 64602 42760 64608
rect 42248 45688 42300 45694
rect 42248 45630 42300 45636
rect 42720 45626 42748 64602
rect 45480 47938 45508 110463
rect 672828 102202 672856 115874
rect 673472 112810 673500 158306
rect 673552 157344 673604 157350
rect 673552 157286 673604 157292
rect 673460 112804 673512 112810
rect 673460 112746 673512 112752
rect 672816 102196 672868 102202
rect 672816 102138 672868 102144
rect 672724 102128 672776 102134
rect 672724 102070 672776 102076
rect 672736 96642 672764 102070
rect 672736 96614 672856 96642
rect 672828 82958 672856 96614
rect 672816 82952 672868 82958
rect 672816 82894 672868 82900
rect 672816 82748 672868 82754
rect 672816 82690 672868 82696
rect 45558 68232 45614 68241
rect 45558 68167 45614 68176
rect 45468 47932 45520 47938
rect 45468 47874 45520 47880
rect 45572 47802 45600 68167
rect 195980 47932 196032 47938
rect 195980 47874 196032 47880
rect 516324 47932 516376 47938
rect 516324 47874 516376 47880
rect 189172 47864 189224 47870
rect 189172 47806 189224 47812
rect 45560 47796 45612 47802
rect 45560 47738 45612 47744
rect 149060 47796 149112 47802
rect 149060 47738 149112 47744
rect 150900 47796 150952 47802
rect 150900 47738 150952 47744
rect 86408 47728 86460 47734
rect 86408 47670 86460 47676
rect 86420 46986 86448 47670
rect 86408 46980 86460 46986
rect 86408 46922 86460 46928
rect 42708 45620 42760 45626
rect 42708 45562 42760 45568
rect 86420 40225 86448 46922
rect 143540 45688 143592 45694
rect 143540 45630 143592 45636
rect 140964 45620 141016 45626
rect 140964 45562 141016 45568
rect 140976 44198 141004 45562
rect 143552 44266 143580 45630
rect 143540 44260 143592 44266
rect 143540 44202 143592 44208
rect 145104 44260 145156 44266
rect 145104 44202 145156 44208
rect 140964 44192 141016 44198
rect 140964 44134 141016 44140
rect 133098 40248 133150 40254
rect 86406 40216 86462 40225
rect 133098 40190 133150 40196
rect 140976 40202 141004 44134
rect 143816 40248 143868 40254
rect 86406 40151 86462 40160
rect 133110 39984 133138 40190
rect 140976 40174 141036 40202
rect 145116 40202 145144 44202
rect 149072 40361 149100 47738
rect 150912 47190 150940 47738
rect 150900 47184 150952 47190
rect 150900 47126 150952 47132
rect 186688 47116 186740 47122
rect 186688 47058 186740 47064
rect 186700 41820 186728 47058
rect 187327 41713 187383 42193
rect 189184 41834 189212 47806
rect 192852 47524 192904 47530
rect 192852 47466 192904 47472
rect 192864 47190 192892 47466
rect 192852 47184 192904 47190
rect 192852 47126 192904 47132
rect 189264 41880 189316 41886
rect 188554 41818 188660 41834
rect 189184 41828 189264 41834
rect 191104 41880 191156 41886
rect 189184 41822 189316 41828
rect 191038 41828 191104 41834
rect 192300 41880 192352 41886
rect 191038 41822 191156 41828
rect 192234 41828 192300 41834
rect 192864 41834 192892 47126
rect 194692 47116 194744 47122
rect 194692 47058 194744 47064
rect 192234 41822 192352 41828
rect 189184 41820 189304 41822
rect 188554 41812 188672 41818
rect 188554 41806 188620 41812
rect 189198 41806 189304 41820
rect 191038 41806 191144 41822
rect 192234 41806 192340 41822
rect 192772 41820 192892 41834
rect 192772 41818 192878 41820
rect 192760 41812 192878 41818
rect 188620 41754 188672 41760
rect 192812 41806 192878 41812
rect 193522 41818 193628 41834
rect 193522 41812 193640 41818
rect 193522 41806 193588 41812
rect 192760 41754 192812 41760
rect 193588 41754 193640 41760
rect 194043 41713 194099 42193
rect 194704 41820 194732 47058
rect 195992 47054 196020 47874
rect 414204 47864 414256 47870
rect 425060 47864 425112 47870
rect 414204 47806 414256 47812
rect 425058 47832 425060 47841
rect 430764 47864 430816 47870
rect 425112 47832 425114 47841
rect 201500 47524 201552 47530
rect 201500 47466 201552 47472
rect 358820 47524 358872 47530
rect 358820 47466 358872 47472
rect 359372 47524 359424 47530
rect 359372 47466 359424 47472
rect 199660 47252 199712 47258
rect 199660 47194 199712 47200
rect 199016 47116 199068 47122
rect 199016 47058 199068 47064
rect 195980 47048 196032 47054
rect 195980 46990 196032 46996
rect 195336 44260 195388 44266
rect 195336 44202 195388 44208
rect 195348 41834 195376 44202
rect 195428 41880 195480 41886
rect 195348 41828 195428 41834
rect 195348 41822 195480 41828
rect 195348 41820 195468 41822
rect 195992 41820 196020 46990
rect 199028 46986 199056 47058
rect 199016 46980 199068 46986
rect 199016 46922 199068 46928
rect 195362 41806 195468 41820
rect 196452 41818 198504 41834
rect 199028 41820 199056 46922
rect 199568 41880 199620 41886
rect 199672 41834 199700 47194
rect 200856 47184 200908 47190
rect 200856 47126 200908 47132
rect 200868 41834 200896 47126
rect 201512 46986 201540 47466
rect 328460 47456 328512 47462
rect 328458 47424 328460 47433
rect 328512 47424 328514 47433
rect 248328 47388 248380 47394
rect 328458 47359 328514 47368
rect 334070 47424 334126 47433
rect 334070 47359 334126 47368
rect 342260 47388 342312 47394
rect 248328 47330 248380 47336
rect 206928 47252 206980 47258
rect 206928 47194 206980 47200
rect 240140 47252 240192 47258
rect 240140 47194 240192 47200
rect 206940 46986 206968 47194
rect 201500 46980 201552 46986
rect 201500 46922 201552 46928
rect 206928 46980 206980 46986
rect 206928 46922 206980 46928
rect 199620 41828 199700 41834
rect 199568 41822 199700 41828
rect 199580 41820 199700 41822
rect 200132 41820 200896 41834
rect 201512 41820 201540 46922
rect 196440 41812 198516 41818
rect 196492 41806 198464 41812
rect 196440 41754 196492 41760
rect 199580 41806 199686 41820
rect 200132 41818 200882 41820
rect 200120 41812 200882 41818
rect 198464 41754 198516 41760
rect 200172 41806 200882 41812
rect 200120 41754 200172 41760
rect 149058 40352 149114 40361
rect 149058 40287 149114 40296
rect 143816 40190 143868 40196
rect 141008 40118 141036 40174
rect 140996 40112 141048 40118
rect 140996 40054 141048 40060
rect 143072 40112 143124 40118
rect 143072 40054 143124 40060
rect 143356 40112 143408 40118
rect 143356 40054 143408 40060
rect 141008 39984 141036 40054
rect 143084 39984 143112 40054
rect 143368 39916 143396 40054
rect 143828 39916 143856 40190
rect 145103 40174 145144 40202
rect 145103 40000 145131 40174
rect 145091 39706 145143 40000
rect 240152 39953 240180 47194
rect 242900 47184 242952 47190
rect 242900 47126 242952 47132
rect 242912 45558 242940 47126
rect 248340 47122 248368 47330
rect 334084 47326 334112 47359
rect 342260 47330 342312 47336
rect 358728 47388 358780 47394
rect 358728 47330 358780 47336
rect 307576 47320 307628 47326
rect 307576 47262 307628 47268
rect 334072 47320 334124 47326
rect 334072 47262 334124 47268
rect 289820 47184 289872 47190
rect 289818 47152 289820 47161
rect 305920 47184 305972 47190
rect 289872 47152 289874 47161
rect 247316 47116 247368 47122
rect 247316 47058 247368 47064
rect 248328 47116 248380 47122
rect 289818 47087 289874 47096
rect 303894 47152 303950 47161
rect 305920 47126 305972 47132
rect 303894 47087 303950 47096
rect 248328 47058 248380 47064
rect 242900 45552 242952 45558
rect 242900 45494 242952 45500
rect 240138 39944 240194 39953
rect 240138 39879 240194 39888
rect 242912 39817 242940 45494
rect 241242 39808 241298 39817
rect 241242 39743 241298 39752
rect 242898 39808 242954 39817
rect 242898 39743 242954 39752
rect 241256 39372 241284 39743
rect 247328 39567 247356 47058
rect 297732 45552 297784 45558
rect 297732 45494 297784 45500
rect 254032 44192 254084 44198
rect 254032 44134 254084 44140
rect 253940 41608 253992 41614
rect 253940 41550 253992 41556
rect 253952 39953 253980 41550
rect 253938 39944 253994 39953
rect 253938 39879 253994 39888
rect 254044 39710 254072 44134
rect 290186 41848 290242 41857
rect 297123 41848 297179 41857
rect 295311 41818 295472 41834
rect 295311 41812 295484 41818
rect 295311 41806 295432 41812
rect 290186 41783 290242 41792
rect 290200 41478 290228 41783
rect 297744 41834 297772 45494
rect 303908 42294 303936 47087
rect 304540 47048 304592 47054
rect 304540 46990 304592 46996
rect 303896 42288 303948 42294
rect 303896 42230 303948 42236
rect 302240 42016 302292 42022
rect 302240 41958 302292 41964
rect 297916 41880 297968 41886
rect 297744 41828 297916 41834
rect 300676 41880 300728 41886
rect 297744 41822 297968 41828
rect 299607 41848 299663 41857
rect 297744 41806 297956 41822
rect 297123 41783 297179 41792
rect 302252 41834 302280 41958
rect 300728 41828 302280 41834
rect 300676 41822 302280 41828
rect 300688 41806 302280 41822
rect 299607 41783 299663 41792
rect 295432 41754 295484 41760
rect 302643 41713 302699 42193
rect 303908 41834 303936 42230
rect 304552 41834 304580 46990
rect 305000 42016 305052 42022
rect 305000 41958 305052 41964
rect 305012 41834 305040 41958
rect 305932 41857 305960 47126
rect 305771 41848 305827 41857
rect 303172 41818 303315 41834
rect 303160 41812 303315 41818
rect 303212 41806 303315 41812
rect 303908 41806 303959 41834
rect 304552 41806 304603 41834
rect 305012 41818 305316 41834
rect 305012 41812 305328 41818
rect 305012 41806 305276 41812
rect 303160 41754 303212 41760
rect 305771 41783 305827 41792
rect 305918 41848 305974 41857
rect 306443 41818 306604 41834
rect 306443 41812 306616 41818
rect 306443 41806 306564 41812
rect 305918 41783 305974 41792
rect 305276 41754 305328 41760
rect 306564 41754 306616 41760
rect 306967 41713 307023 42193
rect 307588 41834 307616 47262
rect 309416 47252 309468 47258
rect 309416 47194 309468 47200
rect 309046 47152 309102 47161
rect 309046 47087 309048 47096
rect 309100 47087 309102 47096
rect 309048 47058 309100 47064
rect 308220 42288 308272 42294
rect 308220 42230 308272 42236
rect 308232 41834 308260 42230
rect 309428 41834 309456 47194
rect 342272 47122 342300 47330
rect 352564 47252 352616 47258
rect 352564 47194 352616 47200
rect 351920 47184 351972 47190
rect 351920 47126 351972 47132
rect 342260 47116 342312 47122
rect 342260 47058 342312 47064
rect 307588 41806 307639 41834
rect 308232 41806 308283 41834
rect 308692 41818 309479 41834
rect 308680 41812 309479 41818
rect 308732 41806 309479 41812
rect 308680 41754 308732 41760
rect 310095 41713 310151 42193
rect 351932 41834 351960 47126
rect 352576 41970 352604 47194
rect 352576 41954 352696 41970
rect 352576 41948 352708 41954
rect 352576 41942 352656 41948
rect 352012 41880 352064 41886
rect 350106 41818 350212 41834
rect 351932 41828 352012 41834
rect 351932 41822 352064 41828
rect 351932 41820 352052 41822
rect 352576 41820 352604 41942
rect 352656 41890 352708 41896
rect 355508 41948 355560 41954
rect 355508 41890 355560 41896
rect 356980 41948 357032 41954
rect 356980 41890 357032 41896
rect 354312 41880 354364 41886
rect 355520 41834 355548 41890
rect 356992 41834 357020 41890
rect 354364 41828 354430 41834
rect 354312 41822 354430 41828
rect 350106 41812 350224 41818
rect 350106 41806 350172 41812
rect 351946 41806 352052 41820
rect 354324 41806 354430 41822
rect 355520 41806 357020 41834
rect 350172 41754 350224 41760
rect 357443 41713 357499 42193
rect 358004 41818 358110 41834
rect 358740 41820 358768 47330
rect 358832 47054 358860 47466
rect 358820 47048 358872 47054
rect 358820 46990 358872 46996
rect 359384 41820 359412 47466
rect 411260 47456 411312 47462
rect 411260 47398 411312 47404
rect 361488 47388 361540 47394
rect 361488 47330 361540 47336
rect 360568 47184 360620 47190
rect 360568 47126 360620 47132
rect 359832 41948 359884 41954
rect 359832 41890 359884 41896
rect 359844 41834 359872 41890
rect 360476 41880 360528 41886
rect 357992 41812 358110 41818
rect 358044 41806 358110 41812
rect 359844 41806 359950 41834
rect 360580 41834 360608 47126
rect 361500 47122 361528 47330
rect 362408 47320 362460 47326
rect 362408 47262 362460 47268
rect 391940 47320 391992 47326
rect 391940 47262 391992 47268
rect 361488 47116 361540 47122
rect 361488 47058 361540 47064
rect 361120 41948 361172 41954
rect 361120 41890 361172 41896
rect 360528 41828 360608 41834
rect 360476 41822 360608 41828
rect 360488 41820 360608 41822
rect 361132 41834 361160 41890
rect 360488 41806 360594 41820
rect 361132 41806 361238 41834
rect 357992 41754 358044 41760
rect 361767 41713 361823 42193
rect 362420 41820 362448 47262
rect 364248 47252 364300 47258
rect 364248 47194 364300 47200
rect 363052 47116 363104 47122
rect 363052 47058 363104 47064
rect 363064 41820 363092 47058
rect 364260 41834 364288 47194
rect 391952 47054 391980 47262
rect 407396 47252 407448 47258
rect 407396 47194 407448 47200
rect 406752 47184 406804 47190
rect 406752 47126 406804 47132
rect 391940 47048 391992 47054
rect 391940 46990 391992 46996
rect 363524 41820 364288 41834
rect 363524 41818 364274 41820
rect 363512 41812 364274 41818
rect 363564 41806 364274 41812
rect 363512 41754 363564 41760
rect 364895 41713 364951 42193
rect 404938 41818 405044 41834
rect 404938 41812 405056 41818
rect 404938 41806 405004 41812
rect 405004 41754 405056 41760
rect 405527 41713 405583 42193
rect 406764 41820 406792 47126
rect 407408 41970 407436 47194
rect 411168 47184 411220 47190
rect 411272 47172 411300 47398
rect 411220 47144 411300 47172
rect 411168 47126 411220 47132
rect 411076 47116 411128 47122
rect 411076 47058 411128 47064
rect 410984 47048 411036 47054
rect 410984 46990 411036 46996
rect 410996 45422 411024 46990
rect 410984 45416 411036 45422
rect 410984 45358 411036 45364
rect 411088 44470 411116 47058
rect 411076 44464 411128 44470
rect 411076 44406 411128 44412
rect 413560 44464 413612 44470
rect 413560 44406 413612 44412
rect 413572 42294 413600 44406
rect 413560 42288 413612 42294
rect 413560 42230 413612 42236
rect 411536 42016 411588 42022
rect 407408 41954 407528 41970
rect 411588 41964 411760 41970
rect 411536 41958 411760 41964
rect 407408 41948 407540 41954
rect 407408 41942 407488 41948
rect 407408 41820 407436 41942
rect 407488 41890 407540 41896
rect 410248 41948 410300 41954
rect 410248 41890 410300 41896
rect 411168 41948 411220 41954
rect 411548 41942 411760 41958
rect 411168 41890 411220 41896
rect 409328 41880 409380 41886
rect 409262 41828 409328 41834
rect 409262 41822 409380 41828
rect 410260 41834 410288 41890
rect 411180 41834 411208 41890
rect 409262 41806 409368 41822
rect 410260 41806 410458 41834
rect 411102 41806 411208 41834
rect 411732 41820 411760 41942
rect 412243 41834 412299 42193
rect 412364 41880 412416 41886
rect 412243 41828 412364 41834
rect 412243 41822 412416 41828
rect 412243 41806 412404 41822
rect 412744 41818 412942 41834
rect 413572 41820 413600 42230
rect 414216 41820 414244 47806
rect 425058 47767 425114 47776
rect 430762 47832 430764 47841
rect 430816 47832 430818 47841
rect 430762 47767 430818 47776
rect 466460 47728 466512 47734
rect 466460 47670 466512 47676
rect 460938 47560 460994 47569
rect 422300 47524 422352 47530
rect 422300 47466 422352 47472
rect 441528 47524 441580 47530
rect 460938 47495 460940 47504
rect 441528 47466 441580 47472
rect 460992 47495 460994 47504
rect 461490 47560 461546 47569
rect 461490 47495 461546 47504
rect 460940 47466 460992 47472
rect 417240 47388 417292 47394
rect 417240 47330 417292 47336
rect 417252 45422 417280 47330
rect 422312 47326 422340 47466
rect 441540 47326 441568 47466
rect 422300 47320 422352 47326
rect 422300 47262 422352 47268
rect 441528 47320 441580 47326
rect 441528 47262 441580 47268
rect 453488 47320 453540 47326
rect 453488 47262 453540 47268
rect 419080 47252 419132 47258
rect 419080 47194 419132 47200
rect 417884 47184 417936 47190
rect 417884 47126 417936 47132
rect 417240 45416 417292 45422
rect 417240 45358 417292 45364
rect 414572 42016 414624 42022
rect 414572 41958 414624 41964
rect 415860 42016 415912 42022
rect 415860 41958 415912 41964
rect 414584 41834 414612 41958
rect 415492 41880 415544 41886
rect 412732 41812 412942 41818
rect 412243 41713 412299 41806
rect 412784 41806 412942 41812
rect 414584 41806 414782 41834
rect 415426 41828 415492 41834
rect 415426 41822 415544 41828
rect 415872 41834 415900 41958
rect 415426 41806 415532 41822
rect 415872 41806 416070 41834
rect 412732 41754 412784 41760
rect 416567 41713 416623 42193
rect 417252 41820 417280 45358
rect 417896 42294 417924 47126
rect 417884 42288 417936 42294
rect 417884 42230 417936 42236
rect 417896 41820 417924 42230
rect 418252 42016 418304 42022
rect 418252 41958 418304 41964
rect 418264 41834 418292 41958
rect 419092 41834 419120 47194
rect 453500 46986 453528 47262
rect 453488 46980 453540 46986
rect 453488 46922 453540 46928
rect 418264 41820 419120 41834
rect 419540 41880 419592 41886
rect 419695 41834 419751 42193
rect 419592 41828 419751 41834
rect 419540 41822 419751 41828
rect 418264 41806 419106 41820
rect 419552 41806 419751 41822
rect 459711 41818 459876 41834
rect 459711 41812 459888 41818
rect 459711 41806 459836 41812
rect 419695 41713 419751 41806
rect 459836 41754 459888 41760
rect 460327 41713 460383 42193
rect 461504 41834 461532 47495
rect 466472 47258 466500 47670
rect 480168 47592 480220 47598
rect 480088 47569 480168 47580
rect 480074 47560 480168 47569
rect 480130 47552 480168 47560
rect 483020 47592 483072 47598
rect 480168 47534 480220 47540
rect 483018 47560 483020 47569
rect 483072 47560 483074 47569
rect 480074 47495 480130 47504
rect 483018 47495 483074 47504
rect 488630 47560 488686 47569
rect 488630 47495 488686 47504
rect 488644 47462 488672 47495
rect 516336 47462 516364 47874
rect 529848 47864 529900 47870
rect 529848 47806 529900 47812
rect 528652 47796 528704 47802
rect 528652 47738 528704 47744
rect 488632 47456 488684 47462
rect 488632 47398 488684 47404
rect 516324 47456 516376 47462
rect 516324 47398 516376 47404
rect 474648 47388 474700 47394
rect 474648 47330 474700 47336
rect 462136 47252 462188 47258
rect 462136 47194 462188 47200
rect 466460 47252 466512 47258
rect 466460 47194 466512 47200
rect 468944 47252 468996 47258
rect 468944 47194 468996 47200
rect 469220 47252 469272 47258
rect 469220 47194 469272 47200
rect 473820 47252 473872 47258
rect 473820 47194 473872 47200
rect 462148 41834 462176 47194
rect 468300 47184 468352 47190
rect 468300 47126 468352 47132
rect 466368 42016 466420 42022
rect 466368 41958 466420 41964
rect 462320 41948 462372 41954
rect 462320 41890 462372 41896
rect 465080 41948 465132 41954
rect 465080 41890 465132 41896
rect 466000 41948 466052 41954
rect 466000 41890 466052 41896
rect 462332 41834 462360 41890
rect 464160 41880 464212 41886
rect 461504 41806 461551 41834
rect 462148 41806 462360 41834
rect 464035 41828 464160 41834
rect 464035 41822 464212 41828
rect 465092 41834 465120 41890
rect 466012 41834 466040 41890
rect 464035 41806 464200 41822
rect 465092 41806 465231 41834
rect 465875 41806 466040 41834
rect 466380 41834 466408 41958
rect 466920 41880 466972 41886
rect 466380 41806 466519 41834
rect 467043 41834 467099 42193
rect 468312 41834 468340 47126
rect 468484 41880 468536 41886
rect 466972 41828 467099 41834
rect 466920 41822 467099 41828
rect 466932 41806 467099 41822
rect 467576 41818 467715 41834
rect 467043 41713 467099 41806
rect 467564 41812 467715 41818
rect 467616 41806 467715 41812
rect 468312 41828 468484 41834
rect 468312 41822 468536 41828
rect 468956 41834 468984 47194
rect 469232 47054 469260 47194
rect 469220 47048 469272 47054
rect 469220 46990 469272 46996
rect 471980 46980 472032 46986
rect 471980 46922 472032 46928
rect 469404 42016 469456 42022
rect 469404 41958 469456 41964
rect 470692 42016 470744 42022
rect 470692 41958 470744 41964
rect 469416 41834 469444 41958
rect 470704 41834 470732 41958
rect 468312 41806 468524 41822
rect 468956 41806 469003 41834
rect 469416 41806 469555 41834
rect 470060 41818 470199 41834
rect 470048 41812 470199 41818
rect 467564 41754 467616 41760
rect 470100 41806 470199 41812
rect 470704 41806 470843 41834
rect 470048 41754 470100 41760
rect 471367 41713 471423 42193
rect 471992 41834 472020 46922
rect 473084 42016 473136 42022
rect 473084 41958 473136 41964
rect 472532 41880 472584 41886
rect 471992 41806 472039 41834
rect 473096 41834 473124 41958
rect 473832 41834 473860 47194
rect 474660 46986 474688 47330
rect 474648 46980 474700 46986
rect 474648 46922 474700 46928
rect 514484 46980 514536 46986
rect 514484 46922 514536 46928
rect 474372 41948 474424 41954
rect 474372 41890 474424 41896
rect 474384 41834 474412 41890
rect 474495 41834 474551 42193
rect 472584 41828 472683 41834
rect 472532 41822 472683 41828
rect 472544 41806 472683 41822
rect 473096 41806 473879 41834
rect 474384 41806 474551 41834
rect 514496 41820 514524 46922
rect 474495 41713 474551 41806
rect 515127 41713 515183 42193
rect 516336 41820 516364 47398
rect 524420 47388 524472 47394
rect 524420 47330 524472 47336
rect 516968 47252 517020 47258
rect 516968 47194 517020 47200
rect 516980 41834 517008 47194
rect 524432 47190 524460 47330
rect 527456 47252 527508 47258
rect 527456 47194 527508 47200
rect 524420 47184 524472 47190
rect 524420 47126 524472 47132
rect 526812 47184 526864 47190
rect 526812 47126 526864 47132
rect 523776 47116 523828 47122
rect 523776 47058 523828 47064
rect 523788 46986 523816 47058
rect 522488 46980 522540 46986
rect 522488 46922 522540 46928
rect 523776 46980 523828 46986
rect 523776 46922 523828 46928
rect 518900 41880 518952 41886
rect 516980 41820 517100 41834
rect 516994 41818 517100 41820
rect 518834 41828 518900 41834
rect 518834 41822 518952 41828
rect 516994 41812 517112 41818
rect 516994 41806 517060 41812
rect 518834 41806 518940 41822
rect 520030 41818 520136 41834
rect 520030 41812 520148 41818
rect 520030 41806 520096 41812
rect 517060 41754 517112 41760
rect 520096 41754 520148 41760
rect 520647 41713 520703 42193
rect 521318 41818 521424 41834
rect 521318 41812 521436 41818
rect 521318 41806 521384 41812
rect 521384 41754 521436 41760
rect 521843 41713 521899 42193
rect 522500 41820 522528 46922
rect 523224 41948 523276 41954
rect 523224 41890 523276 41896
rect 523236 41834 523264 41890
rect 523158 41806 523264 41834
rect 523788 41820 523816 46922
rect 524880 41880 524932 41886
rect 524354 41818 524460 41834
rect 524971 41834 525027 42193
rect 524932 41828 525027 41834
rect 524880 41822 525027 41828
rect 524354 41812 524472 41818
rect 524354 41806 524420 41812
rect 524892 41806 525027 41822
rect 525642 41818 525748 41834
rect 525642 41812 525760 41818
rect 525642 41806 525708 41812
rect 524420 41754 524472 41760
rect 524971 41713 525027 41806
rect 525708 41754 525760 41760
rect 526167 41713 526223 42193
rect 526824 41820 526852 47126
rect 527468 41970 527496 47194
rect 527376 41954 527496 41970
rect 527364 41948 527496 41954
rect 527416 41942 527496 41948
rect 527364 41890 527416 41896
rect 527468 41820 527496 41942
rect 528664 41834 528692 47738
rect 529860 47258 529888 47806
rect 672828 47802 672856 82690
rect 673472 47870 673500 112746
rect 673564 112130 673592 157286
rect 673656 147898 673684 191898
rect 673932 157350 673960 202914
rect 674024 193254 674052 212463
rect 675300 206780 675352 206786
rect 675300 206722 675352 206728
rect 675312 203497 675340 206722
rect 675407 205295 675887 205351
rect 675407 204651 675887 204707
rect 675407 204007 675887 204063
rect 675312 203469 675418 203497
rect 675392 202972 675444 202978
rect 675392 202914 675444 202920
rect 675404 202844 675432 202914
rect 675407 202167 675887 202223
rect 675407 201615 675887 201671
rect 675407 200971 675887 201027
rect 675407 200327 675887 200383
rect 675407 199775 675887 199831
rect 675407 199131 675887 199187
rect 675312 198614 675432 198642
rect 674012 193248 674064 193254
rect 674012 193190 674064 193196
rect 675312 190525 675340 198614
rect 675404 198492 675432 198614
rect 675407 197843 675887 197899
rect 675407 197291 675887 197347
rect 675407 196647 675887 196703
rect 675407 196003 675887 196059
rect 675407 194807 675887 194863
rect 675407 192967 675887 193023
rect 675404 191962 675432 192372
rect 675392 191956 675444 191962
rect 675392 191898 675444 191904
rect 675407 191127 675887 191183
rect 675312 190497 675418 190525
rect 675407 160295 675887 160351
rect 675407 159651 675887 159707
rect 675407 159007 675887 159063
rect 675404 158370 675432 158508
rect 675392 158364 675444 158370
rect 675392 158306 675444 158312
rect 675404 157350 675432 157828
rect 673920 157344 673972 157350
rect 673920 157286 673972 157292
rect 675392 157344 675444 157350
rect 675392 157286 675444 157292
rect 675407 157167 675887 157223
rect 675407 156615 675887 156671
rect 675407 155971 675887 156027
rect 675407 155327 675887 155383
rect 675407 154775 675887 154831
rect 675407 154131 675887 154187
rect 675312 153501 675418 153529
rect 673644 147892 673696 147898
rect 673644 147834 673696 147840
rect 674012 147892 674064 147898
rect 674012 147834 674064 147840
rect 674024 140706 674052 147834
rect 675312 145525 675340 153501
rect 675407 152843 675887 152899
rect 675407 152291 675887 152347
rect 675407 151647 675887 151703
rect 675407 151003 675887 151059
rect 675407 149807 675887 149863
rect 675407 147967 675887 148023
rect 675392 147892 675444 147898
rect 675392 147834 675444 147840
rect 675404 147356 675432 147834
rect 675407 146127 675887 146183
rect 675312 145497 675418 145525
rect 673932 140678 674052 140706
rect 673932 121530 673960 140678
rect 673840 121502 673960 121530
rect 673552 112124 673604 112130
rect 673552 112066 673604 112072
rect 673460 47864 673512 47870
rect 673460 47806 673512 47812
rect 672816 47796 672868 47802
rect 672816 47738 672868 47744
rect 529848 47252 529900 47258
rect 529848 47194 529900 47200
rect 634820 47184 634872 47190
rect 634820 47126 634872 47132
rect 569132 47116 569184 47122
rect 569132 47058 569184 47064
rect 527928 41820 528692 41834
rect 527928 41818 528678 41820
rect 527916 41812 528678 41818
rect 527968 41806 528678 41812
rect 527916 41754 527968 41760
rect 529295 41713 529351 42193
rect 290188 41472 290240 41478
rect 290188 41414 290240 41420
rect 252100 39704 252152 39710
rect 252100 39646 252152 39652
rect 254032 39704 254084 39710
rect 254032 39646 254084 39652
rect 252112 39372 252140 39646
rect 569144 39644 569172 47058
rect 579160 45552 579212 45558
rect 579160 45494 579212 45500
rect 569224 44192 569276 44198
rect 569224 44134 569276 44140
rect 569236 40225 569264 44134
rect 579172 40225 579200 45494
rect 622950 40488 623006 40497
rect 622950 40423 623006 40432
rect 569222 40216 569278 40225
rect 569222 40151 569278 40160
rect 579158 40216 579214 40225
rect 579158 40151 579214 40160
rect 579172 39644 579200 40151
rect 622964 39681 622992 40423
rect 634832 40225 634860 47126
rect 673564 45558 673592 112066
rect 673840 102202 673868 121502
rect 675407 115095 675887 115151
rect 675407 114451 675887 114507
rect 675407 113807 675887 113863
rect 675404 112810 675432 113283
rect 675392 112804 675444 112810
rect 675392 112746 675444 112752
rect 675404 112130 675432 112639
rect 675392 112124 675444 112130
rect 675392 112066 675444 112072
rect 675407 111967 675887 112023
rect 675407 111415 675887 111471
rect 675407 110771 675887 110827
rect 675407 110127 675887 110183
rect 675407 109575 675887 109631
rect 675407 108931 675887 108987
rect 675312 108310 675418 108338
rect 673644 102196 673696 102202
rect 673644 102138 673696 102144
rect 673828 102196 673880 102202
rect 673828 102138 673880 102144
rect 673656 102066 673684 102138
rect 673644 102060 673696 102066
rect 673644 102002 673696 102008
rect 673656 47938 673684 102002
rect 675312 100314 675340 108310
rect 675407 107643 675887 107699
rect 675407 107091 675887 107147
rect 675407 106447 675887 106503
rect 675407 105803 675887 105859
rect 675407 104607 675887 104663
rect 675407 102767 675887 102823
rect 675404 102066 675432 102151
rect 675392 102060 675444 102066
rect 675392 102002 675444 102008
rect 675407 100927 675887 100983
rect 675312 100286 675418 100314
rect 673644 47932 673696 47938
rect 673644 47874 673696 47880
rect 673552 45552 673604 45558
rect 673552 45494 673604 45500
rect 632978 40216 633034 40225
rect 632978 40151 633034 40160
rect 634818 40216 634874 40225
rect 634818 40151 634874 40160
rect 622950 39672 623006 39681
rect 632992 39644 633020 40151
rect 622950 39607 623006 39616
<< via2 >>
rect 328550 997328 328606 997384
rect 39670 922256 39726 922312
rect 45466 990120 45522 990176
rect 39670 920216 39726 920272
rect 39670 908112 39726 908168
rect 40130 877512 40186 877568
rect 41418 875064 41474 875120
rect 40130 870032 40186 870088
rect 40498 830728 40554 830784
rect 39670 827464 39726 827520
rect 40498 811552 40554 811608
rect 42430 866632 42486 866688
rect 42614 885964 42670 886000
rect 42614 885944 42616 885964
rect 42616 885944 42668 885964
rect 42668 885944 42670 885964
rect 42890 885944 42946 886000
rect 44178 870032 44234 870088
rect 42706 866632 42762 866688
rect 39854 778504 39910 778560
rect 39854 772792 39910 772848
rect 40222 550568 40278 550624
rect 40222 546352 40278 546408
rect 39762 492904 39818 492960
rect 39946 455368 40002 455424
rect 39670 451832 39726 451888
rect 39670 440952 39726 441008
rect 41694 275657 41750 275713
rect 42246 275657 42302 275713
rect 41694 184933 41750 184989
rect 42338 184933 42394 184989
rect 39762 120128 39818 120184
rect 41418 115912 41474 115968
rect 42154 115912 42210 115968
rect 39394 84224 39450 84280
rect 44362 917224 44418 917280
rect 45834 877512 45890 877568
rect 77298 990276 77354 990312
rect 77298 990256 77300 990276
rect 77300 990256 77352 990276
rect 77352 990256 77354 990276
rect 132498 990428 132500 990448
rect 132500 990428 132552 990448
rect 132552 990428 132554 990448
rect 132498 990392 132554 990428
rect 140778 990392 140834 990448
rect 347686 997056 347742 997112
rect 672630 996512 672686 996568
rect 585690 996376 585746 996432
rect 672446 996376 672502 996432
rect 82910 990256 82966 990312
rect 328458 990276 328514 990312
rect 328458 990256 328460 990276
rect 328460 990256 328512 990276
rect 328512 990256 328514 990276
rect 44638 835216 44694 835272
rect 44454 828008 44510 828064
rect 672538 828688 672594 828744
rect 673366 908112 673422 908168
rect 672630 826104 672686 826160
rect 673274 826104 673330 826160
rect 672538 823656 672594 823712
rect 673182 823656 673238 823712
rect 672814 792104 672870 792160
rect 672998 792104 673054 792160
rect 673090 721384 673146 721440
rect 672998 714856 673054 714912
rect 672998 514120 673054 514176
rect 673182 514120 673238 514176
rect 673090 511400 673146 511456
rect 673274 511400 673330 511456
rect 672998 509088 673054 509144
rect 44638 493176 44694 493232
rect 44454 488552 44510 488608
rect 672998 463664 673054 463720
rect 44362 448568 44418 448624
rect 677874 918584 677930 918640
rect 677598 915320 677654 915376
rect 677598 912736 677654 912792
rect 677874 912736 677930 912792
rect 677874 908112 677930 908168
rect 677782 907704 677838 907760
rect 673734 850040 673790 850096
rect 673918 850040 673974 850096
rect 673826 772792 673882 772848
rect 675206 772792 675262 772848
rect 673734 685344 673790 685400
rect 675390 685344 675446 685400
rect 673366 467472 673422 467528
rect 673274 463664 673330 463720
rect 678058 480120 678114 480176
rect 677874 469920 677930 469976
rect 673090 427896 673146 427952
rect 673366 420824 673422 420880
rect 672722 391992 672778 392048
rect 672722 386416 672778 386472
rect 677414 427896 677470 427952
rect 677598 425720 677654 425776
rect 673550 338680 673606 338736
rect 672538 295432 672594 295488
rect 672630 295160 672686 295216
rect 675390 338680 675446 338736
rect 673458 292984 673514 293040
rect 675390 292984 675446 293040
rect 673826 212472 673882 212528
rect 674010 212472 674066 212528
rect 672538 193160 672594 193216
rect 672906 193160 672962 193216
rect 44178 120128 44234 120184
rect 44178 110472 44234 110528
rect 45466 110472 45522 110528
rect 44270 75792 44326 75848
rect 44270 73208 44326 73264
rect 44270 68176 44326 68232
rect 45558 68176 45614 68232
rect 86406 40160 86462 40216
rect 425058 47812 425060 47832
rect 425060 47812 425112 47832
rect 425112 47812 425114 47832
rect 328458 47404 328460 47424
rect 328460 47404 328512 47424
rect 328512 47404 328514 47424
rect 328458 47368 328514 47404
rect 334070 47368 334126 47424
rect 149058 40296 149114 40352
rect 289818 47132 289820 47152
rect 289820 47132 289872 47152
rect 289872 47132 289874 47152
rect 289818 47096 289874 47132
rect 303894 47096 303950 47152
rect 240138 39888 240194 39944
rect 241242 39752 241298 39808
rect 242898 39752 242954 39808
rect 253938 39888 253994 39944
rect 290186 41792 290242 41848
rect 297123 41792 297179 41848
rect 299607 41792 299663 41848
rect 305771 41792 305827 41848
rect 305918 41792 305974 41848
rect 309046 47116 309102 47152
rect 309046 47096 309048 47116
rect 309048 47096 309100 47116
rect 309100 47096 309102 47116
rect 425058 47776 425114 47812
rect 430762 47812 430764 47832
rect 430764 47812 430816 47832
rect 430816 47812 430818 47832
rect 430762 47776 430818 47812
rect 460938 47524 460994 47560
rect 460938 47504 460940 47524
rect 460940 47504 460992 47524
rect 460992 47504 460994 47524
rect 461490 47504 461546 47560
rect 480074 47504 480130 47560
rect 483018 47540 483020 47560
rect 483020 47540 483072 47560
rect 483072 47540 483074 47560
rect 483018 47504 483074 47540
rect 488630 47504 488686 47560
rect 622950 40432 623006 40488
rect 569222 40160 569278 40216
rect 579158 40160 579214 40216
rect 632978 40160 633034 40216
rect 634818 40160 634874 40216
rect 622950 39616 623006 39672
<< metal3 >>
rect 328545 997386 328611 997389
rect 338622 997386 338682 997628
rect 341006 997596 341012 997660
rect 341076 997596 341082 997660
rect 343590 997386 343650 997628
rect 580796 997598 581746 997658
rect 581686 997522 581746 997598
rect 585734 997522 585794 997628
rect 581686 997462 585794 997522
rect 328545 997384 343650 997386
rect 328545 997328 328550 997384
rect 328606 997328 343650 997384
rect 328545 997326 343650 997328
rect 328545 997323 328611 997326
rect 343590 997114 343650 997326
rect 347681 997114 347747 997117
rect 343590 997112 347747 997114
rect 343590 997056 347686 997112
rect 347742 997056 347747 997112
rect 343590 997054 347747 997056
rect 585734 997114 585794 997462
rect 585734 997054 585978 997114
rect 347681 997051 347747 997054
rect 585918 996570 585978 997054
rect 672625 996570 672691 996573
rect 585918 996568 672691 996570
rect 585918 996512 672630 996568
rect 672686 996512 672691 996568
rect 585918 996510 672691 996512
rect 672625 996507 672691 996510
rect 585685 996434 585751 996437
rect 672441 996434 672507 996437
rect 585685 996432 672507 996434
rect 585685 996376 585690 996432
rect 585746 996376 672446 996432
rect 672502 996376 672507 996432
rect 585685 996374 672507 996376
rect 585685 996371 585751 996374
rect 672441 996371 672507 996374
rect 132493 990450 132559 990453
rect 140773 990450 140839 990453
rect 132493 990448 140839 990450
rect 132493 990392 132498 990448
rect 132554 990392 140778 990448
rect 140834 990392 140839 990448
rect 132493 990390 140839 990392
rect 132493 990387 132559 990390
rect 140773 990387 140839 990390
rect 77293 990314 77359 990317
rect 82905 990314 82971 990317
rect 77293 990312 82971 990314
rect 77293 990256 77298 990312
rect 77354 990256 82910 990312
rect 82966 990256 82971 990312
rect 77293 990254 82971 990256
rect 77293 990251 77359 990254
rect 82905 990251 82971 990254
rect 328453 990314 328519 990317
rect 341006 990314 341012 990316
rect 328453 990312 341012 990314
rect 328453 990256 328458 990312
rect 328514 990256 341012 990312
rect 328453 990254 341012 990256
rect 328453 990251 328519 990254
rect 341006 990252 341012 990254
rect 341076 990252 341082 990316
rect 45461 990178 45527 990181
rect 676254 990178 676260 990180
rect 45461 990176 676260 990178
rect 45461 990120 45466 990176
rect 45522 990120 676260 990176
rect 45461 990118 676260 990120
rect 45461 990115 45527 990118
rect 676254 990116 676260 990118
rect 676324 990116 676330 990180
rect 39665 922314 39731 922317
rect 39468 922312 39731 922314
rect 39468 922256 39670 922312
rect 39726 922256 39731 922312
rect 39468 922254 39731 922256
rect 39665 922251 39731 922254
rect 39665 920274 39731 920277
rect 39438 920272 39731 920274
rect 39438 920216 39670 920272
rect 39726 920216 39731 920272
rect 39438 920214 39731 920216
rect 39438 919730 39498 920214
rect 39665 920211 39731 920214
rect 39438 919700 39866 919730
rect 39468 919670 39866 919700
rect 39806 919322 39866 919670
rect 39438 919262 39866 919322
rect 39438 917282 39498 919262
rect 677542 918580 677548 918644
rect 677612 918642 677618 918644
rect 677869 918642 677935 918645
rect 677612 918640 677935 918642
rect 677612 918584 677874 918640
rect 677930 918584 677935 918640
rect 677612 918582 677935 918584
rect 677612 918580 677618 918582
rect 677869 918579 677935 918582
rect 44357 917282 44423 917285
rect 39438 917280 44423 917282
rect 39438 917252 44362 917280
rect 39468 917224 44362 917252
rect 44418 917224 44423 917280
rect 39468 917222 44423 917224
rect 44357 917219 44423 917222
rect 677593 915378 677659 915381
rect 677593 915376 678132 915378
rect 677593 915320 677598 915376
rect 677654 915320 678132 915376
rect 677593 915318 678132 915320
rect 677593 915315 677659 915318
rect 677593 912794 677659 912797
rect 677869 912794 677935 912797
rect 677593 912792 678132 912794
rect 677593 912736 677598 912792
rect 677654 912736 677874 912792
rect 677930 912736 678132 912792
rect 677593 912734 678132 912736
rect 677593 912731 677659 912734
rect 677869 912731 677935 912734
rect 39665 908170 39731 908173
rect 40166 908170 40172 908172
rect 39665 908168 40172 908170
rect 39665 908112 39670 908168
rect 39726 908112 40172 908168
rect 39665 908110 40172 908112
rect 39665 908107 39731 908110
rect 40166 908108 40172 908110
rect 40236 908108 40242 908172
rect 673361 908170 673427 908173
rect 677869 908170 677935 908173
rect 673361 908168 678162 908170
rect 673361 908112 673366 908168
rect 673422 908112 677874 908168
rect 677930 908112 678162 908168
rect 673361 908110 678162 908112
rect 673361 908107 673427 908110
rect 677869 908107 677935 908110
rect 676254 907700 676260 907764
rect 676324 907762 676330 907764
rect 677777 907762 677843 907765
rect 676324 907760 677843 907762
rect 676324 907704 677782 907760
rect 677838 907704 677843 907760
rect 678102 907732 678162 908110
rect 676324 907702 677843 907704
rect 676324 907700 676330 907702
rect 677777 907699 677843 907702
rect 42609 886002 42675 886005
rect 42885 886002 42951 886005
rect 42609 886000 42951 886002
rect 42609 885944 42614 886000
rect 42670 885944 42890 886000
rect 42946 885944 42951 886000
rect 42609 885942 42951 885944
rect 42609 885939 42675 885942
rect 42885 885939 42951 885942
rect 40125 877570 40191 877573
rect 45829 877570 45895 877573
rect 39622 877568 45895 877570
rect 39622 877512 40130 877568
rect 40186 877512 45834 877568
rect 45890 877512 45895 877568
rect 39622 877510 45895 877512
rect 39622 877404 39682 877510
rect 40125 877507 40191 877510
rect 45829 877507 45895 877510
rect 41413 875122 41479 875125
rect 39652 875120 41479 875122
rect 39652 875064 41418 875120
rect 41474 875064 41479 875120
rect 39652 875062 41479 875064
rect 41413 875059 41479 875062
rect 40125 870090 40191 870093
rect 44173 870090 44239 870093
rect 39622 870088 44239 870090
rect 39622 870032 40130 870088
rect 40186 870032 44178 870088
rect 44234 870032 44239 870088
rect 39622 870030 44239 870032
rect 39622 869924 39682 870030
rect 40125 870027 40191 870030
rect 44173 870027 44239 870030
rect 42425 866690 42491 866693
rect 42701 866690 42767 866693
rect 42425 866688 42767 866690
rect 42425 866632 42430 866688
rect 42486 866632 42706 866688
rect 42762 866632 42767 866688
rect 42425 866630 42767 866632
rect 42425 866627 42491 866630
rect 42701 866627 42767 866630
rect 673729 850098 673795 850101
rect 673913 850098 673979 850101
rect 673729 850096 673979 850098
rect 673729 850040 673734 850096
rect 673790 850040 673918 850096
rect 673974 850040 673979 850096
rect 673729 850038 673979 850040
rect 673729 850035 673795 850038
rect 673913 850035 673979 850038
rect 44633 835274 44699 835277
rect 39652 835272 44699 835274
rect 39652 835216 44638 835272
rect 44694 835216 44699 835272
rect 39652 835214 44699 835216
rect 44633 835211 44699 835214
rect 40350 830724 40356 830788
rect 40420 830786 40426 830788
rect 40493 830786 40559 830789
rect 40420 830784 40559 830786
rect 40420 830728 40498 830784
rect 40554 830728 40559 830784
rect 40420 830726 40559 830728
rect 40420 830724 40426 830726
rect 40493 830723 40559 830726
rect 672533 828746 672599 828749
rect 672533 828744 677794 828746
rect 672533 828688 672538 828744
rect 672594 828688 677794 828744
rect 672533 828686 677794 828688
rect 672533 828683 672599 828686
rect 677734 828580 677794 828686
rect 44449 828066 44515 828069
rect 39806 828064 44515 828066
rect 39806 828008 44454 828064
rect 44510 828008 44515 828064
rect 39806 828006 44515 828008
rect 39806 827794 39866 828006
rect 44449 828003 44515 828006
rect 39652 827734 39866 827794
rect 39665 827522 39731 827525
rect 39806 827522 39866 827734
rect 39665 827520 39866 827522
rect 39665 827464 39670 827520
rect 39726 827464 39866 827520
rect 39665 827462 39866 827464
rect 39665 827459 39731 827462
rect 672625 826162 672691 826165
rect 673269 826162 673335 826165
rect 672625 826160 677764 826162
rect 672625 826104 672630 826160
rect 672686 826104 673274 826160
rect 673330 826104 677764 826160
rect 672625 826102 677764 826104
rect 672625 826099 672691 826102
rect 673269 826099 673335 826102
rect 672533 823714 672599 823717
rect 673177 823714 673243 823717
rect 672533 823712 677764 823714
rect 672533 823656 672538 823712
rect 672594 823656 673182 823712
rect 673238 823656 677764 823712
rect 672533 823654 677764 823656
rect 672533 823651 672599 823654
rect 673177 823651 673243 823654
rect 40493 811612 40559 811613
rect 40493 811608 40540 811612
rect 40604 811610 40610 811612
rect 40493 811552 40498 811608
rect 40493 811548 40540 811552
rect 40604 811550 40650 811610
rect 40604 811548 40610 811550
rect 40493 811547 40559 811548
rect 40350 811276 40356 811340
rect 40420 811276 40426 811340
rect 40358 811202 40418 811276
rect 40902 811202 40908 811204
rect 40358 811142 40908 811202
rect 40902 811140 40908 811142
rect 40972 811140 40978 811204
rect 40534 792100 40540 792164
rect 40604 792162 40610 792164
rect 40902 792162 40908 792164
rect 40604 792102 40908 792162
rect 40604 792100 40610 792102
rect 40902 792100 40908 792102
rect 40972 792100 40978 792164
rect 672809 792162 672875 792165
rect 672993 792162 673059 792165
rect 672809 792160 673059 792162
rect 672809 792104 672814 792160
rect 672870 792104 672998 792160
rect 673054 792104 673059 792160
rect 672809 792102 673059 792104
rect 672809 792099 672875 792102
rect 672993 792099 673059 792102
rect 39849 778562 39915 778565
rect 40534 778562 40540 778564
rect 39849 778560 40540 778562
rect 39849 778504 39854 778560
rect 39910 778504 40540 778560
rect 39849 778502 40540 778504
rect 39849 778499 39915 778502
rect 40534 778500 40540 778502
rect 40604 778500 40610 778564
rect 39849 772852 39915 772853
rect 39798 772850 39804 772852
rect 39758 772790 39804 772850
rect 39868 772848 39915 772852
rect 39910 772792 39915 772848
rect 39798 772788 39804 772790
rect 39868 772788 39915 772792
rect 39849 772787 39915 772788
rect 673821 772850 673887 772853
rect 675201 772850 675267 772853
rect 673821 772848 675267 772850
rect 673821 772792 673826 772848
rect 673882 772792 675206 772848
rect 675262 772792 675267 772848
rect 673821 772790 675267 772792
rect 673821 772787 673887 772790
rect 675201 772787 675267 772790
rect 39982 769932 39988 769996
rect 40052 769932 40058 769996
rect 39990 769858 40050 769932
rect 40350 769858 40356 769860
rect 39990 769798 40356 769858
rect 40350 769796 40356 769798
rect 40420 769796 40426 769860
rect 40350 761636 40356 761700
rect 40420 761636 40426 761700
rect 40358 761562 40418 761636
rect 41086 761562 41092 761564
rect 40358 761502 41092 761562
rect 41086 761500 41092 761502
rect 41156 761500 41162 761564
rect 41086 758916 41092 758980
rect 41156 758916 41162 758980
rect 40534 758780 40540 758844
rect 40604 758842 40610 758844
rect 41094 758842 41154 758916
rect 40604 758782 41154 758842
rect 40604 758780 40610 758782
rect 40534 739938 40540 739940
rect 40358 739878 40540 739938
rect 40358 739804 40418 739878
rect 40534 739876 40540 739878
rect 40604 739876 40610 739940
rect 40350 739740 40356 739804
rect 40420 739740 40426 739804
rect 672942 721380 672948 721444
rect 673012 721442 673018 721444
rect 673085 721442 673151 721445
rect 673012 721440 673151 721442
rect 673012 721384 673090 721440
rect 673146 721384 673151 721440
rect 673012 721382 673151 721384
rect 673012 721380 673018 721382
rect 673085 721379 673151 721382
rect 40350 720292 40356 720356
rect 40420 720354 40426 720356
rect 40718 720354 40724 720356
rect 40420 720294 40724 720354
rect 40420 720292 40426 720294
rect 40718 720292 40724 720294
rect 40788 720292 40794 720356
rect 672993 714916 673059 714917
rect 672942 714852 672948 714916
rect 673012 714914 673059 714916
rect 673012 714912 673104 714914
rect 673054 714856 673104 714912
rect 673012 714854 673104 714856
rect 673012 714852 673059 714854
rect 672993 714851 673059 714852
rect 40718 701314 40724 701316
rect 40358 701254 40724 701314
rect 40358 701180 40418 701254
rect 40718 701252 40724 701254
rect 40788 701252 40794 701316
rect 40350 701116 40356 701180
rect 40420 701116 40426 701180
rect 673729 685402 673795 685405
rect 675385 685402 675451 685405
rect 673729 685400 675451 685402
rect 673729 685344 673734 685400
rect 673790 685344 675390 685400
rect 675446 685344 675451 685400
rect 673729 685342 675451 685344
rect 673729 685339 673795 685342
rect 675385 685339 675451 685342
rect 40350 681668 40356 681732
rect 40420 681730 40426 681732
rect 40718 681730 40724 681732
rect 40420 681670 40724 681730
rect 40420 681668 40426 681670
rect 40718 681668 40724 681670
rect 40788 681668 40794 681732
rect 40718 662690 40724 662692
rect 40358 662630 40724 662690
rect 40358 662556 40418 662630
rect 40718 662628 40724 662630
rect 40788 662628 40794 662692
rect 40350 662492 40356 662556
rect 40420 662492 40426 662556
rect 40350 598844 40356 598908
rect 40420 598906 40426 598908
rect 40718 598906 40724 598908
rect 40420 598846 40724 598906
rect 40420 598844 40426 598846
rect 40718 598844 40724 598846
rect 40788 598844 40794 598908
rect 40718 579866 40724 579868
rect 40358 579806 40724 579866
rect 40358 579732 40418 579806
rect 40718 579804 40724 579806
rect 40788 579804 40794 579868
rect 40350 579668 40356 579732
rect 40420 579668 40426 579732
rect 40217 550626 40283 550629
rect 40350 550626 40356 550628
rect 40217 550624 40356 550626
rect 40217 550568 40222 550624
rect 40278 550568 40356 550624
rect 40217 550566 40356 550568
rect 40217 550563 40283 550566
rect 40350 550564 40356 550566
rect 40420 550564 40426 550628
rect 40217 546412 40283 546413
rect 40166 546410 40172 546412
rect 40126 546350 40172 546410
rect 40236 546408 40283 546412
rect 40278 546352 40283 546408
rect 40166 546348 40172 546350
rect 40236 546348 40283 546352
rect 40217 546347 40283 546348
rect 40350 540908 40356 540972
rect 40420 540970 40426 540972
rect 40718 540970 40724 540972
rect 40420 540910 40724 540970
rect 40420 540908 40426 540910
rect 40718 540908 40724 540910
rect 40788 540908 40794 540972
rect 40718 521930 40724 521932
rect 40358 521870 40724 521930
rect 40358 521796 40418 521870
rect 40718 521868 40724 521870
rect 40788 521868 40794 521932
rect 40350 521732 40356 521796
rect 40420 521732 40426 521796
rect 672993 514178 673059 514181
rect 673177 514178 673243 514181
rect 672993 514176 677794 514178
rect 672993 514120 672998 514176
rect 673054 514120 673182 514176
rect 673238 514120 677794 514176
rect 672993 514118 677794 514120
rect 672993 514115 673059 514118
rect 673177 514115 673243 514118
rect 677734 514012 677794 514118
rect 673085 511458 673151 511461
rect 673269 511458 673335 511461
rect 673085 511456 677764 511458
rect 673085 511400 673090 511456
rect 673146 511400 673274 511456
rect 673330 511400 677764 511456
rect 673085 511398 677764 511400
rect 673085 511395 673151 511398
rect 673269 511395 673335 511398
rect 672993 509146 673059 509149
rect 672993 509144 677764 509146
rect 672993 509088 672998 509144
rect 673054 509088 677764 509144
rect 672993 509086 677764 509088
rect 672993 509083 673059 509086
rect 40350 508058 40356 508060
rect 39990 507998 40356 508058
rect 39990 507788 40050 507998
rect 40350 507996 40356 507998
rect 40420 507996 40426 508060
rect 39982 507724 39988 507788
rect 40052 507724 40058 507788
rect 44633 493234 44699 493237
rect 39652 493232 44699 493234
rect 39652 493176 44638 493232
rect 44694 493176 44699 493232
rect 39652 493174 44699 493176
rect 39806 492965 39866 493174
rect 44633 493171 44699 493174
rect 39757 492960 39866 492965
rect 39757 492904 39762 492960
rect 39818 492904 39866 492960
rect 39757 492902 39866 492904
rect 39757 492899 39823 492902
rect 44449 488610 44515 488613
rect 39806 488608 44515 488610
rect 39806 488552 44454 488608
rect 44510 488552 44515 488608
rect 39806 488550 44515 488552
rect 39806 488338 39866 488550
rect 44449 488547 44515 488550
rect 39652 488278 39866 488338
rect 677542 480116 677548 480180
rect 677612 480178 677618 480180
rect 678053 480178 678119 480181
rect 677612 480176 678119 480178
rect 677612 480120 678058 480176
rect 678114 480120 678119 480176
rect 677612 480118 678119 480120
rect 677612 480116 677618 480118
rect 678053 480115 678119 480118
rect 677869 469978 677935 469981
rect 677869 469976 678132 469978
rect 677869 469920 677874 469976
rect 677930 469920 678132 469976
rect 677869 469918 678132 469920
rect 677869 469915 677935 469918
rect 673361 467530 673427 467533
rect 673361 467528 678132 467530
rect 673361 467472 673366 467528
rect 673422 467500 678132 467528
rect 673422 467472 678162 467500
rect 673361 467470 678162 467472
rect 673361 467467 673427 467470
rect 678102 465052 678162 467470
rect 672993 463722 673059 463725
rect 673269 463722 673335 463725
rect 672993 463720 673335 463722
rect 672993 463664 672998 463720
rect 673054 463664 673274 463720
rect 673330 463664 673335 463720
rect 672993 463662 673335 463664
rect 672993 463659 673059 463662
rect 673269 463659 673335 463662
rect 39941 455426 40007 455429
rect 40166 455426 40172 455428
rect 39941 455424 40172 455426
rect 39941 455368 39946 455424
rect 40002 455368 40172 455424
rect 39941 455366 40172 455368
rect 39941 455363 40007 455366
rect 40166 455364 40172 455366
rect 40236 455364 40242 455428
rect 39665 451890 39731 451893
rect 40166 451890 40172 451892
rect 39665 451888 40172 451890
rect 39665 451832 39670 451888
rect 39726 451832 40172 451888
rect 39665 451830 40172 451832
rect 39665 451827 39731 451830
rect 40166 451828 40172 451830
rect 40236 451828 40242 451892
rect 44357 448626 44423 448629
rect 39468 448624 44423 448626
rect 39468 448596 44362 448624
rect 39438 448568 44362 448596
rect 44418 448568 44423 448624
rect 39438 448566 44423 448568
rect 39438 446012 39498 448566
rect 44357 448563 44423 448566
rect 39665 441010 39731 441013
rect 39468 441008 39731 441010
rect 39468 440952 39670 441008
rect 39726 440952 39731 441008
rect 39468 440950 39731 440952
rect 39665 440947 39731 440950
rect 673085 427954 673151 427957
rect 677409 427954 677475 427957
rect 673085 427952 677475 427954
rect 673085 427896 673090 427952
rect 673146 427896 677414 427952
rect 677470 427896 677475 427952
rect 673085 427894 677475 427896
rect 673085 427891 673151 427894
rect 677409 427891 677475 427894
rect 677593 425778 677659 425781
rect 677593 425776 677764 425778
rect 677593 425720 677598 425776
rect 677654 425720 677764 425776
rect 677593 425718 677764 425720
rect 677593 425715 677659 425718
rect 673361 420882 673427 420885
rect 673361 420880 677764 420882
rect 673361 420824 673366 420880
rect 673422 420824 677764 420880
rect 673361 420822 677764 420824
rect 673361 420819 673427 420822
rect 672717 392052 672783 392053
rect 672717 392048 672764 392052
rect 672828 392050 672834 392052
rect 672717 391992 672722 392048
rect 672717 391988 672764 391992
rect 672828 391990 672874 392050
rect 672828 391988 672834 391990
rect 672717 391987 672783 391988
rect 672717 386476 672783 386477
rect 672717 386472 672764 386476
rect 672828 386474 672834 386476
rect 672717 386416 672722 386472
rect 672717 386412 672764 386416
rect 672828 386414 672874 386474
rect 672828 386412 672834 386414
rect 672717 386411 672783 386412
rect 673545 338738 673611 338741
rect 675385 338738 675451 338741
rect 673545 338736 675451 338738
rect 673545 338680 673550 338736
rect 673606 338680 675390 338736
rect 675446 338680 675451 338736
rect 673545 338678 675451 338680
rect 673545 338675 673611 338678
rect 675385 338675 675451 338678
rect 672533 295490 672599 295493
rect 672533 295488 672642 295490
rect 672533 295432 672538 295488
rect 672594 295432 672642 295488
rect 672533 295427 672642 295432
rect 672582 295221 672642 295427
rect 672582 295216 672691 295221
rect 672582 295160 672630 295216
rect 672686 295160 672691 295216
rect 672582 295158 672691 295160
rect 672625 295155 672691 295158
rect 673453 293042 673519 293045
rect 675385 293042 675451 293045
rect 673453 293040 675451 293042
rect 673453 292984 673458 293040
rect 673514 292984 675390 293040
rect 675446 292984 675451 293040
rect 673453 292982 675451 292984
rect 673453 292979 673519 292982
rect 675385 292979 675451 292982
rect 41689 275715 41755 275718
rect 42241 275715 42307 275718
rect 41689 275713 42307 275715
rect 41689 275657 41694 275713
rect 41750 275657 42246 275713
rect 42302 275657 42307 275713
rect 41689 275655 42307 275657
rect 41689 275652 41755 275655
rect 42241 275652 42307 275655
rect 673821 212530 673887 212533
rect 674005 212530 674071 212533
rect 673821 212528 674071 212530
rect 673821 212472 673826 212528
rect 673882 212472 674010 212528
rect 674066 212472 674071 212528
rect 673821 212470 674071 212472
rect 673821 212467 673887 212470
rect 674005 212467 674071 212470
rect 672533 193218 672599 193221
rect 672901 193218 672967 193221
rect 672533 193216 672967 193218
rect 672533 193160 672538 193216
rect 672594 193160 672906 193216
rect 672962 193160 672967 193216
rect 672533 193158 672967 193160
rect 672533 193155 672599 193158
rect 672901 193155 672967 193158
rect 41689 184991 41755 184994
rect 42333 184991 42399 184994
rect 41689 184989 42399 184991
rect 41689 184933 41694 184989
rect 41750 184933 42338 184989
rect 42394 184933 42399 184989
rect 41689 184931 42399 184933
rect 41689 184928 41755 184931
rect 42333 184928 42399 184931
rect 39757 120186 39823 120189
rect 44173 120186 44239 120189
rect 39757 120184 44239 120186
rect 39757 120128 39762 120184
rect 39818 120128 44178 120184
rect 44234 120128 44239 120184
rect 39757 120126 44239 120128
rect 39757 120123 39823 120126
rect 44173 120123 44239 120126
rect 41413 115970 41479 115973
rect 42149 115970 42215 115973
rect 39806 115968 42215 115970
rect 39806 115912 41418 115968
rect 41474 115912 42154 115968
rect 42210 115912 42215 115968
rect 39806 115910 42215 115912
rect 39806 115562 39866 115910
rect 41413 115907 41479 115910
rect 42149 115907 42215 115910
rect 39622 115502 39866 115562
rect 39622 115396 39682 115502
rect 44173 110530 44239 110533
rect 45461 110530 45527 110533
rect 39806 110528 45527 110530
rect 39806 110472 44178 110528
rect 44234 110472 45466 110528
rect 45522 110472 45527 110528
rect 39806 110470 45527 110472
rect 39806 110430 39866 110470
rect 44173 110467 44239 110470
rect 45461 110467 45527 110470
rect 39622 110370 39866 110430
rect 39622 110364 39682 110370
rect 39389 84282 39455 84285
rect 40166 84282 40172 84284
rect 39389 84280 40172 84282
rect 39389 84224 39394 84280
rect 39450 84224 40172 84280
rect 39389 84222 40172 84224
rect 39389 84219 39455 84222
rect 40166 84220 40172 84222
rect 40236 84220 40242 84284
rect 44265 75850 44331 75853
rect 39438 75848 44331 75850
rect 39438 75792 44270 75848
rect 44326 75792 44331 75848
rect 39438 75790 44331 75792
rect 39438 75684 39498 75790
rect 44265 75787 44331 75790
rect 44265 73266 44331 73269
rect 39468 73264 44331 73266
rect 39468 73208 44270 73264
rect 44326 73208 44331 73264
rect 39468 73206 44331 73208
rect 44265 73203 44331 73206
rect 44265 68234 44331 68237
rect 45553 68234 45619 68237
rect 39468 68232 45619 68234
rect 39468 68176 44270 68232
rect 44326 68176 45558 68232
rect 45614 68176 45619 68232
rect 39468 68174 45619 68176
rect 44265 68171 44331 68174
rect 45553 68171 45619 68174
rect 425053 47834 425119 47837
rect 430757 47834 430823 47837
rect 425053 47832 430823 47834
rect 425053 47776 425058 47832
rect 425114 47776 430762 47832
rect 430818 47776 430823 47832
rect 425053 47774 430823 47776
rect 425053 47771 425119 47774
rect 430757 47771 430823 47774
rect 460933 47562 460999 47565
rect 461485 47562 461551 47565
rect 480069 47562 480135 47565
rect 460933 47560 480135 47562
rect 460933 47504 460938 47560
rect 460994 47504 461490 47560
rect 461546 47504 480074 47560
rect 480130 47504 480135 47560
rect 460933 47502 480135 47504
rect 460933 47499 460999 47502
rect 461485 47499 461551 47502
rect 480069 47499 480135 47502
rect 483013 47562 483079 47565
rect 488625 47562 488691 47565
rect 483013 47560 488691 47562
rect 483013 47504 483018 47560
rect 483074 47504 488630 47560
rect 488686 47504 488691 47560
rect 483013 47502 488691 47504
rect 483013 47499 483079 47502
rect 488625 47499 488691 47502
rect 328453 47426 328519 47429
rect 334065 47426 334131 47429
rect 328453 47424 334131 47426
rect 328453 47368 328458 47424
rect 328514 47368 334070 47424
rect 334126 47368 334131 47424
rect 328453 47366 334131 47368
rect 328453 47363 328519 47366
rect 334065 47363 334131 47366
rect 289813 47154 289879 47157
rect 303889 47154 303955 47157
rect 309041 47154 309107 47157
rect 289813 47152 309107 47154
rect 289813 47096 289818 47152
rect 289874 47096 303894 47152
rect 303950 47096 309046 47152
rect 309102 47096 309107 47152
rect 289813 47094 309107 47096
rect 289813 47091 289879 47094
rect 303889 47091 303955 47094
rect 309041 47091 309107 47094
rect 290181 41850 290247 41853
rect 297118 41850 297184 41853
rect 299602 41850 299668 41853
rect 305766 41850 305832 41853
rect 305913 41850 305979 41853
rect 290181 41848 300410 41850
rect 290181 41792 290186 41848
rect 290242 41792 297123 41848
rect 297179 41792 299607 41848
rect 299663 41792 300410 41848
rect 290181 41790 300410 41792
rect 290181 41787 290247 41790
rect 297118 41787 297184 41790
rect 299602 41787 299668 41790
rect 300350 41714 300410 41790
rect 305134 41848 305979 41850
rect 305134 41792 305771 41848
rect 305827 41792 305918 41848
rect 305974 41792 305979 41848
rect 305134 41790 305979 41792
rect 305134 41714 305194 41790
rect 305766 41787 305832 41790
rect 305913 41787 305979 41790
rect 300350 41654 305194 41714
rect 622945 40490 623011 40493
rect 84334 40488 623011 40490
rect 84334 40432 622950 40488
rect 623006 40432 623011 40488
rect 84334 40430 623011 40432
rect 84334 40218 84394 40430
rect 622945 40427 623011 40430
rect 149053 40354 149119 40357
rect 145838 40352 149119 40354
rect 145838 40296 149058 40352
rect 149114 40296 149119 40352
rect 145838 40294 149119 40296
rect 84150 40158 84394 40218
rect 86401 40218 86467 40221
rect 86401 40216 86602 40218
rect 86401 40160 86406 40216
rect 86462 40160 86602 40216
rect 86401 40158 86602 40160
rect 84150 39644 84210 40158
rect 86401 40155 86467 40158
rect 86542 39810 86602 40158
rect 86542 39750 88994 39810
rect 86542 39644 86602 39750
rect 88934 39644 88994 39750
rect 141667 38031 141813 39999
rect 145838 39967 145898 40294
rect 149053 40291 149119 40294
rect 569217 40218 569283 40221
rect 579153 40218 579219 40221
rect 569174 40216 579219 40218
rect 569174 40160 569222 40216
rect 569278 40160 579158 40216
rect 579214 40160 579219 40216
rect 569174 40158 579219 40160
rect 569174 40155 569283 40158
rect 579153 40155 579219 40158
rect 632973 40218 633039 40221
rect 634813 40218 634879 40221
rect 632973 40216 634879 40218
rect 632973 40160 632978 40216
rect 633034 40160 634818 40216
rect 634874 40160 634879 40216
rect 632973 40158 634879 40160
rect 632973 40155 633039 40158
rect 634813 40155 634879 40158
rect 240133 39946 240199 39949
rect 253933 39946 253999 39949
rect 240133 39944 246498 39946
rect 240133 39888 240138 39944
rect 240194 39888 246498 39944
rect 240133 39886 246498 39888
rect 240133 39883 240199 39886
rect 241237 39810 241303 39813
rect 242893 39810 242959 39813
rect 241156 39808 242959 39810
rect 241156 39752 241242 39808
rect 241298 39752 242898 39808
rect 242954 39752 242959 39808
rect 241156 39750 242959 39752
rect 241237 39747 241346 39750
rect 242893 39747 242959 39750
rect 241286 39372 241346 39747
rect 246438 39538 246498 39886
rect 248830 39944 253999 39946
rect 248830 39888 253938 39944
rect 253994 39888 253999 39944
rect 248830 39886 253999 39888
rect 248830 39538 248890 39886
rect 253933 39883 253999 39886
rect 569174 39644 569234 40155
rect 622945 39674 623011 39677
rect 622945 39672 623116 39674
rect 622945 39616 622950 39672
rect 623006 39616 623116 39672
rect 622945 39614 623116 39616
rect 622945 39611 623011 39614
rect 246438 39478 248890 39538
rect 246438 39372 246498 39478
rect 248830 39372 248890 39478
<< via3 >>
rect 341012 997596 341076 997660
rect 341012 990252 341076 990316
rect 676260 990116 676324 990180
rect 677548 918580 677612 918644
rect 40172 908108 40236 908172
rect 676260 907700 676324 907764
rect 40356 830724 40420 830788
rect 40540 811608 40604 811612
rect 40540 811552 40554 811608
rect 40554 811552 40604 811608
rect 40540 811548 40604 811552
rect 40356 811276 40420 811340
rect 40908 811140 40972 811204
rect 40540 792100 40604 792164
rect 40908 792100 40972 792164
rect 40540 778500 40604 778564
rect 39804 772848 39868 772852
rect 39804 772792 39854 772848
rect 39854 772792 39868 772848
rect 39804 772788 39868 772792
rect 39988 769932 40052 769996
rect 40356 769796 40420 769860
rect 40356 761636 40420 761700
rect 41092 761500 41156 761564
rect 41092 758916 41156 758980
rect 40540 758780 40604 758844
rect 40540 739876 40604 739940
rect 40356 739740 40420 739804
rect 672948 721380 673012 721444
rect 40356 720292 40420 720356
rect 40724 720292 40788 720356
rect 672948 714912 673012 714916
rect 672948 714856 672998 714912
rect 672998 714856 673012 714912
rect 672948 714852 673012 714856
rect 40724 701252 40788 701316
rect 40356 701116 40420 701180
rect 40356 681668 40420 681732
rect 40724 681668 40788 681732
rect 40724 662628 40788 662692
rect 40356 662492 40420 662556
rect 40356 598844 40420 598908
rect 40724 598844 40788 598908
rect 40724 579804 40788 579868
rect 40356 579668 40420 579732
rect 40356 550564 40420 550628
rect 40172 546408 40236 546412
rect 40172 546352 40222 546408
rect 40222 546352 40236 546408
rect 40172 546348 40236 546352
rect 40356 540908 40420 540972
rect 40724 540908 40788 540972
rect 40724 521868 40788 521932
rect 40356 521732 40420 521796
rect 40356 507996 40420 508060
rect 39988 507724 40052 507788
rect 677548 480116 677612 480180
rect 40172 455364 40236 455428
rect 40172 451828 40236 451892
rect 672764 392048 672828 392052
rect 672764 391992 672778 392048
rect 672778 391992 672828 392048
rect 672764 391988 672828 391992
rect 672764 386472 672828 386476
rect 672764 386416 672778 386472
rect 672778 386416 672828 386472
rect 672764 386412 672828 386416
rect 40172 84220 40236 84284
<< metal4 >>
rect 341011 997660 341077 997661
rect 341011 997596 341012 997660
rect 341076 997596 341077 997660
rect 341011 997595 341077 997596
rect 341014 990317 341074 997595
rect 341011 990316 341077 990317
rect 341011 990252 341012 990316
rect 341076 990252 341077 990316
rect 341011 990251 341077 990252
rect 676259 990180 676325 990181
rect 676259 990116 676260 990180
rect 676324 990116 676325 990180
rect 676259 990115 676325 990116
rect 40171 908172 40237 908173
rect 40171 908108 40172 908172
rect 40236 908108 40237 908172
rect 40171 908107 40237 908108
rect 40174 840170 40234 908107
rect 676262 907765 676322 990115
rect 677547 918644 677613 918645
rect 677547 918580 677548 918644
rect 677612 918580 677613 918644
rect 677547 918579 677613 918580
rect 676259 907764 676325 907765
rect 676259 907700 676260 907764
rect 676324 907700 676325 907764
rect 676259 907699 676325 907700
rect 40174 840110 40418 840170
rect 40358 830789 40418 840110
rect 40355 830788 40421 830789
rect 40355 830724 40356 830788
rect 40420 830724 40421 830788
rect 40355 830723 40421 830724
rect 40539 811612 40605 811613
rect 40539 811610 40540 811612
rect 40358 811550 40540 811610
rect 40358 811341 40418 811550
rect 40539 811548 40540 811550
rect 40604 811548 40605 811612
rect 40539 811547 40605 811548
rect 40355 811340 40421 811341
rect 40355 811276 40356 811340
rect 40420 811276 40421 811340
rect 40355 811275 40421 811276
rect 40907 811204 40973 811205
rect 40907 811140 40908 811204
rect 40972 811140 40973 811204
rect 40907 811139 40973 811140
rect 40910 792165 40970 811139
rect 40539 792164 40605 792165
rect 40539 792100 40540 792164
rect 40604 792100 40605 792164
rect 40539 792099 40605 792100
rect 40907 792164 40973 792165
rect 40907 792100 40908 792164
rect 40972 792100 40973 792164
rect 40907 792099 40973 792100
rect 40542 778565 40602 792099
rect 40539 778564 40605 778565
rect 40539 778500 40540 778564
rect 40604 778500 40605 778564
rect 40539 778499 40605 778500
rect 39803 772852 39869 772853
rect 39803 772788 39804 772852
rect 39868 772850 39869 772852
rect 39868 772790 40050 772850
rect 39868 772788 39869 772790
rect 39803 772787 39869 772788
rect 39990 769997 40050 772790
rect 39987 769996 40053 769997
rect 39987 769932 39988 769996
rect 40052 769932 40053 769996
rect 39987 769931 40053 769932
rect 40355 769860 40421 769861
rect 40355 769796 40356 769860
rect 40420 769796 40421 769860
rect 40355 769795 40421 769796
rect 40358 761701 40418 769795
rect 40355 761700 40421 761701
rect 40355 761636 40356 761700
rect 40420 761636 40421 761700
rect 40355 761635 40421 761636
rect 41091 761564 41157 761565
rect 41091 761500 41092 761564
rect 41156 761500 41157 761564
rect 41091 761499 41157 761500
rect 41094 758981 41154 761499
rect 41091 758980 41157 758981
rect 41091 758916 41092 758980
rect 41156 758916 41157 758980
rect 41091 758915 41157 758916
rect 40539 758844 40605 758845
rect 40539 758780 40540 758844
rect 40604 758780 40605 758844
rect 40539 758779 40605 758780
rect 40542 739941 40602 758779
rect 40539 739940 40605 739941
rect 40539 739876 40540 739940
rect 40604 739876 40605 739940
rect 40539 739875 40605 739876
rect 40355 739804 40421 739805
rect 40355 739740 40356 739804
rect 40420 739740 40421 739804
rect 40355 739739 40421 739740
rect 40358 720357 40418 739739
rect 672947 721444 673013 721445
rect 672947 721380 672948 721444
rect 673012 721380 673013 721444
rect 672947 721379 673013 721380
rect 40355 720356 40421 720357
rect 40355 720292 40356 720356
rect 40420 720292 40421 720356
rect 40355 720291 40421 720292
rect 40723 720356 40789 720357
rect 40723 720292 40724 720356
rect 40788 720292 40789 720356
rect 40723 720291 40789 720292
rect 40726 701317 40786 720291
rect 672950 714917 673010 721379
rect 672947 714916 673013 714917
rect 672947 714852 672948 714916
rect 673012 714852 673013 714916
rect 672947 714851 673013 714852
rect 40723 701316 40789 701317
rect 40723 701252 40724 701316
rect 40788 701252 40789 701316
rect 40723 701251 40789 701252
rect 40355 701180 40421 701181
rect 40355 701116 40356 701180
rect 40420 701116 40421 701180
rect 40355 701115 40421 701116
rect 40358 681733 40418 701115
rect 40355 681732 40421 681733
rect 40355 681668 40356 681732
rect 40420 681668 40421 681732
rect 40355 681667 40421 681668
rect 40723 681732 40789 681733
rect 40723 681668 40724 681732
rect 40788 681668 40789 681732
rect 40723 681667 40789 681668
rect 40726 662693 40786 681667
rect 40723 662692 40789 662693
rect 40723 662628 40724 662692
rect 40788 662628 40789 662692
rect 40723 662627 40789 662628
rect 40355 662556 40421 662557
rect 40355 662492 40356 662556
rect 40420 662492 40421 662556
rect 40355 662491 40421 662492
rect 40358 652490 40418 662491
rect 39990 652430 40418 652490
rect 39990 637530 40050 652430
rect 39990 637470 40418 637530
rect 40358 598909 40418 637470
rect 40355 598908 40421 598909
rect 40355 598844 40356 598908
rect 40420 598844 40421 598908
rect 40355 598843 40421 598844
rect 40723 598908 40789 598909
rect 40723 598844 40724 598908
rect 40788 598844 40789 598908
rect 40723 598843 40789 598844
rect 40726 579869 40786 598843
rect 40723 579868 40789 579869
rect 40723 579804 40724 579868
rect 40788 579804 40789 579868
rect 40723 579803 40789 579804
rect 40355 579732 40421 579733
rect 40355 579668 40356 579732
rect 40420 579668 40421 579732
rect 40355 579667 40421 579668
rect 40358 550629 40418 579667
rect 40355 550628 40421 550629
rect 40355 550564 40356 550628
rect 40420 550564 40421 550628
rect 40355 550563 40421 550564
rect 40171 546412 40237 546413
rect 40171 546348 40172 546412
rect 40236 546348 40237 546412
rect 40171 546347 40237 546348
rect 40174 540970 40234 546347
rect 40355 540972 40421 540973
rect 40355 540970 40356 540972
rect 40174 540910 40356 540970
rect 40355 540908 40356 540910
rect 40420 540908 40421 540972
rect 40355 540907 40421 540908
rect 40723 540972 40789 540973
rect 40723 540908 40724 540972
rect 40788 540908 40789 540972
rect 40723 540907 40789 540908
rect 40726 521933 40786 540907
rect 40723 521932 40789 521933
rect 40723 521868 40724 521932
rect 40788 521868 40789 521932
rect 40723 521867 40789 521868
rect 40355 521796 40421 521797
rect 40355 521732 40356 521796
rect 40420 521732 40421 521796
rect 40355 521731 40421 521732
rect 40358 508061 40418 521731
rect 40355 508060 40421 508061
rect 40355 507996 40356 508060
rect 40420 507996 40421 508060
rect 40355 507995 40421 507996
rect 39987 507788 40053 507789
rect 39987 507724 39988 507788
rect 40052 507724 40053 507788
rect 39987 507723 40053 507724
rect 39990 488610 40050 507723
rect 39990 488550 40234 488610
rect 40174 455429 40234 488550
rect 677550 480181 677610 918579
rect 677547 480180 677613 480181
rect 677547 480116 677548 480180
rect 677612 480116 677613 480180
rect 677547 480115 677613 480116
rect 40171 455428 40237 455429
rect 40171 455364 40172 455428
rect 40236 455364 40237 455428
rect 40171 455363 40237 455364
rect 40171 451892 40237 451893
rect 40171 451828 40172 451892
rect 40236 451828 40237 451892
rect 40171 451827 40237 451828
rect 40174 84285 40234 451827
rect 672763 392052 672829 392053
rect 672763 391988 672764 392052
rect 672828 391988 672829 392052
rect 672763 391987 672829 391988
rect 672766 386477 672826 391987
rect 672763 386476 672829 386477
rect 672763 386412 672764 386476
rect 672828 386412 672829 386476
rect 672763 386411 672829 386412
rect 40171 84284 40237 84285
rect 40171 84220 40172 84284
rect 40236 84220 40237 84284
rect 40171 84219 40237 84220
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334620 1018402 347160 1030924
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 576820 1018402 589360 1030924
rect 628240 1018512 640760 1031002
rect 6598 956440 19088 968960
rect 698512 952840 711002 965360
rect 6086 913863 19572 925191
rect 698028 909409 711514 920737
rect 698512 863640 711002 876160
rect 6675 828820 19197 841360
rect 698402 819640 710924 832180
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 6675 484220 19197 496760
rect 698028 461609 711514 472937
rect 6086 442663 19572 453991
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6675 111420 19197 123960
rect 698512 101240 711002 113760
rect 6086 69863 19572 81191
rect 80040 6675 92580 19197
rect 136713 7143 144149 18309
rect 187640 6598 200160 19088
rect 243009 6086 254337 19572
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 624040 6675 636580 19197
use sky130_ef_io__corner_pad  user1_corner
timestamp 1606493992
transform 1 0 677600 0 1 996800
box -271 -204 40000 40800
use sky130_ef_io__com_bus_slice_5um  FILLER_173
timestamp 1606493992
transform 1 0 676000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_174
timestamp 1606493992
transform 1 0 677000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_175
timestamp 1606493992
transform 1 0 677200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_176
timestamp 1606493992
transform 1 0 677400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_816
timestamp 1606493992
transform 0 1 678007 -1 0 995600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_817
timestamp 1606493992
transform 0 1 678007 -1 0 996600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_818
timestamp 1606493992
transform 0 1 678007 -1 0 996800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_811
timestamp 1606493992
transform 0 1 678007 -1 0 975600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_812
timestamp 1606493992
transform 0 1 678007 -1 0 979600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_813
timestamp 1606493992
transform 0 1 678007 -1 0 983600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_814
timestamp 1606493992
transform 0 1 678007 -1 0 987600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_815
timestamp 1606493992
transform 0 1 678007 -1 0 991600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_164
timestamp 1606493992
transform 1 0 642000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_165
timestamp 1606493992
transform 1 0 646000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_166
timestamp 1606493992
transform 1 0 650000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_167
timestamp 1606493992
transform 1 0 654000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_168
timestamp 1606493992
transform 1 0 658000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_169
timestamp 1606493992
transform 1 0 662000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_170
timestamp 1606493992
transform 1 0 666000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_171
timestamp 1606493992
transform 1 0 670000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_172
timestamp 1606493992
transform 1 0 674000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[15\]
timestamp 1606493992
transform 1 0 626000 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_160
timestamp 1606493992
transform 1 0 624600 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_161
timestamp 1606493992
transform 1 0 625600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_162
timestamp 1606493992
transform 1 0 625800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_156
timestamp 1606493992
transform 1 0 610600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_157
timestamp 1606493992
transform 1 0 614600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_158
timestamp 1606493992
transform 1 0 618600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_159
timestamp 1606493992
transform 1 0 622600 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_152
timestamp 1606493992
transform 1 0 594600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_153
timestamp 1606493992
transform 1 0 598600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_154
timestamp 1606493992
transform 1 0 602600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_155
timestamp 1606493992
transform 1 0 606600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_151
timestamp 1606493992
transform 1 0 590600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_pad  user1_vssa_hvclamp_pad\[0\]
timestamp 1606493992
transform 1 0 575600 0 1 998007
box 0 -434 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_144
timestamp 1606493992
transform 1 0 564200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_145
timestamp 1606493992
transform 1 0 568200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_146
timestamp 1606493992
transform 1 0 572200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_147
timestamp 1606493992
transform 1 0 574200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_148
timestamp 1606493992
transform 1 0 575200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_149
timestamp 1606493992
transform 1 0 575400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_141
timestamp 1606493992
transform 1 0 552200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_142
timestamp 1606493992
transform 1 0 556200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_143
timestamp 1606493992
transform 1 0 560200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_138
timestamp 1606493992
transform 1 0 540200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_139
timestamp 1606493992
transform 1 0 544200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_140
timestamp 1606493992
transform 1 0 548200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[16\]
timestamp 1606493992
transform 1 0 524200 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_134
timestamp 1606493992
transform 1 0 522800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_135
timestamp 1606493992
transform 1 0 523800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_136
timestamp 1606493992
transform 1 0 524000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_130
timestamp 1606493992
transform 1 0 508800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_131
timestamp 1606493992
transform 1 0 512800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_132
timestamp 1606493992
transform 1 0 516800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_133
timestamp 1606493992
transform 1 0 520800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_127
timestamp 1606493992
transform 1 0 496800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_128
timestamp 1606493992
transform 1 0 500800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_129
timestamp 1606493992
transform 1 0 504800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_125
timestamp 1606493992
transform 1 0 488800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_126
timestamp 1606493992
transform 1 0 492800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[17\]
timestamp 1606493992
transform 1 0 472800 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_118
timestamp 1606493992
transform 1 0 465200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_119
timestamp 1606493992
transform 1 0 469200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_120
timestamp 1606493992
transform 1 0 471200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_121
timestamp 1606493992
transform 1 0 472200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_122
timestamp 1606493992
transform 1 0 472400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_123
timestamp 1606493992
transform 1 0 472600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_117
timestamp 1606493992
transform 1 0 461200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_116
timestamp 1606493992
transform 1 0 457200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_115
timestamp 1606493992
transform 1 0 453200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_114
timestamp 1606493992
transform 1 0 449200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_113
timestamp 1606493992
transform 1 0 445200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_112
timestamp 1606493992
transform 1 0 441200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_107
timestamp 1606493992
transform 1 0 434800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_108
timestamp 1606493992
transform 1 0 435000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_0
timestamp 1606493992
transform 1 0 435200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__disconnect_vccd_slice_5um  disconnect_vccd_0
timestamp 1606493992
transform 1 0 436200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_111
timestamp 1606493992
transform 1 0 437200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_105
timestamp 1606493992
transform 1 0 431800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_106
timestamp 1606493992
transform 1 0 433800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_104
timestamp 1606493992
transform 1 0 427800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_103
timestamp 1606493992
transform 1 0 423800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_101
timestamp 1606493992
transform 1 0 415800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_102
timestamp 1606493992
transform 1 0 419800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_97
timestamp 1606493992
transform 1 0 399800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_98
timestamp 1606493992
transform 1 0 403800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_99
timestamp 1606493992
transform 1 0 407800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_100
timestamp 1606493992
transform 1 0 411800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[0\]
timestamp 1606493992
transform 1 0 383800 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_92
timestamp 1606493992
transform 1 0 380400 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_93
timestamp 1606493992
transform 1 0 382400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_94
timestamp 1606493992
transform 1 0 383400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_95
timestamp 1606493992
transform 1 0 383600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_84
timestamp 1606493992
transform 1 0 348400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_85
timestamp 1606493992
transform 1 0 352400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_86
timestamp 1606493992
transform 1 0 356400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_87
timestamp 1606493992
transform 1 0 360400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_88
timestamp 1606493992
transform 1 0 364400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_89
timestamp 1606493992
transform 1 0 368400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_90
timestamp 1606493992
transform 1 0 372400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_91
timestamp 1606493992
transform 1 0 376400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__vssio_hvc_pad  mgmt_vssio_hvclamp_pad\[0\]
timestamp 1606493992
transform 1 0 333400 0 1 998007
box 0 -434 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_78
timestamp 1606493992
transform 1 0 326000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_79
timestamp 1606493992
transform 1 0 330000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_80
timestamp 1606493992
transform 1 0 332000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_81
timestamp 1606493992
transform 1 0 333000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_82
timestamp 1606493992
transform 1 0 333200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_75
timestamp 1606493992
transform 1 0 314000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_76
timestamp 1606493992
transform 1 0 318000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_77
timestamp 1606493992
transform 1 0 322000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_71
timestamp 1606493992
transform 1 0 298000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_72
timestamp 1606493992
transform 1 0 302000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_73
timestamp 1606493992
transform 1 0 306000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_74
timestamp 1606493992
transform 1 0 310000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[1\]
timestamp 1606493992
transform 1 0 282000 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_63
timestamp 1606493992
transform 1 0 270400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_64
timestamp 1606493992
transform 1 0 274400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_65
timestamp 1606493992
transform 1 0 278400 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_66
timestamp 1606493992
transform 1 0 280400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_67
timestamp 1606493992
transform 1 0 281400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_68
timestamp 1606493992
transform 1 0 281600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_69
timestamp 1606493992
transform 1 0 281800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_59
timestamp 1606493992
transform 1 0 254400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_60
timestamp 1606493992
transform 1 0 258400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_61
timestamp 1606493992
transform 1 0 262400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_62
timestamp 1606493992
transform 1 0 266400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_57
timestamp 1606493992
transform 1 0 246400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_58
timestamp 1606493992
transform 1 0 250400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[2\]
timestamp 1606493992
transform 1 0 230400 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_53
timestamp 1606493992
transform 1 0 229000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_54
timestamp 1606493992
transform 1 0 230000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_55
timestamp 1606493992
transform 1 0 230200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_48
timestamp 1606493992
transform 1 0 211000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_49
timestamp 1606493992
transform 1 0 215000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_50
timestamp 1606493992
transform 1 0 219000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_51
timestamp 1606493992
transform 1 0 223000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_52
timestamp 1606493992
transform 1 0 227000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_46
timestamp 1606493992
transform 1 0 203000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_47
timestamp 1606493992
transform 1 0 207000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_44
timestamp 1606493992
transform 1 0 195000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_45
timestamp 1606493992
transform 1 0 199000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[3\]
timestamp 1606493992
transform 1 0 179000 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_38
timestamp 1606493992
transform 1 0 171600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_39
timestamp 1606493992
transform 1 0 175600 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_40
timestamp 1606493992
transform 1 0 177600 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_41
timestamp 1606493992
transform 1 0 178600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_42
timestamp 1606493992
transform 1 0 178800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_35
timestamp 1606493992
transform 1 0 159600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_36
timestamp 1606493992
transform 1 0 163600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_37
timestamp 1606493992
transform 1 0 167600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_31
timestamp 1606493992
transform 1 0 143600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_32
timestamp 1606493992
transform 1 0 147600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_33
timestamp 1606493992
transform 1 0 151600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_34
timestamp 1606493992
transform 1 0 155600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[4\]
timestamp 1606493992
transform 1 0 127600 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_1um  FILLER_28
timestamp 1606493992
transform 1 0 127200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_29
timestamp 1606493992
transform 1 0 127400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_26
timestamp 1606493992
transform 1 0 124200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_27
timestamp 1606493992
transform 1 0 126200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_25
timestamp 1606493992
transform 1 0 120200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_24
timestamp 1606493992
transform 1 0 116200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_23
timestamp 1606493992
transform 1 0 112200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_22
timestamp 1606493992
transform 1 0 108200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_21
timestamp 1606493992
transform 1 0 104200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_20
timestamp 1606493992
transform 1 0 100200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_19
timestamp 1606493992
transform 1 0 96200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_18
timestamp 1606493992
transform 1 0 92200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[5\]
timestamp 1606493992
transform 1 0 76200 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_14
timestamp 1606493992
transform 1 0 74800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_15
timestamp 1606493992
transform 1 0 75800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_16
timestamp 1606493992
transform 1 0 76000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_10
timestamp 1606493992
transform 1 0 60800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_11
timestamp 1606493992
transform 1 0 64800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_12
timestamp 1606493992
transform 1 0 68800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_13
timestamp 1606493992
transform 1 0 72800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_6
timestamp 1606493992
transform 1 0 44800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_7
timestamp 1606493992
transform 1 0 48800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_8
timestamp 1606493992
transform 1 0 52800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_9
timestamp 1606493992
transform 1 0 56800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__corner_pad  user2_corner
timestamp 1606493992
transform 0 -1 40800 1 0 997600
box -271 -204 40000 40800
use sky130_ef_io__com_bus_slice_20um  FILLER_5
timestamp 1606493992
transform 1 0 40800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_608
timestamp 1606493992
transform 0 -1 39593 1 0 994200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_609
timestamp 1606493992
transform 0 -1 39593 1 0 996200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_610
timestamp 1606493992
transform 0 -1 39593 1 0 997200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_611
timestamp 1606493992
transform 0 -1 39593 1 0 997400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_603
timestamp 1606493992
transform 0 -1 39593 1 0 974200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_604
timestamp 1606493992
transform 0 -1 39593 1 0 978200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_605
timestamp 1606493992
transform 0 -1 39593 1 0 982200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_606
timestamp 1606493992
transform 0 -1 39593 1 0 986200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_607
timestamp 1606493992
transform 0 -1 39593 1 0 990200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[14\]
timestamp 1606493992
transform 0 1 675407 -1 0 967600
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_803
timestamp 1606493992
transform 0 1 678007 -1 0 934600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_804
timestamp 1606493992
transform 0 1 678007 -1 0 938600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_805
timestamp 1606493992
transform 0 1 678007 -1 0 942600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_806
timestamp 1606493992
transform 0 1 678007 -1 0 946600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_807
timestamp 1606493992
transform 0 1 678007 -1 0 950600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_808
timestamp 1606493992
transform 0 1 678007 -1 0 951600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_810
timestamp 1606493992
transform 0 1 678007 -1 0 971600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_602
timestamp 1606493992
transform 0 -1 39593 1 0 970200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[6\]
timestamp 1606493992
transform 0 -1 42193 1 0 954200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_597
timestamp 1606493992
transform 0 -1 39593 1 0 947000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_598
timestamp 1606493992
transform 0 -1 39593 1 0 951000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_599
timestamp 1606493992
transform 0 -1 39593 1 0 953000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_600
timestamp 1606493992
transform 0 -1 39593 1 0 954000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_593
timestamp 1606493992
transform 0 -1 39593 1 0 931000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_594
timestamp 1606493992
transform 0 -1 39593 1 0 935000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_595
timestamp 1606493992
transform 0 -1 39593 1 0 939000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_596
timestamp 1606493992
transform 0 -1 39593 1 0 943000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_801
timestamp 1606493992
transform 0 1 678007 -1 0 926600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_802
timestamp 1606493992
transform 0 1 678007 -1 0 930600
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_pad  user1_vccd_lvclamp_pad
timestamp 1606493992
transform 0 1 678007 -1 0 922600
box 0 -46 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_797
timestamp 1606493992
transform 0 1 678007 -1 0 906400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_798
timestamp 1606493992
transform 0 1 678007 -1 0 907400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_799
timestamp 1606493992
transform 0 1 678007 -1 0 907600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_793
timestamp 1606493992
transform 0 1 678007 -1 0 890400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_794
timestamp 1606493992
transform 0 1 678007 -1 0 894400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_795
timestamp 1606493992
transform 0 1 678007 -1 0 898400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_796
timestamp 1606493992
transform 0 1 678007 -1 0 902400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_592
timestamp 1606493992
transform 0 -1 39593 1 0 927000
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_pad  user2_vccd_lvclamp_pad
timestamp 1606493992
transform 0 -1 39593 1 0 912000
box 0 -46 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_587
timestamp 1606493992
transform 0 -1 39593 1 0 904800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_588
timestamp 1606493992
transform 0 -1 39593 1 0 908800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_589
timestamp 1606493992
transform 0 -1 39593 1 0 910800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_590
timestamp 1606493992
transform 0 -1 39593 1 0 911800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_583
timestamp 1606493992
transform 0 -1 39593 1 0 888800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_584
timestamp 1606493992
transform 0 -1 39593 1 0 892800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_585
timestamp 1606493992
transform 0 -1 39593 1 0 896800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_586
timestamp 1606493992
transform 0 -1 39593 1 0 900800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[13\]
timestamp 1606493992
transform 0 1 675407 -1 0 878400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_785
timestamp 1606493992
transform 0 1 678007 -1 0 849400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_786
timestamp 1606493992
transform 0 1 678007 -1 0 853400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_787
timestamp 1606493992
transform 0 1 678007 -1 0 857400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_788
timestamp 1606493992
transform 0 1 678007 -1 0 861400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_789
timestamp 1606493992
transform 0 1 678007 -1 0 862400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_791
timestamp 1606493992
transform 0 1 678007 -1 0 882400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_792
timestamp 1606493992
transform 0 1 678007 -1 0 886400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_582
timestamp 1606493992
transform 0 -1 39593 1 0 884800
box 0 0 4000 39593
use sky130_ef_io__vddio_hvc_pad  mgmt_vddio_hvclamp_pad\[1\]
timestamp 1606493992
transform 0 -1 39593 1 0 869800
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_577
timestamp 1606493992
transform 0 -1 39593 1 0 862600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_578
timestamp 1606493992
transform 0 -1 39593 1 0 866600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_579
timestamp 1606493992
transform 0 -1 39593 1 0 868600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_580
timestamp 1606493992
transform 0 -1 39593 1 0 869600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_573
timestamp 1606493992
transform 0 -1 39593 1 0 846600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_574
timestamp 1606493992
transform 0 -1 39593 1 0 850600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_575
timestamp 1606493992
transform 0 -1 39593 1 0 854600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_576
timestamp 1606493992
transform 0 -1 39593 1 0 858600
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_pad  user1_vdda_hvclamp_pad\[0\]
timestamp 1606493992
transform 0 1 678007 -1 0 833400
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_776
timestamp 1606493992
transform 0 1 678007 -1 0 809200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_777
timestamp 1606493992
transform 0 1 678007 -1 0 813200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_778
timestamp 1606493992
transform 0 1 678007 -1 0 817200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_779
timestamp 1606493992
transform 0 1 678007 -1 0 818200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_780
timestamp 1606493992
transform 0 1 678007 -1 0 818400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_782
timestamp 1606493992
transform 0 1 678007 -1 0 837400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_783
timestamp 1606493992
transform 0 1 678007 -1 0 841400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_784
timestamp 1606493992
transform 0 1 678007 -1 0 845400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_572
timestamp 1606493992
transform 0 -1 39593 1 0 842600
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_pad  user2_vssa_hvclamp_pad
timestamp 1606493992
transform 0 -1 39593 1 0 827600
box 0 -434 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_567
timestamp 1606493992
transform 0 -1 39593 1 0 820400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_568
timestamp 1606493992
transform 0 -1 39593 1 0 824400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_569
timestamp 1606493992
transform 0 -1 39593 1 0 826400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_570
timestamp 1606493992
transform 0 -1 39593 1 0 827400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_563
timestamp 1606493992
transform 0 -1 39593 1 0 804400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_564
timestamp 1606493992
transform 0 -1 39593 1 0 808400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_565
timestamp 1606493992
transform 0 -1 39593 1 0 812400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_566
timestamp 1606493992
transform 0 -1 39593 1 0 816400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[12\]
timestamp 1606493992
transform 0 1 675407 -1 0 789200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_767
timestamp 1606493992
transform 0 1 678007 -1 0 764200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_768
timestamp 1606493992
transform 0 1 678007 -1 0 768200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_769
timestamp 1606493992
transform 0 1 678007 -1 0 772200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_770
timestamp 1606493992
transform 0 1 678007 -1 0 773200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_772
timestamp 1606493992
transform 0 1 678007 -1 0 793200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_773
timestamp 1606493992
transform 0 1 678007 -1 0 797200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_774
timestamp 1606493992
transform 0 1 678007 -1 0 801200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_775
timestamp 1606493992
transform 0 1 678007 -1 0 805200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_562
timestamp 1606493992
transform 0 -1 39593 1 0 800400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[7\]
timestamp 1606493992
transform 0 -1 42193 1 0 784400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_557
timestamp 1606493992
transform 0 -1 39593 1 0 777200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_558
timestamp 1606493992
transform 0 -1 39593 1 0 781200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_559
timestamp 1606493992
transform 0 -1 39593 1 0 783200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_560
timestamp 1606493992
transform 0 -1 39593 1 0 784200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_553
timestamp 1606493992
transform 0 -1 39593 1 0 761200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_554
timestamp 1606493992
transform 0 -1 39593 1 0 765200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_555
timestamp 1606493992
transform 0 -1 39593 1 0 769200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_556
timestamp 1606493992
transform 0 -1 39593 1 0 773200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[11\]
timestamp 1606493992
transform 0 1 675407 -1 0 744200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_759
timestamp 1606493992
transform 0 1 678007 -1 0 723200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_760
timestamp 1606493992
transform 0 1 678007 -1 0 727200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_761
timestamp 1606493992
transform 0 1 678007 -1 0 728200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_763
timestamp 1606493992
transform 0 1 678007 -1 0 748200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_764
timestamp 1606493992
transform 0 1 678007 -1 0 752200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_765
timestamp 1606493992
transform 0 1 678007 -1 0 756200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_766
timestamp 1606493992
transform 0 1 678007 -1 0 760200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_552
timestamp 1606493992
transform 0 -1 39593 1 0 757200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[8\]
timestamp 1606493992
transform 0 -1 42193 1 0 741200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_547
timestamp 1606493992
transform 0 -1 39593 1 0 734000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_548
timestamp 1606493992
transform 0 -1 39593 1 0 738000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_549
timestamp 1606493992
transform 0 -1 39593 1 0 740000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_550
timestamp 1606493992
transform 0 -1 39593 1 0 741000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_543
timestamp 1606493992
transform 0 -1 39593 1 0 718000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_544
timestamp 1606493992
transform 0 -1 39593 1 0 722000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_545
timestamp 1606493992
transform 0 -1 39593 1 0 726000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_546
timestamp 1606493992
transform 0 -1 39593 1 0 730000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[10\]
timestamp 1606493992
transform 0 1 675407 -1 0 699200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_750
timestamp 1606493992
transform 0 1 678007 -1 0 682000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_751
timestamp 1606493992
transform 0 1 678007 -1 0 683000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_752
timestamp 1606493992
transform 0 1 678007 -1 0 683200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_754
timestamp 1606493992
transform 0 1 678007 -1 0 703200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_755
timestamp 1606493992
transform 0 1 678007 -1 0 707200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_756
timestamp 1606493992
transform 0 1 678007 -1 0 711200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_757
timestamp 1606493992
transform 0 1 678007 -1 0 715200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_758
timestamp 1606493992
transform 0 1 678007 -1 0 719200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[9\]
timestamp 1606493992
transform 0 -1 42193 1 0 698000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_534
timestamp 1606493992
transform 0 -1 39593 1 0 678800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_535
timestamp 1606493992
transform 0 -1 39593 1 0 682800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_536
timestamp 1606493992
transform 0 -1 39593 1 0 686800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_537
timestamp 1606493992
transform 0 -1 39593 1 0 690800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_538
timestamp 1606493992
transform 0 -1 39593 1 0 694800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_539
timestamp 1606493992
transform 0 -1 39593 1 0 696800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_540
timestamp 1606493992
transform 0 -1 39593 1 0 697800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_542
timestamp 1606493992
transform 0 -1 39593 1 0 714000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[9\]
timestamp 1606493992
transform 0 1 675407 -1 0 654000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_741
timestamp 1606493992
transform 0 1 678007 -1 0 637000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_742
timestamp 1606493992
transform 0 1 678007 -1 0 638000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_744
timestamp 1606493992
transform 0 1 678007 -1 0 658000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_745
timestamp 1606493992
transform 0 1 678007 -1 0 662000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_746
timestamp 1606493992
transform 0 1 678007 -1 0 666000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_747
timestamp 1606493992
transform 0 1 678007 -1 0 670000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_748
timestamp 1606493992
transform 0 1 678007 -1 0 674000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_749
timestamp 1606493992
transform 0 1 678007 -1 0 678000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_532
timestamp 1606493992
transform 0 -1 39593 1 0 670800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_533
timestamp 1606493992
transform 0 -1 39593 1 0 674800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[10\]
timestamp 1606493992
transform 0 -1 42193 1 0 654800
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_528
timestamp 1606493992
transform 0 -1 39593 1 0 651600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_529
timestamp 1606493992
transform 0 -1 39593 1 0 653600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_530
timestamp 1606493992
transform 0 -1 39593 1 0 654600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_524
timestamp 1606493992
transform 0 -1 39593 1 0 635600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_525
timestamp 1606493992
transform 0 -1 39593 1 0 639600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_526
timestamp 1606493992
transform 0 -1 39593 1 0 643600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_527
timestamp 1606493992
transform 0 -1 39593 1 0 647600
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[8\]
timestamp 1606493992
transform 0 1 675407 -1 0 609000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_732
timestamp 1606493992
transform 0 1 678007 -1 0 592800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_733
timestamp 1606493992
transform 0 1 678007 -1 0 593000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_735
timestamp 1606493992
transform 0 1 678007 -1 0 613000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_736
timestamp 1606493992
transform 0 1 678007 -1 0 617000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_737
timestamp 1606493992
transform 0 1 678007 -1 0 621000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_738
timestamp 1606493992
transform 0 1 678007 -1 0 625000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_739
timestamp 1606493992
transform 0 1 678007 -1 0 629000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_740
timestamp 1606493992
transform 0 1 678007 -1 0 633000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_522
timestamp 1606493992
transform 0 -1 39593 1 0 627600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_523
timestamp 1606493992
transform 0 -1 39593 1 0 631600
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[11\]
timestamp 1606493992
transform 0 -1 42193 1 0 611600
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_518
timestamp 1606493992
transform 0 -1 39593 1 0 608400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_519
timestamp 1606493992
transform 0 -1 39593 1 0 610400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_520
timestamp 1606493992
transform 0 -1 39593 1 0 611400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_514
timestamp 1606493992
transform 0 -1 39593 1 0 592400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_515
timestamp 1606493992
transform 0 -1 39593 1 0 596400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_516
timestamp 1606493992
transform 0 -1 39593 1 0 600400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_517
timestamp 1606493992
transform 0 -1 39593 1 0 604400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_725
timestamp 1606493992
transform 0 1 678007 -1 0 567800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_726
timestamp 1606493992
transform 0 1 678007 -1 0 571800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_727
timestamp 1606493992
transform 0 1 678007 -1 0 575800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_728
timestamp 1606493992
transform 0 1 678007 -1 0 579800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_729
timestamp 1606493992
transform 0 1 678007 -1 0 583800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_730
timestamp 1606493992
transform 0 1 678007 -1 0 587800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_731
timestamp 1606493992
transform 0 1 678007 -1 0 591800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_512
timestamp 1606493992
transform 0 -1 39593 1 0 584400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_513
timestamp 1606493992
transform 0 -1 39593 1 0 588400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[12\]
timestamp 1606493992
transform 0 -1 42193 1 0 568400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_508
timestamp 1606493992
transform 0 -1 39593 1 0 565200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_509
timestamp 1606493992
transform 0 -1 39593 1 0 567200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_510
timestamp 1606493992
transform 0 -1 39593 1 0 568200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_504
timestamp 1606493992
transform 0 -1 39593 1 0 549200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_505
timestamp 1606493992
transform 0 -1 39593 1 0 553200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_506
timestamp 1606493992
transform 0 -1 39593 1 0 557200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_507
timestamp 1606493992
transform 0 -1 39593 1 0 561200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[7\]
timestamp 1606493992
transform 0 1 675407 -1 0 563800
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_716
timestamp 1606493992
transform 0 1 678007 -1 0 522800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_717
timestamp 1606493992
transform 0 1 678007 -1 0 526800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_718
timestamp 1606493992
transform 0 1 678007 -1 0 530800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_719
timestamp 1606493992
transform 0 1 678007 -1 0 534800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_720
timestamp 1606493992
transform 0 1 678007 -1 0 538800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_721
timestamp 1606493992
transform 0 1 678007 -1 0 542800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_722
timestamp 1606493992
transform 0 1 678007 -1 0 546800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_723
timestamp 1606493992
transform 0 1 678007 -1 0 547800
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[13\]
timestamp 1606493992
transform 0 -1 42193 1 0 525200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_495
timestamp 1606493992
transform 0 -1 39593 1 0 510000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_496
timestamp 1606493992
transform 0 -1 39593 1 0 514000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_497
timestamp 1606493992
transform 0 -1 39593 1 0 518000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_498
timestamp 1606493992
transform 0 -1 39593 1 0 522000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_499
timestamp 1606493992
transform 0 -1 39593 1 0 524000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_500
timestamp 1606493992
transform 0 -1 39593 1 0 525000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_502
timestamp 1606493992
transform 0 -1 39593 1 0 541200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_503
timestamp 1606493992
transform 0 -1 39593 1 0 545200
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_pad  user1_vdda_hvclamp_pad\[1\]
timestamp 1606493992
transform 0 1 678007 -1 0 518800
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_707
timestamp 1606493992
transform 0 1 678007 -1 0 478800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_708
timestamp 1606493992
transform 0 1 678007 -1 0 482800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_709
timestamp 1606493992
transform 0 1 678007 -1 0 486800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_710
timestamp 1606493992
transform 0 1 678007 -1 0 490800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_711
timestamp 1606493992
transform 0 1 678007 -1 0 494800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_712
timestamp 1606493992
transform 0 1 678007 -1 0 498800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_713
timestamp 1606493992
transform 0 1 678007 -1 0 502800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_714
timestamp 1606493992
transform 0 1 678007 -1 0 503800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_492
timestamp 1606493992
transform 0 -1 39593 1 0 498000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_493
timestamp 1606493992
transform 0 -1 39593 1 0 502000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_494
timestamp 1606493992
transform 0 -1 39593 1 0 506000
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_pad  user2_vdda_hvclamp_pad
timestamp 1606493992
transform 0 -1 39593 1 0 483000
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_488
timestamp 1606493992
transform 0 -1 39593 1 0 479800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_489
timestamp 1606493992
transform 0 -1 39593 1 0 481800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_490
timestamp 1606493992
transform 0 -1 39593 1 0 482800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_485
timestamp 1606493992
transform 0 -1 39593 1 0 467800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_486
timestamp 1606493992
transform 0 -1 39593 1 0 471800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_487
timestamp 1606493992
transform 0 -1 39593 1 0 475800
box 0 0 4000 39593
use sky130_ef_io__vssd_lvc_pad  user1_vssd_lvclmap_pad
timestamp 1606493992
transform 0 1 678007 -1 0 474800
box 0 -46 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_703
timestamp 1606493992
transform 0 1 678007 -1 0 458600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_704
timestamp 1606493992
transform 0 1 678007 -1 0 459600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_705
timestamp 1606493992
transform 0 1 678007 -1 0 459800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_699
timestamp 1606493992
transform 0 1 678007 -1 0 442600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_700
timestamp 1606493992
transform 0 1 678007 -1 0 446600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_701
timestamp 1606493992
transform 0 1 678007 -1 0 450600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_702
timestamp 1606493992
transform 0 1 678007 -1 0 454600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_697
timestamp 1606493992
transform 0 1 678007 -1 0 434600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_698
timestamp 1606493992
transform 0 1 678007 -1 0 438600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_482
timestamp 1606493992
transform 0 -1 39593 1 0 455800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_483
timestamp 1606493992
transform 0 -1 39593 1 0 459800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_484
timestamp 1606493992
transform 0 -1 39593 1 0 463800
box 0 0 4000 39593
use sky130_ef_io__vssd_lvc_pad  user2_vssd_lvclmap_pad
timestamp 1606493992
transform 0 -1 39593 1 0 440800
box 0 -46 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_478
timestamp 1606493992
transform 0 -1 39593 1 0 437600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_479
timestamp 1606493992
transform 0 -1 39593 1 0 439600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_480
timestamp 1606493992
transform 0 -1 39593 1 0 440600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_475
timestamp 1606493992
transform 0 -1 39593 1 0 425600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_476
timestamp 1606493992
transform 0 -1 39593 1 0 429600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_477
timestamp 1606493992
transform 0 -1 39593 1 0 433600
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_pad  user1_vssa_hvclamp_pad\[1\]
timestamp 1606493992
transform 0 1 678007 -1 0 430600
box 0 -434 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_688
timestamp 1606493992
transform 0 1 678007 -1 0 390600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_689
timestamp 1606493992
transform 0 1 678007 -1 0 394600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_690
timestamp 1606493992
transform 0 1 678007 -1 0 398600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_691
timestamp 1606493992
transform 0 1 678007 -1 0 402600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_692
timestamp 1606493992
transform 0 1 678007 -1 0 406600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_693
timestamp 1606493992
transform 0 1 678007 -1 0 410600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_694
timestamp 1606493992
transform 0 1 678007 -1 0 414600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_695
timestamp 1606493992
transform 0 1 678007 -1 0 415600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_472
timestamp 1606493992
transform 0 -1 39593 1 0 413600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_473
timestamp 1606493992
transform 0 -1 39593 1 0 417600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_474
timestamp 1606493992
transform 0 -1 39593 1 0 421600
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[14\]
timestamp 1606493992
transform 0 -1 42193 1 0 397600
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_469
timestamp 1606493992
transform 0 -1 39593 1 0 396400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_470
timestamp 1606493992
transform 0 -1 39593 1 0 397400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_465
timestamp 1606493992
transform 0 -1 39593 1 0 382400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_466
timestamp 1606493992
transform 0 -1 39593 1 0 386400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_467
timestamp 1606493992
transform 0 -1 39593 1 0 390400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_468
timestamp 1606493992
transform 0 -1 39593 1 0 394400
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[6\]
timestamp 1606493992
transform 0 1 675407 -1 0 386600
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_1um  FILLER_686
timestamp 1606493992
transform 0 1 678007 -1 0 370600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_682
timestamp 1606493992
transform 0 1 678007 -1 0 361400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_683
timestamp 1606493992
transform 0 1 678007 -1 0 365400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_684
timestamp 1606493992
transform 0 1 678007 -1 0 369400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_685
timestamp 1606493992
transform 0 1 678007 -1 0 370400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_678
timestamp 1606493992
transform 0 1 678007 -1 0 345400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_679
timestamp 1606493992
transform 0 1 678007 -1 0 349400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_680
timestamp 1606493992
transform 0 1 678007 -1 0 353400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_681
timestamp 1606493992
transform 0 1 678007 -1 0 357400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_462
timestamp 1606493992
transform 0 -1 39593 1 0 370400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_463
timestamp 1606493992
transform 0 -1 39593 1 0 374400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_464
timestamp 1606493992
transform 0 -1 39593 1 0 378400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[15\]
timestamp 1606493992
transform 0 -1 42193 1 0 354400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_1um  FILLER_460
timestamp 1606493992
transform 0 -1 39593 1 0 354200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_455
timestamp 1606493992
transform 0 -1 39593 1 0 339200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_456
timestamp 1606493992
transform 0 -1 39593 1 0 343200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_457
timestamp 1606493992
transform 0 -1 39593 1 0 347200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_458
timestamp 1606493992
transform 0 -1 39593 1 0 351200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_459
timestamp 1606493992
transform 0 -1 39593 1 0 353200
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[5\]
timestamp 1606493992
transform 0 1 675407 -1 0 341400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_669
timestamp 1606493992
transform 0 1 678007 -1 0 300400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_670
timestamp 1606493992
transform 0 1 678007 -1 0 304400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_671
timestamp 1606493992
transform 0 1 678007 -1 0 308400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_672
timestamp 1606493992
transform 0 1 678007 -1 0 312400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_673
timestamp 1606493992
transform 0 1 678007 -1 0 316400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_674
timestamp 1606493992
transform 0 1 678007 -1 0 320400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_675
timestamp 1606493992
transform 0 1 678007 -1 0 324400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_676
timestamp 1606493992
transform 0 1 678007 -1 0 325400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_453
timestamp 1606493992
transform 0 -1 39593 1 0 331200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_454
timestamp 1606493992
transform 0 -1 39593 1 0 335200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_452
timestamp 1606493992
transform 0 -1 39593 1 0 327200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[16\]
timestamp 1606493992
transform 0 -1 42193 1 0 311200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_445
timestamp 1606493992
transform 0 -1 39593 1 0 296000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_446
timestamp 1606493992
transform 0 -1 39593 1 0 300000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_447
timestamp 1606493992
transform 0 -1 39593 1 0 304000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_448
timestamp 1606493992
transform 0 -1 39593 1 0 308000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_449
timestamp 1606493992
transform 0 -1 39593 1 0 310000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_450
timestamp 1606493992
transform 0 -1 39593 1 0 311000
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[4\]
timestamp 1606493992
transform 0 1 675407 -1 0 296400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_661
timestamp 1606493992
transform 0 1 678007 -1 0 259400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_662
timestamp 1606493992
transform 0 1 678007 -1 0 263400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_663
timestamp 1606493992
transform 0 1 678007 -1 0 267400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_664
timestamp 1606493992
transform 0 1 678007 -1 0 271400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_665
timestamp 1606493992
transform 0 1 678007 -1 0 275400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_666
timestamp 1606493992
transform 0 1 678007 -1 0 279400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_667
timestamp 1606493992
transform 0 1 678007 -1 0 280400
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[17\]
timestamp 1606493992
transform 0 -1 42193 1 0 268000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_436
timestamp 1606493992
transform 0 -1 39593 1 0 256800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_437
timestamp 1606493992
transform 0 -1 39593 1 0 260800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_438
timestamp 1606493992
transform 0 -1 39593 1 0 264800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_439
timestamp 1606493992
transform 0 -1 39593 1 0 266800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_440
timestamp 1606493992
transform 0 -1 39593 1 0 267800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_442
timestamp 1606493992
transform 0 -1 39593 1 0 284000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_443
timestamp 1606493992
transform 0 -1 39593 1 0 288000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_444
timestamp 1606493992
transform 0 -1 39593 1 0 292000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[3\]
timestamp 1606493992
transform 0 1 675407 -1 0 251400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_652
timestamp 1606493992
transform 0 1 678007 -1 0 218200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_653
timestamp 1606493992
transform 0 1 678007 -1 0 222200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_654
timestamp 1606493992
transform 0 1 678007 -1 0 226200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_655
timestamp 1606493992
transform 0 1 678007 -1 0 230200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_656
timestamp 1606493992
transform 0 1 678007 -1 0 234200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_657
timestamp 1606493992
transform 0 1 678007 -1 0 235200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_658
timestamp 1606493992
transform 0 1 678007 -1 0 235400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_660
timestamp 1606493992
transform 0 1 678007 -1 0 255400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_433
timestamp 1606493992
transform 0 -1 39593 1 0 244800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_434
timestamp 1606493992
transform 0 -1 39593 1 0 248800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_435
timestamp 1606493992
transform 0 -1 39593 1 0 252800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_432
timestamp 1606493992
transform 0 -1 39593 1 0 240800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[18\]
timestamp 1606493992
transform 0 -1 42193 1 0 224800
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_426
timestamp 1606493992
transform 0 -1 39593 1 0 213600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_427
timestamp 1606493992
transform 0 -1 39593 1 0 217600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_428
timestamp 1606493992
transform 0 -1 39593 1 0 221600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_429
timestamp 1606493992
transform 0 -1 39593 1 0 223600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_430
timestamp 1606493992
transform 0 -1 39593 1 0 224600
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[2\]
timestamp 1606493992
transform 0 1 675407 -1 0 206200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_643
timestamp 1606493992
transform 0 1 678007 -1 0 173200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_644
timestamp 1606493992
transform 0 1 678007 -1 0 177200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_645
timestamp 1606493992
transform 0 1 678007 -1 0 181200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_646
timestamp 1606493992
transform 0 1 678007 -1 0 185200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_647
timestamp 1606493992
transform 0 1 678007 -1 0 189200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_648
timestamp 1606493992
transform 0 1 678007 -1 0 190200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_650
timestamp 1606493992
transform 0 1 678007 -1 0 210200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_651
timestamp 1606493992
transform 0 1 678007 -1 0 214200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_423
timestamp 1606493992
transform 0 -1 39593 1 0 201600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_424
timestamp 1606493992
transform 0 -1 39593 1 0 205600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_425
timestamp 1606493992
transform 0 -1 39593 1 0 209600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_422
timestamp 1606493992
transform 0 -1 39593 1 0 197600
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[19\]
timestamp 1606493992
transform 0 -1 42193 1 0 181600
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_416
timestamp 1606493992
transform 0 -1 39593 1 0 170400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_417
timestamp 1606493992
transform 0 -1 39593 1 0 174400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_418
timestamp 1606493992
transform 0 -1 39593 1 0 178400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_419
timestamp 1606493992
transform 0 -1 39593 1 0 180400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_420
timestamp 1606493992
transform 0 -1 39593 1 0 181400
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[1\]
timestamp 1606493992
transform 0 1 675407 -1 0 161200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_634
timestamp 1606493992
transform 0 1 678007 -1 0 132000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_635
timestamp 1606493992
transform 0 1 678007 -1 0 136000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_636
timestamp 1606493992
transform 0 1 678007 -1 0 140000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_637
timestamp 1606493992
transform 0 1 678007 -1 0 144000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_638
timestamp 1606493992
transform 0 1 678007 -1 0 145000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_639
timestamp 1606493992
transform 0 1 678007 -1 0 145200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_641
timestamp 1606493992
transform 0 1 678007 -1 0 165200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_642
timestamp 1606493992
transform 0 1 678007 -1 0 169200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_415
timestamp 1606493992
transform 0 -1 39593 1 0 166400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_414
timestamp 1606493992
transform 0 -1 39593 1 0 162400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_413
timestamp 1606493992
transform 0 -1 39593 1 0 158400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_408
timestamp 1606493992
transform 0 -1 39593 1 0 151200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_409
timestamp 1606493992
transform 0 -1 39593 1 0 152200
box 0 0 200 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_2
timestamp 1606493992
transform 0 -1 39593 1 0 152400
box 0 0 1000 39593
use sky130_ef_io__disconnect_vccd_slice_5um  disconnect_vccd_2
timestamp 1606493992
transform 0 -1 39593 1 0 153400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_412
timestamp 1606493992
transform 0 -1 39593 1 0 154400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_407
timestamp 1606493992
transform 0 -1 39593 1 0 149200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_406
timestamp 1606493992
transform 0 -1 39593 1 0 145200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_405
timestamp 1606493992
transform 0 -1 39593 1 0 141200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_404
timestamp 1606493992
transform 0 -1 39593 1 0 137200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_403
timestamp 1606493992
transform 0 -1 39593 1 0 133200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_402
timestamp 1606493992
transform 0 -1 39593 1 0 129200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[0\]
timestamp 1606493992
transform 0 1 675407 -1 0 116000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_626
timestamp 1606493992
transform 0 1 678007 -1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_627
timestamp 1606493992
transform 0 1 678007 -1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_628
timestamp 1606493992
transform 0 1 678007 -1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_629
timestamp 1606493992
transform 0 1 678007 -1 0 100000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_631
timestamp 1606493992
transform 0 1 678007 -1 0 120000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_632
timestamp 1606493992
transform 0 1 678007 -1 0 124000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_633
timestamp 1606493992
transform 0 1 678007 -1 0 128000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_401
timestamp 1606493992
transform 0 -1 39593 1 0 125200
box 0 0 4000 39593
use sky130_ef_io__vddio_hvc_pad  mgmt_vddio_hvclamp_pad\[0\]
timestamp 1606493992
transform 0 -1 39593 1 0 110200
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_396
timestamp 1606493992
transform 0 -1 39593 1 0 103000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_397
timestamp 1606493992
transform 0 -1 39593 1 0 107000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_398
timestamp 1606493992
transform 0 -1 39593 1 0 109000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_399
timestamp 1606493992
transform 0 -1 39593 1 0 110000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_392
timestamp 1606493992
transform 0 -1 39593 1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_393
timestamp 1606493992
transform 0 -1 39593 1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_394
timestamp 1606493992
transform 0 -1 39593 1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_395
timestamp 1606493992
transform 0 -1 39593 1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_625
timestamp 1606493992
transform 0 1 678007 -1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_624
timestamp 1606493992
transform 0 1 678007 -1 0 83000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_623
timestamp 1606493992
transform 0 1 678007 -1 0 79000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_622
timestamp 1606493992
transform 0 1 678007 -1 0 75000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_619
timestamp 1606493992
transform 0 1 678007 -1 0 69000
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_1
timestamp 1606493992
transform 0 1 678007 -1 0 70000
box 0 0 1000 39593
use sky130_ef_io__disconnect_vccd_slice_5um  disconnect_vccd_1
timestamp 1606493992
transform 0 1 678007 -1 0 71000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_618
timestamp 1606493992
transform 0 1 678007 -1 0 68000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_617
timestamp 1606493992
transform 0 1 678007 -1 0 64000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_616
timestamp 1606493992
transform 0 1 678007 -1 0 60000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_615
timestamp 1606493992
transform 0 1 678007 -1 0 56000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_614
timestamp 1606493992
transform 0 1 678007 -1 0 52000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_613
timestamp 1606493992
transform 0 1 678007 -1 0 48000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_391
timestamp 1606493992
transform 0 -1 39593 1 0 83000
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_pad  mgmt_vccd_lvclamp_pad
timestamp 1606493992
transform 0 -1 39593 1 0 68000
box 0 -46 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_386
timestamp 1606493992
transform 0 -1 39593 1 0 60800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_387
timestamp 1606493992
transform 0 -1 39593 1 0 64800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_388
timestamp 1606493992
transform 0 -1 39593 1 0 66800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_389
timestamp 1606493992
transform 0 -1 39593 1 0 67800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_382
timestamp 1606493992
transform 0 -1 39593 1 0 44800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_383
timestamp 1606493992
transform 0 -1 39593 1 0 48800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_384
timestamp 1606493992
transform 0 -1 39593 1 0 52800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_385
timestamp 1606493992
transform 0 -1 39593 1 0 56800
box 0 0 4000 39593
use sky130_ef_io__corner_pad  mgmt_corner\[1\]
timestamp 1606493992
transform 0 1 676800 -1 0 40000
box -271 -204 40000 40800
use sky130_ef_io__com_bus_slice_5um  FILLER_377
timestamp 1606493992
transform -1 0 676200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_378
timestamp 1606493992
transform -1 0 676400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_379
timestamp 1606493992
transform -1 0 676600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_380
timestamp 1606493992
transform -1 0 676800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_612
timestamp 1606493992
transform 0 1 678007 -1 0 44000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_376
timestamp 1606493992
transform -1 0 675200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_375
timestamp 1606493992
transform -1 0 673200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_72
timestamp 1606493992
transform -1 0 669200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_71
timestamp 1606493992
transform -1 0 665200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_70
timestamp 1606493992
transform -1 0 661200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_69
timestamp 1606493992
transform -1 0 657200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_68
timestamp 1606493992
transform -1 0 653200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_368
timestamp 1606493992
transform -1 0 645200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_67
timestamp 1606493992
transform -1 0 649200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_365
timestamp 1606493992
transform -1 0 643800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_366
timestamp 1606493992
transform -1 0 644800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_367
timestamp 1606493992
transform -1 0 645000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_364
timestamp 1606493992
transform -1 0 641800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_pad  mgmt_vdda_hvclamp_pad
timestamp 1606493992
transform -1 0 637800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_360
timestamp 1606493992
transform -1 0 622400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_361
timestamp 1606493992
transform -1 0 622600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_362
timestamp 1606493992
transform -1 0 622800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_65
timestamp 1606493992
transform -1 0 611400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_66
timestamp 1606493992
transform -1 0 615400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_358
timestamp 1606493992
transform -1 0 619400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_359
timestamp 1606493992
transform -1 0 621400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_350
timestamp 1606493992
transform -1 0 591200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_351
timestamp 1606493992
transform -1 0 591400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_61
timestamp 1606493992
transform -1 0 595400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_62
timestamp 1606493992
transform -1 0 599400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_63
timestamp 1606493992
transform -1 0 603400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_64
timestamp 1606493992
transform -1 0 607400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_347
timestamp 1606493992
transform -1 0 588000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_348
timestamp 1606493992
transform -1 0 590000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_349
timestamp 1606493992
transform -1 0 591000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__vssio_hvc_pad  mgmt_vssio_hvclamp_pad\[1\]
timestamp 1606493992
transform -1 0 584000 0 -1 39593
box 0 -434 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_342
timestamp 1606493992
transform -1 0 567600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_343
timestamp 1606493992
transform -1 0 568600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_344
timestamp 1606493992
transform -1 0 568800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_345
timestamp 1606493992
transform -1 0 569000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_58
timestamp 1606493992
transform -1 0 553600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_59
timestamp 1606493992
transform -1 0 557600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_60
timestamp 1606493992
transform -1 0 561600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_341
timestamp 1606493992
transform -1 0 565600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_56
timestamp 1606493992
transform -1 0 545600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_57
timestamp 1606493992
transform -1 0 549600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_330
timestamp 1606493992
transform -1 0 534200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_331
timestamp 1606493992
transform -1 0 536200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_332
timestamp 1606493992
transform -1 0 537200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_333
timestamp 1606493992
transform -1 0 537400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_334
timestamp 1606493992
transform -1 0 537600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_55
timestamp 1606493992
transform -1 0 541600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  gpio_pad
timestamp 1606493992
transform -1 0 530200 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_324
timestamp 1606493992
transform -1 0 510800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_325
timestamp 1606493992
transform -1 0 512800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_326
timestamp 1606493992
transform -1 0 513800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_327
timestamp 1606493992
transform -1 0 514000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_328
timestamp 1606493992
transform -1 0 514200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_54
timestamp 1606493992
transform -1 0 506800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_53
timestamp 1606493992
transform -1 0 502800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_52
timestamp 1606493992
transform -1 0 498800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_51
timestamp 1606493992
transform -1 0 494800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_50
timestamp 1606493992
transform -1 0 490800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_315
timestamp 1606493992
transform -1 0 482400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_316
timestamp 1606493992
transform -1 0 482600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_317
timestamp 1606493992
transform -1 0 482800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_49
timestamp 1606493992
transform -1 0 486800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_314
timestamp 1606493992
transform -1 0 481400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_313
timestamp 1606493992
transform -1 0 479400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_io1_pad
timestamp 1606493992
transform -1 0 475400 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_308
timestamp 1606493992
transform -1 0 458000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_309
timestamp 1606493992
transform -1 0 459000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_310
timestamp 1606493992
transform -1 0 459200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_311
timestamp 1606493992
transform -1 0 459400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_46
timestamp 1606493992
transform -1 0 444000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_47
timestamp 1606493992
transform -1 0 448000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_48
timestamp 1606493992
transform -1 0 452000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_307
timestamp 1606493992
transform -1 0 456000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_297
timestamp 1606493992
transform -1 0 426600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_298
timestamp 1606493992
transform -1 0 427600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_299
timestamp 1606493992
transform -1 0 427800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_300
timestamp 1606493992
transform -1 0 428000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_43
timestamp 1606493992
transform -1 0 432000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_44
timestamp 1606493992
transform -1 0 436000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_45
timestamp 1606493992
transform -1 0 440000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_296
timestamp 1606493992
transform -1 0 424600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_io0_pad
timestamp 1606493992
transform -1 0 420600 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_290
timestamp 1606493992
transform -1 0 401200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_291
timestamp 1606493992
transform -1 0 403200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_292
timestamp 1606493992
transform -1 0 404200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_293
timestamp 1606493992
transform -1 0 404400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_294
timestamp 1606493992
transform -1 0 404600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_39
timestamp 1606493992
transform -1 0 385200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_40
timestamp 1606493992
transform -1 0 389200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_41
timestamp 1606493992
transform -1 0 393200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_42
timestamp 1606493992
transform -1 0 397200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_281
timestamp 1606493992
transform -1 0 372800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_282
timestamp 1606493992
transform -1 0 373000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_283
timestamp 1606493992
transform -1 0 373200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_37
timestamp 1606493992
transform -1 0 377200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_38
timestamp 1606493992
transform -1 0 381200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_279
timestamp 1606493992
transform -1 0 369800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_280
timestamp 1606493992
transform -1 0 371800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_clk_pad
timestamp 1606493992
transform -1 0 365800 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_36
timestamp 1606493992
transform -1 0 342400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_273
timestamp 1606493992
transform -1 0 346400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_274
timestamp 1606493992
transform -1 0 348400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_275
timestamp 1606493992
transform -1 0 349400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_276
timestamp 1606493992
transform -1 0 349600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_277
timestamp 1606493992
transform -1 0 349800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_35
timestamp 1606493992
transform -1 0 338400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_34
timestamp 1606493992
transform -1 0 334400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_33
timestamp 1606493992
transform -1 0 330400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_32
timestamp 1606493992
transform -1 0 326400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_264
timestamp 1606493992
transform -1 0 318000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_265
timestamp 1606493992
transform -1 0 318200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_266
timestamp 1606493992
transform -1 0 318400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_31
timestamp 1606493992
transform -1 0 322400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_263
timestamp 1606493992
transform -1 0 317000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_262
timestamp 1606493992
transform -1 0 315000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_csb_pad
timestamp 1606493992
transform -1 0 311000 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_256
timestamp 1606493992
transform -1 0 291600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_257
timestamp 1606493992
transform -1 0 293600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_258
timestamp 1606493992
transform -1 0 294600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_259
timestamp 1606493992
transform -1 0 294800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_260
timestamp 1606493992
transform -1 0 295000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_27
timestamp 1606493992
transform -1 0 275600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_28
timestamp 1606493992
transform -1 0 279600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_29
timestamp 1606493992
transform -1 0 283600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_30
timestamp 1606493992
transform -1 0 287600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_245
timestamp 1606493992
transform -1 0 260200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_246
timestamp 1606493992
transform -1 0 262200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_247
timestamp 1606493992
transform -1 0 263200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_248
timestamp 1606493992
transform -1 0 263400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_249
timestamp 1606493992
transform -1 0 263600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_25
timestamp 1606493992
transform -1 0 267600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_26
timestamp 1606493992
transform -1 0 271600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__vssd_lvc_pad  mgmt_vssd_lvclmap_pad
timestamp 1606493992
transform -1 0 256200 0 -1 39593
box 0 -46 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_243
timestamp 1606493992
transform -1 0 241200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_24
timestamp 1606493992
transform -1 0 233800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_239
timestamp 1606493992
transform -1 0 237800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_240
timestamp 1606493992
transform -1 0 239800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_241
timestamp 1606493992
transform -1 0 240800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_242
timestamp 1606493992
transform -1 0 241000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_20
timestamp 1606493992
transform -1 0 217800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_21
timestamp 1606493992
transform -1 0 221800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_22
timestamp 1606493992
transform -1 0 225800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_23
timestamp 1606493992
transform -1 0 229800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_228
timestamp 1606493992
transform -1 0 206400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_229
timestamp 1606493992
transform -1 0 208400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_230
timestamp 1606493992
transform -1 0 209400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_231
timestamp 1606493992
transform -1 0 209600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_232
timestamp 1606493992
transform -1 0 209800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_19
timestamp 1606493992
transform -1 0 213800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  clock_pad
timestamp 1606493992
transform -1 0 202400 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_1um  FILLER_225
timestamp 1606493992
transform -1 0 186200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_226
timestamp 1606493992
transform -1 0 186400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_17
timestamp 1606493992
transform -1 0 175000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_18
timestamp 1606493992
transform -1 0 179000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_222
timestamp 1606493992
transform -1 0 183000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_223
timestamp 1606493992
transform -1 0 185000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_224
timestamp 1606493992
transform -1 0 186000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_14
timestamp 1606493992
transform -1 0 163000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_15
timestamp 1606493992
transform -1 0 167000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_16
timestamp 1606493992
transform -1 0 171000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_211
timestamp 1606493992
transform -1 0 151600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_212
timestamp 1606493992
transform -1 0 153600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_213
timestamp 1606493992
transform -1 0 154600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_214
timestamp 1606493992
transform -1 0 154800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_215
timestamp 1606493992
transform -1 0 155000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_13
timestamp 1606493992
transform -1 0 159000 0 -1 39593
box 0 0 4000 39593
use sky130_fd_io__top_xres4v2  resetb_pad
timestamp 1606493992
transform -1 0 147600 0 -1 40000
box -103 0 15124 40000
use sky130_ef_io__com_bus_slice_10um  FILLER_206
timestamp 1606493992
transform -1 0 131200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_207
timestamp 1606493992
transform -1 0 132200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_208
timestamp 1606493992
transform -1 0 132400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_209
timestamp 1606493992
transform -1 0 132600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_205
timestamp 1606493992
transform -1 0 129200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_12
timestamp 1606493992
transform -1 0 125200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_11
timestamp 1606493992
transform -1 0 121200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_10
timestamp 1606493992
transform -1 0 117200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_9
timestamp 1606493992
transform -1 0 113200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_8
timestamp 1606493992
transform -1 0 109200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_197
timestamp 1606493992
transform -1 0 101000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_198
timestamp 1606493992
transform -1 0 101200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_7
timestamp 1606493992
transform -1 0 105200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_195
timestamp 1606493992
transform -1 0 99800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_196
timestamp 1606493992
transform -1 0 100800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_194
timestamp 1606493992
transform -1 0 97800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_pad  mgmt_vssa_hvclamp_pad
timestamp 1606493992
transform -1 0 93800 0 -1 39593
box 0 -434 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_189
timestamp 1606493992
transform -1 0 77400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_190
timestamp 1606493992
transform -1 0 78400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_191
timestamp 1606493992
transform -1 0 78600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_192
timestamp 1606493992
transform -1 0 78800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_4
timestamp 1606493992
transform -1 0 63400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_5
timestamp 1606493992
transform -1 0 67400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_6
timestamp 1606493992
transform -1 0 71400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_188
timestamp 1606493992
transform -1 0 75400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_178
timestamp 1606493992
transform -1 0 46000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_179
timestamp 1606493992
transform -1 0 47000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_180
timestamp 1606493992
transform -1 0 47200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_181
timestamp 1606493992
transform -1 0 47400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_1
timestamp 1606493992
transform -1 0 51400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_2
timestamp 1606493992
transform -1 0 55400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_3
timestamp 1606493992
transform -1 0 59400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__corner_pad  mgmt_corner\[0\]
timestamp 1606493992
transform -1 0 40000 0 -1 40800
box -271 -204 40000 40800
use sky130_ef_io__com_bus_slice_20um  FILLER_177
timestamp 1606493992
transform -1 0 44000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_381
timestamp 1606493992
transform 0 -1 39593 1 0 40800
box 0 0 4000 39593
<< labels >>
rlabel metal5 s 187640 6598 200160 19088 4 clock
port 1 nsew
rlabel metal2 s 187327 41713 187383 42193 4 clock_core
port 2 nsew
rlabel metal2 s 194043 41713 194099 42193 4 por
port 3 nsew
rlabel metal5 s 351040 6598 363560 19088 4 flash_clk
port 4 nsew
rlabel metal2 s 361767 41713 361823 42193 4 flash_clk_core
port 5 nsew
rlabel metal2 s 357443 41713 357499 42193 4 flash_clk_ieb_core
port 6 nsew
rlabel metal2 s 364895 41713 364951 42193 4 flash_clk_oeb_core
port 7 nsew
rlabel metal5 s 296240 6598 308760 19088 4 flash_csb
port 8 nsew
rlabel metal2 s 306967 41713 307023 42193 4 flash_csb_core
port 9 nsew
rlabel metal2 s 302643 41713 302699 42193 4 flash_csb_ieb_core
port 10 nsew
rlabel metal2 s 310095 41713 310151 42193 4 flash_csb_oeb_core
port 11 nsew
rlabel metal5 s 405840 6598 418360 19088 4 flash_io0
port 12 nsew
rlabel metal2 s 405527 41713 405583 42193 4 flash_io0_di_core
port 13 nsew
rlabel metal2 s 416567 41713 416623 42193 4 flash_io0_do_core
port 14 nsew
rlabel metal2 s 412243 41713 412299 42193 4 flash_io0_ieb_core
port 15 nsew
rlabel metal2 s 419695 41713 419751 42193 4 flash_io0_oeb_core
port 16 nsew
rlabel metal5 s 460640 6598 473160 19088 4 flash_io1
port 17 nsew
rlabel metal2 s 460327 41713 460383 42193 4 flash_io1_di_core
port 18 nsew
rlabel metal2 s 471367 41713 471423 42193 4 flash_io1_do_core
port 19 nsew
rlabel metal2 s 467043 41713 467099 42193 4 flash_io1_ieb_core
port 20 nsew
rlabel metal2 s 474495 41713 474551 42193 4 flash_io1_oeb_core
port 21 nsew
rlabel metal5 s 515440 6598 527960 19088 4 gpio
port 22 nsew
rlabel metal2 s 515127 41713 515183 42193 4 gpio_in_core
port 23 nsew
rlabel metal2 s 521843 41713 521899 42193 4 gpio_inenb_core
port 24 nsew
rlabel metal2 s 520647 41713 520703 42193 4 gpio_mode0_core
port 25 nsew
rlabel metal2 s 524971 41713 525027 42193 4 gpio_mode1_core
port 26 nsew
rlabel metal2 s 526167 41713 526223 42193 4 gpio_out_core
port 27 nsew
rlabel metal2 s 529295 41713 529351 42193 4 gpio_outenb_core
port 28 nsew
rlabel metal5 s 6086 69863 19572 81191 4 vccd
port 29 nsew
rlabel metal5 s 624040 6675 636580 19197 4 vdda
port 30 nsew
rlabel metal5 s 6675 111420 19197 123960 4 vddio
port 31 nsew
rlabel metal5 s 80040 6675 92580 19197 4 vssa
port 32 nsew
rlabel metal5 s 243009 6086 254337 19572 4 vssd
port 33 nsew
rlabel metal5 s 334620 1018402 347160 1030924 4 vssio
port 34 nsew
rlabel metal5 s 698512 101240 711002 113760 4 mprj_io[0]
port 35 nsew
rlabel metal2 s 675407 105803 675887 105859 4 mprj_io_analog_en[0]
port 36 nsew
rlabel metal2 s 675407 107091 675887 107147 4 mprj_io_analog_pol[0]
port 37 nsew
rlabel metal2 s 675407 110127 675887 110183 4 mprj_io_analog_sel[0]
port 38 nsew
rlabel metal2 s 675407 106447 675887 106503 4 mprj_io_dm[0]
port 39 nsew
rlabel metal2 s 675407 104607 675887 104663 4 mprj_io_dm[1]
port 40 nsew
rlabel metal2 s 675407 110771 675887 110827 4 mprj_io_dm[2]
port 41 nsew
rlabel metal2 s 675407 108931 675887 108987 4 mprj_io_enh[0]
port 42 nsew
rlabel metal2 s 675407 109575 675887 109631 4 mprj_io_hldh_n[0]
port 43 nsew
rlabel metal2 s 675407 111415 675887 111471 4 mprj_io_holdover[0]
port 44 nsew
rlabel metal2 s 675407 114451 675887 114507 4 mprj_io_ib_mode_sel[0]
port 45 nsew
rlabel metal2 s 675407 107643 675887 107699 4 mprj_io_inp_dis[0]
port 46 nsew
rlabel metal2 s 675407 115095 675887 115151 4 mprj_io_oeb[0]
port 47 nsew
rlabel metal2 s 675407 111967 675887 112023 4 mprj_io_out[0]
port 48 nsew
rlabel metal2 s 675407 102767 675887 102823 4 mprj_io_slow_sel[0]
port 49 nsew
rlabel metal2 s 675407 113807 675887 113863 4 mprj_io_vtrip_sel[0]
port 50 nsew
rlabel metal2 s 675407 100927 675887 100983 4 mprj_io_in[0]
port 51 nsew
rlabel metal2 s 675407 686611 675887 686667 4 mprj_analog_io[3]
port 52 nsew
rlabel metal5 s 698512 684440 711002 696960 4 mprj_io[10]
port 53 nsew
rlabel metal2 s 675407 689003 675887 689059 4 mprj_io_analog_en[10]
port 54 nsew
rlabel metal2 s 675407 690291 675887 690347 4 mprj_io_analog_pol[10]
port 55 nsew
rlabel metal2 s 675407 693327 675887 693383 4 mprj_io_analog_sel[10]
port 56 nsew
rlabel metal2 s 675407 689647 675887 689703 4 mprj_io_dm[30]
port 57 nsew
rlabel metal2 s 675407 687807 675887 687863 4 mprj_io_dm[31]
port 58 nsew
rlabel metal2 s 675407 693971 675887 694027 4 mprj_io_dm[32]
port 59 nsew
rlabel metal2 s 675407 692131 675887 692187 4 mprj_io_enh[10]
port 60 nsew
rlabel metal2 s 675407 692775 675887 692831 4 mprj_io_hldh_n[10]
port 61 nsew
rlabel metal2 s 675407 694615 675887 694671 4 mprj_io_holdover[10]
port 62 nsew
rlabel metal2 s 675407 697651 675887 697707 4 mprj_io_ib_mode_sel[10]
port 63 nsew
rlabel metal2 s 675407 690843 675887 690899 4 mprj_io_inp_dis[10]
port 64 nsew
rlabel metal2 s 675407 698295 675887 698351 4 mprj_io_oeb[10]
port 65 nsew
rlabel metal2 s 675407 695167 675887 695223 4 mprj_io_out[10]
port 66 nsew
rlabel metal2 s 675407 685967 675887 686023 4 mprj_io_slow_sel[10]
port 67 nsew
rlabel metal2 s 675407 697007 675887 697063 4 mprj_io_vtrip_sel[10]
port 68 nsew
rlabel metal2 s 675407 684127 675887 684183 4 mprj_io_in[10]
port 69 nsew
rlabel metal2 s 675407 731611 675887 731667 4 mprj_analog_io[4]
port 70 nsew
rlabel metal5 s 698512 729440 711002 741960 4 mprj_io[11]
port 71 nsew
rlabel metal2 s 675407 734003 675887 734059 4 mprj_io_analog_en[11]
port 72 nsew
rlabel metal2 s 675407 735291 675887 735347 4 mprj_io_analog_pol[11]
port 73 nsew
rlabel metal2 s 675407 738327 675887 738383 4 mprj_io_analog_sel[11]
port 74 nsew
rlabel metal2 s 675407 734647 675887 734703 4 mprj_io_dm[33]
port 75 nsew
rlabel metal2 s 675407 732807 675887 732863 4 mprj_io_dm[34]
port 76 nsew
rlabel metal2 s 675407 738971 675887 739027 4 mprj_io_dm[35]
port 77 nsew
rlabel metal2 s 675407 737131 675887 737187 4 mprj_io_enh[11]
port 78 nsew
rlabel metal2 s 675407 737775 675887 737831 4 mprj_io_hldh_n[11]
port 79 nsew
rlabel metal2 s 675407 739615 675887 739671 4 mprj_io_holdover[11]
port 80 nsew
rlabel metal2 s 675407 742651 675887 742707 4 mprj_io_ib_mode_sel[11]
port 81 nsew
rlabel metal2 s 675407 735843 675887 735899 4 mprj_io_inp_dis[11]
port 82 nsew
rlabel metal2 s 675407 743295 675887 743351 4 mprj_io_oeb[11]
port 83 nsew
rlabel metal2 s 675407 740167 675887 740223 4 mprj_io_out[11]
port 84 nsew
rlabel metal2 s 675407 730967 675887 731023 4 mprj_io_slow_sel[11]
port 85 nsew
rlabel metal2 s 675407 742007 675887 742063 4 mprj_io_vtrip_sel[11]
port 86 nsew
rlabel metal2 s 675407 729127 675887 729183 4 mprj_io_in[11]
port 87 nsew
rlabel metal2 s 675407 776611 675887 776667 4 mprj_analog_io[5]
port 88 nsew
rlabel metal5 s 698512 774440 711002 786960 4 mprj_io[12]
port 89 nsew
rlabel metal2 s 675407 779003 675887 779059 4 mprj_io_analog_en[12]
port 90 nsew
rlabel metal2 s 675407 780291 675887 780347 4 mprj_io_analog_pol[12]
port 91 nsew
rlabel metal2 s 675407 783327 675887 783383 4 mprj_io_analog_sel[12]
port 92 nsew
rlabel metal2 s 675407 779647 675887 779703 4 mprj_io_dm[36]
port 93 nsew
rlabel metal2 s 675407 777807 675887 777863 4 mprj_io_dm[37]
port 94 nsew
rlabel metal2 s 675407 783971 675887 784027 4 mprj_io_dm[38]
port 95 nsew
rlabel metal2 s 675407 782131 675887 782187 4 mprj_io_enh[12]
port 96 nsew
rlabel metal2 s 675407 782775 675887 782831 4 mprj_io_hldh_n[12]
port 97 nsew
rlabel metal2 s 675407 784615 675887 784671 4 mprj_io_holdover[12]
port 98 nsew
rlabel metal2 s 675407 787651 675887 787707 4 mprj_io_ib_mode_sel[12]
port 99 nsew
rlabel metal2 s 675407 780843 675887 780899 4 mprj_io_inp_dis[12]
port 100 nsew
rlabel metal2 s 675407 788295 675887 788351 4 mprj_io_oeb[12]
port 101 nsew
rlabel metal2 s 675407 785167 675887 785223 4 mprj_io_out[12]
port 102 nsew
rlabel metal2 s 675407 775967 675887 776023 4 mprj_io_slow_sel[12]
port 103 nsew
rlabel metal2 s 675407 787007 675887 787063 4 mprj_io_vtrip_sel[12]
port 104 nsew
rlabel metal2 s 675407 774127 675887 774183 4 mprj_io_in[12]
port 105 nsew
rlabel metal2 s 675407 865811 675887 865867 4 mprj_analog_io[6]
port 106 nsew
rlabel metal5 s 698512 863640 711002 876160 4 mprj_io[13]
port 107 nsew
rlabel metal2 s 675407 868203 675887 868259 4 mprj_io_analog_en[13]
port 108 nsew
rlabel metal2 s 675407 869491 675887 869547 4 mprj_io_analog_pol[13]
port 109 nsew
rlabel metal2 s 675407 872527 675887 872583 4 mprj_io_analog_sel[13]
port 110 nsew
rlabel metal2 s 675407 868847 675887 868903 4 mprj_io_dm[39]
port 111 nsew
rlabel metal2 s 675407 867007 675887 867063 4 mprj_io_dm[40]
port 112 nsew
rlabel metal2 s 675407 873171 675887 873227 4 mprj_io_dm[41]
port 113 nsew
rlabel metal2 s 675407 871331 675887 871387 4 mprj_io_enh[13]
port 114 nsew
rlabel metal2 s 675407 871975 675887 872031 4 mprj_io_hldh_n[13]
port 115 nsew
rlabel metal2 s 675407 873815 675887 873871 4 mprj_io_holdover[13]
port 116 nsew
rlabel metal2 s 675407 876851 675887 876907 4 mprj_io_ib_mode_sel[13]
port 117 nsew
rlabel metal2 s 675407 870043 675887 870099 4 mprj_io_inp_dis[13]
port 118 nsew
rlabel metal2 s 675407 877495 675887 877551 4 mprj_io_oeb[13]
port 119 nsew
rlabel metal2 s 675407 874367 675887 874423 4 mprj_io_out[13]
port 120 nsew
rlabel metal2 s 675407 865167 675887 865223 4 mprj_io_slow_sel[13]
port 121 nsew
rlabel metal2 s 675407 876207 675887 876263 4 mprj_io_vtrip_sel[13]
port 122 nsew
rlabel metal2 s 675407 863327 675887 863383 4 mprj_io_in[13]
port 123 nsew
rlabel metal2 s 675407 955011 675887 955067 4 mprj_analog_io[7]
port 124 nsew
rlabel metal5 s 698512 952840 711002 965360 4 mprj_io[14]
port 125 nsew
rlabel metal2 s 675407 957403 675887 957459 4 mprj_io_analog_en[14]
port 126 nsew
rlabel metal2 s 675407 958691 675887 958747 4 mprj_io_analog_pol[14]
port 127 nsew
rlabel metal2 s 675407 961727 675887 961783 4 mprj_io_analog_sel[14]
port 128 nsew
rlabel metal2 s 675407 958047 675887 958103 4 mprj_io_dm[42]
port 129 nsew
rlabel metal2 s 675407 956207 675887 956263 4 mprj_io_dm[43]
port 130 nsew
rlabel metal2 s 675407 962371 675887 962427 4 mprj_io_dm[44]
port 131 nsew
rlabel metal2 s 675407 960531 675887 960587 4 mprj_io_enh[14]
port 132 nsew
rlabel metal2 s 675407 961175 675887 961231 4 mprj_io_hldh_n[14]
port 133 nsew
rlabel metal2 s 675407 963015 675887 963071 4 mprj_io_holdover[14]
port 134 nsew
rlabel metal2 s 675407 966051 675887 966107 4 mprj_io_ib_mode_sel[14]
port 135 nsew
rlabel metal2 s 675407 959243 675887 959299 4 mprj_io_inp_dis[14]
port 136 nsew
rlabel metal2 s 675407 966695 675887 966751 4 mprj_io_oeb[14]
port 137 nsew
rlabel metal2 s 675407 963567 675887 963623 4 mprj_io_out[14]
port 138 nsew
rlabel metal2 s 675407 954367 675887 954423 4 mprj_io_slow_sel[14]
port 139 nsew
rlabel metal2 s 675407 965407 675887 965463 4 mprj_io_vtrip_sel[14]
port 140 nsew
rlabel metal2 s 675407 952527 675887 952583 4 mprj_io_in[14]
port 141 nsew
rlabel metal2 s 638533 995407 638589 995887 4 mprj_analog_io[8]
port 142 nsew
rlabel metal5 s 628240 1018512 640760 1031002 4 mprj_io[15]
port 143 nsew
rlabel metal2 s 636141 995407 636197 995887 4 mprj_io_analog_en[15]
port 144 nsew
rlabel metal2 s 634853 995407 634909 995887 4 mprj_io_analog_pol[15]
port 145 nsew
rlabel metal2 s 631817 995407 631873 995887 4 mprj_io_analog_sel[15]
port 146 nsew
rlabel metal2 s 635497 995407 635553 995887 4 mprj_io_dm[45]
port 147 nsew
rlabel metal2 s 637337 995407 637393 995887 4 mprj_io_dm[46]
port 148 nsew
rlabel metal2 s 631173 995407 631229 995887 4 mprj_io_dm[47]
port 149 nsew
rlabel metal2 s 633013 995407 633069 995887 4 mprj_io_enh[15]
port 150 nsew
rlabel metal2 s 632369 995407 632425 995887 4 mprj_io_hldh_n[15]
port 151 nsew
rlabel metal2 s 630529 995407 630585 995887 4 mprj_io_holdover[15]
port 152 nsew
rlabel metal2 s 627493 995407 627549 995887 4 mprj_io_ib_mode_sel[15]
port 153 nsew
rlabel metal2 s 634301 995407 634357 995887 4 mprj_io_inp_dis[15]
port 154 nsew
rlabel metal2 s 626849 995407 626905 995887 4 mprj_io_oeb[15]
port 155 nsew
rlabel metal2 s 629977 995407 630033 995887 4 mprj_io_out[15]
port 156 nsew
rlabel metal2 s 639177 995407 639233 995887 4 mprj_io_slow_sel[15]
port 157 nsew
rlabel metal2 s 628137 995407 628193 995887 4 mprj_io_vtrip_sel[15]
port 158 nsew
rlabel metal2 s 641017 995407 641073 995887 4 mprj_io_in[15]
port 159 nsew
rlabel metal2 s 536733 995407 536789 995887 4 mprj_analog_io[9]
port 160 nsew
rlabel metal5 s 526440 1018512 538960 1031002 4 mprj_io[16]
port 161 nsew
rlabel metal2 s 534341 995407 534397 995887 4 mprj_io_analog_en[16]
port 162 nsew
rlabel metal2 s 533053 995407 533109 995887 4 mprj_io_analog_pol[16]
port 163 nsew
rlabel metal2 s 530017 995407 530073 995887 4 mprj_io_analog_sel[16]
port 164 nsew
rlabel metal2 s 533697 995407 533753 995887 4 mprj_io_dm[48]
port 165 nsew
rlabel metal2 s 535537 995407 535593 995887 4 mprj_io_dm[49]
port 166 nsew
rlabel metal2 s 529373 995407 529429 995887 4 mprj_io_dm[50]
port 167 nsew
rlabel metal2 s 531213 995407 531269 995887 4 mprj_io_enh[16]
port 168 nsew
rlabel metal2 s 530569 995407 530625 995887 4 mprj_io_hldh_n[16]
port 169 nsew
rlabel metal2 s 528729 995407 528785 995887 4 mprj_io_holdover[16]
port 170 nsew
rlabel metal2 s 525693 995407 525749 995887 4 mprj_io_ib_mode_sel[16]
port 171 nsew
rlabel metal2 s 532501 995407 532557 995887 4 mprj_io_inp_dis[16]
port 172 nsew
rlabel metal2 s 525049 995407 525105 995887 4 mprj_io_oeb[16]
port 173 nsew
rlabel metal2 s 528177 995407 528233 995887 4 mprj_io_out[16]
port 174 nsew
rlabel metal2 s 537377 995407 537433 995887 4 mprj_io_slow_sel[16]
port 175 nsew
rlabel metal2 s 526337 995407 526393 995887 4 mprj_io_vtrip_sel[16]
port 176 nsew
rlabel metal2 s 539217 995407 539273 995887 4 mprj_io_in[16]
port 177 nsew
rlabel metal2 s 485333 995407 485389 995887 4 mprj_analog_io[10]
port 178 nsew
rlabel metal5 s 475040 1018512 487560 1031002 4 mprj_io[17]
port 179 nsew
rlabel metal2 s 482941 995407 482997 995887 4 mprj_io_analog_en[17]
port 180 nsew
rlabel metal2 s 481653 995407 481709 995887 4 mprj_io_analog_pol[17]
port 181 nsew
rlabel metal2 s 478617 995407 478673 995887 4 mprj_io_analog_sel[17]
port 182 nsew
rlabel metal2 s 482297 995407 482353 995887 4 mprj_io_dm[51]
port 183 nsew
rlabel metal2 s 484137 995407 484193 995887 4 mprj_io_dm[52]
port 184 nsew
rlabel metal2 s 477973 995407 478029 995887 4 mprj_io_dm[53]
port 185 nsew
rlabel metal2 s 479813 995407 479869 995887 4 mprj_io_enh[17]
port 186 nsew
rlabel metal2 s 479169 995407 479225 995887 4 mprj_io_hldh_n[17]
port 187 nsew
rlabel metal2 s 477329 995407 477385 995887 4 mprj_io_holdover[17]
port 188 nsew
rlabel metal2 s 474293 995407 474349 995887 4 mprj_io_ib_mode_sel[17]
port 189 nsew
rlabel metal2 s 481101 995407 481157 995887 4 mprj_io_inp_dis[17]
port 190 nsew
rlabel metal2 s 473649 995407 473705 995887 4 mprj_io_oeb[17]
port 191 nsew
rlabel metal2 s 476777 995407 476833 995887 4 mprj_io_out[17]
port 192 nsew
rlabel metal2 s 485977 995407 486033 995887 4 mprj_io_slow_sel[17]
port 193 nsew
rlabel metal2 s 474937 995407 474993 995887 4 mprj_io_vtrip_sel[17]
port 194 nsew
rlabel metal2 s 487817 995407 487873 995887 4 mprj_io_in[17]
port 195 nsew
rlabel metal5 s 698512 146440 711002 158960 4 mprj_io[1]
port 196 nsew
rlabel metal2 s 675407 151003 675887 151059 4 mprj_io_analog_en[1]
port 197 nsew
rlabel metal2 s 675407 152291 675887 152347 4 mprj_io_analog_pol[1]
port 198 nsew
rlabel metal2 s 675407 155327 675887 155383 4 mprj_io_analog_sel[1]
port 199 nsew
rlabel metal2 s 675407 151647 675887 151703 4 mprj_io_dm[3]
port 200 nsew
rlabel metal2 s 675407 149807 675887 149863 4 mprj_io_dm[4]
port 201 nsew
rlabel metal2 s 675407 155971 675887 156027 4 mprj_io_dm[5]
port 202 nsew
rlabel metal2 s 675407 154131 675887 154187 4 mprj_io_enh[1]
port 203 nsew
rlabel metal2 s 675407 154775 675887 154831 4 mprj_io_hldh_n[1]
port 204 nsew
rlabel metal2 s 675407 156615 675887 156671 4 mprj_io_holdover[1]
port 205 nsew
rlabel metal2 s 675407 159651 675887 159707 4 mprj_io_ib_mode_sel[1]
port 206 nsew
rlabel metal2 s 675407 152843 675887 152899 4 mprj_io_inp_dis[1]
port 207 nsew
rlabel metal2 s 675407 160295 675887 160351 4 mprj_io_oeb[1]
port 208 nsew
rlabel metal2 s 675407 157167 675887 157223 4 mprj_io_out[1]
port 209 nsew
rlabel metal2 s 675407 147967 675887 148023 4 mprj_io_slow_sel[1]
port 210 nsew
rlabel metal2 s 675407 159007 675887 159063 4 mprj_io_vtrip_sel[1]
port 211 nsew
rlabel metal2 s 675407 146127 675887 146183 4 mprj_io_in[1]
port 212 nsew
rlabel metal5 s 698512 191440 711002 203960 4 mprj_io[2]
port 213 nsew
rlabel metal2 s 675407 196003 675887 196059 4 mprj_io_analog_en[2]
port 214 nsew
rlabel metal2 s 675407 197291 675887 197347 4 mprj_io_analog_pol[2]
port 215 nsew
rlabel metal2 s 675407 200327 675887 200383 4 mprj_io_analog_sel[2]
port 216 nsew
rlabel metal2 s 675407 196647 675887 196703 4 mprj_io_dm[6]
port 217 nsew
rlabel metal2 s 675407 194807 675887 194863 4 mprj_io_dm[7]
port 218 nsew
rlabel metal2 s 675407 200971 675887 201027 4 mprj_io_dm[8]
port 219 nsew
rlabel metal2 s 675407 199131 675887 199187 4 mprj_io_enh[2]
port 220 nsew
rlabel metal2 s 675407 199775 675887 199831 4 mprj_io_hldh_n[2]
port 221 nsew
rlabel metal2 s 675407 201615 675887 201671 4 mprj_io_holdover[2]
port 222 nsew
rlabel metal2 s 675407 204651 675887 204707 4 mprj_io_ib_mode_sel[2]
port 223 nsew
rlabel metal2 s 675407 197843 675887 197899 4 mprj_io_inp_dis[2]
port 224 nsew
rlabel metal2 s 675407 205295 675887 205351 4 mprj_io_oeb[2]
port 225 nsew
rlabel metal2 s 675407 202167 675887 202223 4 mprj_io_out[2]
port 226 nsew
rlabel metal2 s 675407 192967 675887 193023 4 mprj_io_slow_sel[2]
port 227 nsew
rlabel metal2 s 675407 204007 675887 204063 4 mprj_io_vtrip_sel[2]
port 228 nsew
rlabel metal2 s 675407 191127 675887 191183 4 mprj_io_in[2]
port 229 nsew
rlabel metal5 s 698512 236640 711002 249160 4 mprj_io[3]
port 230 nsew
rlabel metal2 s 675407 241203 675887 241259 4 mprj_io_analog_en[3]
port 231 nsew
rlabel metal2 s 675407 242491 675887 242547 4 mprj_io_analog_pol[3]
port 232 nsew
rlabel metal2 s 675407 245527 675887 245583 4 mprj_io_analog_sel[3]
port 233 nsew
rlabel metal2 s 675407 240007 675887 240063 4 mprj_io_dm[10]
port 234 nsew
rlabel metal2 s 675407 246171 675887 246227 4 mprj_io_dm[11]
port 235 nsew
rlabel metal2 s 675407 241847 675887 241903 4 mprj_io_dm[9]
port 236 nsew
rlabel metal2 s 675407 244331 675887 244387 4 mprj_io_enh[3]
port 237 nsew
rlabel metal2 s 675407 244975 675887 245031 4 mprj_io_hldh_n[3]
port 238 nsew
rlabel metal2 s 675407 246815 675887 246871 4 mprj_io_holdover[3]
port 239 nsew
rlabel metal2 s 675407 249851 675887 249907 4 mprj_io_ib_mode_sel[3]
port 240 nsew
rlabel metal2 s 675407 243043 675887 243099 4 mprj_io_inp_dis[3]
port 241 nsew
rlabel metal2 s 675407 250495 675887 250551 4 mprj_io_oeb[3]
port 242 nsew
rlabel metal2 s 675407 247367 675887 247423 4 mprj_io_out[3]
port 243 nsew
rlabel metal2 s 675407 238167 675887 238223 4 mprj_io_slow_sel[3]
port 244 nsew
rlabel metal2 s 675407 249207 675887 249263 4 mprj_io_vtrip_sel[3]
port 245 nsew
rlabel metal2 s 675407 236327 675887 236383 4 mprj_io_in[3]
port 246 nsew
rlabel metal5 s 698512 281640 711002 294160 4 mprj_io[4]
port 247 nsew
rlabel metal2 s 675407 286203 675887 286259 4 mprj_io_analog_en[4]
port 248 nsew
rlabel metal2 s 675407 287491 675887 287547 4 mprj_io_analog_pol[4]
port 249 nsew
rlabel metal2 s 675407 290527 675887 290583 4 mprj_io_analog_sel[4]
port 250 nsew
rlabel metal2 s 675407 286847 675887 286903 4 mprj_io_dm[12]
port 251 nsew
rlabel metal2 s 675407 285007 675887 285063 4 mprj_io_dm[13]
port 252 nsew
rlabel metal2 s 675407 291171 675887 291227 4 mprj_io_dm[14]
port 253 nsew
rlabel metal2 s 675407 289331 675887 289387 4 mprj_io_enh[4]
port 254 nsew
rlabel metal2 s 675407 289975 675887 290031 4 mprj_io_hldh_n[4]
port 255 nsew
rlabel metal2 s 675407 291815 675887 291871 4 mprj_io_holdover[4]
port 256 nsew
rlabel metal2 s 675407 294851 675887 294907 4 mprj_io_ib_mode_sel[4]
port 257 nsew
rlabel metal2 s 675407 288043 675887 288099 4 mprj_io_inp_dis[4]
port 258 nsew
rlabel metal2 s 675407 295495 675887 295551 4 mprj_io_oeb[4]
port 259 nsew
rlabel metal2 s 675407 292367 675887 292423 4 mprj_io_out[4]
port 260 nsew
rlabel metal2 s 675407 283167 675887 283223 4 mprj_io_slow_sel[4]
port 261 nsew
rlabel metal2 s 675407 294207 675887 294263 4 mprj_io_vtrip_sel[4]
port 262 nsew
rlabel metal2 s 675407 281327 675887 281383 4 mprj_io_in[4]
port 263 nsew
rlabel metal5 s 698512 326640 711002 339160 4 mprj_io[5]
port 264 nsew
rlabel metal2 s 675407 331203 675887 331259 4 mprj_io_analog_en[5]
port 265 nsew
rlabel metal2 s 675407 332491 675887 332547 4 mprj_io_analog_pol[5]
port 266 nsew
rlabel metal2 s 675407 335527 675887 335583 4 mprj_io_analog_sel[5]
port 267 nsew
rlabel metal2 s 675407 331847 675887 331903 4 mprj_io_dm[15]
port 268 nsew
rlabel metal2 s 675407 330007 675887 330063 4 mprj_io_dm[16]
port 269 nsew
rlabel metal2 s 675407 336171 675887 336227 4 mprj_io_dm[17]
port 270 nsew
rlabel metal2 s 675407 334331 675887 334387 4 mprj_io_enh[5]
port 271 nsew
rlabel metal2 s 675407 334975 675887 335031 4 mprj_io_hldh_n[5]
port 272 nsew
rlabel metal2 s 675407 336815 675887 336871 4 mprj_io_holdover[5]
port 273 nsew
rlabel metal2 s 675407 339851 675887 339907 4 mprj_io_ib_mode_sel[5]
port 274 nsew
rlabel metal2 s 675407 333043 675887 333099 4 mprj_io_inp_dis[5]
port 275 nsew
rlabel metal2 s 675407 340495 675887 340551 4 mprj_io_oeb[5]
port 276 nsew
rlabel metal2 s 675407 337367 675887 337423 4 mprj_io_out[5]
port 277 nsew
rlabel metal2 s 675407 328167 675887 328223 4 mprj_io_slow_sel[5]
port 278 nsew
rlabel metal2 s 675407 339207 675887 339263 4 mprj_io_vtrip_sel[5]
port 279 nsew
rlabel metal2 s 675407 326327 675887 326383 4 mprj_io_in[5]
port 280 nsew
rlabel metal5 s 698512 371840 711002 384360 4 mprj_io[6]
port 281 nsew
rlabel metal2 s 675407 376403 675887 376459 4 mprj_io_analog_en[6]
port 282 nsew
rlabel metal2 s 675407 377691 675887 377747 4 mprj_io_analog_pol[6]
port 283 nsew
rlabel metal2 s 675407 380727 675887 380783 4 mprj_io_analog_sel[6]
port 284 nsew
rlabel metal2 s 675407 377047 675887 377103 4 mprj_io_dm[18]
port 285 nsew
rlabel metal2 s 675407 375207 675887 375263 4 mprj_io_dm[19]
port 286 nsew
rlabel metal2 s 675407 381371 675887 381427 4 mprj_io_dm[20]
port 287 nsew
rlabel metal2 s 675407 379531 675887 379587 4 mprj_io_enh[6]
port 288 nsew
rlabel metal2 s 675407 380175 675887 380231 4 mprj_io_hldh_n[6]
port 289 nsew
rlabel metal2 s 675407 382015 675887 382071 4 mprj_io_holdover[6]
port 290 nsew
rlabel metal2 s 675407 385051 675887 385107 4 mprj_io_ib_mode_sel[6]
port 291 nsew
rlabel metal2 s 675407 378243 675887 378299 4 mprj_io_inp_dis[6]
port 292 nsew
rlabel metal2 s 675407 385695 675887 385751 4 mprj_io_oeb[6]
port 293 nsew
rlabel metal2 s 675407 382567 675887 382623 4 mprj_io_out[6]
port 294 nsew
rlabel metal2 s 675407 373367 675887 373423 4 mprj_io_slow_sel[6]
port 295 nsew
rlabel metal2 s 675407 384407 675887 384463 4 mprj_io_vtrip_sel[6]
port 296 nsew
rlabel metal2 s 675407 371527 675887 371583 4 mprj_io_in[6]
port 297 nsew
rlabel metal2 s 675407 551211 675887 551267 4 mprj_analog_io[0]
port 298 nsew
rlabel metal5 s 698512 549040 711002 561560 4 mprj_io[7]
port 299 nsew
rlabel metal2 s 675407 553603 675887 553659 4 mprj_io_analog_en[7]
port 300 nsew
rlabel metal2 s 675407 554891 675887 554947 4 mprj_io_analog_pol[7]
port 301 nsew
rlabel metal2 s 675407 557927 675887 557983 4 mprj_io_analog_sel[7]
port 302 nsew
rlabel metal2 s 675407 554247 675887 554303 4 mprj_io_dm[21]
port 303 nsew
rlabel metal2 s 675407 552407 675887 552463 4 mprj_io_dm[22]
port 304 nsew
rlabel metal2 s 675407 558571 675887 558627 4 mprj_io_dm[23]
port 305 nsew
rlabel metal2 s 675407 556731 675887 556787 4 mprj_io_enh[7]
port 306 nsew
rlabel metal2 s 675407 557375 675887 557431 4 mprj_io_hldh_n[7]
port 307 nsew
rlabel metal2 s 675407 559215 675887 559271 4 mprj_io_holdover[7]
port 308 nsew
rlabel metal2 s 675407 562251 675887 562307 4 mprj_io_ib_mode_sel[7]
port 309 nsew
rlabel metal2 s 675407 555443 675887 555499 4 mprj_io_inp_dis[7]
port 310 nsew
rlabel metal2 s 675407 562895 675887 562951 4 mprj_io_oeb[7]
port 311 nsew
rlabel metal2 s 675407 559767 675887 559823 4 mprj_io_out[7]
port 312 nsew
rlabel metal2 s 675407 550567 675887 550623 4 mprj_io_slow_sel[7]
port 313 nsew
rlabel metal2 s 675407 561607 675887 561663 4 mprj_io_vtrip_sel[7]
port 314 nsew
rlabel metal2 s 675407 548727 675887 548783 4 mprj_io_in[7]
port 315 nsew
rlabel metal2 s 675407 596411 675887 596467 4 mprj_analog_io[1]
port 316 nsew
rlabel metal5 s 698512 594240 711002 606760 4 mprj_io[8]
port 317 nsew
rlabel metal2 s 675407 598803 675887 598859 4 mprj_io_analog_en[8]
port 318 nsew
rlabel metal2 s 675407 600091 675887 600147 4 mprj_io_analog_pol[8]
port 319 nsew
rlabel metal2 s 675407 603127 675887 603183 4 mprj_io_analog_sel[8]
port 320 nsew
rlabel metal2 s 675407 599447 675887 599503 4 mprj_io_dm[24]
port 321 nsew
rlabel metal2 s 675407 597607 675887 597663 4 mprj_io_dm[25]
port 322 nsew
rlabel metal2 s 675407 603771 675887 603827 4 mprj_io_dm[26]
port 323 nsew
rlabel metal2 s 675407 601931 675887 601987 4 mprj_io_enh[8]
port 324 nsew
rlabel metal2 s 675407 602575 675887 602631 4 mprj_io_hldh_n[8]
port 325 nsew
rlabel metal2 s 675407 604415 675887 604471 4 mprj_io_holdover[8]
port 326 nsew
rlabel metal2 s 675407 607451 675887 607507 4 mprj_io_ib_mode_sel[8]
port 327 nsew
rlabel metal2 s 675407 600643 675887 600699 4 mprj_io_inp_dis[8]
port 328 nsew
rlabel metal2 s 675407 608095 675887 608151 4 mprj_io_oeb[8]
port 329 nsew
rlabel metal2 s 675407 604967 675887 605023 4 mprj_io_out[8]
port 330 nsew
rlabel metal2 s 675407 595767 675887 595823 4 mprj_io_slow_sel[8]
port 331 nsew
rlabel metal2 s 675407 606807 675887 606863 4 mprj_io_vtrip_sel[8]
port 332 nsew
rlabel metal2 s 675407 593927 675887 593983 4 mprj_io_in[8]
port 333 nsew
rlabel metal2 s 675407 641411 675887 641467 4 mprj_analog_io[2]
port 334 nsew
rlabel metal5 s 698512 639240 711002 651760 4 mprj_io[9]
port 335 nsew
rlabel metal2 s 675407 643803 675887 643859 4 mprj_io_analog_en[9]
port 336 nsew
rlabel metal2 s 675407 645091 675887 645147 4 mprj_io_analog_pol[9]
port 337 nsew
rlabel metal2 s 675407 648127 675887 648183 4 mprj_io_analog_sel[9]
port 338 nsew
rlabel metal2 s 675407 644447 675887 644503 4 mprj_io_dm[27]
port 339 nsew
rlabel metal2 s 675407 642607 675887 642663 4 mprj_io_dm[28]
port 340 nsew
rlabel metal2 s 675407 648771 675887 648827 4 mprj_io_dm[29]
port 341 nsew
rlabel metal2 s 675407 646931 675887 646987 4 mprj_io_enh[9]
port 342 nsew
rlabel metal2 s 675407 647575 675887 647631 4 mprj_io_hldh_n[9]
port 343 nsew
rlabel metal2 s 675407 649415 675887 649471 4 mprj_io_holdover[9]
port 344 nsew
rlabel metal2 s 675407 652451 675887 652507 4 mprj_io_ib_mode_sel[9]
port 345 nsew
rlabel metal2 s 675407 645643 675887 645699 4 mprj_io_inp_dis[9]
port 346 nsew
rlabel metal2 s 675407 653095 675887 653151 4 mprj_io_oeb[9]
port 347 nsew
rlabel metal2 s 675407 649967 675887 650023 4 mprj_io_out[9]
port 348 nsew
rlabel metal2 s 675407 640767 675887 640823 4 mprj_io_slow_sel[9]
port 349 nsew
rlabel metal2 s 675407 651807 675887 651863 4 mprj_io_vtrip_sel[9]
port 350 nsew
rlabel metal2 s 675407 638927 675887 638983 4 mprj_io_in[9]
port 351 nsew
rlabel metal2 s 396333 995407 396389 995887 4 mprj_analog_io[11]
port 352 nsew
rlabel metal5 s 386040 1018512 398560 1031002 4 mprj_io[18]
port 353 nsew
rlabel metal2 s 393941 995407 393997 995887 4 mprj_io_analog_en[18]
port 354 nsew
rlabel metal2 s 392653 995407 392709 995887 4 mprj_io_analog_pol[18]
port 355 nsew
rlabel metal2 s 389617 995407 389673 995887 4 mprj_io_analog_sel[18]
port 356 nsew
rlabel metal2 s 393297 995407 393353 995887 4 mprj_io_dm[54]
port 357 nsew
rlabel metal2 s 395137 995407 395193 995887 4 mprj_io_dm[55]
port 358 nsew
rlabel metal2 s 388973 995407 389029 995887 4 mprj_io_dm[56]
port 359 nsew
rlabel metal2 s 390813 995407 390869 995887 4 mprj_io_enh[18]
port 360 nsew
rlabel metal2 s 390169 995407 390225 995887 4 mprj_io_hldh_n[18]
port 361 nsew
rlabel metal2 s 388329 995407 388385 995887 4 mprj_io_holdover[18]
port 362 nsew
rlabel metal2 s 385293 995407 385349 995887 4 mprj_io_ib_mode_sel[18]
port 363 nsew
rlabel metal2 s 392101 995407 392157 995887 4 mprj_io_inp_dis[18]
port 364 nsew
rlabel metal2 s 384649 995407 384705 995887 4 mprj_io_oeb[18]
port 365 nsew
rlabel metal2 s 387777 995407 387833 995887 4 mprj_io_out[18]
port 366 nsew
rlabel metal2 s 396977 995407 397033 995887 4 mprj_io_slow_sel[18]
port 367 nsew
rlabel metal2 s 385937 995407 385993 995887 4 mprj_io_vtrip_sel[18]
port 368 nsew
rlabel metal2 s 398817 995407 398873 995887 4 mprj_io_in[18]
port 369 nsew
rlabel metal2 s 41713 667333 42193 667389 4 mprj_analog_io[21]
port 370 nsew
rlabel metal5 s 6598 657040 19088 669560 4 mprj_io[28]
port 371 nsew
rlabel metal2 s 41713 664941 42193 664997 4 mprj_io_analog_en[28]
port 372 nsew
rlabel metal2 s 41713 663653 42193 663709 4 mprj_io_analog_pol[28]
port 373 nsew
rlabel metal2 s 41713 660617 42193 660673 4 mprj_io_analog_sel[28]
port 374 nsew
rlabel metal2 s 41713 664297 42193 664353 4 mprj_io_dm[84]
port 375 nsew
rlabel metal2 s 41713 666137 42193 666193 4 mprj_io_dm[85]
port 376 nsew
rlabel metal2 s 41713 659973 42193 660029 4 mprj_io_dm[86]
port 377 nsew
rlabel metal2 s 41713 661813 42193 661869 4 mprj_io_enh[28]
port 378 nsew
rlabel metal2 s 41713 661169 42193 661225 4 mprj_io_hldh_n[28]
port 379 nsew
rlabel metal2 s 41713 659329 42193 659385 4 mprj_io_holdover[28]
port 380 nsew
rlabel metal2 s 41713 656293 42193 656349 4 mprj_io_ib_mode_sel[28]
port 381 nsew
rlabel metal2 s 41713 663101 42193 663157 4 mprj_io_inp_dis[28]
port 382 nsew
rlabel metal2 s 41713 655649 42193 655705 4 mprj_io_oeb[28]
port 383 nsew
rlabel metal2 s 41713 658777 42193 658833 4 mprj_io_out[28]
port 384 nsew
rlabel metal2 s 41713 667977 42193 668033 4 mprj_io_slow_sel[28]
port 385 nsew
rlabel metal2 s 41713 656937 42193 656993 4 mprj_io_vtrip_sel[28]
port 386 nsew
rlabel metal2 s 41713 669817 42193 669873 4 mprj_io_in[28]
port 387 nsew
rlabel metal2 s 41713 624133 42193 624189 4 mprj_analog_io[22]
port 388 nsew
rlabel metal5 s 6598 613840 19088 626360 4 mprj_io[29]
port 389 nsew
rlabel metal2 s 41713 621741 42193 621797 4 mprj_io_analog_en[29]
port 390 nsew
rlabel metal2 s 41713 620453 42193 620509 4 mprj_io_analog_pol[29]
port 391 nsew
rlabel metal2 s 41713 617417 42193 617473 4 mprj_io_analog_sel[29]
port 392 nsew
rlabel metal2 s 41713 621097 42193 621153 4 mprj_io_dm[87]
port 393 nsew
rlabel metal2 s 41713 622937 42193 622993 4 mprj_io_dm[88]
port 394 nsew
rlabel metal2 s 41713 616773 42193 616829 4 mprj_io_dm[89]
port 395 nsew
rlabel metal2 s 41713 618613 42193 618669 4 mprj_io_enh[29]
port 396 nsew
rlabel metal2 s 41713 617969 42193 618025 4 mprj_io_hldh_n[29]
port 397 nsew
rlabel metal2 s 41713 616129 42193 616185 4 mprj_io_holdover[29]
port 398 nsew
rlabel metal2 s 41713 613093 42193 613149 4 mprj_io_ib_mode_sel[29]
port 399 nsew
rlabel metal2 s 41713 619901 42193 619957 4 mprj_io_inp_dis[29]
port 400 nsew
rlabel metal2 s 41713 612449 42193 612505 4 mprj_io_oeb[29]
port 401 nsew
rlabel metal2 s 41713 615577 42193 615633 4 mprj_io_out[29]
port 402 nsew
rlabel metal2 s 41713 624777 42193 624833 4 mprj_io_slow_sel[29]
port 403 nsew
rlabel metal2 s 41713 613737 42193 613793 4 mprj_io_vtrip_sel[29]
port 404 nsew
rlabel metal2 s 41713 626617 42193 626673 4 mprj_io_in[29]
port 405 nsew
rlabel metal2 s 41713 580933 42193 580989 4 mprj_analog_io[23]
port 406 nsew
rlabel metal5 s 6598 570640 19088 583160 4 mprj_io[30]
port 407 nsew
rlabel metal2 s 41713 578541 42193 578597 4 mprj_io_analog_en[30]
port 408 nsew
rlabel metal2 s 41713 577253 42193 577309 4 mprj_io_analog_pol[30]
port 409 nsew
rlabel metal2 s 41713 574217 42193 574273 4 mprj_io_analog_sel[30]
port 410 nsew
rlabel metal2 s 41713 577897 42193 577953 4 mprj_io_dm[90]
port 411 nsew
rlabel metal2 s 41713 579737 42193 579793 4 mprj_io_dm[91]
port 412 nsew
rlabel metal2 s 41713 573573 42193 573629 4 mprj_io_dm[92]
port 413 nsew
rlabel metal2 s 41713 575413 42193 575469 4 mprj_io_enh[30]
port 414 nsew
rlabel metal2 s 41713 574769 42193 574825 4 mprj_io_hldh_n[30]
port 415 nsew
rlabel metal2 s 41713 572929 42193 572985 4 mprj_io_holdover[30]
port 416 nsew
rlabel metal2 s 41713 569893 42193 569949 4 mprj_io_ib_mode_sel[30]
port 417 nsew
rlabel metal2 s 41713 576701 42193 576757 4 mprj_io_inp_dis[30]
port 418 nsew
rlabel metal2 s 41713 569249 42193 569305 4 mprj_io_oeb[30]
port 419 nsew
rlabel metal2 s 41713 572377 42193 572433 4 mprj_io_out[30]
port 420 nsew
rlabel metal2 s 41713 581577 42193 581633 4 mprj_io_slow_sel[30]
port 421 nsew
rlabel metal2 s 41713 570537 42193 570593 4 mprj_io_vtrip_sel[30]
port 422 nsew
rlabel metal2 s 41713 583417 42193 583473 4 mprj_io_in[30]
port 423 nsew
rlabel metal2 s 41713 537733 42193 537789 4 mprj_analog_io[24]
port 424 nsew
rlabel metal5 s 6598 527440 19088 539960 4 mprj_io[31]
port 425 nsew
rlabel metal2 s 41713 535341 42193 535397 4 mprj_io_analog_en[31]
port 426 nsew
rlabel metal2 s 41713 534053 42193 534109 4 mprj_io_analog_pol[31]
port 427 nsew
rlabel metal2 s 41713 531017 42193 531073 4 mprj_io_analog_sel[31]
port 428 nsew
rlabel metal2 s 41713 534697 42193 534753 4 mprj_io_dm[93]
port 429 nsew
rlabel metal2 s 41713 536537 42193 536593 4 mprj_io_dm[94]
port 430 nsew
rlabel metal2 s 41713 530373 42193 530429 4 mprj_io_dm[95]
port 431 nsew
rlabel metal2 s 41713 532213 42193 532269 4 mprj_io_enh[31]
port 432 nsew
rlabel metal2 s 41713 531569 42193 531625 4 mprj_io_hldh_n[31]
port 433 nsew
rlabel metal2 s 41713 529729 42193 529785 4 mprj_io_holdover[31]
port 434 nsew
rlabel metal2 s 41713 526693 42193 526749 4 mprj_io_ib_mode_sel[31]
port 435 nsew
rlabel metal2 s 41713 533501 42193 533557 4 mprj_io_inp_dis[31]
port 436 nsew
rlabel metal2 s 41713 526049 42193 526105 4 mprj_io_oeb[31]
port 437 nsew
rlabel metal2 s 41713 529177 42193 529233 4 mprj_io_out[31]
port 438 nsew
rlabel metal2 s 41713 538377 42193 538433 4 mprj_io_slow_sel[31]
port 439 nsew
rlabel metal2 s 41713 527337 42193 527393 4 mprj_io_vtrip_sel[31]
port 440 nsew
rlabel metal2 s 41713 540217 42193 540273 4 mprj_io_in[31]
port 441 nsew
rlabel metal2 s 41713 410133 42193 410189 4 mprj_analog_io[25]
port 442 nsew
rlabel metal5 s 6598 399840 19088 412360 4 mprj_io[32]
port 443 nsew
rlabel metal2 s 41713 407741 42193 407797 4 mprj_io_analog_en[32]
port 444 nsew
rlabel metal2 s 41713 406453 42193 406509 4 mprj_io_analog_pol[32]
port 445 nsew
rlabel metal2 s 41713 403417 42193 403473 4 mprj_io_analog_sel[32]
port 446 nsew
rlabel metal2 s 41713 407097 42193 407153 4 mprj_io_dm[96]
port 447 nsew
rlabel metal2 s 41713 408937 42193 408993 4 mprj_io_dm[97]
port 448 nsew
rlabel metal2 s 41713 402773 42193 402829 4 mprj_io_dm[98]
port 449 nsew
rlabel metal2 s 41713 404613 42193 404669 4 mprj_io_enh[32]
port 450 nsew
rlabel metal2 s 41713 403969 42193 404025 4 mprj_io_hldh_n[32]
port 451 nsew
rlabel metal2 s 41713 402129 42193 402185 4 mprj_io_holdover[32]
port 452 nsew
rlabel metal2 s 41713 399093 42193 399149 4 mprj_io_ib_mode_sel[32]
port 453 nsew
rlabel metal2 s 41713 405901 42193 405957 4 mprj_io_inp_dis[32]
port 454 nsew
rlabel metal2 s 41713 398449 42193 398505 4 mprj_io_oeb[32]
port 455 nsew
rlabel metal2 s 41713 401577 42193 401633 4 mprj_io_out[32]
port 456 nsew
rlabel metal2 s 41713 410777 42193 410833 4 mprj_io_slow_sel[32]
port 457 nsew
rlabel metal2 s 41713 399737 42193 399793 4 mprj_io_vtrip_sel[32]
port 458 nsew
rlabel metal2 s 41713 412617 42193 412673 4 mprj_io_in[32]
port 459 nsew
rlabel metal2 s 41713 366933 42193 366989 4 mprj_analog_io[26]
port 460 nsew
rlabel metal5 s 6598 356640 19088 369160 4 mprj_io[33]
port 461 nsew
rlabel metal2 s 41713 364541 42193 364597 4 mprj_io_analog_en[33]
port 462 nsew
rlabel metal2 s 41713 363253 42193 363309 4 mprj_io_analog_pol[33]
port 463 nsew
rlabel metal2 s 41713 360217 42193 360273 4 mprj_io_analog_sel[33]
port 464 nsew
rlabel metal2 s 41713 365737 42193 365793 4 mprj_io_dm[100]
port 465 nsew
rlabel metal2 s 41713 359573 42193 359629 4 mprj_io_dm[101]
port 466 nsew
rlabel metal2 s 41713 363897 42193 363953 4 mprj_io_dm[99]
port 467 nsew
rlabel metal2 s 41713 361413 42193 361469 4 mprj_io_enh[33]
port 468 nsew
rlabel metal2 s 41713 360769 42193 360825 4 mprj_io_hldh_n[33]
port 469 nsew
rlabel metal2 s 41713 358929 42193 358985 4 mprj_io_holdover[33]
port 470 nsew
rlabel metal2 s 41713 355893 42193 355949 4 mprj_io_ib_mode_sel[33]
port 471 nsew
rlabel metal2 s 41713 362701 42193 362757 4 mprj_io_inp_dis[33]
port 472 nsew
rlabel metal2 s 41713 355249 42193 355305 4 mprj_io_oeb[33]
port 473 nsew
rlabel metal2 s 41713 358377 42193 358433 4 mprj_io_out[33]
port 474 nsew
rlabel metal2 s 41713 367577 42193 367633 4 mprj_io_slow_sel[33]
port 475 nsew
rlabel metal2 s 41713 356537 42193 356593 4 mprj_io_vtrip_sel[33]
port 476 nsew
rlabel metal2 s 41713 369417 42193 369473 4 mprj_io_in[33]
port 477 nsew
rlabel metal2 s 41713 323733 42193 323789 4 mprj_analog_io[27]
port 478 nsew
rlabel metal5 s 6598 313440 19088 325960 4 mprj_io[34]
port 479 nsew
rlabel metal2 s 41713 321341 42193 321397 4 mprj_io_analog_en[34]
port 480 nsew
rlabel metal2 s 41713 320053 42193 320109 4 mprj_io_analog_pol[34]
port 481 nsew
rlabel metal2 s 41713 317017 42193 317073 4 mprj_io_analog_sel[34]
port 482 nsew
rlabel metal2 s 41713 320697 42193 320753 4 mprj_io_dm[102]
port 483 nsew
rlabel metal2 s 41713 322537 42193 322593 4 mprj_io_dm[103]
port 484 nsew
rlabel metal2 s 41713 316373 42193 316429 4 mprj_io_dm[104]
port 485 nsew
rlabel metal2 s 41713 318213 42193 318269 4 mprj_io_enh[34]
port 486 nsew
rlabel metal2 s 41713 317569 42193 317625 4 mprj_io_hldh_n[34]
port 487 nsew
rlabel metal2 s 41713 315729 42193 315785 4 mprj_io_holdover[34]
port 488 nsew
rlabel metal2 s 41713 312693 42193 312749 4 mprj_io_ib_mode_sel[34]
port 489 nsew
rlabel metal2 s 41713 319501 42193 319557 4 mprj_io_inp_dis[34]
port 490 nsew
rlabel metal2 s 41713 312049 42193 312105 4 mprj_io_oeb[34]
port 491 nsew
rlabel metal2 s 41713 315177 42193 315233 4 mprj_io_out[34]
port 492 nsew
rlabel metal2 s 41713 324377 42193 324433 4 mprj_io_slow_sel[34]
port 493 nsew
rlabel metal2 s 41713 313337 42193 313393 4 mprj_io_vtrip_sel[34]
port 494 nsew
rlabel metal2 s 41713 326217 42193 326273 4 mprj_io_in[34]
port 495 nsew
rlabel metal2 s 41713 280533 42193 280589 4 mprj_analog_io[28]
port 496 nsew
rlabel metal5 s 6598 270240 19088 282760 4 mprj_io[35]
port 497 nsew
rlabel metal2 s 41713 278141 42193 278197 4 mprj_io_analog_en[35]
port 498 nsew
rlabel metal2 s 41713 276853 42193 276909 4 mprj_io_analog_pol[35]
port 499 nsew
rlabel metal2 s 41713 273817 42193 273873 4 mprj_io_analog_sel[35]
port 500 nsew
rlabel metal2 s 41713 277497 42193 277553 4 mprj_io_dm[105]
port 501 nsew
rlabel metal2 s 41713 279337 42193 279393 4 mprj_io_dm[106]
port 502 nsew
rlabel metal2 s 41713 273173 42193 273229 4 mprj_io_dm[107]
port 503 nsew
rlabel metal2 s 41713 275013 42193 275069 4 mprj_io_enh[35]
port 504 nsew
rlabel metal2 s 41713 274369 42193 274425 4 mprj_io_hldh_n[35]
port 505 nsew
rlabel metal2 s 41713 272529 42193 272585 4 mprj_io_holdover[35]
port 506 nsew
rlabel metal2 s 41713 269493 42193 269549 4 mprj_io_ib_mode_sel[35]
port 507 nsew
rlabel metal2 s 41713 276301 42193 276357 4 mprj_io_inp_dis[35]
port 508 nsew
rlabel metal2 s 41713 268849 42193 268905 4 mprj_io_oeb[35]
port 509 nsew
rlabel metal2 s 41713 271977 42193 272033 4 mprj_io_out[35]
port 510 nsew
rlabel metal2 s 41713 281177 42193 281233 4 mprj_io_slow_sel[35]
port 511 nsew
rlabel metal2 s 41713 270137 42193 270193 4 mprj_io_vtrip_sel[35]
port 512 nsew
rlabel metal2 s 41713 283017 42193 283073 4 mprj_io_in[35]
port 513 nsew
rlabel metal2 s 41713 237333 42193 237389 4 mprj_analog_io[29]
port 514 nsew
rlabel metal5 s 6598 227040 19088 239560 4 mprj_io[36]
port 515 nsew
rlabel metal2 s 41713 234941 42193 234997 4 mprj_io_analog_en[36]
port 516 nsew
rlabel metal2 s 41713 233653 42193 233709 4 mprj_io_analog_pol[36]
port 517 nsew
rlabel metal2 s 41713 230617 42193 230673 4 mprj_io_analog_sel[36]
port 518 nsew
rlabel metal2 s 41713 234297 42193 234353 4 mprj_io_dm[108]
port 519 nsew
rlabel metal2 s 41713 236137 42193 236193 4 mprj_io_dm[109]
port 520 nsew
rlabel metal2 s 41713 229973 42193 230029 4 mprj_io_dm[110]
port 521 nsew
rlabel metal2 s 41713 231813 42193 231869 4 mprj_io_enh[36]
port 522 nsew
rlabel metal2 s 41713 231169 42193 231225 4 mprj_io_hldh_n[36]
port 523 nsew
rlabel metal2 s 41713 229329 42193 229385 4 mprj_io_holdover[36]
port 524 nsew
rlabel metal2 s 41713 226293 42193 226349 4 mprj_io_ib_mode_sel[36]
port 525 nsew
rlabel metal2 s 41713 233101 42193 233157 4 mprj_io_inp_dis[36]
port 526 nsew
rlabel metal2 s 41713 225649 42193 225705 4 mprj_io_oeb[36]
port 527 nsew
rlabel metal2 s 41713 228777 42193 228833 4 mprj_io_out[36]
port 528 nsew
rlabel metal2 s 41713 237977 42193 238033 4 mprj_io_slow_sel[36]
port 529 nsew
rlabel metal2 s 41713 226937 42193 226993 4 mprj_io_vtrip_sel[36]
port 530 nsew
rlabel metal2 s 41713 239817 42193 239873 4 mprj_io_in[36]
port 531 nsew
rlabel metal2 s 41713 194133 42193 194189 4 mprj_analog_io[30]
port 532 nsew
rlabel metal5 s 6598 183840 19088 196360 4 mprj_io[37]
port 533 nsew
rlabel metal2 s 41713 191741 42193 191797 4 mprj_io_analog_en[37]
port 534 nsew
rlabel metal2 s 41713 190453 42193 190509 4 mprj_io_analog_pol[37]
port 535 nsew
rlabel metal2 s 41713 187417 42193 187473 4 mprj_io_analog_sel[37]
port 536 nsew
rlabel metal2 s 41713 191097 42193 191153 4 mprj_io_dm[111]
port 537 nsew
rlabel metal2 s 41713 192937 42193 192993 4 mprj_io_dm[112]
port 538 nsew
rlabel metal2 s 41713 186773 42193 186829 4 mprj_io_dm[113]
port 539 nsew
rlabel metal2 s 41713 188613 42193 188669 4 mprj_io_enh[37]
port 540 nsew
rlabel metal2 s 41713 187969 42193 188025 4 mprj_io_hldh_n[37]
port 541 nsew
rlabel metal2 s 41713 186129 42193 186185 4 mprj_io_holdover[37]
port 542 nsew
rlabel metal2 s 41713 183093 42193 183149 4 mprj_io_ib_mode_sel[37]
port 543 nsew
rlabel metal2 s 41713 189901 42193 189957 4 mprj_io_inp_dis[37]
port 544 nsew
rlabel metal2 s 41713 182449 42193 182505 4 mprj_io_oeb[37]
port 545 nsew
rlabel metal2 s 41713 185577 42193 185633 4 mprj_io_out[37]
port 546 nsew
rlabel metal2 s 41713 194777 42193 194833 4 mprj_io_slow_sel[37]
port 547 nsew
rlabel metal2 s 41713 183737 42193 183793 4 mprj_io_vtrip_sel[37]
port 548 nsew
rlabel metal2 s 41713 196617 42193 196673 4 mprj_io_in[37]
port 549 nsew
rlabel metal2 s 294533 995407 294589 995887 4 mprj_analog_io[12]
port 550 nsew
rlabel metal5 s 284240 1018512 296760 1031002 4 mprj_io[19]
port 551 nsew
rlabel metal2 s 292141 995407 292197 995887 4 mprj_io_analog_en[19]
port 552 nsew
rlabel metal2 s 290853 995407 290909 995887 4 mprj_io_analog_pol[19]
port 553 nsew
rlabel metal2 s 287817 995407 287873 995887 4 mprj_io_analog_sel[19]
port 554 nsew
rlabel metal2 s 291497 995407 291553 995887 4 mprj_io_dm[57]
port 555 nsew
rlabel metal2 s 293337 995407 293393 995887 4 mprj_io_dm[58]
port 556 nsew
rlabel metal2 s 287173 995407 287229 995887 4 mprj_io_dm[59]
port 557 nsew
rlabel metal2 s 289013 995407 289069 995887 4 mprj_io_enh[19]
port 558 nsew
rlabel metal2 s 288369 995407 288425 995887 4 mprj_io_hldh_n[19]
port 559 nsew
rlabel metal2 s 286529 995407 286585 995887 4 mprj_io_holdover[19]
port 560 nsew
rlabel metal2 s 283493 995407 283549 995887 4 mprj_io_ib_mode_sel[19]
port 561 nsew
rlabel metal2 s 290301 995407 290357 995887 4 mprj_io_inp_dis[19]
port 562 nsew
rlabel metal2 s 282849 995407 282905 995887 4 mprj_io_oeb[19]
port 563 nsew
rlabel metal2 s 285977 995407 286033 995887 4 mprj_io_out[19]
port 564 nsew
rlabel metal2 s 295177 995407 295233 995887 4 mprj_io_slow_sel[19]
port 565 nsew
rlabel metal2 s 284137 995407 284193 995887 4 mprj_io_vtrip_sel[19]
port 566 nsew
rlabel metal2 s 297017 995407 297073 995887 4 mprj_io_in[19]
port 567 nsew
rlabel metal2 s 242933 995407 242989 995887 4 mprj_analog_io[13]
port 568 nsew
rlabel metal5 s 232640 1018512 245160 1031002 4 mprj_io[20]
port 569 nsew
rlabel metal2 s 240541 995407 240597 995887 4 mprj_io_analog_en[20]
port 570 nsew
rlabel metal2 s 239253 995407 239309 995887 4 mprj_io_analog_pol[20]
port 571 nsew
rlabel metal2 s 236217 995407 236273 995887 4 mprj_io_analog_sel[20]
port 572 nsew
rlabel metal2 s 239897 995407 239953 995887 4 mprj_io_dm[60]
port 573 nsew
rlabel metal2 s 241737 995407 241793 995887 4 mprj_io_dm[61]
port 574 nsew
rlabel metal2 s 235573 995407 235629 995887 4 mprj_io_dm[62]
port 575 nsew
rlabel metal2 s 237413 995407 237469 995887 4 mprj_io_enh[20]
port 576 nsew
rlabel metal2 s 236769 995407 236825 995887 4 mprj_io_hldh_n[20]
port 577 nsew
rlabel metal2 s 234929 995407 234985 995887 4 mprj_io_holdover[20]
port 578 nsew
rlabel metal2 s 231893 995407 231949 995887 4 mprj_io_ib_mode_sel[20]
port 579 nsew
rlabel metal2 s 238701 995407 238757 995887 4 mprj_io_inp_dis[20]
port 580 nsew
rlabel metal2 s 231249 995407 231305 995887 4 mprj_io_oeb[20]
port 581 nsew
rlabel metal2 s 234377 995407 234433 995887 4 mprj_io_out[20]
port 582 nsew
rlabel metal2 s 243577 995407 243633 995887 4 mprj_io_slow_sel[20]
port 583 nsew
rlabel metal2 s 232537 995407 232593 995887 4 mprj_io_vtrip_sel[20]
port 584 nsew
rlabel metal2 s 245417 995407 245473 995887 4 mprj_io_in[20]
port 585 nsew
rlabel metal2 s 191533 995407 191589 995887 4 mprj_analog_io[14]
port 586 nsew
rlabel metal5 s 181240 1018512 193760 1031002 4 mprj_io[21]
port 587 nsew
rlabel metal2 s 189141 995407 189197 995887 4 mprj_io_analog_en[21]
port 588 nsew
rlabel metal2 s 187853 995407 187909 995887 4 mprj_io_analog_pol[21]
port 589 nsew
rlabel metal2 s 184817 995407 184873 995887 4 mprj_io_analog_sel[21]
port 590 nsew
rlabel metal2 s 188497 995407 188553 995887 4 mprj_io_dm[63]
port 591 nsew
rlabel metal2 s 190337 995407 190393 995887 4 mprj_io_dm[64]
port 592 nsew
rlabel metal2 s 184173 995407 184229 995887 4 mprj_io_dm[65]
port 593 nsew
rlabel metal2 s 186013 995407 186069 995887 4 mprj_io_enh[21]
port 594 nsew
rlabel metal2 s 185369 995407 185425 995887 4 mprj_io_hldh_n[21]
port 595 nsew
rlabel metal2 s 183529 995407 183585 995887 4 mprj_io_holdover[21]
port 596 nsew
rlabel metal2 s 180493 995407 180549 995887 4 mprj_io_ib_mode_sel[21]
port 597 nsew
rlabel metal2 s 187301 995407 187357 995887 4 mprj_io_inp_dis[21]
port 598 nsew
rlabel metal2 s 179849 995407 179905 995887 4 mprj_io_oeb[21]
port 599 nsew
rlabel metal2 s 182977 995407 183033 995887 4 mprj_io_out[21]
port 600 nsew
rlabel metal2 s 192177 995407 192233 995887 4 mprj_io_slow_sel[21]
port 601 nsew
rlabel metal2 s 181137 995407 181193 995887 4 mprj_io_vtrip_sel[21]
port 602 nsew
rlabel metal2 s 194017 995407 194073 995887 4 mprj_io_in[21]
port 603 nsew
rlabel metal2 s 140133 995407 140189 995887 4 mprj_analog_io[15]
port 604 nsew
rlabel metal5 s 129840 1018512 142360 1031002 4 mprj_io[22]
port 605 nsew
rlabel metal2 s 137741 995407 137797 995887 4 mprj_io_analog_en[22]
port 606 nsew
rlabel metal2 s 136453 995407 136509 995887 4 mprj_io_analog_pol[22]
port 607 nsew
rlabel metal2 s 133417 995407 133473 995887 4 mprj_io_analog_sel[22]
port 608 nsew
rlabel metal2 s 137097 995407 137153 995887 4 mprj_io_dm[66]
port 609 nsew
rlabel metal2 s 138937 995407 138993 995887 4 mprj_io_dm[67]
port 610 nsew
rlabel metal2 s 132773 995407 132829 995887 4 mprj_io_dm[68]
port 611 nsew
rlabel metal2 s 134613 995407 134669 995887 4 mprj_io_enh[22]
port 612 nsew
rlabel metal2 s 133969 995407 134025 995887 4 mprj_io_hldh_n[22]
port 613 nsew
rlabel metal2 s 132129 995407 132185 995887 4 mprj_io_holdover[22]
port 614 nsew
rlabel metal2 s 129093 995407 129149 995887 4 mprj_io_ib_mode_sel[22]
port 615 nsew
rlabel metal2 s 135901 995407 135957 995887 4 mprj_io_inp_dis[22]
port 616 nsew
rlabel metal2 s 128449 995407 128505 995887 4 mprj_io_oeb[22]
port 617 nsew
rlabel metal2 s 131577 995407 131633 995887 4 mprj_io_out[22]
port 618 nsew
rlabel metal2 s 140777 995407 140833 995887 4 mprj_io_slow_sel[22]
port 619 nsew
rlabel metal2 s 129737 995407 129793 995887 4 mprj_io_vtrip_sel[22]
port 620 nsew
rlabel metal2 s 142617 995407 142673 995887 4 mprj_io_in[22]
port 621 nsew
rlabel metal2 s 88733 995407 88789 995887 4 mprj_analog_io[16]
port 622 nsew
rlabel metal5 s 78440 1018512 90960 1031002 4 mprj_io[23]
port 623 nsew
rlabel metal2 s 86341 995407 86397 995887 4 mprj_io_analog_en[23]
port 624 nsew
rlabel metal2 s 85053 995407 85109 995887 4 mprj_io_analog_pol[23]
port 625 nsew
rlabel metal2 s 82017 995407 82073 995887 4 mprj_io_analog_sel[23]
port 626 nsew
rlabel metal2 s 85697 995407 85753 995887 4 mprj_io_dm[69]
port 627 nsew
rlabel metal2 s 87537 995407 87593 995887 4 mprj_io_dm[70]
port 628 nsew
rlabel metal2 s 81373 995407 81429 995887 4 mprj_io_dm[71]
port 629 nsew
rlabel metal2 s 83213 995407 83269 995887 4 mprj_io_enh[23]
port 630 nsew
rlabel metal2 s 82569 995407 82625 995887 4 mprj_io_hldh_n[23]
port 631 nsew
rlabel metal2 s 80729 995407 80785 995887 4 mprj_io_holdover[23]
port 632 nsew
rlabel metal2 s 77693 995407 77749 995887 4 mprj_io_ib_mode_sel[23]
port 633 nsew
rlabel metal2 s 84501 995407 84557 995887 4 mprj_io_inp_dis[23]
port 634 nsew
rlabel metal2 s 77049 995407 77105 995887 4 mprj_io_oeb[23]
port 635 nsew
rlabel metal2 s 80177 995407 80233 995887 4 mprj_io_out[23]
port 636 nsew
rlabel metal2 s 89377 995407 89433 995887 4 mprj_io_slow_sel[23]
port 637 nsew
rlabel metal2 s 78337 995407 78393 995887 4 mprj_io_vtrip_sel[23]
port 638 nsew
rlabel metal2 s 91217 995407 91273 995887 4 mprj_io_in[23]
port 639 nsew
rlabel metal2 s 41713 966733 42193 966789 4 mprj_analog_io[17]
port 640 nsew
rlabel metal5 s 6598 956440 19088 968960 4 mprj_io[24]
port 641 nsew
rlabel metal2 s 41713 964341 42193 964397 4 mprj_io_analog_en[24]
port 642 nsew
rlabel metal2 s 41713 963053 42193 963109 4 mprj_io_analog_pol[24]
port 643 nsew
rlabel metal2 s 41713 960017 42193 960073 4 mprj_io_analog_sel[24]
port 644 nsew
rlabel metal2 s 41713 963697 42193 963753 4 mprj_io_dm[72]
port 645 nsew
rlabel metal2 s 41713 965537 42193 965593 4 mprj_io_dm[73]
port 646 nsew
rlabel metal2 s 41713 959373 42193 959429 4 mprj_io_dm[74]
port 647 nsew
rlabel metal2 s 41713 961213 42193 961269 4 mprj_io_enh[24]
port 648 nsew
rlabel metal2 s 41713 960569 42193 960625 4 mprj_io_hldh_n[24]
port 649 nsew
rlabel metal2 s 41713 958729 42193 958785 4 mprj_io_holdover[24]
port 650 nsew
rlabel metal2 s 41713 955693 42193 955749 4 mprj_io_ib_mode_sel[24]
port 651 nsew
rlabel metal2 s 41713 962501 42193 962557 4 mprj_io_inp_dis[24]
port 652 nsew
rlabel metal2 s 41713 955049 42193 955105 4 mprj_io_oeb[24]
port 653 nsew
rlabel metal2 s 41713 958177 42193 958233 4 mprj_io_out[24]
port 654 nsew
rlabel metal2 s 41713 967377 42193 967433 4 mprj_io_slow_sel[24]
port 655 nsew
rlabel metal2 s 41713 956337 42193 956393 4 mprj_io_vtrip_sel[24]
port 656 nsew
rlabel metal2 s 41713 969217 42193 969273 4 mprj_io_in[24]
port 657 nsew
rlabel metal2 s 41713 796933 42193 796989 4 mprj_analog_io[18]
port 658 nsew
rlabel metal5 s 6598 786640 19088 799160 4 mprj_io[25]
port 659 nsew
rlabel metal2 s 41713 794541 42193 794597 4 mprj_io_analog_en[25]
port 660 nsew
rlabel metal2 s 41713 793253 42193 793309 4 mprj_io_analog_pol[25]
port 661 nsew
rlabel metal2 s 41713 790217 42193 790273 4 mprj_io_analog_sel[25]
port 662 nsew
rlabel metal2 s 41713 793897 42193 793953 4 mprj_io_dm[75]
port 663 nsew
rlabel metal2 s 41713 795737 42193 795793 4 mprj_io_dm[76]
port 664 nsew
rlabel metal2 s 41713 789573 42193 789629 4 mprj_io_dm[77]
port 665 nsew
rlabel metal2 s 41713 791413 42193 791469 4 mprj_io_enh[25]
port 666 nsew
rlabel metal2 s 41713 790769 42193 790825 4 mprj_io_hldh_n[25]
port 667 nsew
rlabel metal2 s 41713 788929 42193 788985 4 mprj_io_holdover[25]
port 668 nsew
rlabel metal2 s 41713 785893 42193 785949 4 mprj_io_ib_mode_sel[25]
port 669 nsew
rlabel metal2 s 41713 792701 42193 792757 4 mprj_io_inp_dis[25]
port 670 nsew
rlabel metal2 s 41713 785249 42193 785305 4 mprj_io_oeb[25]
port 671 nsew
rlabel metal2 s 41713 788377 42193 788433 4 mprj_io_out[25]
port 672 nsew
rlabel metal2 s 41713 797577 42193 797633 4 mprj_io_slow_sel[25]
port 673 nsew
rlabel metal2 s 41713 786537 42193 786593 4 mprj_io_vtrip_sel[25]
port 674 nsew
rlabel metal2 s 41713 799417 42193 799473 4 mprj_io_in[25]
port 675 nsew
rlabel metal2 s 41713 753733 42193 753789 4 mprj_analog_io[19]
port 676 nsew
rlabel metal5 s 6598 743440 19088 755960 4 mprj_io[26]
port 677 nsew
rlabel metal2 s 41713 751341 42193 751397 4 mprj_io_analog_en[26]
port 678 nsew
rlabel metal2 s 41713 750053 42193 750109 4 mprj_io_analog_pol[26]
port 679 nsew
rlabel metal2 s 41713 747017 42193 747073 4 mprj_io_analog_sel[26]
port 680 nsew
rlabel metal2 s 41713 750697 42193 750753 4 mprj_io_dm[78]
port 681 nsew
rlabel metal2 s 41713 752537 42193 752593 4 mprj_io_dm[79]
port 682 nsew
rlabel metal2 s 41713 746373 42193 746429 4 mprj_io_dm[80]
port 683 nsew
rlabel metal2 s 41713 748213 42193 748269 4 mprj_io_enh[26]
port 684 nsew
rlabel metal2 s 41713 747569 42193 747625 4 mprj_io_hldh_n[26]
port 685 nsew
rlabel metal2 s 41713 745729 42193 745785 4 mprj_io_holdover[26]
port 686 nsew
rlabel metal2 s 41713 742693 42193 742749 4 mprj_io_ib_mode_sel[26]
port 687 nsew
rlabel metal2 s 41713 749501 42193 749557 4 mprj_io_inp_dis[26]
port 688 nsew
rlabel metal2 s 41713 742049 42193 742105 4 mprj_io_oeb[26]
port 689 nsew
rlabel metal2 s 41713 745177 42193 745233 4 mprj_io_out[26]
port 690 nsew
rlabel metal2 s 41713 754377 42193 754433 4 mprj_io_slow_sel[26]
port 691 nsew
rlabel metal2 s 41713 743337 42193 743393 4 mprj_io_vtrip_sel[26]
port 692 nsew
rlabel metal2 s 41713 756217 42193 756273 4 mprj_io_in[26]
port 693 nsew
rlabel metal2 s 41713 710533 42193 710589 4 mprj_analog_io[20]
port 694 nsew
rlabel metal5 s 6598 700240 19088 712760 4 mprj_io[27]
port 695 nsew
rlabel metal2 s 41713 708141 42193 708197 4 mprj_io_analog_en[27]
port 696 nsew
rlabel metal2 s 41713 706853 42193 706909 4 mprj_io_analog_pol[27]
port 697 nsew
rlabel metal2 s 41713 703817 42193 703873 4 mprj_io_analog_sel[27]
port 698 nsew
rlabel metal2 s 41713 707497 42193 707553 4 mprj_io_dm[81]
port 699 nsew
rlabel metal2 s 41713 709337 42193 709393 4 mprj_io_dm[82]
port 700 nsew
rlabel metal2 s 41713 703173 42193 703229 4 mprj_io_dm[83]
port 701 nsew
rlabel metal2 s 41713 705013 42193 705069 4 mprj_io_enh[27]
port 702 nsew
rlabel metal2 s 41713 704369 42193 704425 4 mprj_io_hldh_n[27]
port 703 nsew
rlabel metal2 s 41713 702529 42193 702585 4 mprj_io_holdover[27]
port 704 nsew
rlabel metal2 s 41713 699493 42193 699549 4 mprj_io_ib_mode_sel[27]
port 705 nsew
rlabel metal2 s 41713 706301 42193 706357 4 mprj_io_inp_dis[27]
port 706 nsew
rlabel metal2 s 41713 698849 42193 698905 4 mprj_io_oeb[27]
port 707 nsew
rlabel metal2 s 41713 701977 42193 702033 4 mprj_io_out[27]
port 708 nsew
rlabel metal2 s 41713 711177 42193 711233 4 mprj_io_slow_sel[27]
port 709 nsew
rlabel metal2 s 41713 700137 42193 700193 4 mprj_io_vtrip_sel[27]
port 710 nsew
rlabel metal2 s 41713 713017 42193 713073 4 mprj_io_in[27]
port 711 nsew
rlabel metal2 s 145091 39706 145143 40000 4 porb_h
port 712 nsew
rlabel metal5 s 136713 7143 144149 18309 4 resetb
port 713 nsew
rlabel metal3 s 141667 38031 141813 39999 4 resetb_core_h
port 714 nsew
rlabel metal5 s 698028 909409 711514 920737 4 vccd1
port 715 nsew
rlabel metal5 s 698402 819640 710924 832180 4 vdda1
port 716 nsew
rlabel metal5 s 576820 1018402 589360 1030924 4 vssa1
port 717 nsew
rlabel metal5 s 698028 461609 711514 472937 4 vssd1
port 718 nsew
rlabel metal5 s 6086 913863 19572 925191 4 vccd2
port 719 nsew
rlabel metal5 s 6675 484220 19197 496760 4 vdda2
port 720 nsew
rlabel metal5 s 6675 828820 19197 841360 4 vssa2
port 721 nsew
rlabel metal5 s 6086 442663 19572 453991 4 vssd2
port 722 nsew
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
string GDS_FILE /project/openlane/chip_io/runs/chip_io/results/magic/chip_io.gds
string GDS_END 35122950
string GDS_START 34578978
<< end >>
