magic
tech sky130A
magscale 1 2
timestamp 1622551585
<< obsli1 >>
rect 1104 1071 72864 3825
<< obsm1 >>
rect 566 1040 72864 4004
<< metal2 >>
rect 570 4000 626 5000
rect 846 4000 902 5000
rect 1122 4000 1178 5000
rect 1398 4000 1454 5000
rect 1674 4000 1730 5000
rect 1950 4000 2006 5000
rect 2226 4000 2282 5000
rect 2502 4000 2558 5000
rect 2778 4000 2834 5000
rect 3054 4000 3110 5000
rect 3330 4000 3386 5000
rect 3606 4000 3662 5000
rect 3882 4000 3938 5000
rect 4158 4000 4214 5000
rect 4434 4000 4490 5000
rect 4710 4000 4766 5000
rect 4986 4000 5042 5000
rect 5262 4000 5318 5000
rect 5538 4000 5594 5000
rect 5814 4000 5870 5000
rect 6090 4000 6146 5000
rect 6366 4000 6422 5000
rect 6642 4000 6698 5000
rect 6918 4000 6974 5000
rect 7194 4000 7250 5000
rect 7470 4000 7526 5000
rect 7746 4000 7802 5000
rect 8022 4000 8078 5000
rect 8298 4000 8354 5000
rect 8574 4000 8630 5000
rect 8850 4000 8906 5000
rect 9126 4000 9182 5000
rect 9402 4000 9458 5000
rect 9678 4000 9734 5000
rect 9954 4000 10010 5000
rect 10230 4000 10286 5000
rect 10506 4000 10562 5000
rect 10782 4000 10838 5000
rect 11058 4000 11114 5000
rect 11334 4000 11390 5000
rect 11610 4000 11666 5000
rect 11886 4000 11942 5000
rect 12162 4000 12218 5000
rect 12438 4000 12494 5000
rect 12714 4000 12770 5000
rect 12990 4000 13046 5000
rect 13266 4000 13322 5000
rect 13542 4000 13598 5000
rect 13818 4000 13874 5000
rect 14094 4000 14150 5000
rect 14370 4000 14426 5000
rect 14646 4000 14702 5000
rect 14922 4000 14978 5000
rect 15198 4000 15254 5000
rect 15474 4000 15530 5000
rect 15750 4000 15806 5000
rect 16026 4000 16082 5000
rect 16302 4000 16358 5000
rect 16578 4000 16634 5000
rect 16854 4000 16910 5000
rect 17130 4000 17186 5000
rect 17406 4000 17462 5000
rect 17682 4000 17738 5000
rect 17958 4000 18014 5000
rect 18234 4000 18290 5000
rect 18510 4000 18566 5000
rect 18786 4000 18842 5000
rect 19062 4000 19118 5000
rect 19338 4000 19394 5000
rect 19614 4000 19670 5000
rect 19890 4000 19946 5000
rect 20166 4000 20222 5000
rect 20442 4000 20498 5000
rect 20718 4000 20774 5000
rect 20994 4000 21050 5000
rect 21270 4000 21326 5000
rect 21546 4000 21602 5000
rect 21822 4000 21878 5000
rect 22098 4000 22154 5000
rect 22374 4000 22430 5000
rect 22650 4000 22706 5000
rect 22926 4000 22982 5000
rect 23202 4000 23258 5000
rect 23478 4000 23534 5000
rect 23754 4000 23810 5000
rect 24030 4000 24086 5000
rect 24306 4000 24362 5000
rect 24582 4000 24638 5000
rect 24858 4000 24914 5000
rect 25134 4000 25190 5000
rect 25410 4000 25466 5000
rect 25686 4000 25742 5000
rect 25962 4000 26018 5000
rect 26238 4000 26294 5000
rect 26514 4000 26570 5000
rect 26790 4000 26846 5000
rect 27066 4000 27122 5000
rect 27342 4000 27398 5000
rect 27618 4000 27674 5000
rect 27894 4000 27950 5000
rect 28170 4000 28226 5000
rect 28446 4000 28502 5000
rect 28722 4000 28778 5000
rect 28998 4000 29054 5000
rect 29274 4000 29330 5000
rect 29550 4000 29606 5000
rect 29826 4000 29882 5000
rect 30102 4000 30158 5000
rect 30378 4000 30434 5000
rect 36174 4000 36230 5000
rect 36450 4000 36506 5000
rect 36726 4000 36782 5000
rect 37002 4000 37058 5000
rect 37278 4000 37334 5000
rect 37554 4000 37610 5000
rect 37830 4000 37886 5000
rect 38106 4000 38162 5000
rect 38382 4000 38438 5000
rect 38658 4000 38714 5000
rect 38934 4000 38990 5000
rect 39210 4000 39266 5000
rect 39486 4000 39542 5000
rect 39762 4000 39818 5000
rect 40038 4000 40094 5000
rect 40314 4000 40370 5000
rect 40590 4000 40646 5000
rect 40866 4000 40922 5000
rect 41142 4000 41198 5000
rect 41418 4000 41474 5000
rect 41694 4000 41750 5000
rect 41970 4000 42026 5000
rect 42246 4000 42302 5000
rect 42522 4000 42578 5000
rect 42798 4000 42854 5000
rect 43074 4000 43130 5000
rect 43350 4000 43406 5000
rect 43626 4000 43682 5000
rect 43902 4000 43958 5000
rect 44178 4000 44234 5000
rect 44454 4000 44510 5000
rect 44730 4000 44786 5000
rect 45006 4000 45062 5000
rect 45282 4000 45338 5000
rect 45558 4000 45614 5000
rect 45834 4000 45890 5000
rect 46110 4000 46166 5000
rect 46386 4000 46442 5000
rect 46662 4000 46718 5000
rect 46938 4000 46994 5000
rect 47214 4000 47270 5000
rect 47490 4000 47546 5000
rect 47766 4000 47822 5000
rect 48042 4000 48098 5000
rect 48318 4000 48374 5000
rect 48594 4000 48650 5000
rect 48870 4000 48926 5000
rect 49146 4000 49202 5000
rect 49422 4000 49478 5000
rect 49698 4000 49754 5000
rect 49974 4000 50030 5000
rect 50250 4000 50306 5000
rect 50526 4000 50582 5000
rect 50802 4000 50858 5000
rect 51078 4000 51134 5000
rect 51354 4000 51410 5000
rect 51630 4000 51686 5000
rect 51906 4000 51962 5000
rect 52182 4000 52238 5000
rect 52458 4000 52514 5000
rect 52734 4000 52790 5000
rect 53010 4000 53066 5000
rect 53286 4000 53342 5000
rect 53562 4000 53618 5000
rect 53838 4000 53894 5000
rect 54114 4000 54170 5000
rect 54390 4000 54446 5000
rect 54666 4000 54722 5000
rect 54942 4000 54998 5000
rect 55218 4000 55274 5000
rect 55494 4000 55550 5000
rect 55770 4000 55826 5000
rect 56046 4000 56102 5000
rect 56322 4000 56378 5000
rect 56598 4000 56654 5000
rect 56874 4000 56930 5000
rect 57150 4000 57206 5000
rect 57426 4000 57482 5000
rect 57702 4000 57758 5000
rect 57978 4000 58034 5000
rect 58254 4000 58310 5000
rect 58530 4000 58586 5000
rect 58806 4000 58862 5000
rect 59082 4000 59138 5000
rect 59358 4000 59414 5000
rect 59634 4000 59690 5000
rect 59910 4000 59966 5000
rect 60186 4000 60242 5000
rect 60462 4000 60518 5000
rect 60738 4000 60794 5000
rect 61014 4000 61070 5000
rect 61290 4000 61346 5000
rect 61566 4000 61622 5000
rect 61842 4000 61898 5000
rect 62118 4000 62174 5000
rect 62394 4000 62450 5000
rect 62670 4000 62726 5000
rect 62946 4000 63002 5000
rect 63222 4000 63278 5000
rect 63498 4000 63554 5000
rect 63774 4000 63830 5000
rect 64050 4000 64106 5000
rect 64326 4000 64382 5000
rect 64602 4000 64658 5000
rect 64878 4000 64934 5000
rect 65154 4000 65210 5000
rect 65430 4000 65486 5000
rect 65706 4000 65762 5000
rect 65982 4000 66038 5000
rect 66258 4000 66314 5000
rect 66534 4000 66590 5000
rect 66810 4000 66866 5000
rect 67086 4000 67142 5000
rect 67362 4000 67418 5000
rect 570 0 626 1000
rect 846 0 902 1000
rect 1122 0 1178 1000
rect 1398 0 1454 1000
rect 1674 0 1730 1000
rect 1950 0 2006 1000
rect 2226 0 2282 1000
rect 2502 0 2558 1000
rect 2778 0 2834 1000
rect 3054 1040 3154 3856
rect 3054 0 3110 1000
rect 3330 0 3386 1000
rect 3606 0 3662 1000
rect 3882 0 3938 1000
rect 4158 0 4214 1000
rect 4434 0 4490 1000
rect 4710 0 4766 1000
rect 4986 0 5042 1000
rect 5262 0 5318 1000
rect 5538 0 5594 1000
rect 5814 0 5870 1000
rect 6090 0 6146 1000
rect 6366 0 6422 1000
rect 6642 0 6698 1000
rect 6918 0 6974 1000
rect 7194 0 7250 1000
rect 7470 0 7526 1000
rect 7746 0 7802 1000
rect 8022 0 8078 1000
rect 8298 0 8354 1000
rect 8574 0 8630 1000
rect 8850 0 8906 1000
rect 9054 1040 9154 3856
rect 9126 0 9182 1000
rect 9402 0 9458 1000
rect 9678 0 9734 1000
rect 9954 0 10010 1000
rect 10230 0 10286 1000
rect 10506 0 10562 1000
rect 10782 0 10838 1000
rect 11058 0 11114 1000
rect 11334 0 11390 1000
rect 11610 0 11666 1000
rect 11886 0 11942 1000
rect 12162 0 12218 1000
rect 12438 0 12494 1000
rect 12714 0 12770 1000
rect 12990 0 13046 1000
rect 13266 0 13322 1000
rect 13542 0 13598 1000
rect 13818 0 13874 1000
rect 14094 0 14150 1000
rect 14370 0 14426 1000
rect 14646 0 14702 1000
rect 15054 1040 15154 3856
rect 14922 0 14978 1000
rect 15198 0 15254 1000
rect 15474 0 15530 1000
rect 15750 0 15806 1000
rect 16026 0 16082 1000
rect 16302 0 16358 1000
rect 16578 0 16634 1000
rect 16854 0 16910 1000
rect 17130 0 17186 1000
rect 17406 0 17462 1000
rect 17682 0 17738 1000
rect 17958 0 18014 1000
rect 18234 0 18290 1000
rect 18510 0 18566 1000
rect 18786 0 18842 1000
rect 19062 0 19118 1000
rect 19338 0 19394 1000
rect 19614 0 19670 1000
rect 19890 0 19946 1000
rect 20166 0 20222 1000
rect 20442 0 20498 1000
rect 20718 0 20774 1000
rect 21054 1040 21154 3856
rect 20994 0 21050 1000
rect 21270 0 21326 1000
rect 21546 0 21602 1000
rect 21822 0 21878 1000
rect 22098 0 22154 1000
rect 22374 0 22430 1000
rect 22650 0 22706 1000
rect 22926 0 22982 1000
rect 23202 0 23258 1000
rect 23478 0 23534 1000
rect 23754 0 23810 1000
rect 24030 0 24086 1000
rect 24306 0 24362 1000
rect 24582 0 24638 1000
rect 24858 0 24914 1000
rect 25134 0 25190 1000
rect 25410 0 25466 1000
rect 25686 0 25742 1000
rect 25962 0 26018 1000
rect 26238 0 26294 1000
rect 26514 0 26570 1000
rect 26790 0 26846 1000
rect 27054 1040 27154 3856
rect 27066 0 27122 1000
rect 27342 0 27398 1000
rect 27618 0 27674 1000
rect 27894 0 27950 1000
rect 28170 0 28226 1000
rect 28446 0 28502 1000
rect 28722 0 28778 1000
rect 28998 0 29054 1000
rect 29274 0 29330 1000
rect 29550 0 29606 1000
rect 29826 0 29882 1000
rect 30102 0 30158 1000
rect 30378 0 30434 1000
rect 30654 0 30710 1000
rect 30930 0 30986 1000
rect 31206 0 31262 1000
rect 31482 0 31538 1000
rect 31758 0 31814 1000
rect 32034 0 32090 1000
rect 32310 0 32366 1000
rect 33054 1040 33154 3856
rect 38106 0 38162 1000
rect 38382 0 38438 1000
rect 38658 0 38714 1000
rect 39054 1040 39154 3856
rect 38934 0 38990 1000
rect 39210 0 39266 1000
rect 39486 0 39542 1000
rect 39762 0 39818 1000
rect 40038 0 40094 1000
rect 40314 0 40370 1000
rect 40590 0 40646 1000
rect 40866 0 40922 1000
rect 41142 0 41198 1000
rect 41418 0 41474 1000
rect 41694 0 41750 1000
rect 41970 0 42026 1000
rect 42246 0 42302 1000
rect 42522 0 42578 1000
rect 42798 0 42854 1000
rect 43074 0 43130 1000
rect 43350 0 43406 1000
rect 43626 0 43682 1000
rect 43902 0 43958 1000
rect 44178 0 44234 1000
rect 44454 0 44510 1000
rect 44730 0 44786 1000
rect 45054 1040 45154 3856
rect 45006 0 45062 1000
rect 45282 0 45338 1000
rect 45558 0 45614 1000
rect 45834 0 45890 1000
rect 46110 0 46166 1000
rect 46386 0 46442 1000
rect 46662 0 46718 1000
rect 46938 0 46994 1000
rect 47214 0 47270 1000
rect 47490 0 47546 1000
rect 47766 0 47822 1000
rect 48042 0 48098 1000
rect 48318 0 48374 1000
rect 48594 0 48650 1000
rect 48870 0 48926 1000
rect 49146 0 49202 1000
rect 49422 0 49478 1000
rect 49698 0 49754 1000
rect 49974 0 50030 1000
rect 50250 0 50306 1000
rect 50526 0 50582 1000
rect 50802 0 50858 1000
rect 51054 1040 51154 3856
rect 51078 0 51134 1000
rect 51354 0 51410 1000
rect 51630 0 51686 1000
rect 51906 0 51962 1000
rect 52182 0 52238 1000
rect 52458 0 52514 1000
rect 52734 0 52790 1000
rect 53010 0 53066 1000
rect 53286 0 53342 1000
rect 53562 0 53618 1000
rect 53838 0 53894 1000
rect 54114 0 54170 1000
rect 54390 0 54446 1000
rect 54666 0 54722 1000
rect 54942 0 54998 1000
rect 55218 0 55274 1000
rect 55494 0 55550 1000
rect 55770 0 55826 1000
rect 56046 0 56102 1000
rect 56322 0 56378 1000
rect 56598 0 56654 1000
rect 56874 0 56930 1000
rect 57054 1040 57154 3856
rect 57150 0 57206 1000
rect 57426 0 57482 1000
rect 57702 0 57758 1000
rect 57978 0 58034 1000
rect 58254 0 58310 1000
rect 58530 0 58586 1000
rect 58806 0 58862 1000
rect 59082 0 59138 1000
rect 59358 0 59414 1000
rect 59634 0 59690 1000
rect 59910 0 59966 1000
rect 60186 0 60242 1000
rect 60462 0 60518 1000
rect 60738 0 60794 1000
rect 61014 0 61070 1000
rect 61290 0 61346 1000
rect 61566 0 61622 1000
rect 61842 0 61898 1000
rect 62118 0 62174 1000
rect 62394 0 62450 1000
rect 62670 0 62726 1000
rect 63054 1040 63154 3856
rect 62946 0 63002 1000
rect 63222 0 63278 1000
rect 63498 0 63554 1000
rect 63774 0 63830 1000
rect 64050 0 64106 1000
rect 64326 0 64382 1000
rect 64602 0 64658 1000
rect 64878 0 64934 1000
rect 65154 0 65210 1000
rect 65430 0 65486 1000
rect 65706 0 65762 1000
rect 65982 0 66038 1000
rect 66258 0 66314 1000
rect 66534 0 66590 1000
rect 66810 0 66866 1000
rect 67086 0 67142 1000
rect 67362 0 67418 1000
rect 67638 0 67694 1000
rect 67914 0 67970 1000
rect 68190 0 68246 1000
rect 68466 0 68522 1000
rect 68742 0 68798 1000
rect 69054 1040 69154 3856
rect 69018 0 69074 1000
rect 69294 0 69350 1000
rect 69570 0 69626 1000
rect 69846 0 69902 1000
<< obsm2 >>
rect 682 3944 790 4010
rect 958 3944 1066 4010
rect 1234 3944 1342 4010
rect 1510 3944 1618 4010
rect 1786 3944 1894 4010
rect 2062 3944 2170 4010
rect 2338 3944 2446 4010
rect 2614 3944 2722 4010
rect 2890 3944 2998 4010
rect 3166 3944 3274 4010
rect 3442 3944 3550 4010
rect 3718 3944 3826 4010
rect 3994 3944 4102 4010
rect 4270 3944 4378 4010
rect 4546 3944 4654 4010
rect 4822 3944 4930 4010
rect 5098 3944 5206 4010
rect 5374 3944 5482 4010
rect 5650 3944 5758 4010
rect 5926 3944 6034 4010
rect 6202 3944 6310 4010
rect 6478 3944 6586 4010
rect 6754 3944 6862 4010
rect 7030 3944 7138 4010
rect 7306 3944 7414 4010
rect 7582 3944 7690 4010
rect 7858 3944 7966 4010
rect 8134 3944 8242 4010
rect 8410 3944 8518 4010
rect 8686 3944 8794 4010
rect 8962 3944 9070 4010
rect 9238 3944 9346 4010
rect 9514 3944 9622 4010
rect 9790 3944 9898 4010
rect 10066 3944 10174 4010
rect 10342 3944 10450 4010
rect 10618 3944 10726 4010
rect 10894 3944 11002 4010
rect 11170 3944 11278 4010
rect 11446 3944 11554 4010
rect 11722 3944 11830 4010
rect 11998 3944 12106 4010
rect 12274 3944 12382 4010
rect 12550 3944 12658 4010
rect 12826 3944 12934 4010
rect 13102 3944 13210 4010
rect 13378 3944 13486 4010
rect 13654 3944 13762 4010
rect 13930 3944 14038 4010
rect 14206 3944 14314 4010
rect 14482 3944 14590 4010
rect 14758 3944 14866 4010
rect 15034 3944 15142 4010
rect 15310 3944 15418 4010
rect 15586 3944 15694 4010
rect 15862 3944 15970 4010
rect 16138 3944 16246 4010
rect 16414 3944 16522 4010
rect 16690 3944 16798 4010
rect 16966 3944 17074 4010
rect 17242 3944 17350 4010
rect 17518 3944 17626 4010
rect 17794 3944 17902 4010
rect 18070 3944 18178 4010
rect 18346 3944 18454 4010
rect 18622 3944 18730 4010
rect 18898 3944 19006 4010
rect 19174 3944 19282 4010
rect 19450 3944 19558 4010
rect 19726 3944 19834 4010
rect 20002 3944 20110 4010
rect 20278 3944 20386 4010
rect 20554 3944 20662 4010
rect 20830 3944 20938 4010
rect 21106 3944 21214 4010
rect 21382 3944 21490 4010
rect 21658 3944 21766 4010
rect 21934 3944 22042 4010
rect 22210 3944 22318 4010
rect 22486 3944 22594 4010
rect 22762 3944 22870 4010
rect 23038 3944 23146 4010
rect 23314 3944 23422 4010
rect 23590 3944 23698 4010
rect 23866 3944 23974 4010
rect 24142 3944 24250 4010
rect 24418 3944 24526 4010
rect 24694 3944 24802 4010
rect 24970 3944 25078 4010
rect 25246 3944 25354 4010
rect 25522 3944 25630 4010
rect 25798 3944 25906 4010
rect 26074 3944 26182 4010
rect 26350 3944 26458 4010
rect 26626 3944 26734 4010
rect 26902 3944 27010 4010
rect 27178 3944 27286 4010
rect 27454 3944 27562 4010
rect 27730 3944 27838 4010
rect 28006 3944 28114 4010
rect 28282 3944 28390 4010
rect 28558 3944 28666 4010
rect 28834 3944 28942 4010
rect 29110 3944 29218 4010
rect 29386 3944 29494 4010
rect 29662 3944 29770 4010
rect 29938 3944 30046 4010
rect 30214 3944 30322 4010
rect 30490 3944 36118 4010
rect 36286 3944 36394 4010
rect 36562 3944 36670 4010
rect 36838 3944 36946 4010
rect 37114 3944 37222 4010
rect 37390 3944 37498 4010
rect 37666 3944 37774 4010
rect 37942 3944 38050 4010
rect 38218 3944 38326 4010
rect 38494 3944 38602 4010
rect 38770 3944 38878 4010
rect 39046 3944 39154 4010
rect 39322 3944 39430 4010
rect 39598 3944 39706 4010
rect 39874 3944 39982 4010
rect 40150 3944 40258 4010
rect 40426 3944 40534 4010
rect 40702 3944 40810 4010
rect 40978 3944 41086 4010
rect 41254 3944 41362 4010
rect 41530 3944 41638 4010
rect 41806 3944 41914 4010
rect 42082 3944 42190 4010
rect 42358 3944 42466 4010
rect 42634 3944 42742 4010
rect 42910 3944 43018 4010
rect 43186 3944 43294 4010
rect 43462 3944 43570 4010
rect 43738 3944 43846 4010
rect 44014 3944 44122 4010
rect 44290 3944 44398 4010
rect 44566 3944 44674 4010
rect 44842 3944 44950 4010
rect 45118 3944 45226 4010
rect 45394 3944 45502 4010
rect 45670 3944 45778 4010
rect 45946 3944 46054 4010
rect 46222 3944 46330 4010
rect 46498 3944 46606 4010
rect 46774 3944 46882 4010
rect 47050 3944 47158 4010
rect 47326 3944 47434 4010
rect 47602 3944 47710 4010
rect 47878 3944 47986 4010
rect 48154 3944 48262 4010
rect 48430 3944 48538 4010
rect 48706 3944 48814 4010
rect 48982 3944 49090 4010
rect 49258 3944 49366 4010
rect 49534 3944 49642 4010
rect 49810 3944 49918 4010
rect 50086 3944 50194 4010
rect 50362 3944 50470 4010
rect 50638 3944 50746 4010
rect 50914 3944 51022 4010
rect 51190 3944 51298 4010
rect 51466 3944 51574 4010
rect 51742 3944 51850 4010
rect 52018 3944 52126 4010
rect 52294 3944 52402 4010
rect 52570 3944 52678 4010
rect 52846 3944 52954 4010
rect 53122 3944 53230 4010
rect 53398 3944 53506 4010
rect 53674 3944 53782 4010
rect 53950 3944 54058 4010
rect 54226 3944 54334 4010
rect 54502 3944 54610 4010
rect 54778 3944 54886 4010
rect 55054 3944 55162 4010
rect 55330 3944 55438 4010
rect 55606 3944 55714 4010
rect 55882 3944 55990 4010
rect 56158 3944 56266 4010
rect 56434 3944 56542 4010
rect 56710 3944 56818 4010
rect 56986 3944 57094 4010
rect 57262 3944 57370 4010
rect 57538 3944 57646 4010
rect 57814 3944 57922 4010
rect 58090 3944 58198 4010
rect 58366 3944 58474 4010
rect 58642 3944 58750 4010
rect 58918 3944 59026 4010
rect 59194 3944 59302 4010
rect 59470 3944 59578 4010
rect 59746 3944 59854 4010
rect 60022 3944 60130 4010
rect 60298 3944 60406 4010
rect 60574 3944 60682 4010
rect 60850 3944 60958 4010
rect 61126 3944 61234 4010
rect 61402 3944 61510 4010
rect 61678 3944 61786 4010
rect 61954 3944 62062 4010
rect 62230 3944 62338 4010
rect 62506 3944 62614 4010
rect 62782 3944 62890 4010
rect 63058 3944 63166 4010
rect 63334 3944 63442 4010
rect 63610 3944 63718 4010
rect 63886 3944 63994 4010
rect 64162 3944 64270 4010
rect 64438 3944 64546 4010
rect 64714 3944 64822 4010
rect 64990 3944 65098 4010
rect 65266 3944 65374 4010
rect 65542 3944 65650 4010
rect 65818 3944 65926 4010
rect 66094 3944 66202 4010
rect 66370 3944 66478 4010
rect 66646 3944 66754 4010
rect 66922 3944 67030 4010
rect 67198 3944 67306 4010
rect 67474 3944 69900 4010
rect 572 3912 69900 3944
rect 572 1056 2998 3912
rect 682 870 790 1056
rect 958 870 1066 1056
rect 1234 870 1342 1056
rect 1510 870 1618 1056
rect 1786 870 1894 1056
rect 2062 870 2170 1056
rect 2338 870 2446 1056
rect 2614 870 2722 1056
rect 2890 870 2998 1056
rect 3210 1056 8998 3912
rect 3210 984 3274 1056
rect 3166 870 3274 984
rect 3442 870 3550 1056
rect 3718 870 3826 1056
rect 3994 870 4102 1056
rect 4270 870 4378 1056
rect 4546 870 4654 1056
rect 4822 870 4930 1056
rect 5098 870 5206 1056
rect 5374 870 5482 1056
rect 5650 870 5758 1056
rect 5926 870 6034 1056
rect 6202 870 6310 1056
rect 6478 870 6586 1056
rect 6754 870 6862 1056
rect 7030 870 7138 1056
rect 7306 870 7414 1056
rect 7582 870 7690 1056
rect 7858 870 7966 1056
rect 8134 870 8242 1056
rect 8410 870 8518 1056
rect 8686 870 8794 1056
rect 8962 984 8998 1056
rect 9210 1056 14998 3912
rect 8962 870 9070 984
rect 9238 870 9346 1056
rect 9514 870 9622 1056
rect 9790 870 9898 1056
rect 10066 870 10174 1056
rect 10342 870 10450 1056
rect 10618 870 10726 1056
rect 10894 870 11002 1056
rect 11170 870 11278 1056
rect 11446 870 11554 1056
rect 11722 870 11830 1056
rect 11998 870 12106 1056
rect 12274 870 12382 1056
rect 12550 870 12658 1056
rect 12826 870 12934 1056
rect 13102 870 13210 1056
rect 13378 870 13486 1056
rect 13654 870 13762 1056
rect 13930 870 14038 1056
rect 14206 870 14314 1056
rect 14482 870 14590 1056
rect 14758 870 14866 1056
rect 15210 1056 20998 3912
rect 15034 870 15142 984
rect 15310 870 15418 1056
rect 15586 870 15694 1056
rect 15862 870 15970 1056
rect 16138 870 16246 1056
rect 16414 870 16522 1056
rect 16690 870 16798 1056
rect 16966 870 17074 1056
rect 17242 870 17350 1056
rect 17518 870 17626 1056
rect 17794 870 17902 1056
rect 18070 870 18178 1056
rect 18346 870 18454 1056
rect 18622 870 18730 1056
rect 18898 870 19006 1056
rect 19174 870 19282 1056
rect 19450 870 19558 1056
rect 19726 870 19834 1056
rect 20002 870 20110 1056
rect 20278 870 20386 1056
rect 20554 870 20662 1056
rect 20830 870 20938 1056
rect 21210 1056 26998 3912
rect 21210 984 21214 1056
rect 21106 870 21214 984
rect 21382 870 21490 1056
rect 21658 870 21766 1056
rect 21934 870 22042 1056
rect 22210 870 22318 1056
rect 22486 870 22594 1056
rect 22762 870 22870 1056
rect 23038 870 23146 1056
rect 23314 870 23422 1056
rect 23590 870 23698 1056
rect 23866 870 23974 1056
rect 24142 870 24250 1056
rect 24418 870 24526 1056
rect 24694 870 24802 1056
rect 24970 870 25078 1056
rect 25246 870 25354 1056
rect 25522 870 25630 1056
rect 25798 870 25906 1056
rect 26074 870 26182 1056
rect 26350 870 26458 1056
rect 26626 870 26734 1056
rect 26902 984 26998 1056
rect 27210 1056 32998 3912
rect 26902 870 27010 984
rect 27210 984 27286 1056
rect 27178 870 27286 984
rect 27454 870 27562 1056
rect 27730 870 27838 1056
rect 28006 870 28114 1056
rect 28282 870 28390 1056
rect 28558 870 28666 1056
rect 28834 870 28942 1056
rect 29110 870 29218 1056
rect 29386 870 29494 1056
rect 29662 870 29770 1056
rect 29938 870 30046 1056
rect 30214 870 30322 1056
rect 30490 870 30598 1056
rect 30766 870 30874 1056
rect 31042 870 31150 1056
rect 31318 870 31426 1056
rect 31594 870 31702 1056
rect 31870 870 31978 1056
rect 32146 870 32254 1056
rect 32422 984 32998 1056
rect 33210 1056 38998 3912
rect 33210 984 38050 1056
rect 32422 870 38050 984
rect 38218 870 38326 1056
rect 38494 870 38602 1056
rect 38770 870 38878 1056
rect 39210 1056 44998 3912
rect 39046 870 39154 984
rect 39322 870 39430 1056
rect 39598 870 39706 1056
rect 39874 870 39982 1056
rect 40150 870 40258 1056
rect 40426 870 40534 1056
rect 40702 870 40810 1056
rect 40978 870 41086 1056
rect 41254 870 41362 1056
rect 41530 870 41638 1056
rect 41806 870 41914 1056
rect 42082 870 42190 1056
rect 42358 870 42466 1056
rect 42634 870 42742 1056
rect 42910 870 43018 1056
rect 43186 870 43294 1056
rect 43462 870 43570 1056
rect 43738 870 43846 1056
rect 44014 870 44122 1056
rect 44290 870 44398 1056
rect 44566 870 44674 1056
rect 44842 870 44950 1056
rect 45210 1056 50998 3912
rect 45210 984 45226 1056
rect 45118 870 45226 984
rect 45394 870 45502 1056
rect 45670 870 45778 1056
rect 45946 870 46054 1056
rect 46222 870 46330 1056
rect 46498 870 46606 1056
rect 46774 870 46882 1056
rect 47050 870 47158 1056
rect 47326 870 47434 1056
rect 47602 870 47710 1056
rect 47878 870 47986 1056
rect 48154 870 48262 1056
rect 48430 870 48538 1056
rect 48706 870 48814 1056
rect 48982 870 49090 1056
rect 49258 870 49366 1056
rect 49534 870 49642 1056
rect 49810 870 49918 1056
rect 50086 870 50194 1056
rect 50362 870 50470 1056
rect 50638 870 50746 1056
rect 50914 984 50998 1056
rect 51210 1056 56998 3912
rect 50914 870 51022 984
rect 51210 984 51298 1056
rect 51190 870 51298 984
rect 51466 870 51574 1056
rect 51742 870 51850 1056
rect 52018 870 52126 1056
rect 52294 870 52402 1056
rect 52570 870 52678 1056
rect 52846 870 52954 1056
rect 53122 870 53230 1056
rect 53398 870 53506 1056
rect 53674 870 53782 1056
rect 53950 870 54058 1056
rect 54226 870 54334 1056
rect 54502 870 54610 1056
rect 54778 870 54886 1056
rect 55054 870 55162 1056
rect 55330 870 55438 1056
rect 55606 870 55714 1056
rect 55882 870 55990 1056
rect 56158 870 56266 1056
rect 56434 870 56542 1056
rect 56710 870 56818 1056
rect 56986 984 56998 1056
rect 57210 1056 62998 3912
rect 56986 870 57094 984
rect 57262 870 57370 1056
rect 57538 870 57646 1056
rect 57814 870 57922 1056
rect 58090 870 58198 1056
rect 58366 870 58474 1056
rect 58642 870 58750 1056
rect 58918 870 59026 1056
rect 59194 870 59302 1056
rect 59470 870 59578 1056
rect 59746 870 59854 1056
rect 60022 870 60130 1056
rect 60298 870 60406 1056
rect 60574 870 60682 1056
rect 60850 870 60958 1056
rect 61126 870 61234 1056
rect 61402 870 61510 1056
rect 61678 870 61786 1056
rect 61954 870 62062 1056
rect 62230 870 62338 1056
rect 62506 870 62614 1056
rect 62782 870 62890 1056
rect 63210 1056 68998 3912
rect 63058 870 63166 984
rect 63334 870 63442 1056
rect 63610 870 63718 1056
rect 63886 870 63994 1056
rect 64162 870 64270 1056
rect 64438 870 64546 1056
rect 64714 870 64822 1056
rect 64990 870 65098 1056
rect 65266 870 65374 1056
rect 65542 870 65650 1056
rect 65818 870 65926 1056
rect 66094 870 66202 1056
rect 66370 870 66478 1056
rect 66646 870 66754 1056
rect 66922 870 67030 1056
rect 67198 870 67306 1056
rect 67474 870 67582 1056
rect 67750 870 67858 1056
rect 68026 870 68134 1056
rect 68302 870 68410 1056
rect 68578 870 68686 1056
rect 68854 870 68962 1056
rect 69210 1056 69900 3912
rect 69210 984 69238 1056
rect 69130 870 69238 984
rect 69406 870 69514 1056
rect 69682 870 69790 1056
<< metal3 >>
rect 0 3680 1000 3800
rect 0 3272 1000 3392
rect 1104 3350 72864 3450
rect 0 2864 1000 2984
rect 0 2456 1000 2576
rect 1104 2270 72864 2370
rect 0 2048 1000 2168
rect 0 1640 1000 1760
rect 0 1232 1000 1352
rect 1104 1190 72864 1290
<< obsm3 >>
rect 1080 3600 28599 3773
rect 982 3530 28599 3600
rect 982 3472 1024 3530
rect 1080 3192 28599 3270
rect 982 3064 28599 3192
rect 1080 2784 28599 3064
rect 982 2656 28599 2784
rect 1080 2450 28599 2656
rect 982 2248 1024 2376
rect 1080 1968 28599 2190
rect 982 1840 28599 1968
rect 1080 1560 28599 1840
rect 982 1432 28599 1560
rect 1080 1370 28599 1432
<< labels >>
rlabel metal2 s 32310 0 32366 1000 6 HI[0]
port 1 nsew signal output
rlabel metal2 s 20994 0 21050 1000 6 HI[100]
port 2 nsew signal output
rlabel metal2 s 30378 0 30434 1000 6 HI[101]
port 3 nsew signal output
rlabel metal2 s 10230 0 10286 1000 6 HI[102]
port 4 nsew signal output
rlabel metal2 s 846 0 902 1000 6 HI[103]
port 5 nsew signal output
rlabel metal2 s 26238 0 26294 1000 6 HI[104]
port 6 nsew signal output
rlabel metal2 s 32034 0 32090 1000 6 HI[105]
port 7 nsew signal output
rlabel metal2 s 8298 0 8354 1000 6 HI[106]
port 8 nsew signal output
rlabel metal2 s 31758 0 31814 1000 6 HI[107]
port 9 nsew signal output
rlabel metal2 s 26514 0 26570 1000 6 HI[108]
port 10 nsew signal output
rlabel metal2 s 9954 0 10010 1000 6 HI[109]
port 11 nsew signal output
rlabel metal2 s 17406 0 17462 1000 6 HI[10]
port 12 nsew signal output
rlabel metal2 s 5814 0 5870 1000 6 HI[110]
port 13 nsew signal output
rlabel metal2 s 26790 0 26846 1000 6 HI[111]
port 14 nsew signal output
rlabel metal2 s 17682 0 17738 1000 6 HI[112]
port 15 nsew signal output
rlabel metal2 s 27618 0 27674 1000 6 HI[113]
port 16 nsew signal output
rlabel metal2 s 1122 0 1178 1000 6 HI[114]
port 17 nsew signal output
rlabel metal2 s 27066 0 27122 1000 6 HI[115]
port 18 nsew signal output
rlabel metal2 s 14646 0 14702 1000 6 HI[116]
port 19 nsew signal output
rlabel metal2 s 5262 0 5318 1000 6 HI[117]
port 20 nsew signal output
rlabel metal2 s 18234 0 18290 1000 6 HI[118]
port 21 nsew signal output
rlabel metal2 s 11886 0 11942 1000 6 HI[119]
port 22 nsew signal output
rlabel metal2 s 27342 0 27398 1000 6 HI[11]
port 23 nsew signal output
rlabel metal2 s 18510 0 18566 1000 6 HI[120]
port 24 nsew signal output
rlabel metal2 s 1674 0 1730 1000 6 HI[121]
port 25 nsew signal output
rlabel metal2 s 11334 0 11390 1000 6 HI[122]
port 26 nsew signal output
rlabel metal2 s 30654 0 30710 1000 6 HI[123]
port 27 nsew signal output
rlabel metal2 s 12438 0 12494 1000 6 HI[124]
port 28 nsew signal output
rlabel metal2 s 6918 0 6974 1000 6 HI[125]
port 29 nsew signal output
rlabel metal2 s 19062 0 19118 1000 6 HI[126]
port 30 nsew signal output
rlabel metal2 s 27894 0 27950 1000 6 HI[127]
port 31 nsew signal output
rlabel metal2 s 15474 0 15530 1000 6 HI[128]
port 32 nsew signal output
rlabel metal2 s 19338 0 19394 1000 6 HI[129]
port 33 nsew signal output
rlabel metal2 s 17958 0 18014 1000 6 HI[12]
port 34 nsew signal output
rlabel metal2 s 28170 0 28226 1000 6 HI[130]
port 35 nsew signal output
rlabel metal2 s 19614 0 19670 1000 6 HI[131]
port 36 nsew signal output
rlabel metal2 s 4710 0 4766 1000 6 HI[132]
port 37 nsew signal output
rlabel metal2 s 10782 0 10838 1000 6 HI[133]
port 38 nsew signal output
rlabel metal2 s 28446 0 28502 1000 6 HI[134]
port 39 nsew signal output
rlabel metal2 s 13542 0 13598 1000 6 HI[135]
port 40 nsew signal output
rlabel metal2 s 30930 0 30986 1000 6 HI[136]
port 41 nsew signal output
rlabel metal2 s 20442 0 20498 1000 6 HI[137]
port 42 nsew signal output
rlabel metal2 s 7194 0 7250 1000 6 HI[138]
port 43 nsew signal output
rlabel metal2 s 6366 0 6422 1000 6 HI[139]
port 44 nsew signal output
rlabel metal2 s 21270 0 21326 1000 6 HI[13]
port 45 nsew signal output
rlabel metal2 s 28722 0 28778 1000 6 HI[140]
port 46 nsew signal output
rlabel metal2 s 3606 0 3662 1000 6 HI[141]
port 47 nsew signal output
rlabel metal2 s 20718 0 20774 1000 6 HI[142]
port 48 nsew signal output
rlabel metal2 s 4434 0 4490 1000 6 HI[143]
port 49 nsew signal output
rlabel metal2 s 28998 0 29054 1000 6 HI[144]
port 50 nsew signal output
rlabel metal2 s 31206 0 31262 1000 6 HI[145]
port 51 nsew signal output
rlabel metal2 s 18786 0 18842 1000 6 HI[146]
port 52 nsew signal output
rlabel metal2 s 16578 0 16634 1000 6 HI[147]
port 53 nsew signal output
rlabel metal2 s 23202 0 23258 1000 6 HI[148]
port 54 nsew signal output
rlabel metal2 s 17130 0 17186 1000 6 HI[149]
port 55 nsew signal output
rlabel metal2 s 8022 0 8078 1000 6 HI[14]
port 56 nsew signal output
rlabel metal2 s 21546 0 21602 1000 6 HI[150]
port 57 nsew signal output
rlabel metal2 s 15198 0 15254 1000 6 HI[151]
port 58 nsew signal output
rlabel metal2 s 7470 0 7526 1000 6 HI[152]
port 59 nsew signal output
rlabel metal2 s 21822 0 21878 1000 6 HI[153]
port 60 nsew signal output
rlabel metal2 s 12714 0 12770 1000 6 HI[154]
port 61 nsew signal output
rlabel metal2 s 8850 0 8906 1000 6 HI[155]
port 62 nsew signal output
rlabel metal2 s 22098 0 22154 1000 6 HI[156]
port 63 nsew signal output
rlabel metal2 s 9126 0 9182 1000 6 HI[157]
port 64 nsew signal output
rlabel metal2 s 1950 0 2006 1000 6 HI[158]
port 65 nsew signal output
rlabel metal2 s 22374 0 22430 1000 6 HI[159]
port 66 nsew signal output
rlabel metal2 s 2226 0 2282 1000 6 HI[15]
port 67 nsew signal output
rlabel metal2 s 9678 0 9734 1000 6 HI[160]
port 68 nsew signal output
rlabel metal2 s 22650 0 22706 1000 6 HI[161]
port 69 nsew signal output
rlabel metal2 s 16302 0 16358 1000 6 HI[162]
port 70 nsew signal output
rlabel metal2 s 3330 0 3386 1000 6 HI[163]
port 71 nsew signal output
rlabel metal2 s 22926 0 22982 1000 6 HI[164]
port 72 nsew signal output
rlabel metal2 s 4158 0 4214 1000 6 HI[165]
port 73 nsew signal output
rlabel metal2 s 10506 0 10562 1000 6 HI[166]
port 74 nsew signal output
rlabel metal2 s 3882 0 3938 1000 6 HI[167]
port 75 nsew signal output
rlabel metal2 s 29274 0 29330 1000 6 HI[168]
port 76 nsew signal output
rlabel metal2 s 16854 0 16910 1000 6 HI[169]
port 77 nsew signal output
rlabel metal2 s 11058 0 11114 1000 6 HI[16]
port 78 nsew signal output
rlabel metal2 s 13266 0 13322 1000 6 HI[170]
port 79 nsew signal output
rlabel metal2 s 23478 0 23534 1000 6 HI[171]
port 80 nsew signal output
rlabel metal2 s 6090 0 6146 1000 6 HI[172]
port 81 nsew signal output
rlabel metal2 s 11610 0 11666 1000 6 HI[173]
port 82 nsew signal output
rlabel metal2 s 570 0 626 1000 6 HI[174]
port 83 nsew signal output
rlabel metal2 s 23754 0 23810 1000 6 HI[175]
port 84 nsew signal output
rlabel metal2 s 4986 0 5042 1000 6 HI[176]
port 85 nsew signal output
rlabel metal2 s 12162 0 12218 1000 6 HI[177]
port 86 nsew signal output
rlabel metal2 s 14094 0 14150 1000 6 HI[178]
port 87 nsew signal output
rlabel metal2 s 24030 0 24086 1000 6 HI[179]
port 88 nsew signal output
rlabel metal2 s 7746 0 7802 1000 6 HI[17]
port 89 nsew signal output
rlabel metal2 s 29550 0 29606 1000 6 HI[180]
port 90 nsew signal output
rlabel metal2 s 2778 0 2834 1000 6 HI[181]
port 91 nsew signal output
rlabel metal2 s 24306 0 24362 1000 6 HI[182]
port 92 nsew signal output
rlabel metal2 s 2502 0 2558 1000 6 HI[183]
port 93 nsew signal output
rlabel metal2 s 16026 0 16082 1000 6 HI[184]
port 94 nsew signal output
rlabel metal2 s 31482 0 31538 1000 6 HI[185]
port 95 nsew signal output
rlabel metal2 s 24582 0 24638 1000 6 HI[186]
port 96 nsew signal output
rlabel metal2 s 6642 0 6698 1000 6 HI[187]
port 97 nsew signal output
rlabel metal2 s 13818 0 13874 1000 6 HI[188]
port 98 nsew signal output
rlabel metal2 s 8574 0 8630 1000 6 HI[189]
port 99 nsew signal output
rlabel metal2 s 24858 0 24914 1000 6 HI[18]
port 100 nsew signal output
rlabel metal2 s 29826 0 29882 1000 6 HI[190]
port 101 nsew signal output
rlabel metal2 s 14370 0 14426 1000 6 HI[191]
port 102 nsew signal output
rlabel metal2 s 5538 0 5594 1000 6 HI[192]
port 103 nsew signal output
rlabel metal2 s 25134 0 25190 1000 6 HI[193]
port 104 nsew signal output
rlabel metal2 s 20166 0 20222 1000 6 HI[194]
port 105 nsew signal output
rlabel metal2 s 14922 0 14978 1000 6 HI[195]
port 106 nsew signal output
rlabel metal2 s 1398 0 1454 1000 6 HI[196]
port 107 nsew signal output
rlabel metal2 s 25410 0 25466 1000 6 HI[197]
port 108 nsew signal output
rlabel metal2 s 9402 0 9458 1000 6 HI[198]
port 109 nsew signal output
rlabel metal2 s 30102 0 30158 1000 6 HI[199]
port 110 nsew signal output
rlabel metal2 s 3054 0 3110 1000 6 HI[19]
port 111 nsew signal output
rlabel metal2 s 15750 0 15806 1000 6 HI[1]
port 112 nsew signal output
rlabel metal2 s 25686 0 25742 1000 6 HI[200]
port 113 nsew signal output
rlabel metal2 s 19890 0 19946 1000 6 HI[201]
port 114 nsew signal output
rlabel metal2 s 12990 0 13046 1000 6 HI[202]
port 115 nsew signal output
rlabel metal2 s 25962 0 26018 1000 6 HI[203]
port 116 nsew signal output
rlabel metal2 s 30378 4000 30434 5000 6 HI[204]
port 117 nsew signal output
rlabel metal3 s 0 1232 1000 1352 6 HI[205]
port 118 nsew signal output
rlabel metal3 s 0 1640 1000 1760 6 HI[206]
port 119 nsew signal output
rlabel metal3 s 0 2048 1000 2168 6 HI[207]
port 120 nsew signal output
rlabel metal3 s 0 2456 1000 2576 6 HI[208]
port 121 nsew signal output
rlabel metal3 s 0 2864 1000 2984 6 HI[209]
port 122 nsew signal output
rlabel metal3 s 0 3272 1000 3392 6 HI[20]
port 123 nsew signal output
rlabel metal3 s 0 3680 1000 3800 6 HI[210]
port 124 nsew signal output
rlabel metal2 s 570 4000 626 5000 6 HI[211]
port 125 nsew signal output
rlabel metal2 s 846 4000 902 5000 6 HI[212]
port 126 nsew signal output
rlabel metal2 s 1122 4000 1178 5000 6 HI[213]
port 127 nsew signal output
rlabel metal2 s 1398 4000 1454 5000 6 HI[214]
port 128 nsew signal output
rlabel metal2 s 1674 4000 1730 5000 6 HI[215]
port 129 nsew signal output
rlabel metal2 s 1950 4000 2006 5000 6 HI[216]
port 130 nsew signal output
rlabel metal2 s 2226 4000 2282 5000 6 HI[217]
port 131 nsew signal output
rlabel metal2 s 2502 4000 2558 5000 6 HI[218]
port 132 nsew signal output
rlabel metal2 s 2778 4000 2834 5000 6 HI[219]
port 133 nsew signal output
rlabel metal2 s 3054 4000 3110 5000 6 HI[21]
port 134 nsew signal output
rlabel metal2 s 3330 4000 3386 5000 6 HI[220]
port 135 nsew signal output
rlabel metal2 s 3606 4000 3662 5000 6 HI[221]
port 136 nsew signal output
rlabel metal2 s 3882 4000 3938 5000 6 HI[222]
port 137 nsew signal output
rlabel metal2 s 4158 4000 4214 5000 6 HI[223]
port 138 nsew signal output
rlabel metal2 s 4434 4000 4490 5000 6 HI[224]
port 139 nsew signal output
rlabel metal2 s 4710 4000 4766 5000 6 HI[225]
port 140 nsew signal output
rlabel metal2 s 4986 4000 5042 5000 6 HI[226]
port 141 nsew signal output
rlabel metal2 s 5262 4000 5318 5000 6 HI[227]
port 142 nsew signal output
rlabel metal2 s 5538 4000 5594 5000 6 HI[228]
port 143 nsew signal output
rlabel metal2 s 5814 4000 5870 5000 6 HI[229]
port 144 nsew signal output
rlabel metal2 s 6090 4000 6146 5000 6 HI[22]
port 145 nsew signal output
rlabel metal2 s 6366 4000 6422 5000 6 HI[230]
port 146 nsew signal output
rlabel metal2 s 6642 4000 6698 5000 6 HI[231]
port 147 nsew signal output
rlabel metal2 s 6918 4000 6974 5000 6 HI[232]
port 148 nsew signal output
rlabel metal2 s 7194 4000 7250 5000 6 HI[233]
port 149 nsew signal output
rlabel metal2 s 7470 4000 7526 5000 6 HI[234]
port 150 nsew signal output
rlabel metal2 s 7746 4000 7802 5000 6 HI[235]
port 151 nsew signal output
rlabel metal2 s 8022 4000 8078 5000 6 HI[236]
port 152 nsew signal output
rlabel metal2 s 8298 4000 8354 5000 6 HI[237]
port 153 nsew signal output
rlabel metal2 s 8574 4000 8630 5000 6 HI[238]
port 154 nsew signal output
rlabel metal2 s 8850 4000 8906 5000 6 HI[239]
port 155 nsew signal output
rlabel metal2 s 9126 4000 9182 5000 6 HI[23]
port 156 nsew signal output
rlabel metal2 s 9402 4000 9458 5000 6 HI[240]
port 157 nsew signal output
rlabel metal2 s 9678 4000 9734 5000 6 HI[241]
port 158 nsew signal output
rlabel metal2 s 9954 4000 10010 5000 6 HI[242]
port 159 nsew signal output
rlabel metal2 s 10230 4000 10286 5000 6 HI[243]
port 160 nsew signal output
rlabel metal2 s 10506 4000 10562 5000 6 HI[244]
port 161 nsew signal output
rlabel metal2 s 10782 4000 10838 5000 6 HI[245]
port 162 nsew signal output
rlabel metal2 s 11058 4000 11114 5000 6 HI[246]
port 163 nsew signal output
rlabel metal2 s 11334 4000 11390 5000 6 HI[247]
port 164 nsew signal output
rlabel metal2 s 11610 4000 11666 5000 6 HI[248]
port 165 nsew signal output
rlabel metal2 s 11886 4000 11942 5000 6 HI[249]
port 166 nsew signal output
rlabel metal2 s 12162 4000 12218 5000 6 HI[24]
port 167 nsew signal output
rlabel metal2 s 12438 4000 12494 5000 6 HI[250]
port 168 nsew signal output
rlabel metal2 s 12714 4000 12770 5000 6 HI[251]
port 169 nsew signal output
rlabel metal2 s 12990 4000 13046 5000 6 HI[252]
port 170 nsew signal output
rlabel metal2 s 13266 4000 13322 5000 6 HI[253]
port 171 nsew signal output
rlabel metal2 s 13542 4000 13598 5000 6 HI[254]
port 172 nsew signal output
rlabel metal2 s 13818 4000 13874 5000 6 HI[255]
port 173 nsew signal output
rlabel metal2 s 14094 4000 14150 5000 6 HI[256]
port 174 nsew signal output
rlabel metal2 s 14370 4000 14426 5000 6 HI[257]
port 175 nsew signal output
rlabel metal2 s 14646 4000 14702 5000 6 HI[258]
port 176 nsew signal output
rlabel metal2 s 14922 4000 14978 5000 6 HI[259]
port 177 nsew signal output
rlabel metal2 s 15198 4000 15254 5000 6 HI[25]
port 178 nsew signal output
rlabel metal2 s 15474 4000 15530 5000 6 HI[260]
port 179 nsew signal output
rlabel metal2 s 15750 4000 15806 5000 6 HI[261]
port 180 nsew signal output
rlabel metal2 s 16026 4000 16082 5000 6 HI[262]
port 181 nsew signal output
rlabel metal2 s 16302 4000 16358 5000 6 HI[263]
port 182 nsew signal output
rlabel metal2 s 16578 4000 16634 5000 6 HI[264]
port 183 nsew signal output
rlabel metal2 s 16854 4000 16910 5000 6 HI[265]
port 184 nsew signal output
rlabel metal2 s 17130 4000 17186 5000 6 HI[266]
port 185 nsew signal output
rlabel metal2 s 17406 4000 17462 5000 6 HI[267]
port 186 nsew signal output
rlabel metal2 s 17682 4000 17738 5000 6 HI[268]
port 187 nsew signal output
rlabel metal2 s 17958 4000 18014 5000 6 HI[269]
port 188 nsew signal output
rlabel metal2 s 18234 4000 18290 5000 6 HI[26]
port 189 nsew signal output
rlabel metal2 s 18510 4000 18566 5000 6 HI[270]
port 190 nsew signal output
rlabel metal2 s 18786 4000 18842 5000 6 HI[271]
port 191 nsew signal output
rlabel metal2 s 19062 4000 19118 5000 6 HI[272]
port 192 nsew signal output
rlabel metal2 s 19338 4000 19394 5000 6 HI[273]
port 193 nsew signal output
rlabel metal2 s 19614 4000 19670 5000 6 HI[274]
port 194 nsew signal output
rlabel metal2 s 19890 4000 19946 5000 6 HI[275]
port 195 nsew signal output
rlabel metal2 s 20166 4000 20222 5000 6 HI[276]
port 196 nsew signal output
rlabel metal2 s 20442 4000 20498 5000 6 HI[277]
port 197 nsew signal output
rlabel metal2 s 20718 4000 20774 5000 6 HI[278]
port 198 nsew signal output
rlabel metal2 s 20994 4000 21050 5000 6 HI[279]
port 199 nsew signal output
rlabel metal2 s 21270 4000 21326 5000 6 HI[27]
port 200 nsew signal output
rlabel metal2 s 21546 4000 21602 5000 6 HI[280]
port 201 nsew signal output
rlabel metal2 s 21822 4000 21878 5000 6 HI[281]
port 202 nsew signal output
rlabel metal2 s 22098 4000 22154 5000 6 HI[282]
port 203 nsew signal output
rlabel metal2 s 22374 4000 22430 5000 6 HI[283]
port 204 nsew signal output
rlabel metal2 s 22650 4000 22706 5000 6 HI[284]
port 205 nsew signal output
rlabel metal2 s 22926 4000 22982 5000 6 HI[285]
port 206 nsew signal output
rlabel metal2 s 23202 4000 23258 5000 6 HI[286]
port 207 nsew signal output
rlabel metal2 s 23478 4000 23534 5000 6 HI[287]
port 208 nsew signal output
rlabel metal2 s 23754 4000 23810 5000 6 HI[288]
port 209 nsew signal output
rlabel metal2 s 24030 4000 24086 5000 6 HI[289]
port 210 nsew signal output
rlabel metal2 s 24306 4000 24362 5000 6 HI[28]
port 211 nsew signal output
rlabel metal2 s 24582 4000 24638 5000 6 HI[290]
port 212 nsew signal output
rlabel metal2 s 24858 4000 24914 5000 6 HI[291]
port 213 nsew signal output
rlabel metal2 s 25134 4000 25190 5000 6 HI[292]
port 214 nsew signal output
rlabel metal2 s 25410 4000 25466 5000 6 HI[293]
port 215 nsew signal output
rlabel metal2 s 25686 4000 25742 5000 6 HI[294]
port 216 nsew signal output
rlabel metal2 s 25962 4000 26018 5000 6 HI[295]
port 217 nsew signal output
rlabel metal2 s 26238 4000 26294 5000 6 HI[296]
port 218 nsew signal output
rlabel metal2 s 26514 4000 26570 5000 6 HI[297]
port 219 nsew signal output
rlabel metal2 s 26790 4000 26846 5000 6 HI[298]
port 220 nsew signal output
rlabel metal2 s 27066 4000 27122 5000 6 HI[299]
port 221 nsew signal output
rlabel metal2 s 27342 4000 27398 5000 6 HI[29]
port 222 nsew signal output
rlabel metal2 s 27618 4000 27674 5000 6 HI[2]
port 223 nsew signal output
rlabel metal2 s 27894 4000 27950 5000 6 HI[300]
port 224 nsew signal output
rlabel metal2 s 28170 4000 28226 5000 6 HI[301]
port 225 nsew signal output
rlabel metal2 s 28446 4000 28502 5000 6 HI[302]
port 226 nsew signal output
rlabel metal2 s 28722 4000 28778 5000 6 HI[303]
port 227 nsew signal output
rlabel metal2 s 28998 4000 29054 5000 6 HI[304]
port 228 nsew signal output
rlabel metal2 s 29274 4000 29330 5000 6 HI[305]
port 229 nsew signal output
rlabel metal2 s 29550 4000 29606 5000 6 HI[306]
port 230 nsew signal output
rlabel metal2 s 29826 4000 29882 5000 6 HI[307]
port 231 nsew signal output
rlabel metal2 s 30102 4000 30158 5000 6 HI[308]
port 232 nsew signal output
rlabel metal2 s 69846 0 69902 1000 6 HI[309]
port 233 nsew signal output
rlabel metal2 s 58530 0 58586 1000 6 HI[30]
port 234 nsew signal output
rlabel metal2 s 67914 0 67970 1000 6 HI[310]
port 235 nsew signal output
rlabel metal2 s 47766 0 47822 1000 6 HI[311]
port 236 nsew signal output
rlabel metal2 s 38382 0 38438 1000 6 HI[312]
port 237 nsew signal output
rlabel metal2 s 63774 0 63830 1000 6 HI[313]
port 238 nsew signal output
rlabel metal2 s 69570 0 69626 1000 6 HI[314]
port 239 nsew signal output
rlabel metal2 s 45834 0 45890 1000 6 HI[315]
port 240 nsew signal output
rlabel metal2 s 69294 0 69350 1000 6 HI[316]
port 241 nsew signal output
rlabel metal2 s 64050 0 64106 1000 6 HI[317]
port 242 nsew signal output
rlabel metal2 s 47490 0 47546 1000 6 HI[318]
port 243 nsew signal output
rlabel metal2 s 54942 0 54998 1000 6 HI[319]
port 244 nsew signal output
rlabel metal2 s 43350 0 43406 1000 6 HI[31]
port 245 nsew signal output
rlabel metal2 s 64326 0 64382 1000 6 HI[320]
port 246 nsew signal output
rlabel metal2 s 55218 0 55274 1000 6 HI[321]
port 247 nsew signal output
rlabel metal2 s 65154 0 65210 1000 6 HI[322]
port 248 nsew signal output
rlabel metal2 s 38658 0 38714 1000 6 HI[323]
port 249 nsew signal output
rlabel metal2 s 64602 0 64658 1000 6 HI[324]
port 250 nsew signal output
rlabel metal2 s 52182 0 52238 1000 6 HI[325]
port 251 nsew signal output
rlabel metal2 s 42798 0 42854 1000 6 HI[326]
port 252 nsew signal output
rlabel metal2 s 55770 0 55826 1000 6 HI[327]
port 253 nsew signal output
rlabel metal2 s 49422 0 49478 1000 6 HI[328]
port 254 nsew signal output
rlabel metal2 s 64878 0 64934 1000 6 HI[329]
port 255 nsew signal output
rlabel metal2 s 56046 0 56102 1000 6 HI[32]
port 256 nsew signal output
rlabel metal2 s 39210 0 39266 1000 6 HI[330]
port 257 nsew signal output
rlabel metal2 s 48870 0 48926 1000 6 HI[331]
port 258 nsew signal output
rlabel metal2 s 68190 0 68246 1000 6 HI[332]
port 259 nsew signal output
rlabel metal2 s 49974 0 50030 1000 6 HI[333]
port 260 nsew signal output
rlabel metal2 s 44454 0 44510 1000 6 HI[334]
port 261 nsew signal output
rlabel metal2 s 56598 0 56654 1000 6 HI[335]
port 262 nsew signal output
rlabel metal2 s 65430 0 65486 1000 6 HI[336]
port 263 nsew signal output
rlabel metal2 s 53010 0 53066 1000 6 HI[337]
port 264 nsew signal output
rlabel metal2 s 56874 0 56930 1000 6 HI[338]
port 265 nsew signal output
rlabel metal2 s 55494 0 55550 1000 6 HI[339]
port 266 nsew signal output
rlabel metal2 s 65706 0 65762 1000 6 HI[33]
port 267 nsew signal output
rlabel metal2 s 57150 0 57206 1000 6 HI[340]
port 268 nsew signal output
rlabel metal2 s 42246 0 42302 1000 6 HI[341]
port 269 nsew signal output
rlabel metal2 s 48318 0 48374 1000 6 HI[342]
port 270 nsew signal output
rlabel metal2 s 65982 0 66038 1000 6 HI[343]
port 271 nsew signal output
rlabel metal2 s 51078 0 51134 1000 6 HI[344]
port 272 nsew signal output
rlabel metal2 s 68466 0 68522 1000 6 HI[345]
port 273 nsew signal output
rlabel metal2 s 57978 0 58034 1000 6 HI[346]
port 274 nsew signal output
rlabel metal2 s 44730 0 44786 1000 6 HI[347]
port 275 nsew signal output
rlabel metal2 s 43902 0 43958 1000 6 HI[348]
port 276 nsew signal output
rlabel metal2 s 58806 0 58862 1000 6 HI[349]
port 277 nsew signal output
rlabel metal2 s 66258 0 66314 1000 6 HI[34]
port 278 nsew signal output
rlabel metal2 s 41142 0 41198 1000 6 HI[350]
port 279 nsew signal output
rlabel metal2 s 58254 0 58310 1000 6 HI[351]
port 280 nsew signal output
rlabel metal2 s 41970 0 42026 1000 6 HI[352]
port 281 nsew signal output
rlabel metal2 s 66534 0 66590 1000 6 HI[353]
port 282 nsew signal output
rlabel metal2 s 68742 0 68798 1000 6 HI[354]
port 283 nsew signal output
rlabel metal2 s 56322 0 56378 1000 6 HI[355]
port 284 nsew signal output
rlabel metal2 s 54114 0 54170 1000 6 HI[356]
port 285 nsew signal output
rlabel metal2 s 60738 0 60794 1000 6 HI[357]
port 286 nsew signal output
rlabel metal2 s 54666 0 54722 1000 6 HI[358]
port 287 nsew signal output
rlabel metal2 s 45558 0 45614 1000 6 HI[359]
port 288 nsew signal output
rlabel metal2 s 59082 0 59138 1000 6 HI[35]
port 289 nsew signal output
rlabel metal2 s 52734 0 52790 1000 6 HI[360]
port 290 nsew signal output
rlabel metal2 s 45006 0 45062 1000 6 HI[361]
port 291 nsew signal output
rlabel metal2 s 59358 0 59414 1000 6 HI[362]
port 292 nsew signal output
rlabel metal2 s 50250 0 50306 1000 6 HI[363]
port 293 nsew signal output
rlabel metal2 s 46386 0 46442 1000 6 HI[364]
port 294 nsew signal output
rlabel metal2 s 59634 0 59690 1000 6 HI[365]
port 295 nsew signal output
rlabel metal2 s 46662 0 46718 1000 6 HI[366]
port 296 nsew signal output
rlabel metal2 s 39486 0 39542 1000 6 HI[367]
port 297 nsew signal output
rlabel metal2 s 59910 0 59966 1000 6 HI[368]
port 298 nsew signal output
rlabel metal2 s 39762 0 39818 1000 6 HI[369]
port 299 nsew signal output
rlabel metal2 s 47214 0 47270 1000 6 HI[36]
port 300 nsew signal output
rlabel metal2 s 60186 0 60242 1000 6 HI[370]
port 301 nsew signal output
rlabel metal2 s 53838 0 53894 1000 6 HI[371]
port 302 nsew signal output
rlabel metal2 s 40866 0 40922 1000 6 HI[372]
port 303 nsew signal output
rlabel metal2 s 60462 0 60518 1000 6 HI[373]
port 304 nsew signal output
rlabel metal2 s 41694 0 41750 1000 6 HI[374]
port 305 nsew signal output
rlabel metal2 s 48042 0 48098 1000 6 HI[375]
port 306 nsew signal output
rlabel metal2 s 41418 0 41474 1000 6 HI[376]
port 307 nsew signal output
rlabel metal2 s 66810 0 66866 1000 6 HI[377]
port 308 nsew signal output
rlabel metal2 s 54390 0 54446 1000 6 HI[378]
port 309 nsew signal output
rlabel metal2 s 48594 0 48650 1000 6 HI[379]
port 310 nsew signal output
rlabel metal2 s 50802 0 50858 1000 6 HI[37]
port 311 nsew signal output
rlabel metal2 s 61014 0 61070 1000 6 HI[380]
port 312 nsew signal output
rlabel metal2 s 43626 0 43682 1000 6 HI[381]
port 313 nsew signal output
rlabel metal2 s 49146 0 49202 1000 6 HI[382]
port 314 nsew signal output
rlabel metal2 s 38106 0 38162 1000 6 HI[383]
port 315 nsew signal output
rlabel metal2 s 61290 0 61346 1000 6 HI[384]
port 316 nsew signal output
rlabel metal2 s 42522 0 42578 1000 6 HI[385]
port 317 nsew signal output
rlabel metal2 s 49698 0 49754 1000 6 HI[386]
port 318 nsew signal output
rlabel metal2 s 51630 0 51686 1000 6 HI[387]
port 319 nsew signal output
rlabel metal2 s 61566 0 61622 1000 6 HI[388]
port 320 nsew signal output
rlabel metal2 s 45282 0 45338 1000 6 HI[389]
port 321 nsew signal output
rlabel metal2 s 67086 0 67142 1000 6 HI[38]
port 322 nsew signal output
rlabel metal2 s 40314 0 40370 1000 6 HI[390]
port 323 nsew signal output
rlabel metal2 s 61842 0 61898 1000 6 HI[391]
port 324 nsew signal output
rlabel metal2 s 40038 0 40094 1000 6 HI[392]
port 325 nsew signal output
rlabel metal2 s 53562 0 53618 1000 6 HI[393]
port 326 nsew signal output
rlabel metal2 s 69018 0 69074 1000 6 HI[394]
port 327 nsew signal output
rlabel metal2 s 62118 0 62174 1000 6 HI[395]
port 328 nsew signal output
rlabel metal2 s 44178 0 44234 1000 6 HI[396]
port 329 nsew signal output
rlabel metal2 s 51354 0 51410 1000 6 HI[397]
port 330 nsew signal output
rlabel metal2 s 46110 0 46166 1000 6 HI[398]
port 331 nsew signal output
rlabel metal2 s 62394 0 62450 1000 6 HI[399]
port 332 nsew signal output
rlabel metal2 s 67362 0 67418 1000 6 HI[39]
port 333 nsew signal output
rlabel metal2 s 51906 0 51962 1000 6 HI[3]
port 334 nsew signal output
rlabel metal2 s 43074 0 43130 1000 6 HI[400]
port 335 nsew signal output
rlabel metal2 s 62670 0 62726 1000 6 HI[401]
port 336 nsew signal output
rlabel metal2 s 57702 0 57758 1000 6 HI[402]
port 337 nsew signal output
rlabel metal2 s 52458 0 52514 1000 6 HI[403]
port 338 nsew signal output
rlabel metal2 s 38934 0 38990 1000 6 HI[404]
port 339 nsew signal output
rlabel metal2 s 62946 0 63002 1000 6 HI[405]
port 340 nsew signal output
rlabel metal2 s 46938 0 46994 1000 6 HI[406]
port 341 nsew signal output
rlabel metal2 s 67638 0 67694 1000 6 HI[407]
port 342 nsew signal output
rlabel metal2 s 40590 0 40646 1000 6 HI[408]
port 343 nsew signal output
rlabel metal2 s 53286 0 53342 1000 6 HI[409]
port 344 nsew signal output
rlabel metal2 s 63222 0 63278 1000 6 HI[40]
port 345 nsew signal output
rlabel metal2 s 57426 0 57482 1000 6 HI[410]
port 346 nsew signal output
rlabel metal2 s 50526 0 50582 1000 6 HI[411]
port 347 nsew signal output
rlabel metal2 s 63498 0 63554 1000 6 HI[412]
port 348 nsew signal output
rlabel metal2 s 67362 4000 67418 5000 6 HI[413]
port 349 nsew signal output
rlabel metal2 s 36174 4000 36230 5000 6 HI[414]
port 350 nsew signal output
rlabel metal2 s 36450 4000 36506 5000 6 HI[415]
port 351 nsew signal output
rlabel metal2 s 36726 4000 36782 5000 6 HI[416]
port 352 nsew signal output
rlabel metal2 s 37002 4000 37058 5000 6 HI[417]
port 353 nsew signal output
rlabel metal2 s 37278 4000 37334 5000 6 HI[418]
port 354 nsew signal output
rlabel metal2 s 37554 4000 37610 5000 6 HI[419]
port 355 nsew signal output
rlabel metal2 s 37830 4000 37886 5000 6 HI[41]
port 356 nsew signal output
rlabel metal2 s 38106 4000 38162 5000 6 HI[420]
port 357 nsew signal output
rlabel metal2 s 38382 4000 38438 5000 6 HI[421]
port 358 nsew signal output
rlabel metal2 s 38658 4000 38714 5000 6 HI[422]
port 359 nsew signal output
rlabel metal2 s 38934 4000 38990 5000 6 HI[423]
port 360 nsew signal output
rlabel metal2 s 39210 4000 39266 5000 6 HI[424]
port 361 nsew signal output
rlabel metal2 s 39486 4000 39542 5000 6 HI[425]
port 362 nsew signal output
rlabel metal2 s 39762 4000 39818 5000 6 HI[426]
port 363 nsew signal output
rlabel metal2 s 40038 4000 40094 5000 6 HI[427]
port 364 nsew signal output
rlabel metal2 s 40314 4000 40370 5000 6 HI[428]
port 365 nsew signal output
rlabel metal2 s 40590 4000 40646 5000 6 HI[429]
port 366 nsew signal output
rlabel metal2 s 40866 4000 40922 5000 6 HI[42]
port 367 nsew signal output
rlabel metal2 s 41142 4000 41198 5000 6 HI[430]
port 368 nsew signal output
rlabel metal2 s 41418 4000 41474 5000 6 HI[431]
port 369 nsew signal output
rlabel metal2 s 41694 4000 41750 5000 6 HI[432]
port 370 nsew signal output
rlabel metal2 s 41970 4000 42026 5000 6 HI[433]
port 371 nsew signal output
rlabel metal2 s 42246 4000 42302 5000 6 HI[434]
port 372 nsew signal output
rlabel metal2 s 42522 4000 42578 5000 6 HI[435]
port 373 nsew signal output
rlabel metal2 s 42798 4000 42854 5000 6 HI[436]
port 374 nsew signal output
rlabel metal2 s 43074 4000 43130 5000 6 HI[437]
port 375 nsew signal output
rlabel metal2 s 43350 4000 43406 5000 6 HI[438]
port 376 nsew signal output
rlabel metal2 s 43626 4000 43682 5000 6 HI[439]
port 377 nsew signal output
rlabel metal2 s 43902 4000 43958 5000 6 HI[43]
port 378 nsew signal output
rlabel metal2 s 44178 4000 44234 5000 6 HI[440]
port 379 nsew signal output
rlabel metal2 s 44454 4000 44510 5000 6 HI[441]
port 380 nsew signal output
rlabel metal2 s 44730 4000 44786 5000 6 HI[442]
port 381 nsew signal output
rlabel metal2 s 45006 4000 45062 5000 6 HI[443]
port 382 nsew signal output
rlabel metal2 s 45282 4000 45338 5000 6 HI[444]
port 383 nsew signal output
rlabel metal2 s 45558 4000 45614 5000 6 HI[445]
port 384 nsew signal output
rlabel metal2 s 45834 4000 45890 5000 6 HI[446]
port 385 nsew signal output
rlabel metal2 s 46110 4000 46166 5000 6 HI[447]
port 386 nsew signal output
rlabel metal2 s 46386 4000 46442 5000 6 HI[448]
port 387 nsew signal output
rlabel metal2 s 46662 4000 46718 5000 6 HI[449]
port 388 nsew signal output
rlabel metal2 s 46938 4000 46994 5000 6 HI[44]
port 389 nsew signal output
rlabel metal2 s 47214 4000 47270 5000 6 HI[450]
port 390 nsew signal output
rlabel metal2 s 47490 4000 47546 5000 6 HI[451]
port 391 nsew signal output
rlabel metal2 s 47766 4000 47822 5000 6 HI[452]
port 392 nsew signal output
rlabel metal2 s 48042 4000 48098 5000 6 HI[453]
port 393 nsew signal output
rlabel metal2 s 48318 4000 48374 5000 6 HI[454]
port 394 nsew signal output
rlabel metal2 s 48594 4000 48650 5000 6 HI[455]
port 395 nsew signal output
rlabel metal2 s 48870 4000 48926 5000 6 HI[456]
port 396 nsew signal output
rlabel metal2 s 49146 4000 49202 5000 6 HI[457]
port 397 nsew signal output
rlabel metal2 s 49422 4000 49478 5000 6 HI[458]
port 398 nsew signal output
rlabel metal2 s 49698 4000 49754 5000 6 HI[459]
port 399 nsew signal output
rlabel metal2 s 49974 4000 50030 5000 6 HI[45]
port 400 nsew signal output
rlabel metal2 s 50250 4000 50306 5000 6 HI[460]
port 401 nsew signal output
rlabel metal2 s 50526 4000 50582 5000 6 HI[461]
port 402 nsew signal output
rlabel metal2 s 50802 4000 50858 5000 6 HI[46]
port 403 nsew signal output
rlabel metal2 s 51078 4000 51134 5000 6 HI[47]
port 404 nsew signal output
rlabel metal2 s 51354 4000 51410 5000 6 HI[48]
port 405 nsew signal output
rlabel metal2 s 51630 4000 51686 5000 6 HI[49]
port 406 nsew signal output
rlabel metal2 s 51906 4000 51962 5000 6 HI[4]
port 407 nsew signal output
rlabel metal2 s 52182 4000 52238 5000 6 HI[50]
port 408 nsew signal output
rlabel metal2 s 52458 4000 52514 5000 6 HI[51]
port 409 nsew signal output
rlabel metal2 s 52734 4000 52790 5000 6 HI[52]
port 410 nsew signal output
rlabel metal2 s 53010 4000 53066 5000 6 HI[53]
port 411 nsew signal output
rlabel metal2 s 53286 4000 53342 5000 6 HI[54]
port 412 nsew signal output
rlabel metal2 s 53562 4000 53618 5000 6 HI[55]
port 413 nsew signal output
rlabel metal2 s 53838 4000 53894 5000 6 HI[56]
port 414 nsew signal output
rlabel metal2 s 54114 4000 54170 5000 6 HI[57]
port 415 nsew signal output
rlabel metal2 s 54390 4000 54446 5000 6 HI[58]
port 416 nsew signal output
rlabel metal2 s 54666 4000 54722 5000 6 HI[59]
port 417 nsew signal output
rlabel metal2 s 54942 4000 54998 5000 6 HI[5]
port 418 nsew signal output
rlabel metal2 s 55218 4000 55274 5000 6 HI[60]
port 419 nsew signal output
rlabel metal2 s 55494 4000 55550 5000 6 HI[61]
port 420 nsew signal output
rlabel metal2 s 55770 4000 55826 5000 6 HI[62]
port 421 nsew signal output
rlabel metal2 s 56046 4000 56102 5000 6 HI[63]
port 422 nsew signal output
rlabel metal2 s 56322 4000 56378 5000 6 HI[64]
port 423 nsew signal output
rlabel metal2 s 56598 4000 56654 5000 6 HI[65]
port 424 nsew signal output
rlabel metal2 s 56874 4000 56930 5000 6 HI[66]
port 425 nsew signal output
rlabel metal2 s 57150 4000 57206 5000 6 HI[67]
port 426 nsew signal output
rlabel metal2 s 57426 4000 57482 5000 6 HI[68]
port 427 nsew signal output
rlabel metal2 s 57702 4000 57758 5000 6 HI[69]
port 428 nsew signal output
rlabel metal2 s 57978 4000 58034 5000 6 HI[6]
port 429 nsew signal output
rlabel metal2 s 58254 4000 58310 5000 6 HI[70]
port 430 nsew signal output
rlabel metal2 s 58530 4000 58586 5000 6 HI[71]
port 431 nsew signal output
rlabel metal2 s 58806 4000 58862 5000 6 HI[72]
port 432 nsew signal output
rlabel metal2 s 59082 4000 59138 5000 6 HI[73]
port 433 nsew signal output
rlabel metal2 s 59358 4000 59414 5000 6 HI[74]
port 434 nsew signal output
rlabel metal2 s 59634 4000 59690 5000 6 HI[75]
port 435 nsew signal output
rlabel metal2 s 59910 4000 59966 5000 6 HI[76]
port 436 nsew signal output
rlabel metal2 s 60186 4000 60242 5000 6 HI[77]
port 437 nsew signal output
rlabel metal2 s 60462 4000 60518 5000 6 HI[78]
port 438 nsew signal output
rlabel metal2 s 60738 4000 60794 5000 6 HI[79]
port 439 nsew signal output
rlabel metal2 s 61014 4000 61070 5000 6 HI[7]
port 440 nsew signal output
rlabel metal2 s 61290 4000 61346 5000 6 HI[80]
port 441 nsew signal output
rlabel metal2 s 61566 4000 61622 5000 6 HI[81]
port 442 nsew signal output
rlabel metal2 s 61842 4000 61898 5000 6 HI[82]
port 443 nsew signal output
rlabel metal2 s 62118 4000 62174 5000 6 HI[83]
port 444 nsew signal output
rlabel metal2 s 62394 4000 62450 5000 6 HI[84]
port 445 nsew signal output
rlabel metal2 s 62670 4000 62726 5000 6 HI[85]
port 446 nsew signal output
rlabel metal2 s 62946 4000 63002 5000 6 HI[86]
port 447 nsew signal output
rlabel metal2 s 63222 4000 63278 5000 6 HI[87]
port 448 nsew signal output
rlabel metal2 s 63498 4000 63554 5000 6 HI[88]
port 449 nsew signal output
rlabel metal2 s 63774 4000 63830 5000 6 HI[89]
port 450 nsew signal output
rlabel metal2 s 64050 4000 64106 5000 6 HI[8]
port 451 nsew signal output
rlabel metal2 s 64326 4000 64382 5000 6 HI[90]
port 452 nsew signal output
rlabel metal2 s 64602 4000 64658 5000 6 HI[91]
port 453 nsew signal output
rlabel metal2 s 64878 4000 64934 5000 6 HI[92]
port 454 nsew signal output
rlabel metal2 s 65154 4000 65210 5000 6 HI[93]
port 455 nsew signal output
rlabel metal2 s 65430 4000 65486 5000 6 HI[94]
port 456 nsew signal output
rlabel metal2 s 65706 4000 65762 5000 6 HI[95]
port 457 nsew signal output
rlabel metal2 s 65982 4000 66038 5000 6 HI[96]
port 458 nsew signal output
rlabel metal2 s 66258 4000 66314 5000 6 HI[97]
port 459 nsew signal output
rlabel metal2 s 66534 4000 66590 5000 6 HI[98]
port 460 nsew signal output
rlabel metal2 s 66810 4000 66866 5000 6 HI[99]
port 461 nsew signal output
rlabel metal2 s 67086 4000 67142 5000 6 HI[9]
port 462 nsew signal output
rlabel metal2 s 63054 1040 63154 3856 6 vccd1
port 463 nsew power bidirectional
rlabel metal2 s 51054 1040 51154 3856 6 vccd1
port 464 nsew power bidirectional
rlabel metal2 s 39054 1040 39154 3856 6 vccd1
port 465 nsew power bidirectional
rlabel metal2 s 27054 1040 27154 3856 6 vccd1
port 466 nsew power bidirectional
rlabel metal2 s 15054 1040 15154 3856 6 vccd1
port 467 nsew power bidirectional
rlabel metal2 s 3054 1040 3154 3856 6 vccd1
port 468 nsew power bidirectional
rlabel metal3 s 1104 3350 72864 3450 6 vccd1
port 469 nsew power bidirectional
rlabel metal3 s 1104 1190 72864 1290 6 vccd1
port 470 nsew power bidirectional
rlabel metal2 s 69054 1040 69154 3856 6 vssd1
port 471 nsew ground bidirectional
rlabel metal2 s 57054 1040 57154 3856 6 vssd1
port 472 nsew ground bidirectional
rlabel metal2 s 45054 1040 45154 3856 6 vssd1
port 473 nsew ground bidirectional
rlabel metal2 s 33054 1040 33154 3856 6 vssd1
port 474 nsew ground bidirectional
rlabel metal2 s 21054 1040 21154 3856 6 vssd1
port 475 nsew ground bidirectional
rlabel metal2 s 9054 1040 9154 3856 6 vssd1
port 476 nsew ground bidirectional
rlabel metal3 s 1104 2270 72864 2370 6 vssd1
port 477 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 74000 5000
string LEFview TRUE
string GDS_FILE /project/openlane/mprj_logic_high/runs/mprj_logic_high/results/magic/mprj_logic_high.gds
string GDS_END 505678
string GDS_START 24116
<< end >>

