.subckt sky130_fd_pr__model__parasitic__diode_ps2nw A C a=1 p=1
D A C  sky130_fd_pr__model__parasitic__diode_ps2nw area={a}
.ends
