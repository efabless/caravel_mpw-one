magic
tech sky130A
magscale 12 1
timestamp 1598763107
<< metal5 >>
rect 10 100 35 105
rect 5 95 40 100
rect 0 85 45 95
rect 0 45 15 85
rect 30 45 45 85
rect 0 30 45 45
rect 0 0 15 30
rect 30 0 45 30
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
