magic
tech sky130A
magscale 1 2
timestamp 1606435979
<< error_s >>
rect 12547 2767 12605 2773
rect 12665 2767 12723 2773
rect 12783 2767 12841 2773
rect 12901 2767 12959 2773
rect 13019 2767 13077 2773
rect 13137 2767 13195 2773
rect 13255 2767 13313 2773
rect 13373 2767 13431 2773
rect 13491 2767 13549 2773
rect 13609 2767 13667 2773
rect 13727 2767 13785 2773
rect 13845 2767 13903 2773
rect 13963 2767 14021 2773
rect 14081 2767 14139 2773
rect 14199 2767 14257 2773
rect 14317 2767 14375 2773
rect 14435 2767 14493 2773
rect 14553 2767 14611 2773
rect 14671 2767 14729 2773
rect 14789 2767 14847 2773
rect 14907 2767 14965 2773
rect 15025 2767 15083 2773
rect 15143 2767 15201 2773
rect 15261 2767 15319 2773
rect 15379 2767 15437 2773
rect 15497 2767 15555 2773
rect 15615 2767 15673 2773
rect 15733 2767 15791 2773
rect 15851 2767 15909 2773
rect 15969 2767 16027 2773
rect 16087 2767 16145 2773
rect 16205 2767 16263 2773
rect 16323 2767 16381 2773
rect 16441 2767 16499 2773
rect 16559 2767 16617 2773
rect 16677 2767 16735 2773
rect 16795 2767 16853 2773
rect 16913 2767 16971 2773
rect 17031 2767 17089 2773
rect 17149 2767 17207 2773
rect 17267 2767 17325 2773
rect 17385 2767 17443 2773
rect 17503 2767 17561 2773
rect 17621 2767 17679 2773
rect 17739 2767 17797 2773
rect 17857 2767 17915 2773
rect 17975 2767 18033 2773
rect 18093 2767 18151 2773
rect 18211 2767 18269 2773
rect 18329 2767 18387 2773
rect 18447 2767 18505 2773
rect 18565 2767 18623 2773
rect 18683 2767 18741 2773
rect 18801 2767 18859 2773
rect 18919 2767 18977 2773
rect 19037 2767 19095 2773
rect 19155 2767 19213 2773
rect 19273 2767 19331 2773
rect 19391 2767 19449 2773
rect 19509 2767 19567 2773
rect 19627 2767 19685 2773
rect 19745 2767 19803 2773
rect 19863 2767 19921 2773
rect 19981 2767 20039 2773
rect 20099 2767 20157 2773
rect 20217 2767 20275 2773
rect 20335 2767 20393 2773
rect 20453 2767 20511 2773
rect 20571 2767 20629 2773
rect 20689 2767 20747 2773
rect 20807 2767 20865 2773
rect 20925 2767 20983 2773
rect 21043 2767 21101 2773
rect 21161 2767 21219 2773
rect 21279 2767 21337 2773
rect 12547 2733 12559 2767
rect 12665 2733 12677 2767
rect 12783 2733 12795 2767
rect 12901 2733 12913 2767
rect 13019 2733 13031 2767
rect 13137 2733 13149 2767
rect 13255 2733 13267 2767
rect 13373 2733 13385 2767
rect 13491 2733 13503 2767
rect 13609 2733 13621 2767
rect 13727 2733 13739 2767
rect 13845 2733 13857 2767
rect 13963 2733 13975 2767
rect 14081 2733 14093 2767
rect 14199 2733 14211 2767
rect 14317 2733 14329 2767
rect 14435 2733 14447 2767
rect 14553 2733 14565 2767
rect 14671 2733 14683 2767
rect 14789 2733 14801 2767
rect 14907 2733 14919 2767
rect 15025 2733 15037 2767
rect 15143 2733 15155 2767
rect 15261 2733 15273 2767
rect 15379 2733 15391 2767
rect 15497 2733 15509 2767
rect 15615 2733 15627 2767
rect 15733 2733 15745 2767
rect 15851 2733 15863 2767
rect 15969 2733 15981 2767
rect 16087 2733 16099 2767
rect 16205 2733 16217 2767
rect 16323 2733 16335 2767
rect 16441 2733 16453 2767
rect 16559 2733 16571 2767
rect 16677 2733 16689 2767
rect 16795 2733 16807 2767
rect 16913 2733 16925 2767
rect 17031 2733 17043 2767
rect 17149 2733 17161 2767
rect 17267 2733 17279 2767
rect 17385 2733 17397 2767
rect 17503 2733 17515 2767
rect 17621 2733 17633 2767
rect 17739 2733 17751 2767
rect 17857 2733 17869 2767
rect 17975 2733 17987 2767
rect 18093 2733 18105 2767
rect 18211 2733 18223 2767
rect 18329 2733 18341 2767
rect 18447 2733 18459 2767
rect 18565 2733 18577 2767
rect 18683 2733 18695 2767
rect 18801 2733 18813 2767
rect 18919 2733 18931 2767
rect 19037 2733 19049 2767
rect 19155 2733 19167 2767
rect 19273 2733 19285 2767
rect 19391 2733 19403 2767
rect 19509 2733 19521 2767
rect 19627 2733 19639 2767
rect 19745 2733 19757 2767
rect 19863 2733 19875 2767
rect 19981 2733 19993 2767
rect 20099 2733 20111 2767
rect 20217 2733 20229 2767
rect 20335 2733 20347 2767
rect 20453 2733 20465 2767
rect 20571 2733 20583 2767
rect 20689 2733 20701 2767
rect 20807 2733 20819 2767
rect 20925 2733 20937 2767
rect 21043 2733 21055 2767
rect 21161 2733 21173 2767
rect 21279 2733 21291 2767
rect 12547 2727 12605 2733
rect 12665 2727 12723 2733
rect 12783 2727 12841 2733
rect 12901 2727 12959 2733
rect 13019 2727 13077 2733
rect 13137 2727 13195 2733
rect 13255 2727 13313 2733
rect 13373 2727 13431 2733
rect 13491 2727 13549 2733
rect 13609 2727 13667 2733
rect 13727 2727 13785 2733
rect 13845 2727 13903 2733
rect 13963 2727 14021 2733
rect 14081 2727 14139 2733
rect 14199 2727 14257 2733
rect 14317 2727 14375 2733
rect 14435 2727 14493 2733
rect 14553 2727 14611 2733
rect 14671 2727 14729 2733
rect 14789 2727 14847 2733
rect 14907 2727 14965 2733
rect 15025 2727 15083 2733
rect 15143 2727 15201 2733
rect 15261 2727 15319 2733
rect 15379 2727 15437 2733
rect 15497 2727 15555 2733
rect 15615 2727 15673 2733
rect 15733 2727 15791 2733
rect 15851 2727 15909 2733
rect 15969 2727 16027 2733
rect 16087 2727 16145 2733
rect 16205 2727 16263 2733
rect 16323 2727 16381 2733
rect 16441 2727 16499 2733
rect 16559 2727 16617 2733
rect 16677 2727 16735 2733
rect 16795 2727 16853 2733
rect 16913 2727 16971 2733
rect 17031 2727 17089 2733
rect 17149 2727 17207 2733
rect 17267 2727 17325 2733
rect 17385 2727 17443 2733
rect 17503 2727 17561 2733
rect 17621 2727 17679 2733
rect 17739 2727 17797 2733
rect 17857 2727 17915 2733
rect 17975 2727 18033 2733
rect 18093 2727 18151 2733
rect 18211 2727 18269 2733
rect 18329 2727 18387 2733
rect 18447 2727 18505 2733
rect 18565 2727 18623 2733
rect 18683 2727 18741 2733
rect 18801 2727 18859 2733
rect 18919 2727 18977 2733
rect 19037 2727 19095 2733
rect 19155 2727 19213 2733
rect 19273 2727 19331 2733
rect 19391 2727 19449 2733
rect 19509 2727 19567 2733
rect 19627 2727 19685 2733
rect 19745 2727 19803 2733
rect 19863 2727 19921 2733
rect 19981 2727 20039 2733
rect 20099 2727 20157 2733
rect 20217 2727 20275 2733
rect 20335 2727 20393 2733
rect 20453 2727 20511 2733
rect 20571 2727 20629 2733
rect 20689 2727 20747 2733
rect 20807 2727 20865 2733
rect 20925 2727 20983 2733
rect 21043 2727 21101 2733
rect 21161 2727 21219 2733
rect 21279 2727 21337 2733
rect 717 2139 775 2145
rect 835 2139 893 2145
rect 953 2139 1011 2145
rect 1071 2139 1129 2145
rect 1189 2139 1247 2145
rect 1307 2139 1365 2145
rect 1425 2139 1483 2145
rect 1543 2139 1601 2145
rect 1661 2139 1719 2145
rect 1779 2139 1837 2145
rect 1897 2139 1955 2145
rect 2015 2139 2073 2145
rect 2133 2139 2191 2145
rect 2251 2139 2309 2145
rect 2369 2139 2427 2145
rect 717 2105 729 2139
rect 835 2105 847 2139
rect 953 2105 965 2139
rect 1071 2105 1083 2139
rect 1189 2105 1201 2139
rect 1307 2105 1319 2139
rect 1425 2105 1437 2139
rect 1543 2105 1555 2139
rect 1661 2105 1673 2139
rect 1779 2105 1791 2139
rect 1897 2105 1909 2139
rect 2015 2105 2027 2139
rect 2133 2105 2145 2139
rect 2251 2105 2263 2139
rect 2369 2105 2381 2139
rect 717 2099 775 2105
rect 835 2099 893 2105
rect 953 2099 1011 2105
rect 1071 2099 1129 2105
rect 1189 2099 1247 2105
rect 1307 2099 1365 2105
rect 1425 2099 1483 2105
rect 1543 2099 1601 2105
rect 1661 2099 1719 2105
rect 1779 2099 1837 2105
rect 1897 2099 1955 2105
rect 2015 2099 2073 2105
rect 2133 2099 2191 2105
rect 2251 2099 2309 2105
rect 2369 2099 2427 2105
rect 717 1411 775 1417
rect 835 1411 893 1417
rect 953 1411 1011 1417
rect 1071 1411 1129 1417
rect 1189 1411 1247 1417
rect 1307 1411 1365 1417
rect 1425 1411 1483 1417
rect 1543 1411 1601 1417
rect 1661 1411 1719 1417
rect 1779 1411 1837 1417
rect 1897 1411 1955 1417
rect 2015 1411 2073 1417
rect 2133 1411 2191 1417
rect 2251 1411 2309 1417
rect 2369 1411 2427 1417
rect 717 1377 729 1411
rect 835 1377 847 1411
rect 953 1377 965 1411
rect 1071 1377 1083 1411
rect 1189 1377 1201 1411
rect 1307 1377 1319 1411
rect 1425 1377 1437 1411
rect 1543 1377 1555 1411
rect 1661 1377 1673 1411
rect 1779 1377 1791 1411
rect 1897 1377 1909 1411
rect 2015 1377 2027 1411
rect 2133 1377 2145 1411
rect 2251 1377 2263 1411
rect 2369 1377 2381 1411
rect 717 1371 775 1377
rect 835 1371 893 1377
rect 953 1371 1011 1377
rect 1071 1371 1129 1377
rect 1189 1371 1247 1377
rect 1307 1371 1365 1377
rect 1425 1371 1483 1377
rect 1543 1371 1601 1377
rect 1661 1371 1719 1377
rect 1779 1371 1837 1377
rect 1897 1371 1955 1377
rect 2015 1371 2073 1377
rect 2133 1371 2191 1377
rect 2251 1371 2309 1377
rect 2369 1371 2427 1377
rect 2819 1239 2878 2277
rect 4958 2145 5177 2277
rect 3016 2139 3074 2145
rect 3134 2139 3192 2145
rect 3252 2139 3310 2145
rect 3370 2139 3428 2145
rect 3488 2139 3546 2145
rect 3606 2139 3664 2145
rect 3724 2139 3782 2145
rect 3842 2139 3900 2145
rect 3960 2139 4018 2145
rect 4078 2139 4136 2145
rect 4196 2139 4254 2145
rect 4314 2139 4372 2145
rect 4432 2139 4490 2145
rect 4550 2139 4608 2145
rect 4668 2139 4726 2145
rect 4958 2139 5213 2145
rect 5273 2139 5331 2145
rect 5391 2139 5449 2145
rect 5509 2139 5567 2145
rect 5627 2139 5685 2145
rect 5745 2139 5803 2145
rect 5863 2139 5921 2145
rect 5981 2139 6039 2145
rect 6099 2139 6157 2145
rect 6217 2139 6275 2145
rect 6335 2139 6393 2145
rect 6453 2139 6511 2145
rect 6571 2139 6629 2145
rect 6689 2139 6747 2145
rect 6807 2139 6865 2145
rect 3016 2105 3028 2139
rect 3134 2105 3146 2139
rect 3252 2105 3264 2139
rect 3370 2105 3382 2139
rect 3488 2105 3500 2139
rect 3606 2105 3618 2139
rect 3724 2105 3736 2139
rect 3842 2105 3854 2139
rect 3960 2105 3972 2139
rect 4078 2105 4090 2139
rect 4196 2105 4208 2139
rect 4314 2105 4326 2139
rect 4432 2105 4444 2139
rect 4550 2105 4562 2139
rect 4668 2105 4680 2139
rect 4958 2105 5177 2139
rect 5273 2105 5285 2139
rect 5391 2105 5403 2139
rect 5509 2105 5521 2139
rect 5627 2105 5639 2139
rect 5745 2105 5757 2139
rect 5863 2105 5875 2139
rect 5981 2105 5993 2139
rect 6099 2105 6111 2139
rect 6217 2105 6229 2139
rect 6335 2105 6347 2139
rect 6453 2105 6465 2139
rect 6571 2105 6583 2139
rect 6689 2105 6701 2139
rect 6807 2105 6819 2139
rect 3016 2099 3074 2105
rect 3134 2099 3192 2105
rect 3252 2099 3310 2105
rect 3370 2099 3428 2105
rect 3488 2099 3546 2105
rect 3606 2099 3664 2105
rect 3724 2099 3782 2105
rect 3842 2099 3900 2105
rect 3960 2099 4018 2105
rect 4078 2099 4136 2105
rect 4196 2099 4254 2105
rect 4314 2099 4372 2105
rect 4432 2099 4490 2105
rect 4550 2099 4608 2105
rect 4668 2099 4726 2105
rect 4958 2099 5213 2105
rect 5273 2099 5331 2105
rect 5391 2099 5449 2105
rect 5509 2099 5567 2105
rect 5627 2099 5685 2105
rect 5745 2099 5803 2105
rect 5863 2099 5921 2105
rect 5981 2099 6039 2105
rect 6099 2099 6157 2105
rect 6217 2099 6275 2105
rect 6335 2099 6393 2105
rect 6453 2099 6511 2105
rect 6571 2099 6629 2105
rect 6689 2099 6747 2105
rect 6807 2099 6865 2105
rect 4958 1417 5177 2099
rect 3016 1411 3074 1417
rect 3134 1411 3192 1417
rect 3252 1411 3310 1417
rect 3370 1411 3428 1417
rect 3488 1411 3546 1417
rect 3606 1411 3664 1417
rect 3724 1411 3782 1417
rect 3842 1411 3900 1417
rect 3960 1411 4018 1417
rect 4078 1411 4136 1417
rect 4196 1411 4254 1417
rect 4314 1411 4372 1417
rect 4432 1411 4490 1417
rect 4550 1411 4608 1417
rect 4668 1411 4726 1417
rect 4958 1411 5213 1417
rect 5273 1411 5331 1417
rect 5391 1411 5449 1417
rect 5509 1411 5567 1417
rect 5627 1411 5685 1417
rect 5745 1411 5803 1417
rect 5863 1411 5921 1417
rect 5981 1411 6039 1417
rect 6099 1411 6157 1417
rect 6217 1411 6275 1417
rect 6335 1411 6393 1417
rect 6453 1411 6511 1417
rect 6571 1411 6629 1417
rect 6689 1411 6747 1417
rect 6807 1411 6865 1417
rect 3016 1377 3028 1411
rect 3134 1377 3146 1411
rect 3252 1377 3264 1411
rect 3370 1377 3382 1411
rect 3488 1377 3500 1411
rect 3606 1377 3618 1411
rect 3724 1377 3736 1411
rect 3842 1377 3854 1411
rect 3960 1377 3972 1411
rect 4078 1377 4090 1411
rect 4196 1377 4208 1411
rect 4314 1377 4326 1411
rect 4432 1377 4444 1411
rect 4550 1377 4562 1411
rect 4668 1377 4680 1411
rect 4958 1377 5177 1411
rect 5273 1377 5285 1411
rect 5391 1377 5403 1411
rect 5509 1377 5521 1411
rect 5627 1377 5639 1411
rect 5745 1377 5757 1411
rect 5863 1377 5875 1411
rect 5981 1377 5993 1411
rect 6099 1377 6111 1411
rect 6217 1377 6229 1411
rect 6335 1377 6347 1411
rect 6453 1377 6465 1411
rect 6571 1377 6583 1411
rect 6689 1377 6701 1411
rect 6807 1377 6819 1411
rect 3016 1371 3074 1377
rect 3134 1371 3192 1377
rect 3252 1371 3310 1377
rect 3370 1371 3428 1377
rect 3488 1371 3546 1377
rect 3606 1371 3664 1377
rect 3724 1371 3782 1377
rect 3842 1371 3900 1377
rect 3960 1371 4018 1377
rect 4078 1371 4136 1377
rect 4196 1371 4254 1377
rect 4314 1371 4372 1377
rect 4432 1371 4490 1377
rect 4550 1371 4608 1377
rect 4668 1371 4726 1377
rect 4958 1371 5213 1377
rect 5273 1371 5331 1377
rect 5391 1371 5449 1377
rect 5509 1371 5567 1377
rect 5627 1371 5685 1377
rect 5745 1371 5803 1377
rect 5863 1371 5921 1377
rect 5981 1371 6039 1377
rect 6099 1371 6157 1377
rect 6217 1371 6275 1377
rect 6335 1371 6393 1377
rect 6453 1371 6511 1377
rect 6571 1371 6629 1377
rect 6689 1371 6747 1377
rect 6807 1371 6865 1377
rect 4958 1239 5177 1371
rect 12547 1203 12605 1209
rect 12665 1203 12723 1209
rect 12783 1203 12841 1209
rect 12901 1203 12959 1209
rect 13019 1203 13077 1209
rect 13137 1203 13195 1209
rect 13255 1203 13313 1209
rect 13373 1203 13431 1209
rect 13491 1203 13549 1209
rect 13609 1203 13667 1209
rect 13727 1203 13785 1209
rect 13845 1203 13903 1209
rect 13963 1203 14021 1209
rect 14081 1203 14139 1209
rect 14199 1203 14257 1209
rect 14317 1203 14375 1209
rect 14435 1203 14493 1209
rect 14553 1203 14611 1209
rect 14671 1203 14729 1209
rect 14789 1203 14847 1209
rect 14907 1203 14965 1209
rect 15025 1203 15083 1209
rect 15143 1203 15201 1209
rect 15261 1203 15319 1209
rect 15379 1203 15437 1209
rect 15497 1203 15555 1209
rect 15615 1203 15673 1209
rect 15733 1203 15791 1209
rect 15851 1203 15909 1209
rect 15969 1203 16027 1209
rect 16087 1203 16145 1209
rect 16205 1203 16263 1209
rect 16323 1203 16381 1209
rect 16441 1203 16499 1209
rect 16559 1203 16617 1209
rect 16677 1203 16735 1209
rect 16795 1203 16853 1209
rect 16913 1203 16971 1209
rect 17031 1203 17089 1209
rect 17149 1203 17207 1209
rect 17267 1203 17325 1209
rect 17385 1203 17443 1209
rect 17503 1203 17561 1209
rect 17621 1203 17679 1209
rect 17739 1203 17797 1209
rect 17857 1203 17915 1209
rect 17975 1203 18033 1209
rect 18093 1203 18151 1209
rect 18211 1203 18269 1209
rect 18329 1203 18387 1209
rect 18447 1203 18505 1209
rect 18565 1203 18623 1209
rect 18683 1203 18741 1209
rect 18801 1203 18859 1209
rect 18919 1203 18977 1209
rect 19037 1203 19095 1209
rect 19155 1203 19213 1209
rect 19273 1203 19331 1209
rect 19391 1203 19449 1209
rect 19509 1203 19567 1209
rect 19627 1203 19685 1209
rect 19745 1203 19803 1209
rect 19863 1203 19921 1209
rect 19981 1203 20039 1209
rect 20099 1203 20157 1209
rect 20217 1203 20275 1209
rect 20335 1203 20393 1209
rect 20453 1203 20511 1209
rect 20571 1203 20629 1209
rect 20689 1203 20747 1209
rect 20807 1203 20865 1209
rect 20925 1203 20983 1209
rect 21043 1203 21101 1209
rect 21161 1203 21219 1209
rect 21279 1203 21337 1209
rect 12547 1169 12559 1203
rect 12665 1169 12677 1203
rect 12783 1169 12795 1203
rect 12901 1169 12913 1203
rect 13019 1169 13031 1203
rect 13137 1169 13149 1203
rect 13255 1169 13267 1203
rect 13373 1169 13385 1203
rect 13491 1169 13503 1203
rect 13609 1169 13621 1203
rect 13727 1169 13739 1203
rect 13845 1169 13857 1203
rect 13963 1169 13975 1203
rect 14081 1169 14093 1203
rect 14199 1169 14211 1203
rect 14317 1169 14329 1203
rect 14435 1169 14447 1203
rect 14553 1169 14565 1203
rect 14671 1169 14683 1203
rect 14789 1169 14801 1203
rect 14907 1169 14919 1203
rect 15025 1169 15037 1203
rect 15143 1169 15155 1203
rect 15261 1169 15273 1203
rect 15379 1169 15391 1203
rect 15497 1169 15509 1203
rect 15615 1169 15627 1203
rect 15733 1169 15745 1203
rect 15851 1169 15863 1203
rect 15969 1169 15981 1203
rect 16087 1169 16099 1203
rect 16205 1169 16217 1203
rect 16323 1169 16335 1203
rect 16441 1169 16453 1203
rect 16559 1169 16571 1203
rect 16677 1169 16689 1203
rect 16795 1169 16807 1203
rect 16913 1169 16925 1203
rect 17031 1169 17043 1203
rect 17149 1169 17161 1203
rect 17267 1169 17279 1203
rect 17385 1169 17397 1203
rect 17503 1169 17515 1203
rect 17621 1169 17633 1203
rect 17739 1169 17751 1203
rect 17857 1169 17869 1203
rect 17975 1169 17987 1203
rect 18093 1169 18105 1203
rect 18211 1169 18223 1203
rect 18329 1169 18341 1203
rect 18447 1169 18459 1203
rect 18565 1169 18577 1203
rect 18683 1169 18695 1203
rect 18801 1169 18813 1203
rect 18919 1169 18931 1203
rect 19037 1169 19049 1203
rect 19155 1169 19167 1203
rect 19273 1169 19285 1203
rect 19391 1169 19403 1203
rect 19509 1169 19521 1203
rect 19627 1169 19639 1203
rect 19745 1169 19757 1203
rect 19863 1169 19875 1203
rect 19981 1169 19993 1203
rect 20099 1169 20111 1203
rect 20217 1169 20229 1203
rect 20335 1169 20347 1203
rect 20453 1169 20465 1203
rect 20571 1169 20583 1203
rect 20689 1169 20701 1203
rect 20807 1169 20819 1203
rect 20925 1169 20937 1203
rect 21043 1169 21055 1203
rect 21161 1169 21173 1203
rect 21279 1169 21291 1203
rect 12547 1163 12605 1169
rect 12665 1163 12723 1169
rect 12783 1163 12841 1169
rect 12901 1163 12959 1169
rect 13019 1163 13077 1169
rect 13137 1163 13195 1169
rect 13255 1163 13313 1169
rect 13373 1163 13431 1169
rect 13491 1163 13549 1169
rect 13609 1163 13667 1169
rect 13727 1163 13785 1169
rect 13845 1163 13903 1169
rect 13963 1163 14021 1169
rect 14081 1163 14139 1169
rect 14199 1163 14257 1169
rect 14317 1163 14375 1169
rect 14435 1163 14493 1169
rect 14553 1163 14611 1169
rect 14671 1163 14729 1169
rect 14789 1163 14847 1169
rect 14907 1163 14965 1169
rect 15025 1163 15083 1169
rect 15143 1163 15201 1169
rect 15261 1163 15319 1169
rect 15379 1163 15437 1169
rect 15497 1163 15555 1169
rect 15615 1163 15673 1169
rect 15733 1163 15791 1169
rect 15851 1163 15909 1169
rect 15969 1163 16027 1169
rect 16087 1163 16145 1169
rect 16205 1163 16263 1169
rect 16323 1163 16381 1169
rect 16441 1163 16499 1169
rect 16559 1163 16617 1169
rect 16677 1163 16735 1169
rect 16795 1163 16853 1169
rect 16913 1163 16971 1169
rect 17031 1163 17089 1169
rect 17149 1163 17207 1169
rect 17267 1163 17325 1169
rect 17385 1163 17443 1169
rect 17503 1163 17561 1169
rect 17621 1163 17679 1169
rect 17739 1163 17797 1169
rect 17857 1163 17915 1169
rect 17975 1163 18033 1169
rect 18093 1163 18151 1169
rect 18211 1163 18269 1169
rect 18329 1163 18387 1169
rect 18447 1163 18505 1169
rect 18565 1163 18623 1169
rect 18683 1163 18741 1169
rect 18801 1163 18859 1169
rect 18919 1163 18977 1169
rect 19037 1163 19095 1169
rect 19155 1163 19213 1169
rect 19273 1163 19331 1169
rect 19391 1163 19449 1169
rect 19509 1163 19567 1169
rect 19627 1163 19685 1169
rect 19745 1163 19803 1169
rect 19863 1163 19921 1169
rect 19981 1163 20039 1169
rect 20099 1163 20157 1169
rect 20217 1163 20275 1169
rect 20335 1163 20393 1169
rect 20453 1163 20511 1169
rect 20571 1163 20629 1169
rect 20689 1163 20747 1169
rect 20807 1163 20865 1169
rect 20925 1163 20983 1169
rect 21043 1163 21101 1169
rect 21161 1163 21219 1169
rect 21279 1163 21337 1169
rect 1383 583 1441 589
rect 1501 583 1559 589
rect 1619 583 1677 589
rect 1737 583 1795 589
rect 1855 583 1913 589
rect 1973 583 2031 589
rect 2091 583 2149 589
rect 2209 583 2267 589
rect 2327 583 2385 589
rect 2445 583 2503 589
rect 2563 583 2621 589
rect 2681 583 2739 589
rect 2799 583 2857 589
rect 2917 583 2975 589
rect 3035 583 3093 589
rect 3153 583 3211 589
rect 3271 583 3329 589
rect 3389 583 3447 589
rect 3507 583 3565 589
rect 3625 583 3683 589
rect 3743 583 3801 589
rect 3861 583 3919 589
rect 3979 583 4037 589
rect 4097 583 4155 589
rect 4215 583 4273 589
rect 4333 583 4391 589
rect 4451 583 4509 589
rect 4569 583 4627 589
rect 4687 583 4745 589
rect 4805 583 4863 589
rect 4923 583 4981 589
rect 5041 583 5099 589
rect 5159 583 5217 589
rect 5277 583 5335 589
rect 5395 583 5453 589
rect 5513 583 5571 589
rect 5631 583 5689 589
rect 5749 583 5807 589
rect 5867 583 5925 589
rect 5985 583 6043 589
rect 6103 583 6161 589
rect 6221 583 6279 589
rect 6339 583 6397 589
rect 6457 583 6515 589
rect 6575 583 6633 589
rect 6693 583 6751 589
rect 6811 583 6869 589
rect 6929 583 6987 589
rect 7047 583 7105 589
rect 7165 583 7223 589
rect 1383 549 1395 583
rect 1501 549 1513 583
rect 1619 549 1631 583
rect 1737 549 1749 583
rect 1855 549 1867 583
rect 1973 549 1985 583
rect 2091 549 2103 583
rect 2209 549 2221 583
rect 2327 549 2339 583
rect 2445 549 2457 583
rect 2563 549 2575 583
rect 2681 549 2693 583
rect 2799 549 2811 583
rect 2917 549 2929 583
rect 3035 549 3047 583
rect 3153 549 3165 583
rect 3271 549 3283 583
rect 3389 549 3401 583
rect 3507 549 3519 583
rect 3625 549 3637 583
rect 3743 549 3755 583
rect 3861 549 3873 583
rect 3979 549 3991 583
rect 4097 549 4109 583
rect 4215 549 4227 583
rect 4333 549 4345 583
rect 4451 549 4463 583
rect 4569 549 4581 583
rect 4687 549 4699 583
rect 4805 549 4817 583
rect 4923 549 4935 583
rect 5041 549 5053 583
rect 5159 549 5171 583
rect 5277 549 5289 583
rect 5395 549 5407 583
rect 5513 549 5525 583
rect 5631 549 5643 583
rect 5749 549 5761 583
rect 5867 549 5879 583
rect 5985 549 5997 583
rect 6103 549 6115 583
rect 6221 549 6233 583
rect 6339 549 6351 583
rect 6457 549 6469 583
rect 6575 549 6587 583
rect 6693 549 6705 583
rect 6811 549 6823 583
rect 6929 549 6941 583
rect 7047 549 7059 583
rect 7165 549 7177 583
rect 1383 543 1441 549
rect 1501 543 1559 549
rect 1619 543 1677 549
rect 1737 543 1795 549
rect 1855 543 1913 549
rect 1973 543 2031 549
rect 2091 543 2149 549
rect 2209 543 2267 549
rect 2327 543 2385 549
rect 2445 543 2503 549
rect 2563 543 2621 549
rect 2681 543 2739 549
rect 2799 543 2857 549
rect 2917 543 2975 549
rect 3035 543 3093 549
rect 3153 543 3211 549
rect 3271 543 3329 549
rect 3389 543 3447 549
rect 3507 543 3565 549
rect 3625 543 3683 549
rect 3743 543 3801 549
rect 3861 543 3919 549
rect 3979 543 4037 549
rect 4097 543 4155 549
rect 4215 543 4273 549
rect 4333 543 4391 549
rect 4451 543 4509 549
rect 4569 543 4627 549
rect 4687 543 4745 549
rect 4805 543 4863 549
rect 4923 543 4981 549
rect 5041 543 5099 549
rect 5159 543 5217 549
rect 5277 543 5335 549
rect 5395 543 5453 549
rect 5513 543 5571 549
rect 5631 543 5689 549
rect 5749 543 5807 549
rect 5867 543 5925 549
rect 5985 543 6043 549
rect 6103 543 6161 549
rect 6221 543 6279 549
rect 6339 543 6397 549
rect 6457 543 6515 549
rect 6575 543 6633 549
rect 6693 543 6751 549
rect 6811 543 6869 549
rect 6929 543 6987 549
rect 7047 543 7105 549
rect 7165 543 7223 549
rect 1383 -145 1441 -139
rect 1501 -145 1559 -139
rect 1619 -145 1677 -139
rect 1737 -145 1795 -139
rect 1855 -145 1913 -139
rect 1973 -145 2031 -139
rect 2091 -145 2149 -139
rect 2209 -145 2267 -139
rect 2327 -145 2385 -139
rect 2445 -145 2503 -139
rect 2563 -145 2621 -139
rect 2681 -145 2739 -139
rect 2799 -145 2857 -139
rect 2917 -145 2975 -139
rect 3035 -145 3093 -139
rect 3153 -145 3211 -139
rect 3271 -145 3329 -139
rect 3389 -145 3447 -139
rect 3507 -145 3565 -139
rect 3625 -145 3683 -139
rect 3743 -145 3801 -139
rect 3861 -145 3919 -139
rect 3979 -145 4037 -139
rect 4097 -145 4155 -139
rect 4215 -145 4273 -139
rect 4333 -145 4391 -139
rect 4451 -145 4509 -139
rect 4569 -145 4627 -139
rect 4687 -145 4745 -139
rect 4805 -145 4863 -139
rect 4923 -145 4981 -139
rect 5041 -145 5099 -139
rect 5159 -145 5217 -139
rect 5277 -145 5335 -139
rect 5395 -145 5453 -139
rect 5513 -145 5571 -139
rect 5631 -145 5689 -139
rect 5749 -145 5807 -139
rect 5867 -145 5925 -139
rect 5985 -145 6043 -139
rect 6103 -145 6161 -139
rect 6221 -145 6279 -139
rect 6339 -145 6397 -139
rect 6457 -145 6515 -139
rect 6575 -145 6633 -139
rect 6693 -145 6751 -139
rect 6811 -145 6869 -139
rect 6929 -145 6987 -139
rect 7047 -145 7105 -139
rect 7165 -145 7223 -139
rect 1383 -179 1395 -145
rect 1501 -179 1513 -145
rect 1619 -179 1631 -145
rect 1737 -179 1749 -145
rect 1855 -179 1867 -145
rect 1973 -179 1985 -145
rect 2091 -179 2103 -145
rect 2209 -179 2221 -145
rect 2327 -179 2339 -145
rect 2445 -179 2457 -145
rect 2563 -179 2575 -145
rect 2681 -179 2693 -145
rect 2799 -179 2811 -145
rect 2917 -179 2929 -145
rect 3035 -179 3047 -145
rect 3153 -179 3165 -145
rect 3271 -179 3283 -145
rect 3389 -179 3401 -145
rect 3507 -179 3519 -145
rect 3625 -179 3637 -145
rect 3743 -179 3755 -145
rect 3861 -179 3873 -145
rect 3979 -179 3991 -145
rect 4097 -179 4109 -145
rect 4215 -179 4227 -145
rect 4333 -179 4345 -145
rect 4451 -179 4463 -145
rect 4569 -179 4581 -145
rect 4687 -179 4699 -145
rect 4805 -179 4817 -145
rect 4923 -179 4935 -145
rect 5041 -179 5053 -145
rect 5159 -179 5171 -145
rect 5277 -179 5289 -145
rect 5395 -179 5407 -145
rect 5513 -179 5525 -145
rect 5631 -179 5643 -145
rect 5749 -179 5761 -145
rect 5867 -179 5879 -145
rect 5985 -179 5997 -145
rect 6103 -179 6115 -145
rect 6221 -179 6233 -145
rect 6339 -179 6351 -145
rect 6457 -179 6469 -145
rect 6575 -179 6587 -145
rect 6693 -179 6705 -145
rect 6811 -179 6823 -145
rect 6929 -179 6941 -145
rect 7047 -179 7059 -145
rect 7165 -179 7177 -145
rect 1383 -185 1441 -179
rect 1501 -185 1559 -179
rect 1619 -185 1677 -179
rect 1737 -185 1795 -179
rect 1855 -185 1913 -179
rect 1973 -185 2031 -179
rect 2091 -185 2149 -179
rect 2209 -185 2267 -179
rect 2327 -185 2385 -179
rect 2445 -185 2503 -179
rect 2563 -185 2621 -179
rect 2681 -185 2739 -179
rect 2799 -185 2857 -179
rect 2917 -185 2975 -179
rect 3035 -185 3093 -179
rect 3153 -185 3211 -179
rect 3271 -185 3329 -179
rect 3389 -185 3447 -179
rect 3507 -185 3565 -179
rect 3625 -185 3683 -179
rect 3743 -185 3801 -179
rect 3861 -185 3919 -179
rect 3979 -185 4037 -179
rect 4097 -185 4155 -179
rect 4215 -185 4273 -179
rect 4333 -185 4391 -179
rect 4451 -185 4509 -179
rect 4569 -185 4627 -179
rect 4687 -185 4745 -179
rect 4805 -185 4863 -179
rect 4923 -185 4981 -179
rect 5041 -185 5099 -179
rect 5159 -185 5217 -179
rect 5277 -185 5335 -179
rect 5395 -185 5453 -179
rect 5513 -185 5571 -179
rect 5631 -185 5689 -179
rect 5749 -185 5807 -179
rect 5867 -185 5925 -179
rect 5985 -185 6043 -179
rect 6103 -185 6161 -179
rect 6221 -185 6279 -179
rect 6339 -185 6397 -179
rect 6457 -185 6515 -179
rect 6575 -185 6633 -179
rect 6693 -185 6751 -179
rect 6811 -185 6869 -179
rect 6929 -185 6987 -179
rect 7047 -185 7105 -179
rect 7165 -185 7223 -179
rect 1383 -253 1441 -247
rect 1501 -253 1559 -247
rect 1619 -253 1677 -247
rect 1737 -253 1795 -247
rect 1855 -253 1913 -247
rect 1973 -253 2031 -247
rect 2091 -253 2149 -247
rect 2209 -253 2267 -247
rect 2327 -253 2385 -247
rect 2445 -253 2503 -247
rect 2563 -253 2621 -247
rect 2681 -253 2739 -247
rect 2799 -253 2857 -247
rect 2917 -253 2975 -247
rect 3035 -253 3093 -247
rect 3153 -253 3211 -247
rect 3271 -253 3329 -247
rect 3389 -253 3447 -247
rect 3507 -253 3565 -247
rect 3625 -253 3683 -247
rect 3743 -253 3801 -247
rect 3861 -253 3919 -247
rect 3979 -253 4037 -247
rect 4097 -253 4155 -247
rect 4215 -253 4273 -247
rect 4333 -253 4391 -247
rect 4451 -253 4509 -247
rect 4569 -253 4627 -247
rect 4687 -253 4745 -247
rect 4805 -253 4863 -247
rect 4923 -253 4981 -247
rect 5041 -253 5099 -247
rect 5159 -253 5217 -247
rect 5277 -253 5335 -247
rect 5395 -253 5453 -247
rect 5513 -253 5571 -247
rect 5631 -253 5689 -247
rect 5749 -253 5807 -247
rect 5867 -253 5925 -247
rect 5985 -253 6043 -247
rect 6103 -253 6161 -247
rect 6221 -253 6279 -247
rect 6339 -253 6397 -247
rect 6457 -253 6515 -247
rect 6575 -253 6633 -247
rect 6693 -253 6751 -247
rect 6811 -253 6869 -247
rect 6929 -253 6987 -247
rect 7047 -253 7105 -247
rect 7165 -253 7223 -247
rect 1383 -287 1395 -253
rect 1501 -287 1513 -253
rect 1619 -287 1631 -253
rect 1737 -287 1749 -253
rect 1855 -287 1867 -253
rect 1973 -287 1985 -253
rect 2091 -287 2103 -253
rect 2209 -287 2221 -253
rect 2327 -287 2339 -253
rect 2445 -287 2457 -253
rect 2563 -287 2575 -253
rect 2681 -287 2693 -253
rect 2799 -287 2811 -253
rect 2917 -287 2929 -253
rect 3035 -287 3047 -253
rect 3153 -287 3165 -253
rect 3271 -287 3283 -253
rect 3389 -287 3401 -253
rect 3507 -287 3519 -253
rect 3625 -287 3637 -253
rect 3743 -287 3755 -253
rect 3861 -287 3873 -253
rect 3979 -287 3991 -253
rect 4097 -287 4109 -253
rect 4215 -287 4227 -253
rect 4333 -287 4345 -253
rect 4451 -287 4463 -253
rect 4569 -287 4581 -253
rect 4687 -287 4699 -253
rect 4805 -287 4817 -253
rect 4923 -287 4935 -253
rect 5041 -287 5053 -253
rect 5159 -287 5171 -253
rect 5277 -287 5289 -253
rect 5395 -287 5407 -253
rect 5513 -287 5525 -253
rect 5631 -287 5643 -253
rect 5749 -287 5761 -253
rect 5867 -287 5879 -253
rect 5985 -287 5997 -253
rect 6103 -287 6115 -253
rect 6221 -287 6233 -253
rect 6339 -287 6351 -253
rect 6457 -287 6469 -253
rect 6575 -287 6587 -253
rect 6693 -287 6705 -253
rect 6811 -287 6823 -253
rect 6929 -287 6941 -253
rect 7047 -287 7059 -253
rect 7165 -287 7177 -253
rect 1383 -293 1441 -287
rect 1501 -293 1559 -287
rect 1619 -293 1677 -287
rect 1737 -293 1795 -287
rect 1855 -293 1913 -287
rect 1973 -293 2031 -287
rect 2091 -293 2149 -287
rect 2209 -293 2267 -287
rect 2327 -293 2385 -287
rect 2445 -293 2503 -287
rect 2563 -293 2621 -287
rect 2681 -293 2739 -287
rect 2799 -293 2857 -287
rect 2917 -293 2975 -287
rect 3035 -293 3093 -287
rect 3153 -293 3211 -287
rect 3271 -293 3329 -287
rect 3389 -293 3447 -287
rect 3507 -293 3565 -287
rect 3625 -293 3683 -287
rect 3743 -293 3801 -287
rect 3861 -293 3919 -287
rect 3979 -293 4037 -287
rect 4097 -293 4155 -287
rect 4215 -293 4273 -287
rect 4333 -293 4391 -287
rect 4451 -293 4509 -287
rect 4569 -293 4627 -287
rect 4687 -293 4745 -287
rect 4805 -293 4863 -287
rect 4923 -293 4981 -287
rect 5041 -293 5099 -287
rect 5159 -293 5217 -287
rect 5277 -293 5335 -287
rect 5395 -293 5453 -287
rect 5513 -293 5571 -287
rect 5631 -293 5689 -287
rect 5749 -293 5807 -287
rect 5867 -293 5925 -287
rect 5985 -293 6043 -287
rect 6103 -293 6161 -287
rect 6221 -293 6279 -287
rect 6339 -293 6397 -287
rect 6457 -293 6515 -287
rect 6575 -293 6633 -287
rect 6693 -293 6751 -287
rect 6811 -293 6869 -287
rect 6929 -293 6987 -287
rect 7047 -293 7105 -287
rect 7165 -293 7223 -287
rect 1383 -981 1441 -975
rect 1501 -981 1559 -975
rect 1619 -981 1677 -975
rect 1737 -981 1795 -975
rect 1855 -981 1913 -975
rect 1973 -981 2031 -975
rect 2091 -981 2149 -975
rect 2209 -981 2267 -975
rect 2327 -981 2385 -975
rect 2445 -981 2503 -975
rect 2563 -981 2621 -975
rect 2681 -981 2739 -975
rect 2799 -981 2857 -975
rect 2917 -981 2975 -975
rect 3035 -981 3093 -975
rect 3153 -981 3211 -975
rect 3271 -981 3329 -975
rect 3389 -981 3447 -975
rect 3507 -981 3565 -975
rect 3625 -981 3683 -975
rect 3743 -981 3801 -975
rect 3861 -981 3919 -975
rect 3979 -981 4037 -975
rect 4097 -981 4155 -975
rect 4215 -981 4273 -975
rect 4333 -981 4391 -975
rect 4451 -981 4509 -975
rect 4569 -981 4627 -975
rect 4687 -981 4745 -975
rect 4805 -981 4863 -975
rect 4923 -981 4981 -975
rect 5041 -981 5099 -975
rect 5159 -981 5217 -975
rect 5277 -981 5335 -975
rect 5395 -981 5453 -975
rect 5513 -981 5571 -975
rect 5631 -981 5689 -975
rect 5749 -981 5807 -975
rect 5867 -981 5925 -975
rect 5985 -981 6043 -975
rect 6103 -981 6161 -975
rect 6221 -981 6279 -975
rect 6339 -981 6397 -975
rect 6457 -981 6515 -975
rect 6575 -981 6633 -975
rect 6693 -981 6751 -975
rect 6811 -981 6869 -975
rect 6929 -981 6987 -975
rect 7047 -981 7105 -975
rect 7165 -981 7223 -975
rect 1383 -1015 1395 -981
rect 1501 -1015 1513 -981
rect 1619 -1015 1631 -981
rect 1737 -1015 1749 -981
rect 1855 -1015 1867 -981
rect 1973 -1015 1985 -981
rect 2091 -1015 2103 -981
rect 2209 -1015 2221 -981
rect 2327 -1015 2339 -981
rect 2445 -1015 2457 -981
rect 2563 -1015 2575 -981
rect 2681 -1015 2693 -981
rect 2799 -1015 2811 -981
rect 2917 -1015 2929 -981
rect 3035 -1015 3047 -981
rect 3153 -1015 3165 -981
rect 3271 -1015 3283 -981
rect 3389 -1015 3401 -981
rect 3507 -1015 3519 -981
rect 3625 -1015 3637 -981
rect 3743 -1015 3755 -981
rect 3861 -1015 3873 -981
rect 3979 -1015 3991 -981
rect 4097 -1015 4109 -981
rect 4215 -1015 4227 -981
rect 4333 -1015 4345 -981
rect 4451 -1015 4463 -981
rect 4569 -1015 4581 -981
rect 4687 -1015 4699 -981
rect 4805 -1015 4817 -981
rect 4923 -1015 4935 -981
rect 5041 -1015 5053 -981
rect 5159 -1015 5171 -981
rect 5277 -1015 5289 -981
rect 5395 -1015 5407 -981
rect 5513 -1015 5525 -981
rect 5631 -1015 5643 -981
rect 5749 -1015 5761 -981
rect 5867 -1015 5879 -981
rect 5985 -1015 5997 -981
rect 6103 -1015 6115 -981
rect 6221 -1015 6233 -981
rect 6339 -1015 6351 -981
rect 6457 -1015 6469 -981
rect 6575 -1015 6587 -981
rect 6693 -1015 6705 -981
rect 6811 -1015 6823 -981
rect 6929 -1015 6941 -981
rect 7047 -1015 7059 -981
rect 7165 -1015 7177 -981
rect 1383 -1021 1441 -1015
rect 1501 -1021 1559 -1015
rect 1619 -1021 1677 -1015
rect 1737 -1021 1795 -1015
rect 1855 -1021 1913 -1015
rect 1973 -1021 2031 -1015
rect 2091 -1021 2149 -1015
rect 2209 -1021 2267 -1015
rect 2327 -1021 2385 -1015
rect 2445 -1021 2503 -1015
rect 2563 -1021 2621 -1015
rect 2681 -1021 2739 -1015
rect 2799 -1021 2857 -1015
rect 2917 -1021 2975 -1015
rect 3035 -1021 3093 -1015
rect 3153 -1021 3211 -1015
rect 3271 -1021 3329 -1015
rect 3389 -1021 3447 -1015
rect 3507 -1021 3565 -1015
rect 3625 -1021 3683 -1015
rect 3743 -1021 3801 -1015
rect 3861 -1021 3919 -1015
rect 3979 -1021 4037 -1015
rect 4097 -1021 4155 -1015
rect 4215 -1021 4273 -1015
rect 4333 -1021 4391 -1015
rect 4451 -1021 4509 -1015
rect 4569 -1021 4627 -1015
rect 4687 -1021 4745 -1015
rect 4805 -1021 4863 -1015
rect 4923 -1021 4981 -1015
rect 5041 -1021 5099 -1015
rect 5159 -1021 5217 -1015
rect 5277 -1021 5335 -1015
rect 5395 -1021 5453 -1015
rect 5513 -1021 5571 -1015
rect 5631 -1021 5689 -1015
rect 5749 -1021 5807 -1015
rect 5867 -1021 5925 -1015
rect 5985 -1021 6043 -1015
rect 6103 -1021 6161 -1015
rect 6221 -1021 6279 -1015
rect 6339 -1021 6397 -1015
rect 6457 -1021 6515 -1015
rect 6575 -1021 6633 -1015
rect 6693 -1021 6751 -1015
rect 6811 -1021 6869 -1015
rect 6929 -1021 6987 -1015
rect 7047 -1021 7105 -1015
rect 7165 -1021 7223 -1015
rect 1318 -1086 7288 -1083
rect 1272 -1117 7288 -1086
rect 1272 -1120 7242 -1117
rect 1337 -1188 1395 -1182
rect 1455 -1188 1513 -1182
rect 1573 -1188 1631 -1182
rect 1691 -1188 1749 -1182
rect 1809 -1188 1867 -1182
rect 1927 -1188 1985 -1182
rect 2045 -1188 2103 -1182
rect 2163 -1188 2221 -1182
rect 2281 -1188 2339 -1182
rect 2399 -1188 2457 -1182
rect 2517 -1188 2575 -1182
rect 2635 -1188 2693 -1182
rect 2753 -1188 2811 -1182
rect 2871 -1188 2929 -1182
rect 2989 -1188 3047 -1182
rect 3107 -1188 3165 -1182
rect 3225 -1188 3283 -1182
rect 3343 -1188 3401 -1182
rect 3461 -1188 3519 -1182
rect 3579 -1188 3637 -1182
rect 3697 -1188 3755 -1182
rect 3815 -1188 3873 -1182
rect 3933 -1188 3991 -1182
rect 4051 -1188 4109 -1182
rect 4169 -1188 4227 -1182
rect 4287 -1188 4345 -1182
rect 4405 -1188 4463 -1182
rect 4523 -1188 4581 -1182
rect 4641 -1188 4699 -1182
rect 4759 -1188 4817 -1182
rect 4877 -1188 4935 -1182
rect 4995 -1188 5053 -1182
rect 5113 -1188 5171 -1182
rect 5231 -1188 5289 -1182
rect 5349 -1188 5407 -1182
rect 5467 -1188 5525 -1182
rect 5585 -1188 5643 -1182
rect 5703 -1188 5761 -1182
rect 5821 -1188 5879 -1182
rect 5939 -1188 5997 -1182
rect 6057 -1188 6115 -1182
rect 6175 -1188 6233 -1182
rect 6293 -1188 6351 -1182
rect 6411 -1188 6469 -1182
rect 6529 -1188 6587 -1182
rect 6647 -1188 6705 -1182
rect 6765 -1188 6823 -1182
rect 6883 -1188 6941 -1182
rect 7001 -1188 7059 -1182
rect 7119 -1188 7177 -1182
rect 1337 -1222 1349 -1188
rect 1455 -1222 1467 -1188
rect 1573 -1222 1585 -1188
rect 1691 -1222 1703 -1188
rect 1809 -1222 1821 -1188
rect 1927 -1222 1939 -1188
rect 2045 -1222 2057 -1188
rect 2163 -1222 2175 -1188
rect 2281 -1222 2293 -1188
rect 2399 -1222 2411 -1188
rect 2517 -1222 2529 -1188
rect 2635 -1222 2647 -1188
rect 2753 -1222 2765 -1188
rect 2871 -1222 2883 -1188
rect 2989 -1222 3001 -1188
rect 3107 -1222 3119 -1188
rect 3225 -1222 3237 -1188
rect 3343 -1222 3355 -1188
rect 3461 -1222 3473 -1188
rect 3579 -1222 3591 -1188
rect 3697 -1222 3709 -1188
rect 3815 -1222 3827 -1188
rect 3933 -1222 3945 -1188
rect 4051 -1222 4063 -1188
rect 4169 -1222 4181 -1188
rect 4287 -1222 4299 -1188
rect 4405 -1222 4417 -1188
rect 4523 -1222 4535 -1188
rect 4641 -1222 4653 -1188
rect 4759 -1222 4771 -1188
rect 4877 -1222 4889 -1188
rect 4995 -1222 5007 -1188
rect 5113 -1222 5125 -1188
rect 5231 -1222 5243 -1188
rect 5349 -1222 5361 -1188
rect 5467 -1222 5479 -1188
rect 5585 -1222 5597 -1188
rect 5703 -1222 5715 -1188
rect 5821 -1222 5833 -1188
rect 5939 -1222 5951 -1188
rect 6057 -1222 6069 -1188
rect 6175 -1222 6187 -1188
rect 6293 -1222 6305 -1188
rect 6411 -1222 6423 -1188
rect 6529 -1222 6541 -1188
rect 6647 -1222 6659 -1188
rect 6765 -1222 6777 -1188
rect 6883 -1222 6895 -1188
rect 7001 -1222 7013 -1188
rect 7119 -1222 7131 -1188
rect 1337 -1228 1395 -1222
rect 1455 -1228 1513 -1222
rect 1573 -1228 1631 -1222
rect 1691 -1228 1749 -1222
rect 1809 -1228 1867 -1222
rect 1927 -1228 1985 -1222
rect 2045 -1228 2103 -1222
rect 2163 -1228 2221 -1222
rect 2281 -1228 2339 -1222
rect 2399 -1228 2457 -1222
rect 2517 -1228 2575 -1222
rect 2635 -1228 2693 -1222
rect 2753 -1228 2811 -1222
rect 2871 -1228 2929 -1222
rect 2989 -1228 3047 -1222
rect 3107 -1228 3165 -1222
rect 3225 -1228 3283 -1222
rect 3343 -1228 3401 -1222
rect 3461 -1228 3519 -1222
rect 3579 -1228 3637 -1222
rect 3697 -1228 3755 -1222
rect 3815 -1228 3873 -1222
rect 3933 -1228 3991 -1222
rect 4051 -1228 4109 -1222
rect 4169 -1228 4227 -1222
rect 4287 -1228 4345 -1222
rect 4405 -1228 4463 -1222
rect 4523 -1228 4581 -1222
rect 4641 -1228 4699 -1222
rect 4759 -1228 4817 -1222
rect 4877 -1228 4935 -1222
rect 4995 -1228 5053 -1222
rect 5113 -1228 5171 -1222
rect 5231 -1228 5289 -1222
rect 5349 -1228 5407 -1222
rect 5467 -1228 5525 -1222
rect 5585 -1228 5643 -1222
rect 5703 -1228 5761 -1222
rect 5821 -1228 5879 -1222
rect 5939 -1228 5997 -1222
rect 6057 -1228 6115 -1222
rect 6175 -1228 6233 -1222
rect 6293 -1228 6351 -1222
rect 6411 -1228 6469 -1222
rect 6529 -1228 6587 -1222
rect 6647 -1228 6705 -1222
rect 6765 -1228 6823 -1222
rect 6883 -1228 6941 -1222
rect 7001 -1228 7059 -1222
rect 7119 -1228 7177 -1222
rect 1337 -1916 1395 -1910
rect 1455 -1916 1513 -1910
rect 1573 -1916 1631 -1910
rect 1691 -1916 1749 -1910
rect 1809 -1916 1867 -1910
rect 1927 -1916 1985 -1910
rect 2045 -1916 2103 -1910
rect 2163 -1916 2221 -1910
rect 2281 -1916 2339 -1910
rect 2399 -1916 2457 -1910
rect 2517 -1916 2575 -1910
rect 2635 -1916 2693 -1910
rect 2753 -1916 2811 -1910
rect 2871 -1916 2929 -1910
rect 2989 -1916 3047 -1910
rect 3107 -1916 3165 -1910
rect 3225 -1916 3283 -1910
rect 3343 -1916 3401 -1910
rect 3461 -1916 3519 -1910
rect 3579 -1916 3637 -1910
rect 3697 -1916 3755 -1910
rect 3815 -1916 3873 -1910
rect 3933 -1916 3991 -1910
rect 4051 -1916 4109 -1910
rect 4169 -1916 4227 -1910
rect 4287 -1916 4345 -1910
rect 4405 -1916 4463 -1910
rect 4523 -1916 4581 -1910
rect 4641 -1916 4699 -1910
rect 4759 -1916 4817 -1910
rect 4877 -1916 4935 -1910
rect 4995 -1916 5053 -1910
rect 5113 -1916 5171 -1910
rect 5231 -1916 5289 -1910
rect 5349 -1916 5407 -1910
rect 5467 -1916 5525 -1910
rect 5585 -1916 5643 -1910
rect 5703 -1916 5761 -1910
rect 5821 -1916 5879 -1910
rect 5939 -1916 5997 -1910
rect 6057 -1916 6115 -1910
rect 6175 -1916 6233 -1910
rect 6293 -1916 6351 -1910
rect 6411 -1916 6469 -1910
rect 6529 -1916 6587 -1910
rect 6647 -1916 6705 -1910
rect 6765 -1916 6823 -1910
rect 6883 -1916 6941 -1910
rect 7001 -1916 7059 -1910
rect 7119 -1916 7177 -1910
rect 1337 -1950 1349 -1916
rect 1455 -1950 1467 -1916
rect 1573 -1950 1585 -1916
rect 1691 -1950 1703 -1916
rect 1809 -1950 1821 -1916
rect 1927 -1950 1939 -1916
rect 2045 -1950 2057 -1916
rect 2163 -1950 2175 -1916
rect 2281 -1950 2293 -1916
rect 2399 -1950 2411 -1916
rect 2517 -1950 2529 -1916
rect 2635 -1950 2647 -1916
rect 2753 -1950 2765 -1916
rect 2871 -1950 2883 -1916
rect 2989 -1950 3001 -1916
rect 3107 -1950 3119 -1916
rect 3225 -1950 3237 -1916
rect 3343 -1950 3355 -1916
rect 3461 -1950 3473 -1916
rect 3579 -1950 3591 -1916
rect 3697 -1950 3709 -1916
rect 3815 -1950 3827 -1916
rect 3933 -1950 3945 -1916
rect 4051 -1950 4063 -1916
rect 4169 -1950 4181 -1916
rect 4287 -1950 4299 -1916
rect 4405 -1950 4417 -1916
rect 4523 -1950 4535 -1916
rect 4641 -1950 4653 -1916
rect 4759 -1950 4771 -1916
rect 4877 -1950 4889 -1916
rect 4995 -1950 5007 -1916
rect 5113 -1950 5125 -1916
rect 5231 -1950 5243 -1916
rect 5349 -1950 5361 -1916
rect 5467 -1950 5479 -1916
rect 5585 -1950 5597 -1916
rect 5703 -1950 5715 -1916
rect 5821 -1950 5833 -1916
rect 5939 -1950 5951 -1916
rect 6057 -1950 6069 -1916
rect 6175 -1950 6187 -1916
rect 6293 -1950 6305 -1916
rect 6411 -1950 6423 -1916
rect 6529 -1950 6541 -1916
rect 6647 -1950 6659 -1916
rect 6765 -1950 6777 -1916
rect 6883 -1950 6895 -1916
rect 7001 -1950 7013 -1916
rect 7119 -1950 7131 -1916
rect 1337 -1956 1395 -1950
rect 1455 -1956 1513 -1950
rect 1573 -1956 1631 -1950
rect 1691 -1956 1749 -1950
rect 1809 -1956 1867 -1950
rect 1927 -1956 1985 -1950
rect 2045 -1956 2103 -1950
rect 2163 -1956 2221 -1950
rect 2281 -1956 2339 -1950
rect 2399 -1956 2457 -1950
rect 2517 -1956 2575 -1950
rect 2635 -1956 2693 -1950
rect 2753 -1956 2811 -1950
rect 2871 -1956 2929 -1950
rect 2989 -1956 3047 -1950
rect 3107 -1956 3165 -1950
rect 3225 -1956 3283 -1950
rect 3343 -1956 3401 -1950
rect 3461 -1956 3519 -1950
rect 3579 -1956 3637 -1950
rect 3697 -1956 3755 -1950
rect 3815 -1956 3873 -1950
rect 3933 -1956 3991 -1950
rect 4051 -1956 4109 -1950
rect 4169 -1956 4227 -1950
rect 4287 -1956 4345 -1950
rect 4405 -1956 4463 -1950
rect 4523 -1956 4581 -1950
rect 4641 -1956 4699 -1950
rect 4759 -1956 4817 -1950
rect 4877 -1956 4935 -1950
rect 4995 -1956 5053 -1950
rect 5113 -1956 5171 -1950
rect 5231 -1956 5289 -1950
rect 5349 -1956 5407 -1950
rect 5467 -1956 5525 -1950
rect 5585 -1956 5643 -1950
rect 5703 -1956 5761 -1950
rect 5821 -1956 5879 -1950
rect 5939 -1956 5997 -1950
rect 6057 -1956 6115 -1950
rect 6175 -1956 6233 -1950
rect 6293 -1956 6351 -1950
rect 6411 -1956 6469 -1950
rect 6529 -1956 6587 -1950
rect 6647 -1956 6705 -1950
rect 6765 -1956 6823 -1950
rect 6883 -1956 6941 -1950
rect 7001 -1956 7059 -1950
rect 7119 -1956 7177 -1950
rect 1337 -2024 1395 -2018
rect 1455 -2024 1513 -2018
rect 1573 -2024 1631 -2018
rect 1691 -2024 1749 -2018
rect 1809 -2024 1867 -2018
rect 1927 -2024 1985 -2018
rect 2045 -2024 2103 -2018
rect 2163 -2024 2221 -2018
rect 2281 -2024 2339 -2018
rect 2399 -2024 2457 -2018
rect 2517 -2024 2575 -2018
rect 2635 -2024 2693 -2018
rect 2753 -2024 2811 -2018
rect 2871 -2024 2929 -2018
rect 2989 -2024 3047 -2018
rect 3107 -2024 3165 -2018
rect 3225 -2024 3283 -2018
rect 3343 -2024 3401 -2018
rect 3461 -2024 3519 -2018
rect 3579 -2024 3637 -2018
rect 3697 -2024 3755 -2018
rect 3815 -2024 3873 -2018
rect 3933 -2024 3991 -2018
rect 4051 -2024 4109 -2018
rect 4169 -2024 4227 -2018
rect 4287 -2024 4345 -2018
rect 4405 -2024 4463 -2018
rect 4523 -2024 4581 -2018
rect 4641 -2024 4699 -2018
rect 4759 -2024 4817 -2018
rect 4877 -2024 4935 -2018
rect 4995 -2024 5053 -2018
rect 5113 -2024 5171 -2018
rect 5231 -2024 5289 -2018
rect 5349 -2024 5407 -2018
rect 5467 -2024 5525 -2018
rect 5585 -2024 5643 -2018
rect 5703 -2024 5761 -2018
rect 5821 -2024 5879 -2018
rect 5939 -2024 5997 -2018
rect 6057 -2024 6115 -2018
rect 6175 -2024 6233 -2018
rect 6293 -2024 6351 -2018
rect 6411 -2024 6469 -2018
rect 6529 -2024 6587 -2018
rect 6647 -2024 6705 -2018
rect 6765 -2024 6823 -2018
rect 6883 -2024 6941 -2018
rect 7001 -2024 7059 -2018
rect 7119 -2024 7177 -2018
rect 1337 -2058 1349 -2024
rect 1455 -2058 1467 -2024
rect 1573 -2058 1585 -2024
rect 1691 -2058 1703 -2024
rect 1809 -2058 1821 -2024
rect 1927 -2058 1939 -2024
rect 2045 -2058 2057 -2024
rect 2163 -2058 2175 -2024
rect 2281 -2058 2293 -2024
rect 2399 -2058 2411 -2024
rect 2517 -2058 2529 -2024
rect 2635 -2058 2647 -2024
rect 2753 -2058 2765 -2024
rect 2871 -2058 2883 -2024
rect 2989 -2058 3001 -2024
rect 3107 -2058 3119 -2024
rect 3225 -2058 3237 -2024
rect 3343 -2058 3355 -2024
rect 3461 -2058 3473 -2024
rect 3579 -2058 3591 -2024
rect 3697 -2058 3709 -2024
rect 3815 -2058 3827 -2024
rect 3933 -2058 3945 -2024
rect 4051 -2058 4063 -2024
rect 4169 -2058 4181 -2024
rect 4287 -2058 4299 -2024
rect 4405 -2058 4417 -2024
rect 4523 -2058 4535 -2024
rect 4641 -2058 4653 -2024
rect 4759 -2058 4771 -2024
rect 4877 -2058 4889 -2024
rect 4995 -2058 5007 -2024
rect 5113 -2058 5125 -2024
rect 5231 -2058 5243 -2024
rect 5349 -2058 5361 -2024
rect 5467 -2058 5479 -2024
rect 5585 -2058 5597 -2024
rect 5703 -2058 5715 -2024
rect 5821 -2058 5833 -2024
rect 5939 -2058 5951 -2024
rect 6057 -2058 6069 -2024
rect 6175 -2058 6187 -2024
rect 6293 -2058 6305 -2024
rect 6411 -2058 6423 -2024
rect 6529 -2058 6541 -2024
rect 6647 -2058 6659 -2024
rect 6765 -2058 6777 -2024
rect 6883 -2058 6895 -2024
rect 7001 -2058 7013 -2024
rect 7119 -2058 7131 -2024
rect 1337 -2064 1395 -2058
rect 1455 -2064 1513 -2058
rect 1573 -2064 1631 -2058
rect 1691 -2064 1749 -2058
rect 1809 -2064 1867 -2058
rect 1927 -2064 1985 -2058
rect 2045 -2064 2103 -2058
rect 2163 -2064 2221 -2058
rect 2281 -2064 2339 -2058
rect 2399 -2064 2457 -2058
rect 2517 -2064 2575 -2058
rect 2635 -2064 2693 -2058
rect 2753 -2064 2811 -2058
rect 2871 -2064 2929 -2058
rect 2989 -2064 3047 -2058
rect 3107 -2064 3165 -2058
rect 3225 -2064 3283 -2058
rect 3343 -2064 3401 -2058
rect 3461 -2064 3519 -2058
rect 3579 -2064 3637 -2058
rect 3697 -2064 3755 -2058
rect 3815 -2064 3873 -2058
rect 3933 -2064 3991 -2058
rect 4051 -2064 4109 -2058
rect 4169 -2064 4227 -2058
rect 4287 -2064 4345 -2058
rect 4405 -2064 4463 -2058
rect 4523 -2064 4581 -2058
rect 4641 -2064 4699 -2058
rect 4759 -2064 4817 -2058
rect 4877 -2064 4935 -2058
rect 4995 -2064 5053 -2058
rect 5113 -2064 5171 -2058
rect 5231 -2064 5289 -2058
rect 5349 -2064 5407 -2058
rect 5467 -2064 5525 -2058
rect 5585 -2064 5643 -2058
rect 5703 -2064 5761 -2058
rect 5821 -2064 5879 -2058
rect 5939 -2064 5997 -2058
rect 6057 -2064 6115 -2058
rect 6175 -2064 6233 -2058
rect 6293 -2064 6351 -2058
rect 6411 -2064 6469 -2058
rect 6529 -2064 6587 -2058
rect 6647 -2064 6705 -2058
rect 6765 -2064 6823 -2058
rect 6883 -2064 6941 -2058
rect 7001 -2064 7059 -2058
rect 7119 -2064 7177 -2058
rect 1176 -2758 1210 -2520
rect 1290 -2693 1324 -2661
rect 1408 -2693 1442 -2661
rect 1526 -2693 1560 -2661
rect 1644 -2693 1678 -2661
rect 1762 -2693 1796 -2661
rect 1880 -2693 1914 -2661
rect 1998 -2693 2032 -2661
rect 2116 -2693 2150 -2661
rect 2234 -2693 2268 -2661
rect 2352 -2693 2386 -2661
rect 2470 -2693 2504 -2661
rect 2588 -2693 2622 -2661
rect 2706 -2693 2740 -2661
rect 2824 -2693 2858 -2661
rect 2942 -2693 2976 -2661
rect 3060 -2693 3094 -2661
rect 3178 -2693 3212 -2661
rect 3296 -2693 3330 -2661
rect 3414 -2693 3448 -2661
rect 3532 -2693 3566 -2661
rect 3650 -2693 3684 -2661
rect 3768 -2693 3802 -2661
rect 3886 -2693 3920 -2661
rect 4004 -2693 4038 -2661
rect 4122 -2693 4156 -2661
rect 4240 -2693 4274 -2661
rect 4358 -2693 4392 -2661
rect 4476 -2693 4510 -2661
rect 4594 -2693 4628 -2661
rect 4712 -2693 4746 -2661
rect 4830 -2693 4864 -2661
rect 4948 -2693 4982 -2661
rect 5066 -2693 5100 -2661
rect 5184 -2693 5218 -2661
rect 5302 -2693 5336 -2661
rect 5420 -2693 5454 -2661
rect 5538 -2693 5572 -2661
rect 5656 -2693 5690 -2661
rect 5774 -2693 5808 -2661
rect 5892 -2693 5926 -2661
rect 6010 -2693 6044 -2661
rect 6128 -2693 6162 -2661
rect 6246 -2693 6280 -2661
rect 6364 -2693 6398 -2661
rect 6482 -2693 6516 -2661
rect 6600 -2693 6634 -2661
rect 6718 -2693 6752 -2661
rect 6836 -2693 6870 -2661
rect 6954 -2693 6988 -2661
rect 7072 -2693 7106 -2661
rect 7190 -2693 7224 -2661
rect 1278 -2705 7236 -2695
rect 1336 -2714 1396 -2705
rect 1454 -2714 1514 -2705
rect 1572 -2714 1632 -2705
rect 1690 -2714 1750 -2705
rect 1808 -2714 1868 -2705
rect 1926 -2714 1986 -2705
rect 2044 -2714 2104 -2705
rect 2162 -2714 2222 -2705
rect 2280 -2714 2340 -2705
rect 2398 -2714 2458 -2705
rect 2516 -2714 2576 -2705
rect 2634 -2714 2694 -2705
rect 2752 -2714 2812 -2705
rect 2870 -2714 2930 -2705
rect 2988 -2714 3048 -2705
rect 3106 -2714 3166 -2705
rect 3224 -2714 3284 -2705
rect 3342 -2714 3402 -2705
rect 3460 -2714 3520 -2705
rect 3578 -2714 3638 -2705
rect 3696 -2714 3756 -2705
rect 3814 -2714 3874 -2705
rect 3932 -2714 3992 -2705
rect 4050 -2714 4110 -2705
rect 4168 -2714 4228 -2705
rect 4286 -2714 4346 -2705
rect 4404 -2714 4464 -2705
rect 4522 -2714 4582 -2705
rect 4640 -2714 4700 -2705
rect 4758 -2714 4818 -2705
rect 4876 -2714 4936 -2705
rect 4994 -2714 5054 -2705
rect 5112 -2714 5172 -2705
rect 5230 -2714 5290 -2705
rect 5348 -2714 5408 -2705
rect 5466 -2714 5526 -2705
rect 5584 -2714 5644 -2705
rect 5702 -2714 5762 -2705
rect 5820 -2714 5880 -2705
rect 5938 -2714 5998 -2705
rect 6056 -2714 6116 -2705
rect 6174 -2714 6234 -2705
rect 6292 -2714 6352 -2705
rect 6410 -2714 6470 -2705
rect 6528 -2714 6588 -2705
rect 6646 -2714 6706 -2705
rect 6764 -2714 6824 -2705
rect 6882 -2714 6942 -2705
rect 7000 -2714 7060 -2705
rect 7118 -2714 7178 -2705
rect 1311 -2718 1421 -2714
rect 1429 -2718 1539 -2714
rect 1547 -2718 1657 -2714
rect 1665 -2718 1775 -2714
rect 1783 -2718 1893 -2714
rect 1901 -2718 2011 -2714
rect 2019 -2718 2129 -2714
rect 2137 -2718 2247 -2714
rect 2255 -2718 2365 -2714
rect 2373 -2718 2483 -2714
rect 2491 -2718 2601 -2714
rect 2609 -2718 2719 -2714
rect 2727 -2718 2837 -2714
rect 2845 -2718 2955 -2714
rect 2963 -2718 3073 -2714
rect 3081 -2718 3191 -2714
rect 3199 -2718 3309 -2714
rect 3317 -2718 3427 -2714
rect 3435 -2718 3545 -2714
rect 3553 -2718 3663 -2714
rect 3671 -2718 3781 -2714
rect 3789 -2718 3899 -2714
rect 3907 -2718 4017 -2714
rect 4025 -2718 4135 -2714
rect 4143 -2718 4253 -2714
rect 4261 -2718 4371 -2714
rect 4379 -2718 4489 -2714
rect 4497 -2718 4607 -2714
rect 4615 -2718 4725 -2714
rect 4733 -2718 4843 -2714
rect 4851 -2718 4961 -2714
rect 4969 -2718 5079 -2714
rect 5087 -2718 5197 -2714
rect 5205 -2718 5315 -2714
rect 5323 -2718 5433 -2714
rect 5441 -2718 5551 -2714
rect 5559 -2718 5669 -2714
rect 5677 -2718 5787 -2714
rect 5795 -2718 5905 -2714
rect 5913 -2718 6023 -2714
rect 6031 -2718 6141 -2714
rect 6149 -2718 6259 -2714
rect 6267 -2718 6377 -2714
rect 6385 -2718 6495 -2714
rect 6503 -2718 6613 -2714
rect 6621 -2718 6731 -2714
rect 6739 -2718 6849 -2714
rect 6857 -2718 6967 -2714
rect 6975 -2718 7085 -2714
rect 7093 -2718 7203 -2714
rect 1299 -2729 7215 -2718
rect 1386 -2752 1399 -2739
rect 1504 -2752 1517 -2739
rect 1622 -2752 1635 -2739
rect 1740 -2752 1753 -2739
rect 1858 -2752 1871 -2739
rect 1976 -2752 1989 -2739
rect 2094 -2752 2107 -2739
rect 2212 -2752 2225 -2739
rect 2330 -2752 2343 -2739
rect 2448 -2752 2461 -2739
rect 2566 -2752 2579 -2739
rect 2684 -2752 2697 -2739
rect 2802 -2752 2815 -2739
rect 2920 -2752 2933 -2739
rect 3038 -2752 3051 -2739
rect 3156 -2752 3169 -2739
rect 3274 -2752 3287 -2739
rect 3392 -2752 3405 -2739
rect 3510 -2752 3523 -2739
rect 3628 -2752 3641 -2739
rect 3746 -2752 3759 -2739
rect 3864 -2752 3877 -2739
rect 3982 -2752 3995 -2739
rect 4100 -2752 4113 -2739
rect 4218 -2752 4231 -2739
rect 4336 -2752 4349 -2739
rect 4454 -2752 4467 -2739
rect 4572 -2752 4585 -2739
rect 4690 -2752 4703 -2739
rect 4808 -2752 4821 -2739
rect 4926 -2752 4939 -2739
rect 5044 -2752 5057 -2739
rect 5162 -2752 5175 -2739
rect 5280 -2752 5293 -2739
rect 5398 -2752 5411 -2739
rect 5516 -2752 5529 -2739
rect 5634 -2752 5647 -2739
rect 5752 -2752 5765 -2739
rect 5870 -2752 5883 -2739
rect 5988 -2752 6001 -2739
rect 6106 -2752 6119 -2739
rect 6224 -2752 6237 -2739
rect 6342 -2752 6355 -2739
rect 6460 -2752 6473 -2739
rect 6578 -2752 6591 -2739
rect 6696 -2752 6709 -2739
rect 6814 -2752 6827 -2739
rect 6932 -2752 6945 -2739
rect 7050 -2752 7063 -2739
rect 1153 -2792 1210 -2758
rect 1333 -2786 1399 -2752
rect 1153 -4401 1187 -2792
rect 1428 -2797 1441 -2781
rect 1451 -2786 1517 -2752
rect 1546 -2797 1559 -2781
rect 1569 -2786 1635 -2752
rect 1664 -2797 1677 -2781
rect 1687 -2786 1753 -2752
rect 1782 -2797 1795 -2781
rect 1805 -2786 1871 -2752
rect 1900 -2797 1913 -2781
rect 1923 -2786 1989 -2752
rect 2018 -2797 2031 -2781
rect 2041 -2786 2107 -2752
rect 2136 -2797 2149 -2781
rect 2159 -2786 2225 -2752
rect 2254 -2797 2267 -2781
rect 2277 -2786 2343 -2752
rect 2372 -2797 2385 -2781
rect 2395 -2786 2461 -2752
rect 2490 -2797 2503 -2781
rect 2513 -2786 2579 -2752
rect 2608 -2797 2621 -2781
rect 2631 -2786 2697 -2752
rect 2726 -2797 2739 -2781
rect 2749 -2786 2815 -2752
rect 2844 -2797 2857 -2781
rect 2867 -2786 2933 -2752
rect 2962 -2797 2975 -2781
rect 2985 -2786 3051 -2752
rect 3080 -2797 3093 -2781
rect 3103 -2786 3169 -2752
rect 3198 -2797 3211 -2781
rect 3221 -2786 3287 -2752
rect 3316 -2797 3329 -2781
rect 3339 -2786 3405 -2752
rect 3434 -2797 3447 -2781
rect 3457 -2786 3523 -2752
rect 3552 -2797 3565 -2781
rect 3575 -2786 3641 -2752
rect 3670 -2797 3683 -2781
rect 3693 -2786 3759 -2752
rect 3788 -2797 3801 -2781
rect 3811 -2786 3877 -2752
rect 3906 -2797 3919 -2781
rect 3929 -2786 3995 -2752
rect 4024 -2797 4037 -2781
rect 4047 -2786 4113 -2752
rect 4142 -2797 4155 -2781
rect 4165 -2786 4231 -2752
rect 4260 -2797 4273 -2781
rect 4283 -2786 4349 -2752
rect 4378 -2797 4391 -2781
rect 4401 -2786 4467 -2752
rect 4496 -2797 4509 -2781
rect 4519 -2786 4585 -2752
rect 4614 -2797 4627 -2781
rect 4637 -2786 4703 -2752
rect 4732 -2797 4745 -2781
rect 4755 -2786 4821 -2752
rect 4850 -2797 4863 -2781
rect 4873 -2786 4939 -2752
rect 4968 -2797 4981 -2781
rect 4991 -2786 5057 -2752
rect 5086 -2797 5099 -2781
rect 5109 -2786 5175 -2752
rect 5204 -2797 5217 -2781
rect 5227 -2786 5293 -2752
rect 5322 -2797 5335 -2781
rect 5345 -2786 5411 -2752
rect 5440 -2797 5453 -2781
rect 5463 -2786 5529 -2752
rect 5558 -2797 5571 -2781
rect 5581 -2786 5647 -2752
rect 5676 -2797 5689 -2781
rect 5699 -2786 5765 -2752
rect 5794 -2797 5807 -2781
rect 5817 -2786 5883 -2752
rect 5912 -2797 5925 -2781
rect 5935 -2786 6001 -2752
rect 6030 -2797 6043 -2781
rect 6053 -2786 6119 -2752
rect 6148 -2797 6161 -2781
rect 6171 -2786 6237 -2752
rect 6266 -2797 6279 -2781
rect 6289 -2786 6355 -2752
rect 6384 -2797 6397 -2781
rect 6407 -2786 6473 -2752
rect 6502 -2797 6515 -2781
rect 6525 -2786 6591 -2752
rect 6620 -2797 6633 -2781
rect 6643 -2786 6709 -2752
rect 6738 -2797 6751 -2781
rect 6761 -2786 6827 -2752
rect 6856 -2797 6869 -2781
rect 6879 -2786 6945 -2752
rect 6974 -2797 6987 -2781
rect 6997 -2786 7063 -2752
rect 7092 -2797 7105 -2781
rect 7115 -2786 7181 -2752
rect 7304 -2758 7338 -1182
rect 9491 -2006 9549 -2000
rect 9491 -2040 9503 -2006
rect 9491 -2046 9549 -2040
rect 9491 -2434 9549 -2428
rect 9491 -2468 9503 -2434
rect 9491 -2474 9549 -2468
rect 9491 -2542 9549 -2536
rect 9491 -2576 9503 -2542
rect 9491 -2582 9549 -2576
rect 7281 -2792 7338 -2758
rect 1310 -2831 1376 -2797
rect 1428 -2831 1494 -2797
rect 1546 -2831 1612 -2797
rect 1664 -2831 1730 -2797
rect 1782 -2831 1848 -2797
rect 1900 -2831 1966 -2797
rect 2018 -2831 2084 -2797
rect 2136 -2831 2202 -2797
rect 2254 -2831 2320 -2797
rect 2372 -2831 2438 -2797
rect 2490 -2831 2556 -2797
rect 2608 -2831 2674 -2797
rect 2726 -2831 2792 -2797
rect 2844 -2831 2910 -2797
rect 2962 -2831 3028 -2797
rect 3080 -2831 3146 -2797
rect 3198 -2831 3264 -2797
rect 3316 -2831 3382 -2797
rect 3434 -2831 3500 -2797
rect 3552 -2831 3618 -2797
rect 3670 -2831 3736 -2797
rect 3788 -2831 3854 -2797
rect 3906 -2831 3972 -2797
rect 4024 -2831 4090 -2797
rect 4142 -2831 4208 -2797
rect 4260 -2831 4326 -2797
rect 4378 -2831 4444 -2797
rect 4496 -2831 4562 -2797
rect 4614 -2831 4680 -2797
rect 4732 -2831 4798 -2797
rect 4850 -2831 4916 -2797
rect 4968 -2831 5034 -2797
rect 5086 -2831 5152 -2797
rect 5204 -2831 5270 -2797
rect 5322 -2831 5388 -2797
rect 5440 -2831 5506 -2797
rect 5558 -2831 5624 -2797
rect 5676 -2831 5742 -2797
rect 5794 -2831 5860 -2797
rect 5912 -2831 5978 -2797
rect 6030 -2831 6096 -2797
rect 6148 -2831 6214 -2797
rect 6266 -2831 6332 -2797
rect 6384 -2831 6450 -2797
rect 6502 -2831 6568 -2797
rect 6620 -2831 6686 -2797
rect 6738 -2831 6804 -2797
rect 6856 -2831 6922 -2797
rect 6974 -2831 7040 -2797
rect 7092 -2831 7158 -2797
rect 1276 -2856 7192 -2854
rect 1272 -2878 7235 -2856
rect 1255 -2888 7235 -2878
rect 1314 -3525 1372 -3519
rect 1432 -3525 1490 -3519
rect 1550 -3525 1608 -3519
rect 1668 -3525 1726 -3519
rect 1786 -3525 1844 -3519
rect 1904 -3525 1962 -3519
rect 2022 -3525 2080 -3519
rect 2140 -3525 2198 -3519
rect 2258 -3525 2316 -3519
rect 2376 -3525 2434 -3519
rect 2494 -3525 2552 -3519
rect 2612 -3525 2670 -3519
rect 2730 -3525 2788 -3519
rect 2848 -3525 2906 -3519
rect 2966 -3525 3024 -3519
rect 3084 -3525 3142 -3519
rect 3202 -3525 3260 -3519
rect 3320 -3525 3378 -3519
rect 3438 -3525 3496 -3519
rect 3556 -3525 3614 -3519
rect 3674 -3525 3732 -3519
rect 3792 -3525 3850 -3519
rect 3910 -3525 3968 -3519
rect 4028 -3525 4086 -3519
rect 4146 -3525 4204 -3519
rect 4264 -3525 4322 -3519
rect 4382 -3525 4440 -3519
rect 4500 -3525 4558 -3519
rect 4618 -3525 4676 -3519
rect 4736 -3525 4794 -3519
rect 4854 -3525 4912 -3519
rect 4972 -3525 5030 -3519
rect 5090 -3525 5148 -3519
rect 5208 -3525 5266 -3519
rect 5326 -3525 5384 -3519
rect 5444 -3525 5502 -3519
rect 5562 -3525 5620 -3519
rect 5680 -3525 5738 -3519
rect 5798 -3525 5856 -3519
rect 5916 -3525 5974 -3519
rect 6034 -3525 6092 -3519
rect 6152 -3525 6210 -3519
rect 6270 -3525 6328 -3519
rect 6388 -3525 6446 -3519
rect 6506 -3525 6564 -3519
rect 6624 -3525 6682 -3519
rect 6742 -3525 6800 -3519
rect 6860 -3525 6918 -3519
rect 6978 -3525 7036 -3519
rect 7096 -3525 7154 -3519
rect 1314 -3559 1326 -3525
rect 1432 -3559 1444 -3525
rect 1550 -3559 1562 -3525
rect 1668 -3559 1680 -3525
rect 1786 -3559 1798 -3525
rect 1904 -3559 1916 -3525
rect 2022 -3559 2034 -3525
rect 2140 -3559 2152 -3525
rect 2258 -3559 2270 -3525
rect 2376 -3559 2388 -3525
rect 2494 -3559 2506 -3525
rect 2612 -3559 2624 -3525
rect 2730 -3559 2742 -3525
rect 2848 -3559 2860 -3525
rect 2966 -3559 2978 -3525
rect 3084 -3559 3096 -3525
rect 3202 -3559 3214 -3525
rect 3320 -3559 3332 -3525
rect 3438 -3559 3450 -3525
rect 3556 -3559 3568 -3525
rect 3674 -3559 3686 -3525
rect 3792 -3559 3804 -3525
rect 3910 -3559 3922 -3525
rect 4028 -3559 4040 -3525
rect 4146 -3559 4158 -3525
rect 4264 -3559 4276 -3525
rect 4382 -3559 4394 -3525
rect 4500 -3559 4512 -3525
rect 4618 -3559 4630 -3525
rect 4736 -3559 4748 -3525
rect 4854 -3559 4866 -3525
rect 4972 -3559 4984 -3525
rect 5090 -3559 5102 -3525
rect 5208 -3559 5220 -3525
rect 5326 -3559 5338 -3525
rect 5444 -3559 5456 -3525
rect 5562 -3559 5574 -3525
rect 5680 -3559 5692 -3525
rect 5798 -3559 5810 -3525
rect 5916 -3559 5928 -3525
rect 6034 -3559 6046 -3525
rect 6152 -3559 6164 -3525
rect 6270 -3559 6282 -3525
rect 6388 -3559 6400 -3525
rect 6506 -3559 6518 -3525
rect 6624 -3559 6636 -3525
rect 6742 -3559 6754 -3525
rect 6860 -3559 6872 -3525
rect 6978 -3559 6990 -3525
rect 7096 -3559 7108 -3525
rect 1314 -3565 1372 -3559
rect 1432 -3565 1490 -3559
rect 1550 -3565 1608 -3559
rect 1668 -3565 1726 -3559
rect 1786 -3565 1844 -3559
rect 1904 -3565 1962 -3559
rect 2022 -3565 2080 -3559
rect 2140 -3565 2198 -3559
rect 2258 -3565 2316 -3559
rect 2376 -3565 2434 -3559
rect 2494 -3565 2552 -3559
rect 2612 -3565 2670 -3559
rect 2730 -3565 2788 -3559
rect 2848 -3565 2906 -3559
rect 2966 -3565 3024 -3559
rect 3084 -3565 3142 -3559
rect 3202 -3565 3260 -3559
rect 3320 -3565 3378 -3559
rect 3438 -3565 3496 -3559
rect 3556 -3565 3614 -3559
rect 3674 -3565 3732 -3559
rect 3792 -3565 3850 -3559
rect 3910 -3565 3968 -3559
rect 4028 -3565 4086 -3559
rect 4146 -3565 4204 -3559
rect 4264 -3565 4322 -3559
rect 4382 -3565 4440 -3559
rect 4500 -3565 4558 -3559
rect 4618 -3565 4676 -3559
rect 4736 -3565 4794 -3559
rect 4854 -3565 4912 -3559
rect 4972 -3565 5030 -3559
rect 5090 -3565 5148 -3559
rect 5208 -3565 5266 -3559
rect 5326 -3565 5384 -3559
rect 5444 -3565 5502 -3559
rect 5562 -3565 5620 -3559
rect 5680 -3565 5738 -3559
rect 5798 -3565 5856 -3559
rect 5916 -3565 5974 -3559
rect 6034 -3565 6092 -3559
rect 6152 -3565 6210 -3559
rect 6270 -3565 6328 -3559
rect 6388 -3565 6446 -3559
rect 6506 -3565 6564 -3559
rect 6624 -3565 6682 -3559
rect 6742 -3565 6800 -3559
rect 6860 -3565 6918 -3559
rect 6978 -3565 7036 -3559
rect 7096 -3565 7154 -3559
rect 1314 -3633 1372 -3627
rect 1432 -3633 1490 -3627
rect 1550 -3633 1608 -3627
rect 1668 -3633 1726 -3627
rect 1786 -3633 1844 -3627
rect 1904 -3633 1962 -3627
rect 2022 -3633 2080 -3627
rect 2140 -3633 2198 -3627
rect 2258 -3633 2316 -3627
rect 2376 -3633 2434 -3627
rect 2494 -3633 2552 -3627
rect 2612 -3633 2670 -3627
rect 2730 -3633 2788 -3627
rect 2848 -3633 2906 -3627
rect 2966 -3633 3024 -3627
rect 3084 -3633 3142 -3627
rect 3202 -3633 3260 -3627
rect 3320 -3633 3378 -3627
rect 3438 -3633 3496 -3627
rect 3556 -3633 3614 -3627
rect 3674 -3633 3732 -3627
rect 3792 -3633 3850 -3627
rect 3910 -3633 3968 -3627
rect 4028 -3633 4086 -3627
rect 4146 -3633 4204 -3627
rect 4264 -3633 4322 -3627
rect 4382 -3633 4440 -3627
rect 4500 -3633 4558 -3627
rect 4618 -3633 4676 -3627
rect 4736 -3633 4794 -3627
rect 4854 -3633 4912 -3627
rect 4972 -3633 5030 -3627
rect 5090 -3633 5148 -3627
rect 5208 -3633 5266 -3627
rect 5326 -3633 5384 -3627
rect 5444 -3633 5502 -3627
rect 5562 -3633 5620 -3627
rect 5680 -3633 5738 -3627
rect 5798 -3633 5856 -3627
rect 5916 -3633 5974 -3627
rect 6034 -3633 6092 -3627
rect 6152 -3633 6210 -3627
rect 6270 -3633 6328 -3627
rect 6388 -3633 6446 -3627
rect 6506 -3633 6564 -3627
rect 6624 -3633 6682 -3627
rect 6742 -3633 6800 -3627
rect 6860 -3633 6918 -3627
rect 6978 -3633 7036 -3627
rect 7096 -3633 7154 -3627
rect 1314 -3667 1326 -3633
rect 1432 -3667 1444 -3633
rect 1550 -3667 1562 -3633
rect 1668 -3667 1680 -3633
rect 1786 -3667 1798 -3633
rect 1904 -3667 1916 -3633
rect 2022 -3667 2034 -3633
rect 2140 -3667 2152 -3633
rect 2258 -3667 2270 -3633
rect 2376 -3667 2388 -3633
rect 2494 -3667 2506 -3633
rect 2612 -3667 2624 -3633
rect 2730 -3667 2742 -3633
rect 2848 -3667 2860 -3633
rect 2966 -3667 2978 -3633
rect 3084 -3667 3096 -3633
rect 3202 -3667 3214 -3633
rect 3320 -3667 3332 -3633
rect 3438 -3667 3450 -3633
rect 3556 -3667 3568 -3633
rect 3674 -3667 3686 -3633
rect 3792 -3667 3804 -3633
rect 3910 -3667 3922 -3633
rect 4028 -3667 4040 -3633
rect 4146 -3667 4158 -3633
rect 4264 -3667 4276 -3633
rect 4382 -3667 4394 -3633
rect 4500 -3667 4512 -3633
rect 4618 -3667 4630 -3633
rect 4736 -3667 4748 -3633
rect 4854 -3667 4866 -3633
rect 4972 -3667 4984 -3633
rect 5090 -3667 5102 -3633
rect 5208 -3667 5220 -3633
rect 5326 -3667 5338 -3633
rect 5444 -3667 5456 -3633
rect 5562 -3667 5574 -3633
rect 5680 -3667 5692 -3633
rect 5798 -3667 5810 -3633
rect 5916 -3667 5928 -3633
rect 6034 -3667 6046 -3633
rect 6152 -3667 6164 -3633
rect 6270 -3667 6282 -3633
rect 6388 -3667 6400 -3633
rect 6506 -3667 6518 -3633
rect 6624 -3667 6636 -3633
rect 6742 -3667 6754 -3633
rect 6860 -3667 6872 -3633
rect 6978 -3667 6990 -3633
rect 7096 -3667 7108 -3633
rect 1314 -3673 1372 -3667
rect 1432 -3673 1490 -3667
rect 1550 -3673 1608 -3667
rect 1668 -3673 1726 -3667
rect 1786 -3673 1844 -3667
rect 1904 -3673 1962 -3667
rect 2022 -3673 2080 -3667
rect 2140 -3673 2198 -3667
rect 2258 -3673 2316 -3667
rect 2376 -3673 2434 -3667
rect 2494 -3673 2552 -3667
rect 2612 -3673 2670 -3667
rect 2730 -3673 2788 -3667
rect 2848 -3673 2906 -3667
rect 2966 -3673 3024 -3667
rect 3084 -3673 3142 -3667
rect 3202 -3673 3260 -3667
rect 3320 -3673 3378 -3667
rect 3438 -3673 3496 -3667
rect 3556 -3673 3614 -3667
rect 3674 -3673 3732 -3667
rect 3792 -3673 3850 -3667
rect 3910 -3673 3968 -3667
rect 4028 -3673 4086 -3667
rect 4146 -3673 4204 -3667
rect 4264 -3673 4322 -3667
rect 4382 -3673 4440 -3667
rect 4500 -3673 4558 -3667
rect 4618 -3673 4676 -3667
rect 4736 -3673 4794 -3667
rect 4854 -3673 4912 -3667
rect 4972 -3673 5030 -3667
rect 5090 -3673 5148 -3667
rect 5208 -3673 5266 -3667
rect 5326 -3673 5384 -3667
rect 5444 -3673 5502 -3667
rect 5562 -3673 5620 -3667
rect 5680 -3673 5738 -3667
rect 5798 -3673 5856 -3667
rect 5916 -3673 5974 -3667
rect 6034 -3673 6092 -3667
rect 6152 -3673 6210 -3667
rect 6270 -3673 6328 -3667
rect 6388 -3673 6446 -3667
rect 6506 -3673 6564 -3667
rect 6624 -3673 6682 -3667
rect 6742 -3673 6800 -3667
rect 6860 -3673 6918 -3667
rect 6978 -3673 7036 -3667
rect 7096 -3673 7154 -3667
rect 1314 -4361 1372 -4355
rect 1432 -4361 1490 -4355
rect 1550 -4361 1608 -4355
rect 1668 -4361 1726 -4355
rect 1786 -4361 1844 -4355
rect 1904 -4361 1962 -4355
rect 2022 -4361 2080 -4355
rect 2140 -4361 2198 -4355
rect 2258 -4361 2316 -4355
rect 2376 -4361 2434 -4355
rect 2494 -4361 2552 -4355
rect 2612 -4361 2670 -4355
rect 2730 -4361 2788 -4355
rect 2848 -4361 2906 -4355
rect 2966 -4361 3024 -4355
rect 3084 -4361 3142 -4355
rect 3202 -4361 3260 -4355
rect 3320 -4361 3378 -4355
rect 3438 -4361 3496 -4355
rect 3556 -4361 3614 -4355
rect 3674 -4361 3732 -4355
rect 3792 -4361 3850 -4355
rect 3910 -4361 3968 -4355
rect 4028 -4361 4086 -4355
rect 4146 -4361 4204 -4355
rect 4264 -4361 4322 -4355
rect 4382 -4361 4440 -4355
rect 4500 -4361 4558 -4355
rect 4618 -4361 4676 -4355
rect 4736 -4361 4794 -4355
rect 4854 -4361 4912 -4355
rect 4972 -4361 5030 -4355
rect 5090 -4361 5148 -4355
rect 5208 -4361 5266 -4355
rect 5326 -4361 5384 -4355
rect 5444 -4361 5502 -4355
rect 5562 -4361 5620 -4355
rect 5680 -4361 5738 -4355
rect 5798 -4361 5856 -4355
rect 5916 -4361 5974 -4355
rect 6034 -4361 6092 -4355
rect 6152 -4361 6210 -4355
rect 6270 -4361 6328 -4355
rect 6388 -4361 6446 -4355
rect 6506 -4361 6564 -4355
rect 6624 -4361 6682 -4355
rect 6742 -4361 6800 -4355
rect 6860 -4361 6918 -4355
rect 6978 -4361 7036 -4355
rect 7096 -4361 7154 -4355
rect 1314 -4395 1326 -4361
rect 1432 -4395 1444 -4361
rect 1550 -4395 1562 -4361
rect 1668 -4395 1680 -4361
rect 1786 -4395 1798 -4361
rect 1904 -4395 1916 -4361
rect 2022 -4395 2034 -4361
rect 2140 -4395 2152 -4361
rect 2258 -4395 2270 -4361
rect 2376 -4395 2388 -4361
rect 2494 -4395 2506 -4361
rect 2612 -4395 2624 -4361
rect 2730 -4395 2742 -4361
rect 2848 -4395 2860 -4361
rect 2966 -4395 2978 -4361
rect 3084 -4395 3096 -4361
rect 3202 -4395 3214 -4361
rect 3320 -4395 3332 -4361
rect 3438 -4395 3450 -4361
rect 3556 -4395 3568 -4361
rect 3674 -4395 3686 -4361
rect 3792 -4395 3804 -4361
rect 3910 -4395 3922 -4361
rect 4028 -4395 4040 -4361
rect 4146 -4395 4158 -4361
rect 4264 -4395 4276 -4361
rect 4382 -4395 4394 -4361
rect 4500 -4395 4512 -4361
rect 4618 -4395 4630 -4361
rect 4736 -4395 4748 -4361
rect 4854 -4395 4866 -4361
rect 4972 -4395 4984 -4361
rect 5090 -4395 5102 -4361
rect 5208 -4395 5220 -4361
rect 5326 -4395 5338 -4361
rect 5444 -4395 5456 -4361
rect 5562 -4395 5574 -4361
rect 5680 -4395 5692 -4361
rect 5798 -4395 5810 -4361
rect 5916 -4395 5928 -4361
rect 6034 -4395 6046 -4361
rect 6152 -4395 6164 -4361
rect 6270 -4395 6282 -4361
rect 6388 -4395 6400 -4361
rect 6506 -4395 6518 -4361
rect 6624 -4395 6636 -4361
rect 6742 -4395 6754 -4361
rect 6860 -4395 6872 -4361
rect 6978 -4395 6990 -4361
rect 7096 -4395 7108 -4361
rect 1314 -4401 1372 -4395
rect 1432 -4401 1490 -4395
rect 1550 -4401 1608 -4395
rect 1668 -4401 1726 -4395
rect 1786 -4401 1844 -4395
rect 1904 -4401 1962 -4395
rect 2022 -4401 2080 -4395
rect 2140 -4401 2198 -4395
rect 2258 -4401 2316 -4395
rect 2376 -4401 2434 -4395
rect 2494 -4401 2552 -4395
rect 2612 -4401 2670 -4395
rect 2730 -4401 2788 -4395
rect 2848 -4401 2906 -4395
rect 2966 -4401 3024 -4395
rect 3084 -4401 3142 -4395
rect 3202 -4401 3260 -4395
rect 3320 -4401 3378 -4395
rect 3438 -4401 3496 -4395
rect 3556 -4401 3614 -4395
rect 3674 -4401 3732 -4395
rect 3792 -4401 3850 -4395
rect 3910 -4401 3968 -4395
rect 4028 -4401 4086 -4395
rect 4146 -4401 4204 -4395
rect 4264 -4401 4322 -4395
rect 4382 -4401 4440 -4395
rect 4500 -4401 4558 -4395
rect 4618 -4401 4676 -4395
rect 4736 -4401 4794 -4395
rect 4854 -4401 4912 -4395
rect 4972 -4401 5030 -4395
rect 5090 -4401 5148 -4395
rect 5208 -4401 5266 -4395
rect 5326 -4401 5384 -4395
rect 5444 -4401 5502 -4395
rect 5562 -4401 5620 -4395
rect 5680 -4401 5738 -4395
rect 5798 -4401 5856 -4395
rect 5916 -4401 5974 -4395
rect 6034 -4401 6092 -4395
rect 6152 -4401 6210 -4395
rect 6270 -4401 6328 -4395
rect 6388 -4401 6446 -4395
rect 6506 -4401 6564 -4395
rect 6624 -4401 6682 -4395
rect 6742 -4401 6800 -4395
rect 6860 -4401 6918 -4395
rect 6978 -4401 7036 -4395
rect 7096 -4401 7154 -4395
rect 7281 -4401 7315 -2792
rect 9491 -2970 9549 -2964
rect 9491 -3004 9503 -2970
rect 9491 -3010 9549 -3004
rect 1249 -4497 7219 -4443
rect 1314 -4545 1372 -4539
rect 1432 -4545 1490 -4539
rect 1550 -4545 1608 -4539
rect 1668 -4545 1726 -4539
rect 1786 -4545 1844 -4539
rect 1904 -4545 1962 -4539
rect 2022 -4545 2080 -4539
rect 2140 -4545 2198 -4539
rect 2258 -4545 2316 -4539
rect 2376 -4545 2434 -4539
rect 2494 -4545 2552 -4539
rect 2612 -4545 2670 -4539
rect 2730 -4545 2788 -4539
rect 2848 -4545 2906 -4539
rect 2966 -4545 3024 -4539
rect 3084 -4545 3142 -4539
rect 3202 -4545 3260 -4539
rect 3320 -4545 3378 -4539
rect 3438 -4545 3496 -4539
rect 3556 -4545 3614 -4539
rect 3674 -4545 3732 -4539
rect 3792 -4545 3850 -4539
rect 3910 -4545 3968 -4539
rect 4028 -4545 4086 -4539
rect 4146 -4545 4204 -4539
rect 4264 -4545 4322 -4539
rect 4382 -4545 4440 -4539
rect 4500 -4545 4558 -4539
rect 4618 -4545 4676 -4539
rect 4736 -4545 4794 -4539
rect 4854 -4545 4912 -4539
rect 4972 -4545 5030 -4539
rect 5090 -4545 5148 -4539
rect 5208 -4545 5266 -4539
rect 5326 -4545 5384 -4539
rect 5444 -4545 5502 -4539
rect 5562 -4545 5620 -4539
rect 5680 -4545 5738 -4539
rect 5798 -4545 5856 -4539
rect 5916 -4545 5974 -4539
rect 6034 -4545 6092 -4539
rect 6152 -4545 6210 -4539
rect 6270 -4545 6328 -4539
rect 6388 -4545 6446 -4539
rect 6506 -4545 6564 -4539
rect 6624 -4545 6682 -4539
rect 6742 -4545 6800 -4539
rect 6860 -4545 6918 -4539
rect 6978 -4545 7036 -4539
rect 7096 -4545 7154 -4539
rect 1314 -4579 1326 -4545
rect 1432 -4579 1444 -4545
rect 1550 -4579 1562 -4545
rect 1668 -4579 1680 -4545
rect 1786 -4579 1798 -4545
rect 1904 -4579 1916 -4545
rect 2022 -4579 2034 -4545
rect 2140 -4579 2152 -4545
rect 2258 -4579 2270 -4545
rect 2376 -4579 2388 -4545
rect 2494 -4579 2506 -4545
rect 2612 -4579 2624 -4545
rect 2730 -4579 2742 -4545
rect 2848 -4579 2860 -4545
rect 2966 -4579 2978 -4545
rect 3084 -4579 3096 -4545
rect 3202 -4579 3214 -4545
rect 3320 -4579 3332 -4545
rect 3438 -4579 3450 -4545
rect 3556 -4579 3568 -4545
rect 3674 -4579 3686 -4545
rect 3792 -4579 3804 -4545
rect 3910 -4579 3922 -4545
rect 4028 -4579 4040 -4545
rect 4146 -4579 4158 -4545
rect 4264 -4579 4276 -4545
rect 4382 -4579 4394 -4545
rect 4500 -4579 4512 -4545
rect 4618 -4579 4630 -4545
rect 4736 -4579 4748 -4545
rect 4854 -4579 4866 -4545
rect 4972 -4579 4984 -4545
rect 5090 -4579 5102 -4545
rect 5208 -4579 5220 -4545
rect 5326 -4579 5338 -4545
rect 5444 -4579 5456 -4545
rect 5562 -4579 5574 -4545
rect 5680 -4579 5692 -4545
rect 5798 -4579 5810 -4545
rect 5916 -4579 5928 -4545
rect 6034 -4579 6046 -4545
rect 6152 -4579 6164 -4545
rect 6270 -4579 6282 -4545
rect 6388 -4579 6400 -4545
rect 6506 -4579 6518 -4545
rect 6624 -4579 6636 -4545
rect 6742 -4579 6754 -4545
rect 6860 -4579 6872 -4545
rect 6978 -4579 6990 -4545
rect 7096 -4579 7108 -4545
rect 1314 -4585 1372 -4579
rect 1432 -4585 1490 -4579
rect 1550 -4585 1608 -4579
rect 1668 -4585 1726 -4579
rect 1786 -4585 1844 -4579
rect 1904 -4585 1962 -4579
rect 2022 -4585 2080 -4579
rect 2140 -4585 2198 -4579
rect 2258 -4585 2316 -4579
rect 2376 -4585 2434 -4579
rect 2494 -4585 2552 -4579
rect 2612 -4585 2670 -4579
rect 2730 -4585 2788 -4579
rect 2848 -4585 2906 -4579
rect 2966 -4585 3024 -4579
rect 3084 -4585 3142 -4579
rect 3202 -4585 3260 -4579
rect 3320 -4585 3378 -4579
rect 3438 -4585 3496 -4579
rect 3556 -4585 3614 -4579
rect 3674 -4585 3732 -4579
rect 3792 -4585 3850 -4579
rect 3910 -4585 3968 -4579
rect 4028 -4585 4086 -4579
rect 4146 -4585 4204 -4579
rect 4264 -4585 4322 -4579
rect 4382 -4585 4440 -4579
rect 4500 -4585 4558 -4579
rect 4618 -4585 4676 -4579
rect 4736 -4585 4794 -4579
rect 4854 -4585 4912 -4579
rect 4972 -4585 5030 -4579
rect 5090 -4585 5148 -4579
rect 5208 -4585 5266 -4579
rect 5326 -4585 5384 -4579
rect 5444 -4585 5502 -4579
rect 5562 -4585 5620 -4579
rect 5680 -4585 5738 -4579
rect 5798 -4585 5856 -4579
rect 5916 -4585 5974 -4579
rect 6034 -4585 6092 -4579
rect 6152 -4585 6210 -4579
rect 6270 -4585 6328 -4579
rect 6388 -4585 6446 -4579
rect 6506 -4585 6564 -4579
rect 6624 -4585 6682 -4579
rect 6742 -4585 6800 -4579
rect 6860 -4585 6918 -4579
rect 6978 -4585 7036 -4579
rect 7096 -4585 7154 -4579
rect 1314 -5273 1372 -5267
rect 1432 -5273 1490 -5267
rect 1550 -5273 1608 -5267
rect 1668 -5273 1726 -5267
rect 1786 -5273 1844 -5267
rect 1904 -5273 1962 -5267
rect 2022 -5273 2080 -5267
rect 2140 -5273 2198 -5267
rect 2258 -5273 2316 -5267
rect 2376 -5273 2434 -5267
rect 2494 -5273 2552 -5267
rect 2612 -5273 2670 -5267
rect 2730 -5273 2788 -5267
rect 2848 -5273 2906 -5267
rect 2966 -5273 3024 -5267
rect 3084 -5273 3142 -5267
rect 3202 -5273 3260 -5267
rect 3320 -5273 3378 -5267
rect 3438 -5273 3496 -5267
rect 3556 -5273 3614 -5267
rect 3674 -5273 3732 -5267
rect 3792 -5273 3850 -5267
rect 3910 -5273 3968 -5267
rect 4028 -5273 4086 -5267
rect 4146 -5273 4204 -5267
rect 4264 -5273 4322 -5267
rect 4382 -5273 4440 -5267
rect 4500 -5273 4558 -5267
rect 4618 -5273 4676 -5267
rect 4736 -5273 4794 -5267
rect 4854 -5273 4912 -5267
rect 4972 -5273 5030 -5267
rect 5090 -5273 5148 -5267
rect 5208 -5273 5266 -5267
rect 5326 -5273 5384 -5267
rect 5444 -5273 5502 -5267
rect 5562 -5273 5620 -5267
rect 5680 -5273 5738 -5267
rect 5798 -5273 5856 -5267
rect 5916 -5273 5974 -5267
rect 6034 -5273 6092 -5267
rect 6152 -5273 6210 -5267
rect 6270 -5273 6328 -5267
rect 6388 -5273 6446 -5267
rect 6506 -5273 6564 -5267
rect 6624 -5273 6682 -5267
rect 6742 -5273 6800 -5267
rect 6860 -5273 6918 -5267
rect 6978 -5273 7036 -5267
rect 7096 -5273 7154 -5267
rect 1314 -5307 1326 -5273
rect 1432 -5307 1444 -5273
rect 1550 -5307 1562 -5273
rect 1668 -5307 1680 -5273
rect 1786 -5307 1798 -5273
rect 1904 -5307 1916 -5273
rect 2022 -5307 2034 -5273
rect 2140 -5307 2152 -5273
rect 2258 -5307 2270 -5273
rect 2376 -5307 2388 -5273
rect 2494 -5307 2506 -5273
rect 2612 -5307 2624 -5273
rect 2730 -5307 2742 -5273
rect 2848 -5307 2860 -5273
rect 2966 -5307 2978 -5273
rect 3084 -5307 3096 -5273
rect 3202 -5307 3214 -5273
rect 3320 -5307 3332 -5273
rect 3438 -5307 3450 -5273
rect 3556 -5307 3568 -5273
rect 3674 -5307 3686 -5273
rect 3792 -5307 3804 -5273
rect 3910 -5307 3922 -5273
rect 4028 -5307 4040 -5273
rect 4146 -5307 4158 -5273
rect 4264 -5307 4276 -5273
rect 4382 -5307 4394 -5273
rect 4500 -5307 4512 -5273
rect 4618 -5307 4630 -5273
rect 4736 -5307 4748 -5273
rect 4854 -5307 4866 -5273
rect 4972 -5307 4984 -5273
rect 5090 -5307 5102 -5273
rect 5208 -5307 5220 -5273
rect 5326 -5307 5338 -5273
rect 5444 -5307 5456 -5273
rect 5562 -5307 5574 -5273
rect 5680 -5307 5692 -5273
rect 5798 -5307 5810 -5273
rect 5916 -5307 5928 -5273
rect 6034 -5307 6046 -5273
rect 6152 -5307 6164 -5273
rect 6270 -5307 6282 -5273
rect 6388 -5307 6400 -5273
rect 6506 -5307 6518 -5273
rect 6624 -5307 6636 -5273
rect 6742 -5307 6754 -5273
rect 6860 -5307 6872 -5273
rect 6978 -5307 6990 -5273
rect 7096 -5307 7108 -5273
rect 1314 -5313 1372 -5307
rect 1432 -5313 1490 -5307
rect 1550 -5313 1608 -5307
rect 1668 -5313 1726 -5307
rect 1786 -5313 1844 -5307
rect 1904 -5313 1962 -5307
rect 2022 -5313 2080 -5307
rect 2140 -5313 2198 -5307
rect 2258 -5313 2316 -5307
rect 2376 -5313 2434 -5307
rect 2494 -5313 2552 -5307
rect 2612 -5313 2670 -5307
rect 2730 -5313 2788 -5307
rect 2848 -5313 2906 -5307
rect 2966 -5313 3024 -5307
rect 3084 -5313 3142 -5307
rect 3202 -5313 3260 -5307
rect 3320 -5313 3378 -5307
rect 3438 -5313 3496 -5307
rect 3556 -5313 3614 -5307
rect 3674 -5313 3732 -5307
rect 3792 -5313 3850 -5307
rect 3910 -5313 3968 -5307
rect 4028 -5313 4086 -5307
rect 4146 -5313 4204 -5307
rect 4264 -5313 4322 -5307
rect 4382 -5313 4440 -5307
rect 4500 -5313 4558 -5307
rect 4618 -5313 4676 -5307
rect 4736 -5313 4794 -5307
rect 4854 -5313 4912 -5307
rect 4972 -5313 5030 -5307
rect 5090 -5313 5148 -5307
rect 5208 -5313 5266 -5307
rect 5326 -5313 5384 -5307
rect 5444 -5313 5502 -5307
rect 5562 -5313 5620 -5307
rect 5680 -5313 5738 -5307
rect 5798 -5313 5856 -5307
rect 5916 -5313 5974 -5307
rect 6034 -5313 6092 -5307
rect 6152 -5313 6210 -5307
rect 6270 -5313 6328 -5307
rect 6388 -5313 6446 -5307
rect 6506 -5313 6564 -5307
rect 6624 -5313 6682 -5307
rect 6742 -5313 6800 -5307
rect 6860 -5313 6918 -5307
rect 6978 -5313 7036 -5307
rect 7096 -5313 7154 -5307
rect 1314 -5381 1372 -5375
rect 1432 -5381 1490 -5375
rect 1550 -5381 1608 -5375
rect 1668 -5381 1726 -5375
rect 1786 -5381 1844 -5375
rect 1904 -5381 1962 -5375
rect 2022 -5381 2080 -5375
rect 2140 -5381 2198 -5375
rect 2258 -5381 2316 -5375
rect 2376 -5381 2434 -5375
rect 2494 -5381 2552 -5375
rect 2612 -5381 2670 -5375
rect 2730 -5381 2788 -5375
rect 2848 -5381 2906 -5375
rect 2966 -5381 3024 -5375
rect 3084 -5381 3142 -5375
rect 3202 -5381 3260 -5375
rect 3320 -5381 3378 -5375
rect 3438 -5381 3496 -5375
rect 3556 -5381 3614 -5375
rect 3674 -5381 3732 -5375
rect 3792 -5381 3850 -5375
rect 3910 -5381 3968 -5375
rect 4028 -5381 4086 -5375
rect 4146 -5381 4204 -5375
rect 4264 -5381 4322 -5375
rect 4382 -5381 4440 -5375
rect 4500 -5381 4558 -5375
rect 4618 -5381 4676 -5375
rect 4736 -5381 4794 -5375
rect 4854 -5381 4912 -5375
rect 4972 -5381 5030 -5375
rect 5090 -5381 5148 -5375
rect 5208 -5381 5266 -5375
rect 5326 -5381 5384 -5375
rect 5444 -5381 5502 -5375
rect 5562 -5381 5620 -5375
rect 5680 -5381 5738 -5375
rect 5798 -5381 5856 -5375
rect 5916 -5381 5974 -5375
rect 6034 -5381 6092 -5375
rect 6152 -5381 6210 -5375
rect 6270 -5381 6328 -5375
rect 6388 -5381 6446 -5375
rect 6506 -5381 6564 -5375
rect 6624 -5381 6682 -5375
rect 6742 -5381 6800 -5375
rect 6860 -5381 6918 -5375
rect 6978 -5381 7036 -5375
rect 7096 -5381 7154 -5375
rect 1314 -5415 1326 -5381
rect 1432 -5415 1444 -5381
rect 1550 -5415 1562 -5381
rect 1668 -5415 1680 -5381
rect 1786 -5415 1798 -5381
rect 1904 -5415 1916 -5381
rect 2022 -5415 2034 -5381
rect 2140 -5415 2152 -5381
rect 2258 -5415 2270 -5381
rect 2376 -5415 2388 -5381
rect 2494 -5415 2506 -5381
rect 2612 -5415 2624 -5381
rect 2730 -5415 2742 -5381
rect 2848 -5415 2860 -5381
rect 2966 -5415 2978 -5381
rect 3084 -5415 3096 -5381
rect 3202 -5415 3214 -5381
rect 3320 -5415 3332 -5381
rect 3438 -5415 3450 -5381
rect 3556 -5415 3568 -5381
rect 3674 -5415 3686 -5381
rect 3792 -5415 3804 -5381
rect 3910 -5415 3922 -5381
rect 4028 -5415 4040 -5381
rect 4146 -5415 4158 -5381
rect 4264 -5415 4276 -5381
rect 4382 -5415 4394 -5381
rect 4500 -5415 4512 -5381
rect 4618 -5415 4630 -5381
rect 4736 -5415 4748 -5381
rect 4854 -5415 4866 -5381
rect 4972 -5415 4984 -5381
rect 5090 -5415 5102 -5381
rect 5208 -5415 5220 -5381
rect 5326 -5415 5338 -5381
rect 5444 -5415 5456 -5381
rect 5562 -5415 5574 -5381
rect 5680 -5415 5692 -5381
rect 5798 -5415 5810 -5381
rect 5916 -5415 5928 -5381
rect 6034 -5415 6046 -5381
rect 6152 -5415 6164 -5381
rect 6270 -5415 6282 -5381
rect 6388 -5415 6400 -5381
rect 6506 -5415 6518 -5381
rect 6624 -5415 6636 -5381
rect 6742 -5415 6754 -5381
rect 6860 -5415 6872 -5381
rect 6978 -5415 6990 -5381
rect 7096 -5415 7108 -5381
rect 1314 -5421 1372 -5415
rect 1432 -5421 1490 -5415
rect 1550 -5421 1608 -5415
rect 1668 -5421 1726 -5415
rect 1786 -5421 1844 -5415
rect 1904 -5421 1962 -5415
rect 2022 -5421 2080 -5415
rect 2140 -5421 2198 -5415
rect 2258 -5421 2316 -5415
rect 2376 -5421 2434 -5415
rect 2494 -5421 2552 -5415
rect 2612 -5421 2670 -5415
rect 2730 -5421 2788 -5415
rect 2848 -5421 2906 -5415
rect 2966 -5421 3024 -5415
rect 3084 -5421 3142 -5415
rect 3202 -5421 3260 -5415
rect 3320 -5421 3378 -5415
rect 3438 -5421 3496 -5415
rect 3556 -5421 3614 -5415
rect 3674 -5421 3732 -5415
rect 3792 -5421 3850 -5415
rect 3910 -5421 3968 -5415
rect 4028 -5421 4086 -5415
rect 4146 -5421 4204 -5415
rect 4264 -5421 4322 -5415
rect 4382 -5421 4440 -5415
rect 4500 -5421 4558 -5415
rect 4618 -5421 4676 -5415
rect 4736 -5421 4794 -5415
rect 4854 -5421 4912 -5415
rect 4972 -5421 5030 -5415
rect 5090 -5421 5148 -5415
rect 5208 -5421 5266 -5415
rect 5326 -5421 5384 -5415
rect 5444 -5421 5502 -5415
rect 5562 -5421 5620 -5415
rect 5680 -5421 5738 -5415
rect 5798 -5421 5856 -5415
rect 5916 -5421 5974 -5415
rect 6034 -5421 6092 -5415
rect 6152 -5421 6210 -5415
rect 6270 -5421 6328 -5415
rect 6388 -5421 6446 -5415
rect 6506 -5421 6564 -5415
rect 6624 -5421 6682 -5415
rect 6742 -5421 6800 -5415
rect 6860 -5421 6918 -5415
rect 6978 -5421 7036 -5415
rect 7096 -5421 7154 -5415
rect 1314 -6109 1372 -6103
rect 1432 -6109 1490 -6103
rect 1550 -6109 1608 -6103
rect 1668 -6109 1726 -6103
rect 1786 -6109 1844 -6103
rect 1904 -6109 1962 -6103
rect 2022 -6109 2080 -6103
rect 2140 -6109 2198 -6103
rect 2258 -6109 2316 -6103
rect 2376 -6109 2434 -6103
rect 2494 -6109 2552 -6103
rect 2612 -6109 2670 -6103
rect 2730 -6109 2788 -6103
rect 2848 -6109 2906 -6103
rect 2966 -6109 3024 -6103
rect 3084 -6109 3142 -6103
rect 3202 -6109 3260 -6103
rect 3320 -6109 3378 -6103
rect 3438 -6109 3496 -6103
rect 3556 -6109 3614 -6103
rect 3674 -6109 3732 -6103
rect 3792 -6109 3850 -6103
rect 3910 -6109 3968 -6103
rect 4028 -6109 4086 -6103
rect 4146 -6109 4204 -6103
rect 4264 -6109 4322 -6103
rect 4382 -6109 4440 -6103
rect 4500 -6109 4558 -6103
rect 4618 -6109 4676 -6103
rect 4736 -6109 4794 -6103
rect 4854 -6109 4912 -6103
rect 4972 -6109 5030 -6103
rect 5090 -6109 5148 -6103
rect 5208 -6109 5266 -6103
rect 5326 -6109 5384 -6103
rect 5444 -6109 5502 -6103
rect 5562 -6109 5620 -6103
rect 5680 -6109 5738 -6103
rect 5798 -6109 5856 -6103
rect 5916 -6109 5974 -6103
rect 6034 -6109 6092 -6103
rect 6152 -6109 6210 -6103
rect 6270 -6109 6328 -6103
rect 6388 -6109 6446 -6103
rect 6506 -6109 6564 -6103
rect 6624 -6109 6682 -6103
rect 6742 -6109 6800 -6103
rect 6860 -6109 6918 -6103
rect 6978 -6109 7036 -6103
rect 7096 -6109 7154 -6103
rect 1314 -6143 1326 -6109
rect 1432 -6143 1444 -6109
rect 1550 -6143 1562 -6109
rect 1668 -6143 1680 -6109
rect 1786 -6143 1798 -6109
rect 1904 -6143 1916 -6109
rect 2022 -6143 2034 -6109
rect 2140 -6143 2152 -6109
rect 2258 -6143 2270 -6109
rect 2376 -6143 2388 -6109
rect 2494 -6143 2506 -6109
rect 2612 -6143 2624 -6109
rect 2730 -6143 2742 -6109
rect 2848 -6143 2860 -6109
rect 2966 -6143 2978 -6109
rect 3084 -6143 3096 -6109
rect 3202 -6143 3214 -6109
rect 3320 -6143 3332 -6109
rect 3438 -6143 3450 -6109
rect 3556 -6143 3568 -6109
rect 3674 -6143 3686 -6109
rect 3792 -6143 3804 -6109
rect 3910 -6143 3922 -6109
rect 4028 -6143 4040 -6109
rect 4146 -6143 4158 -6109
rect 4264 -6143 4276 -6109
rect 4382 -6143 4394 -6109
rect 4500 -6143 4512 -6109
rect 4618 -6143 4630 -6109
rect 4736 -6143 4748 -6109
rect 4854 -6143 4866 -6109
rect 4972 -6143 4984 -6109
rect 5090 -6143 5102 -6109
rect 5208 -6143 5220 -6109
rect 5326 -6143 5338 -6109
rect 5444 -6143 5456 -6109
rect 5562 -6143 5574 -6109
rect 5680 -6143 5692 -6109
rect 5798 -6143 5810 -6109
rect 5916 -6143 5928 -6109
rect 6034 -6143 6046 -6109
rect 6152 -6143 6164 -6109
rect 6270 -6143 6282 -6109
rect 6388 -6143 6400 -6109
rect 6506 -6143 6518 -6109
rect 6624 -6143 6636 -6109
rect 6742 -6143 6754 -6109
rect 6860 -6143 6872 -6109
rect 6978 -6143 6990 -6109
rect 7096 -6143 7108 -6109
rect 1314 -6149 1372 -6143
rect 1432 -6149 1490 -6143
rect 1550 -6149 1608 -6143
rect 1668 -6149 1726 -6143
rect 1786 -6149 1844 -6143
rect 1904 -6149 1962 -6143
rect 2022 -6149 2080 -6143
rect 2140 -6149 2198 -6143
rect 2258 -6149 2316 -6143
rect 2376 -6149 2434 -6143
rect 2494 -6149 2552 -6143
rect 2612 -6149 2670 -6143
rect 2730 -6149 2788 -6143
rect 2848 -6149 2906 -6143
rect 2966 -6149 3024 -6143
rect 3084 -6149 3142 -6143
rect 3202 -6149 3260 -6143
rect 3320 -6149 3378 -6143
rect 3438 -6149 3496 -6143
rect 3556 -6149 3614 -6143
rect 3674 -6149 3732 -6143
rect 3792 -6149 3850 -6143
rect 3910 -6149 3968 -6143
rect 4028 -6149 4086 -6143
rect 4146 -6149 4204 -6143
rect 4264 -6149 4322 -6143
rect 4382 -6149 4440 -6143
rect 4500 -6149 4558 -6143
rect 4618 -6149 4676 -6143
rect 4736 -6149 4794 -6143
rect 4854 -6149 4912 -6143
rect 4972 -6149 5030 -6143
rect 5090 -6149 5148 -6143
rect 5208 -6149 5266 -6143
rect 5326 -6149 5384 -6143
rect 5444 -6149 5502 -6143
rect 5562 -6149 5620 -6143
rect 5680 -6149 5738 -6143
rect 5798 -6149 5856 -6143
rect 5916 -6149 5974 -6143
rect 6034 -6149 6092 -6143
rect 6152 -6149 6210 -6143
rect 6270 -6149 6328 -6143
rect 6388 -6149 6446 -6143
rect 6506 -6149 6564 -6143
rect 6624 -6149 6682 -6143
rect 6742 -6149 6800 -6143
rect 6860 -6149 6918 -6143
rect 6978 -6149 7036 -6143
rect 7096 -6149 7154 -6143
rect 4741 -6535 4799 -6529
rect 4859 -6535 4917 -6529
rect 4977 -6535 5035 -6529
rect 5095 -6535 5153 -6529
rect 5213 -6535 5271 -6529
rect 5331 -6535 5389 -6529
rect 5449 -6535 5507 -6529
rect 5567 -6535 5625 -6529
rect 5685 -6535 5743 -6529
rect 5803 -6535 5861 -6529
rect 5921 -6535 5979 -6529
rect 6039 -6535 6097 -6529
rect 6157 -6535 6215 -6529
rect 6275 -6535 6333 -6529
rect 6393 -6535 6451 -6529
rect 4741 -6569 4753 -6535
rect 4859 -6569 4871 -6535
rect 4977 -6569 4989 -6535
rect 5095 -6569 5107 -6535
rect 5213 -6569 5225 -6535
rect 5331 -6569 5343 -6535
rect 5449 -6569 5461 -6535
rect 5567 -6569 5579 -6535
rect 5685 -6569 5697 -6535
rect 5803 -6569 5815 -6535
rect 5921 -6569 5933 -6535
rect 6039 -6569 6051 -6535
rect 6157 -6569 6169 -6535
rect 6275 -6569 6287 -6535
rect 6393 -6569 6405 -6535
rect 4741 -6575 4799 -6569
rect 4859 -6575 4917 -6569
rect 4977 -6575 5035 -6569
rect 5095 -6575 5153 -6569
rect 5213 -6575 5271 -6569
rect 5331 -6575 5389 -6569
rect 5449 -6575 5507 -6569
rect 5567 -6575 5625 -6569
rect 5685 -6575 5743 -6569
rect 5803 -6575 5861 -6569
rect 5921 -6575 5979 -6569
rect 6039 -6575 6097 -6569
rect 6157 -6575 6215 -6569
rect 6275 -6575 6333 -6569
rect 6393 -6575 6451 -6569
rect 2648 -6581 2706 -6575
rect 2766 -6581 2824 -6575
rect 2884 -6581 2942 -6575
rect 3002 -6581 3060 -6575
rect 3120 -6581 3178 -6575
rect 3238 -6581 3296 -6575
rect 3356 -6581 3414 -6575
rect 3474 -6581 3532 -6575
rect 3592 -6581 3650 -6575
rect 3710 -6581 3768 -6575
rect 3828 -6581 3886 -6575
rect 3946 -6581 4004 -6575
rect 4064 -6581 4122 -6575
rect 4182 -6581 4240 -6575
rect 4300 -6581 4358 -6575
rect 2648 -6615 2660 -6581
rect 2766 -6615 2778 -6581
rect 2884 -6615 2896 -6581
rect 3002 -6615 3014 -6581
rect 3120 -6615 3132 -6581
rect 3238 -6615 3250 -6581
rect 3356 -6615 3368 -6581
rect 3474 -6615 3486 -6581
rect 3592 -6615 3604 -6581
rect 3710 -6615 3722 -6581
rect 3828 -6615 3840 -6581
rect 3946 -6615 3958 -6581
rect 4064 -6615 4076 -6581
rect 4182 -6615 4194 -6581
rect 4300 -6615 4312 -6581
rect 2648 -6621 2706 -6615
rect 2766 -6621 2824 -6615
rect 2884 -6621 2942 -6615
rect 3002 -6621 3060 -6615
rect 3120 -6621 3178 -6615
rect 3238 -6621 3296 -6615
rect 3356 -6621 3414 -6615
rect 3474 -6621 3532 -6615
rect 3592 -6621 3650 -6615
rect 3710 -6621 3768 -6615
rect 3828 -6621 3886 -6615
rect 3946 -6621 4004 -6615
rect 4064 -6621 4122 -6615
rect 4182 -6621 4240 -6615
rect 4300 -6621 4358 -6615
rect 4741 -7245 4799 -7239
rect 4859 -7245 4917 -7239
rect 4977 -7245 5035 -7239
rect 5095 -7245 5153 -7239
rect 5213 -7245 5271 -7239
rect 5331 -7245 5389 -7239
rect 5449 -7245 5507 -7239
rect 5567 -7245 5625 -7239
rect 5685 -7245 5743 -7239
rect 5803 -7245 5861 -7239
rect 5921 -7245 5979 -7239
rect 6039 -7245 6097 -7239
rect 6157 -7245 6215 -7239
rect 6275 -7245 6333 -7239
rect 6393 -7245 6451 -7239
rect 4741 -7279 4753 -7245
rect 4859 -7279 4871 -7245
rect 4977 -7279 4989 -7245
rect 5095 -7279 5107 -7245
rect 5213 -7279 5225 -7245
rect 5331 -7279 5343 -7245
rect 5449 -7279 5461 -7245
rect 5567 -7279 5579 -7245
rect 5685 -7279 5697 -7245
rect 5803 -7279 5815 -7245
rect 5921 -7279 5933 -7245
rect 6039 -7279 6051 -7245
rect 6157 -7279 6169 -7245
rect 6275 -7279 6287 -7245
rect 6393 -7279 6405 -7245
rect 4741 -7285 4799 -7279
rect 4859 -7285 4917 -7279
rect 4977 -7285 5035 -7279
rect 5095 -7285 5153 -7279
rect 5213 -7285 5271 -7279
rect 5331 -7285 5389 -7279
rect 5449 -7285 5507 -7279
rect 5567 -7285 5625 -7279
rect 5685 -7285 5743 -7279
rect 5803 -7285 5861 -7279
rect 5921 -7285 5979 -7279
rect 6039 -7285 6097 -7279
rect 6157 -7285 6215 -7279
rect 6275 -7285 6333 -7279
rect 6393 -7285 6451 -7279
rect 2648 -7291 2706 -7285
rect 2766 -7291 2824 -7285
rect 2884 -7291 2942 -7285
rect 3002 -7291 3060 -7285
rect 3120 -7291 3178 -7285
rect 3238 -7291 3296 -7285
rect 3356 -7291 3414 -7285
rect 3474 -7291 3532 -7285
rect 3592 -7291 3650 -7285
rect 3710 -7291 3768 -7285
rect 3828 -7291 3886 -7285
rect 3946 -7291 4004 -7285
rect 4064 -7291 4122 -7285
rect 4182 -7291 4240 -7285
rect 4300 -7291 4358 -7285
rect 2648 -7325 2660 -7291
rect 2766 -7325 2778 -7291
rect 2884 -7325 2896 -7291
rect 3002 -7325 3014 -7291
rect 3120 -7325 3132 -7291
rect 3238 -7325 3250 -7291
rect 3356 -7325 3368 -7291
rect 3474 -7325 3486 -7291
rect 3592 -7325 3604 -7291
rect 3710 -7325 3722 -7291
rect 3828 -7325 3840 -7291
rect 3946 -7325 3958 -7291
rect 4064 -7325 4076 -7291
rect 4182 -7325 4194 -7291
rect 4300 -7325 4312 -7291
rect 2648 -7331 2706 -7325
rect 2766 -7331 2824 -7325
rect 2884 -7331 2942 -7325
rect 3002 -7331 3060 -7325
rect 3120 -7331 3178 -7325
rect 3238 -7331 3296 -7325
rect 3356 -7331 3414 -7325
rect 3474 -7331 3532 -7325
rect 3592 -7331 3650 -7325
rect 3710 -7331 3768 -7325
rect 3828 -7331 3886 -7325
rect 3946 -7331 4004 -7325
rect 4064 -7331 4122 -7325
rect 4182 -7331 4240 -7325
rect 4300 -7331 4358 -7325
rect 4741 -7353 4799 -7347
rect 4859 -7353 4917 -7347
rect 4977 -7353 5035 -7347
rect 5095 -7353 5153 -7347
rect 5213 -7353 5271 -7347
rect 5331 -7353 5389 -7347
rect 5449 -7353 5507 -7347
rect 5567 -7353 5625 -7347
rect 5685 -7353 5743 -7347
rect 5803 -7353 5861 -7347
rect 5921 -7353 5979 -7347
rect 6039 -7353 6097 -7347
rect 6157 -7353 6215 -7347
rect 6275 -7353 6333 -7347
rect 6393 -7353 6451 -7347
rect 4741 -7387 4753 -7353
rect 4859 -7387 4871 -7353
rect 4977 -7387 4989 -7353
rect 5095 -7387 5107 -7353
rect 5213 -7387 5225 -7353
rect 5331 -7387 5343 -7353
rect 5449 -7387 5461 -7353
rect 5567 -7387 5579 -7353
rect 5685 -7387 5697 -7353
rect 5803 -7387 5815 -7353
rect 5921 -7387 5933 -7353
rect 6039 -7387 6051 -7353
rect 6157 -7387 6169 -7353
rect 6275 -7387 6287 -7353
rect 6393 -7387 6405 -7353
rect 4741 -7393 4799 -7387
rect 4859 -7393 4917 -7387
rect 4977 -7393 5035 -7387
rect 5095 -7393 5153 -7387
rect 5213 -7393 5271 -7387
rect 5331 -7393 5389 -7387
rect 5449 -7393 5507 -7387
rect 5567 -7393 5625 -7387
rect 5685 -7393 5743 -7387
rect 5803 -7393 5861 -7387
rect 5921 -7393 5979 -7387
rect 6039 -7393 6097 -7387
rect 6157 -7393 6215 -7387
rect 6275 -7393 6333 -7387
rect 6393 -7393 6451 -7387
rect 2648 -7399 2706 -7393
rect 2766 -7399 2824 -7393
rect 2884 -7399 2942 -7393
rect 3002 -7399 3060 -7393
rect 3120 -7399 3178 -7393
rect 3238 -7399 3296 -7393
rect 3356 -7399 3414 -7393
rect 3474 -7399 3532 -7393
rect 3592 -7399 3650 -7393
rect 3710 -7399 3768 -7393
rect 3828 -7399 3886 -7393
rect 3946 -7399 4004 -7393
rect 4064 -7399 4122 -7393
rect 4182 -7399 4240 -7393
rect 4300 -7399 4358 -7393
rect 2648 -7433 2660 -7399
rect 2766 -7433 2778 -7399
rect 2884 -7433 2896 -7399
rect 3002 -7433 3014 -7399
rect 3120 -7433 3132 -7399
rect 3238 -7433 3250 -7399
rect 3356 -7433 3368 -7399
rect 3474 -7433 3486 -7399
rect 3592 -7433 3604 -7399
rect 3710 -7433 3722 -7399
rect 3828 -7433 3840 -7399
rect 3946 -7433 3958 -7399
rect 4064 -7433 4076 -7399
rect 4182 -7433 4194 -7399
rect 4300 -7433 4312 -7399
rect 2648 -7439 2706 -7433
rect 2766 -7439 2824 -7433
rect 2884 -7439 2942 -7433
rect 3002 -7439 3060 -7433
rect 3120 -7439 3178 -7433
rect 3238 -7439 3296 -7433
rect 3356 -7439 3414 -7433
rect 3474 -7439 3532 -7433
rect 3592 -7439 3650 -7433
rect 3710 -7439 3768 -7433
rect 3828 -7439 3886 -7433
rect 3946 -7439 4004 -7433
rect 4064 -7439 4122 -7433
rect 4182 -7439 4240 -7433
rect 4300 -7439 4358 -7433
rect 4741 -8063 4799 -8057
rect 4859 -8063 4917 -8057
rect 4977 -8063 5035 -8057
rect 5095 -8063 5153 -8057
rect 5213 -8063 5271 -8057
rect 5331 -8063 5389 -8057
rect 5449 -8063 5507 -8057
rect 5567 -8063 5625 -8057
rect 5685 -8063 5743 -8057
rect 5803 -8063 5861 -8057
rect 5921 -8063 5979 -8057
rect 6039 -8063 6097 -8057
rect 6157 -8063 6215 -8057
rect 6275 -8063 6333 -8057
rect 6393 -8063 6451 -8057
rect 4741 -8097 4753 -8063
rect 4859 -8097 4871 -8063
rect 4977 -8097 4989 -8063
rect 5095 -8097 5107 -8063
rect 5213 -8097 5225 -8063
rect 5331 -8097 5343 -8063
rect 5449 -8097 5461 -8063
rect 5567 -8097 5579 -8063
rect 5685 -8097 5697 -8063
rect 5803 -8097 5815 -8063
rect 5921 -8097 5933 -8063
rect 6039 -8097 6051 -8063
rect 6157 -8097 6169 -8063
rect 6275 -8097 6287 -8063
rect 6393 -8097 6405 -8063
rect 4741 -8103 4799 -8097
rect 4859 -8103 4917 -8097
rect 4977 -8103 5035 -8097
rect 5095 -8103 5153 -8097
rect 5213 -8103 5271 -8097
rect 5331 -8103 5389 -8097
rect 5449 -8103 5507 -8097
rect 5567 -8103 5625 -8097
rect 5685 -8103 5743 -8097
rect 5803 -8103 5861 -8097
rect 5921 -8103 5979 -8097
rect 6039 -8103 6097 -8097
rect 6157 -8103 6215 -8097
rect 6275 -8103 6333 -8097
rect 6393 -8103 6451 -8097
rect 2648 -8109 2706 -8103
rect 2766 -8109 2824 -8103
rect 2884 -8109 2942 -8103
rect 3002 -8109 3060 -8103
rect 3120 -8109 3178 -8103
rect 3238 -8109 3296 -8103
rect 3356 -8109 3414 -8103
rect 3474 -8109 3532 -8103
rect 3592 -8109 3650 -8103
rect 3710 -8109 3768 -8103
rect 3828 -8109 3886 -8103
rect 3946 -8109 4004 -8103
rect 4064 -8109 4122 -8103
rect 4182 -8109 4240 -8103
rect 4300 -8109 4358 -8103
rect 2648 -8143 2660 -8109
rect 2766 -8143 2778 -8109
rect 2884 -8143 2896 -8109
rect 3002 -8143 3014 -8109
rect 3120 -8143 3132 -8109
rect 3238 -8143 3250 -8109
rect 3356 -8143 3368 -8109
rect 3474 -8143 3486 -8109
rect 3592 -8143 3604 -8109
rect 3710 -8143 3722 -8109
rect 3828 -8143 3840 -8109
rect 3946 -8143 3958 -8109
rect 4064 -8143 4076 -8109
rect 4182 -8143 4194 -8109
rect 4300 -8143 4312 -8109
rect 2648 -8149 2706 -8143
rect 2766 -8149 2824 -8143
rect 2884 -8149 2942 -8143
rect 3002 -8149 3060 -8143
rect 3120 -8149 3178 -8143
rect 3238 -8149 3296 -8143
rect 3356 -8149 3414 -8143
rect 3474 -8149 3532 -8143
rect 3592 -8149 3650 -8143
rect 3710 -8149 3768 -8143
rect 3828 -8149 3886 -8143
rect 3946 -8149 4004 -8143
rect 4064 -8149 4122 -8143
rect 4182 -8149 4240 -8143
rect 4300 -8149 4358 -8143
<< nwell >>
rect 12783 1936 12959 1999
rect 13019 1937 13431 1999
rect 13491 1937 14375 1999
rect 14435 1937 16263 1999
rect 16323 1937 18151 1999
rect 18211 1937 20039 1999
rect 20099 1937 21376 1999
<< pwell >>
rect 22030 -8266 22330 -8220
<< poly >>
rect 12783 1989 12845 1999
rect 12897 1989 12959 1999
rect 13019 1989 13081 1999
rect 13133 1989 13199 1999
rect 13251 1989 13317 1999
rect 13369 1989 13431 1999
rect 13491 1989 13553 1999
rect 13605 1989 13671 1999
rect 13723 1989 13789 1999
rect 13841 1989 13907 1999
rect 13959 1989 14025 1999
rect 14077 1989 14143 1999
rect 14195 1989 14261 1999
rect 14313 1989 14375 1999
rect 14435 1989 14497 1999
rect 14549 1989 14615 1999
rect 14667 1989 14733 1999
rect 14785 1989 14851 1999
rect 14903 1989 14969 1999
rect 15021 1989 15087 1999
rect 15139 1989 15205 1999
rect 15257 1989 15323 1999
rect 15375 1989 15441 1999
rect 15493 1989 15559 1999
rect 15611 1989 15677 1999
rect 15729 1989 15795 1999
rect 15847 1989 15913 1999
rect 15965 1989 16031 1999
rect 16083 1989 16149 1999
rect 16201 1989 16263 1999
rect 16323 1989 16385 1999
rect 16437 1989 16503 1999
rect 16555 1989 16621 1999
rect 16673 1989 16739 1999
rect 16791 1989 16857 1999
rect 16909 1989 16975 1999
rect 17027 1989 17093 1999
rect 17145 1989 17211 1999
rect 17263 1989 17329 1999
rect 17381 1989 17447 1999
rect 17499 1989 17565 1999
rect 17617 1989 17683 1999
rect 17735 1989 17801 1999
rect 17853 1989 17919 1999
rect 17971 1989 18037 1999
rect 18089 1989 18151 1999
rect 18211 1989 18273 1999
rect 18325 1989 18391 1999
rect 18443 1989 18509 1999
rect 18561 1989 18627 1999
rect 18679 1989 18745 1999
rect 18797 1989 18863 1999
rect 18915 1989 18981 1999
rect 19033 1989 19099 1999
rect 19151 1989 19217 1999
rect 19269 1989 19335 1999
rect 19387 1989 19453 1999
rect 19505 1989 19571 1999
rect 19623 1989 19689 1999
rect 19741 1989 19807 1999
rect 19859 1989 19925 1999
rect 19977 1989 20039 1999
rect 20099 1989 20161 1999
rect 20213 1989 20279 1999
rect 20331 1989 20397 1999
rect 20449 1989 20515 1999
rect 20567 1989 20633 1999
rect 20685 1989 20751 1999
rect 20803 1989 20869 1999
rect 20921 1989 20987 1999
rect 21039 1989 21105 1999
rect 21157 1989 21223 1999
rect 21275 1989 21341 1999
rect 12783 1936 12845 1947
rect 12897 1936 12959 1947
rect 13019 1937 13081 1947
rect 13133 1937 13199 1947
rect 13251 1937 13317 1947
rect 13369 1937 13431 1947
rect 13491 1937 13553 1947
rect 13605 1937 13671 1947
rect 13723 1937 13789 1947
rect 13841 1937 13907 1947
rect 13959 1937 14025 1947
rect 14077 1937 14143 1947
rect 14195 1937 14261 1947
rect 14313 1937 14375 1947
rect 14435 1937 14497 1947
rect 14549 1937 14615 1947
rect 14667 1937 14733 1947
rect 14785 1937 14851 1947
rect 14903 1937 14969 1947
rect 15021 1937 15087 1947
rect 15139 1937 15205 1947
rect 15257 1937 15323 1947
rect 15375 1937 15441 1947
rect 15493 1937 15559 1947
rect 15611 1937 15677 1947
rect 15729 1937 15795 1947
rect 15847 1937 15913 1947
rect 15965 1937 16031 1947
rect 16083 1937 16149 1947
rect 16201 1937 16263 1947
rect 16323 1937 16385 1947
rect 16437 1937 16503 1947
rect 16555 1937 16621 1947
rect 16673 1937 16739 1947
rect 16791 1937 16857 1947
rect 16909 1937 16975 1947
rect 17027 1937 17093 1947
rect 17145 1937 17211 1947
rect 17263 1937 17329 1947
rect 17381 1937 17447 1947
rect 17499 1937 17565 1947
rect 17617 1937 17683 1947
rect 17735 1937 17801 1947
rect 17853 1937 17919 1947
rect 17971 1937 18037 1947
rect 18089 1937 18151 1947
rect 18211 1937 18273 1947
rect 18325 1937 18391 1947
rect 18443 1937 18509 1947
rect 18561 1937 18627 1947
rect 18679 1937 18745 1947
rect 18797 1937 18863 1947
rect 18915 1937 18981 1947
rect 19033 1937 19099 1947
rect 19151 1937 19217 1947
rect 19269 1937 19335 1947
rect 19387 1937 19453 1947
rect 19505 1937 19571 1947
rect 19623 1937 19689 1947
rect 19741 1937 19807 1947
rect 19859 1937 19925 1947
rect 19977 1937 20039 1947
rect 20099 1937 20161 1947
rect 20213 1937 20279 1947
rect 20331 1937 20397 1947
rect 20449 1937 20515 1947
rect 20567 1937 20633 1947
rect 20685 1937 20751 1947
rect 20803 1937 20869 1947
rect 20921 1937 20987 1947
rect 21039 1937 21105 1947
rect 21157 1937 21223 1947
rect 21275 1937 21341 1947
rect 22030 -8266 22038 -8220
rect 22096 -8226 22186 -8220
rect 22096 -8260 22112 -8226
rect 22170 -8260 22186 -8226
rect 22096 -8266 22186 -8260
rect 22244 -8226 22330 -8220
rect 22244 -8260 22260 -8226
rect 22318 -8260 22330 -8226
rect 22244 -8266 22330 -8260
<< polycont >>
rect 22112 -8260 22170 -8226
rect 22260 -8260 22318 -8226
<< locali >>
rect 22030 -8260 22038 -8226
rect 22096 -8260 22112 -8226
rect 22170 -8260 22186 -8226
rect 22244 -8260 22260 -8226
rect 22318 -8260 22330 -8226
<< viali >>
rect 22112 -8260 22170 -8226
rect 22260 -8260 22318 -8226
<< metal1 >>
rect 12547 1936 12605 2000
rect 12665 1935 12723 1999
rect 12783 1936 12841 1999
rect 12901 1936 12959 1999
rect 13019 1937 13077 1999
rect 13137 1937 13195 1999
rect 13255 1937 13313 1999
rect 13373 1937 13431 1999
rect 13491 1937 13549 1999
rect 13609 1937 13667 1999
rect 13727 1937 13785 1999
rect 13845 1937 13903 1999
rect 13963 1937 14021 1999
rect 14081 1937 14139 1999
rect 14199 1937 14257 1999
rect 14317 1937 14375 1999
rect 14435 1937 14493 1999
rect 14553 1937 14611 1999
rect 14671 1937 14729 1999
rect 14789 1937 14847 1999
rect 14907 1937 14965 1999
rect 15025 1937 15083 1999
rect 15143 1937 15201 1999
rect 15261 1937 15319 1999
rect 15379 1937 15437 1999
rect 15497 1937 15555 1999
rect 15615 1937 15673 1999
rect 15733 1937 15791 1999
rect 15851 1937 15909 1999
rect 15969 1937 16027 1999
rect 16087 1937 16145 1999
rect 16205 1937 16263 1999
rect 16323 1937 16381 1999
rect 16441 1937 16499 1999
rect 16559 1937 16617 1999
rect 16677 1937 16735 1999
rect 16795 1937 16853 1999
rect 16913 1937 16971 1999
rect 17031 1937 17089 1999
rect 17149 1937 17207 1999
rect 17267 1937 17325 1999
rect 17385 1937 17443 1999
rect 17503 1937 17561 1999
rect 17621 1937 17679 1999
rect 17739 1937 17797 1999
rect 17857 1937 17915 1999
rect 17975 1937 18033 1999
rect 18093 1937 18151 1999
rect 18211 1937 18269 1999
rect 18329 1937 18387 1999
rect 18447 1937 18505 1999
rect 18565 1937 18623 1999
rect 18683 1937 18741 1999
rect 18801 1937 18859 1999
rect 18919 1937 18977 1999
rect 19037 1937 19095 1999
rect 19155 1937 19213 1999
rect 19273 1937 19331 1999
rect 19391 1937 19449 1999
rect 19509 1937 19567 1999
rect 19627 1937 19685 1999
rect 19745 1937 19803 1999
rect 19863 1937 19921 1999
rect 19981 1937 20039 1999
rect 20099 1937 20157 1999
rect 20217 1937 20275 1999
rect 20335 1937 20393 1999
rect 20453 1937 20511 1999
rect 20571 1937 20629 1999
rect 20689 1937 20747 1999
rect 20807 1937 20865 1999
rect 20925 1937 20983 1999
rect 21043 1937 21101 1999
rect 21161 1937 21219 1999
rect 21279 1937 21337 1999
rect 11378 -8266 21212 -8220
rect 21293 -8266 21952 -8220
rect 22030 -8226 22330 -8220
rect 22030 -8260 22112 -8226
rect 22170 -8260 22260 -8226
rect 22318 -8260 22330 -8226
rect 22030 -8266 22330 -8260
use sky130_fd_pr__nfet_01v8_8HUREQ  sky130_fd_pr__nfet_01v8_8HUREQ_0
timestamp 1606416512
transform 1 0 3503 0 1 -7362
box -1052 -919 1052 919
use sky130_fd_pr__nfet_01v8_8HUREQ  sky130_fd_pr__nfet_01v8_8HUREQ_1
timestamp 1606416512
transform 1 0 5596 0 1 -7316
box -1052 -919 1052 919
use sky130_fd_pr__pfet_01v8_YCMRKB  sky130_fd_pr__pfet_01v8_YCMRKB_3
timestamp 1606426375
transform 1 0 4234 0 1 -5344
box -3117 -937 3117 937
use sky130_fd_pr__pfet_01v8_YCMRKB  sky130_fd_pr__pfet_01v8_YCMRKB_2
timestamp 1606426375
transform 1 0 4234 0 1 -3596
box -3117 -937 3117 937
use sky130_fd_pr__pfet_01v8_QCPMCH  sky130_fd_pr__pfet_01v8_QCPMCH_0
timestamp 1606424343
transform 1 0 9520 0 1 -2505
box -211 -637 211 637
use sky130_fd_pr__pfet_01v8_YCMRKB  sky130_fd_pr__pfet_01v8_YCMRKB_0
timestamp 1606426375
transform 1 0 4257 0 1 -1987
box -3117 -937 3117 937
use sky130_fd_pr__pfet_01v8_YCMRKB  sky130_fd_pr__pfet_01v8_YCMRKB_1
timestamp 1606426375
transform 1 0 4303 0 1 -216
box -3117 -937 3117 937
use sky130_fd_pr__pfet_01v8_YC9MKB  sky130_fd_pr__pfet_01v8_YC9MKB_0
timestamp 1606426375
transform 1 0 1572 0 1 1758
box -1052 -519 1052 519
use sky130_fd_pr__pfet_01v8_YC9MKB  sky130_fd_pr__pfet_01v8_YC9MKB_1
timestamp 1606426375
transform 1 0 3871 0 1 1758
box -1052 -519 1052 519
use sky130_fd_pr__pfet_01v8_YC9MKB  sky130_fd_pr__pfet_01v8_YC9MKB_2
timestamp 1606426375
transform 1 0 6010 0 1 1758
box -1052 -519 1052 519
use sky130_fd_pr__pfet_01v8_YC99EG  sky130_fd_pr__pfet_01v8_YC99EG_0
timestamp 1606426095
transform 1 0 16942 0 1 1968
box -4592 -937 4592 937
use sky130_fd_pr__cap_mim_m3_1_BLS9ZS  sky130_fd_pr__cap_mim_m3_1_BLS9ZS_0
timestamp 1606431493
transform -1 0 16853 0 1 -2470
box -5943 -3300 5943 3300
use sky130_fd_pr__nfet_01v8_8JUMX6  sky130_fd_pr__nfet_01v8_8JUMX6_0
timestamp 1606424956
transform 1 0 16813 0 1 -7179
box -5717 -1219 5717 1219
<< end >>
