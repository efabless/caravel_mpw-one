magic
tech sky130A
magscale 1 2
timestamp 1622551583
<< locali >>
rect 21925 2839 21959 2941
<< viali >>
rect 2513 3689 2547 3723
rect 2789 3621 2823 3655
rect 3065 3553 3099 3587
rect 3341 3485 3375 3519
rect 2237 3009 2271 3043
rect 2513 3009 2547 3043
rect 2789 3009 2823 3043
rect 4445 3009 4479 3043
rect 4997 3009 5031 3043
rect 5825 3009 5859 3043
rect 6101 3009 6135 3043
rect 7021 3009 7055 3043
rect 7297 3009 7331 3043
rect 8401 3009 8435 3043
rect 9229 3009 9263 3043
rect 10057 3009 10091 3043
rect 10333 3009 10367 3043
rect 11713 3009 11747 3043
rect 12541 3009 12575 3043
rect 14197 3009 14231 3043
rect 14473 3009 14507 3043
rect 15577 3009 15611 3043
rect 17233 3009 17267 3043
rect 17785 3009 17819 3043
rect 18337 3009 18371 3043
rect 19165 3009 19199 3043
rect 19441 3009 19475 3043
rect 19993 3009 20027 3043
rect 20821 3009 20855 3043
rect 21373 3009 21407 3043
rect 21649 3009 21683 3043
rect 22201 3009 22235 3043
rect 23305 3009 23339 3043
rect 23581 3009 23615 3043
rect 23857 3009 23891 3043
rect 24685 3009 24719 3043
rect 25237 3009 25271 3043
rect 26065 3009 26099 3043
rect 26341 3009 26375 3043
rect 26617 3009 26651 3043
rect 26893 3009 26927 3043
rect 27445 3009 27479 3043
rect 28273 3009 28307 3043
rect 28825 3009 28859 3043
rect 29101 3009 29135 3043
rect 29929 3009 29963 3043
rect 30205 3009 30239 3043
rect 32045 3009 32079 3043
rect 32321 3009 32355 3043
rect 36277 3009 36311 3043
rect 36553 3009 36587 3043
rect 37105 3009 37139 3043
rect 37381 3009 37415 3043
rect 37933 3009 37967 3043
rect 38485 3009 38519 3043
rect 39037 3009 39071 3043
rect 39589 3009 39623 3043
rect 40141 3009 40175 3043
rect 40693 3009 40727 3043
rect 41245 3009 41279 3043
rect 41797 3009 41831 3043
rect 42349 3009 42383 3043
rect 43177 3009 43211 3043
rect 44005 3009 44039 3043
rect 44833 3009 44867 3043
rect 45661 3009 45695 3043
rect 46489 3009 46523 3043
rect 47317 3009 47351 3043
rect 48973 3009 49007 3043
rect 49249 3009 49283 3043
rect 50353 3009 50387 3043
rect 51181 3009 51215 3043
rect 52009 3009 52043 3043
rect 52561 3009 52595 3043
rect 53941 3009 53975 3043
rect 54493 3009 54527 3043
rect 55597 3009 55631 3043
rect 56701 3009 56735 3043
rect 56977 3009 57011 3043
rect 58081 3009 58115 3043
rect 59461 3009 59495 3043
rect 59737 3009 59771 3043
rect 60289 3009 60323 3043
rect 61393 3009 61427 3043
rect 61669 3009 61703 3043
rect 62497 3009 62531 3043
rect 62773 3009 62807 3043
rect 63049 3009 63083 3043
rect 64705 3009 64739 3043
rect 64981 3009 65015 3043
rect 65809 3009 65843 3043
rect 66361 3009 66395 3043
rect 67189 3009 67223 3043
rect 68753 3009 68787 3043
rect 69029 3009 69063 3043
rect 2145 2941 2179 2975
rect 4721 2941 4755 2975
rect 6469 2941 6503 2975
rect 7573 2941 7607 2975
rect 8677 2941 8711 2975
rect 9781 2941 9815 2975
rect 10885 2941 10919 2975
rect 12265 2941 12299 2975
rect 13645 2941 13679 2975
rect 15025 2941 15059 2975
rect 16957 2941 16991 2975
rect 18613 2941 18647 2975
rect 20269 2941 20303 2975
rect 21925 2941 21959 2975
rect 22753 2941 22787 2975
rect 24133 2941 24167 2975
rect 25513 2941 25547 2975
rect 27997 2941 28031 2975
rect 29377 2941 29411 2975
rect 32689 2941 32723 2975
rect 38209 2941 38243 2975
rect 38761 2941 38795 2975
rect 39313 2941 39347 2975
rect 39865 2941 39899 2975
rect 40417 2941 40451 2975
rect 40969 2941 41003 2975
rect 41521 2941 41555 2975
rect 42073 2941 42107 2975
rect 42625 2941 42659 2975
rect 43453 2941 43487 2975
rect 44281 2941 44315 2975
rect 45109 2941 45143 2975
rect 45937 2941 45971 2975
rect 46765 2941 46799 2975
rect 47593 2941 47627 2975
rect 49525 2941 49559 2975
rect 50629 2941 50663 2975
rect 51733 2941 51767 2975
rect 52837 2941 52871 2975
rect 54217 2941 54251 2975
rect 55321 2941 55355 2975
rect 55873 2941 55907 2975
rect 58357 2941 58391 2975
rect 60013 2941 60047 2975
rect 61117 2941 61151 2975
rect 61945 2941 61979 2975
rect 64153 2941 64187 2975
rect 65533 2941 65567 2975
rect 66637 2941 66671 2975
rect 69397 2941 69431 2975
rect 3065 2873 3099 2907
rect 4169 2873 4203 2907
rect 5273 2873 5307 2907
rect 6745 2873 6779 2907
rect 8125 2873 8159 2907
rect 9505 2873 9539 2907
rect 10609 2873 10643 2907
rect 11989 2873 12023 2907
rect 13369 2873 13403 2907
rect 14749 2873 14783 2907
rect 16405 2873 16439 2907
rect 18061 2873 18095 2907
rect 18889 2873 18923 2907
rect 20545 2873 20579 2907
rect 22477 2873 22511 2907
rect 24409 2873 24443 2907
rect 25789 2873 25823 2907
rect 27721 2873 27755 2907
rect 31585 2873 31619 2907
rect 36829 2873 36863 2907
rect 43729 2873 43763 2907
rect 44557 2873 44591 2907
rect 45385 2873 45419 2907
rect 46213 2873 46247 2907
rect 47041 2873 47075 2907
rect 47869 2873 47903 2907
rect 48697 2873 48731 2907
rect 49801 2873 49835 2907
rect 50905 2873 50939 2907
rect 52285 2873 52319 2907
rect 53665 2873 53699 2907
rect 55045 2873 55079 2907
rect 56425 2873 56459 2907
rect 57805 2873 57839 2907
rect 60841 2873 60875 2907
rect 63325 2873 63359 2907
rect 66085 2873 66119 2907
rect 67465 2873 67499 2907
rect 67741 2873 67775 2907
rect 68017 2873 68051 2907
rect 3341 2805 3375 2839
rect 3617 2805 3651 2839
rect 3893 2805 3927 2839
rect 5549 2805 5583 2839
rect 7849 2805 7883 2839
rect 8953 2805 8987 2839
rect 11161 2805 11195 2839
rect 12817 2805 12851 2839
rect 13093 2805 13127 2839
rect 13921 2805 13955 2839
rect 15301 2805 15335 2839
rect 15853 2805 15887 2839
rect 16129 2805 16163 2839
rect 17509 2805 17543 2839
rect 19717 2805 19751 2839
rect 21097 2805 21131 2839
rect 21925 2805 21959 2839
rect 23029 2805 23063 2839
rect 24961 2805 24995 2839
rect 28549 2805 28583 2839
rect 29653 2805 29687 2839
rect 30481 2805 30515 2839
rect 30757 2805 30791 2839
rect 31033 2805 31067 2839
rect 31309 2805 31343 2839
rect 48421 2805 48455 2839
rect 50077 2805 50111 2839
rect 51457 2805 51491 2839
rect 53113 2805 53147 2839
rect 54769 2805 54803 2839
rect 56149 2805 56183 2839
rect 57253 2805 57287 2839
rect 57529 2805 57563 2839
rect 58909 2805 58943 2839
rect 59185 2805 59219 2839
rect 60565 2805 60599 2839
rect 62221 2805 62255 2839
rect 63601 2805 63635 2839
rect 64429 2805 64463 2839
rect 65257 2805 65291 2839
rect 66913 2805 66947 2839
rect 68293 2805 68327 2839
rect 3065 2601 3099 2635
rect 2789 2465 2823 2499
rect 2513 2397 2547 2431
rect 3157 1853 3191 1887
rect 31033 1785 31067 1819
rect 2237 1717 2271 1751
rect 2513 1717 2547 1751
rect 2881 1717 2915 1751
rect 3433 1717 3467 1751
rect 4077 1717 4111 1751
rect 7021 1717 7055 1751
rect 8953 1717 8987 1751
rect 9873 1717 9907 1751
rect 11897 1717 11931 1751
rect 13277 1717 13311 1751
rect 15209 1717 15243 1751
rect 16129 1717 16163 1751
rect 20361 1717 20395 1751
rect 26709 1717 26743 1751
rect 30757 1717 30791 1751
rect 32689 1717 32723 1751
rect 38577 1717 38611 1751
rect 44005 1717 44039 1751
rect 46857 1717 46891 1751
rect 50537 1717 50571 1751
rect 52561 1717 52595 1751
rect 54401 1717 54435 1751
rect 57529 1717 57563 1751
rect 64153 1717 64187 1751
rect 68201 1717 68235 1751
rect 69581 1717 69615 1751
rect 2789 1513 2823 1547
rect 24869 1513 24903 1547
rect 26341 1513 26375 1547
rect 28733 1513 28767 1547
rect 30849 1513 30883 1547
rect 32137 1513 32171 1547
rect 2145 1445 2179 1479
rect 4169 1445 4203 1479
rect 4721 1445 4755 1479
rect 5365 1445 5399 1479
rect 8125 1445 8159 1479
rect 9597 1445 9631 1479
rect 10333 1445 10367 1479
rect 12265 1445 12299 1479
rect 13001 1445 13035 1479
rect 13829 1445 13863 1479
rect 14565 1445 14599 1479
rect 15577 1445 15611 1479
rect 16589 1445 16623 1479
rect 17509 1445 17543 1479
rect 18337 1445 18371 1479
rect 19165 1445 19199 1479
rect 20637 1445 20671 1479
rect 21465 1445 21499 1479
rect 23397 1445 23431 1479
rect 24317 1445 24351 1479
rect 25513 1445 25547 1479
rect 27353 1445 27387 1479
rect 29009 1445 29043 1479
rect 30573 1445 30607 1479
rect 31585 1445 31619 1479
rect 32873 1445 32907 1479
rect 37841 1445 37875 1479
rect 39129 1445 39163 1479
rect 40233 1445 40267 1479
rect 41429 1445 41463 1479
rect 41981 1445 42015 1479
rect 42533 1445 42567 1479
rect 43085 1445 43119 1479
rect 60197 1445 60231 1479
rect 61025 1445 61059 1479
rect 61577 1445 61611 1479
rect 62129 1445 62163 1479
rect 65257 1445 65291 1479
rect 66453 1445 66487 1479
rect 67281 1445 67315 1479
rect 68477 1445 68511 1479
rect 69305 1445 69339 1479
rect 70041 1445 70075 1479
rect 1685 1377 1719 1411
rect 3065 1377 3099 1411
rect 5641 1377 5675 1411
rect 6193 1377 6227 1411
rect 6837 1377 6871 1411
rect 7573 1377 7607 1411
rect 8401 1377 8435 1411
rect 10609 1377 10643 1411
rect 11253 1377 11287 1411
rect 13277 1377 13311 1411
rect 15853 1377 15887 1411
rect 17785 1377 17819 1411
rect 18613 1377 18647 1411
rect 19441 1377 19475 1411
rect 21189 1377 21223 1411
rect 22109 1377 22143 1411
rect 23121 1377 23155 1411
rect 23765 1377 23799 1411
rect 25237 1377 25271 1411
rect 25789 1377 25823 1411
rect 26985 1377 27019 1411
rect 28457 1377 28491 1411
rect 29837 1377 29871 1411
rect 31309 1377 31343 1411
rect 33241 1377 33275 1411
rect 38853 1377 38887 1411
rect 39405 1377 39439 1411
rect 39957 1377 39991 1411
rect 40785 1377 40819 1411
rect 49525 1377 49559 1411
rect 50353 1377 50387 1411
rect 52377 1377 52411 1411
rect 62865 1377 62899 1411
rect 63417 1377 63451 1411
rect 64429 1377 64463 1411
rect 66177 1377 66211 1411
rect 67005 1377 67039 1411
rect 68201 1377 68235 1411
rect 70593 1377 70627 1411
rect 2237 1309 2271 1343
rect 2513 1309 2547 1343
rect 3341 1309 3375 1343
rect 3893 1309 3927 1343
rect 4445 1309 4479 1343
rect 5089 1309 5123 1343
rect 5917 1309 5951 1343
rect 6561 1309 6595 1343
rect 7297 1309 7331 1343
rect 7849 1309 7883 1343
rect 8769 1309 8803 1343
rect 9321 1309 9355 1343
rect 10057 1309 10091 1343
rect 10977 1309 11011 1343
rect 11529 1309 11563 1343
rect 11897 1309 11931 1343
rect 12725 1309 12759 1343
rect 13553 1309 13587 1343
rect 14105 1309 14139 1343
rect 14933 1309 14967 1343
rect 15209 1309 15243 1343
rect 16313 1309 16347 1343
rect 16865 1309 16899 1343
rect 17233 1309 17267 1343
rect 18061 1309 18095 1343
rect 18889 1309 18923 1343
rect 19901 1309 19935 1343
rect 20177 1309 20211 1343
rect 20913 1309 20947 1343
rect 21741 1309 21775 1343
rect 22569 1309 22603 1343
rect 22845 1309 22879 1343
rect 24041 1309 24075 1343
rect 24593 1309 24627 1343
rect 26065 1309 26099 1343
rect 26617 1309 26651 1343
rect 27905 1309 27939 1343
rect 28181 1309 28215 1343
rect 29285 1309 29319 1343
rect 29561 1309 29595 1343
rect 30113 1309 30147 1343
rect 31861 1309 31895 1343
rect 32597 1309 32631 1343
rect 38117 1309 38151 1343
rect 38393 1309 38427 1343
rect 39681 1309 39715 1343
rect 40509 1309 40543 1343
rect 41061 1309 41095 1343
rect 41705 1309 41739 1343
rect 42257 1309 42291 1343
rect 42809 1309 42843 1343
rect 43361 1309 43395 1343
rect 43729 1309 43763 1343
rect 44281 1309 44315 1343
rect 44557 1309 44591 1343
rect 44833 1309 44867 1343
rect 45109 1309 45143 1343
rect 45385 1309 45419 1343
rect 45661 1309 45695 1343
rect 45937 1309 45971 1343
rect 46305 1309 46339 1343
rect 46765 1309 46799 1343
rect 47133 1309 47167 1343
rect 47409 1309 47443 1343
rect 47685 1309 47719 1343
rect 47961 1309 47995 1343
rect 48237 1309 48271 1343
rect 48605 1309 48639 1343
rect 48881 1309 48915 1343
rect 49433 1309 49467 1343
rect 49985 1309 50019 1343
rect 50261 1309 50295 1343
rect 50905 1309 50939 1343
rect 51181 1309 51215 1343
rect 51457 1309 51491 1343
rect 51733 1309 51767 1343
rect 52285 1309 52319 1343
rect 52837 1309 52871 1343
rect 53021 1309 53055 1343
rect 53297 1309 53331 1343
rect 53573 1309 53607 1343
rect 53849 1309 53883 1343
rect 54125 1309 54159 1343
rect 54677 1309 54711 1343
rect 54953 1309 54987 1343
rect 55229 1309 55263 1343
rect 55597 1309 55631 1343
rect 55873 1309 55907 1343
rect 56149 1309 56183 1343
rect 56425 1309 56459 1343
rect 56701 1309 56735 1343
rect 57253 1309 57287 1343
rect 57529 1309 57563 1343
rect 57805 1309 57839 1343
rect 58081 1309 58115 1343
rect 58449 1309 58483 1343
rect 58725 1309 58759 1343
rect 59001 1309 59035 1343
rect 59277 1309 59311 1343
rect 59553 1309 59587 1343
rect 59921 1309 59955 1343
rect 60473 1309 60507 1343
rect 60749 1309 60783 1343
rect 61301 1309 61335 1343
rect 61853 1309 61887 1343
rect 62589 1309 62623 1343
rect 63141 1309 63175 1343
rect 63693 1309 63727 1343
rect 64153 1309 64187 1343
rect 64705 1309 64739 1343
rect 65625 1309 65659 1343
rect 65901 1309 65935 1343
rect 66729 1309 66763 1343
rect 67557 1309 67591 1343
rect 67925 1309 67959 1343
rect 68753 1309 68787 1343
rect 69029 1309 69063 1343
rect 69765 1309 69799 1343
<< metal1 >>
rect 3050 3952 3056 4004
rect 3108 3992 3114 4004
rect 3786 3992 3792 4004
rect 3108 3964 3792 3992
rect 3108 3952 3114 3964
rect 3786 3952 3792 3964
rect 3844 3952 3850 4004
rect 9122 3952 9128 4004
rect 9180 3992 9186 4004
rect 10042 3992 10048 4004
rect 9180 3964 10048 3992
rect 9180 3952 9186 3964
rect 10042 3952 10048 3964
rect 10100 3952 10106 4004
rect 20990 3952 20996 4004
rect 21048 3992 21054 4004
rect 22738 3992 22744 4004
rect 21048 3964 22744 3992
rect 21048 3952 21054 3964
rect 22738 3952 22744 3964
rect 22796 3952 22802 4004
rect 27062 3952 27068 4004
rect 27120 3992 27126 4004
rect 29086 3992 29092 4004
rect 27120 3964 29092 3992
rect 27120 3952 27126 3964
rect 29086 3952 29092 3964
rect 29144 3952 29150 4004
rect 45002 3952 45008 4004
rect 45060 3992 45066 4004
rect 45646 3992 45652 4004
rect 45060 3964 45652 3992
rect 45060 3952 45066 3964
rect 45646 3952 45652 3964
rect 45704 3952 45710 4004
rect 51074 3952 51080 4004
rect 51132 3992 51138 4004
rect 51994 3992 52000 4004
rect 51132 3964 52000 3992
rect 51132 3952 51138 3964
rect 51994 3952 52000 3964
rect 52052 3952 52058 4004
rect 57146 3952 57152 4004
rect 57204 3992 57210 4004
rect 57330 3992 57336 4004
rect 57204 3964 57336 3992
rect 57204 3952 57210 3964
rect 57330 3952 57336 3964
rect 57388 3952 57394 4004
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 3510 3924 3516 3936
rect 2832 3896 3516 3924
rect 2832 3884 2838 3896
rect 3510 3884 3516 3896
rect 3568 3884 3574 3936
rect 1104 3834 72864 3856
rect 1104 3782 9078 3834
rect 9130 3782 21078 3834
rect 21130 3782 33078 3834
rect 33130 3782 45078 3834
rect 45130 3782 57078 3834
rect 57130 3782 69078 3834
rect 69130 3782 72864 3834
rect 1104 3760 72864 3782
rect 1118 3680 1124 3732
rect 1176 3720 1182 3732
rect 2501 3723 2559 3729
rect 2501 3720 2513 3723
rect 1176 3692 2513 3720
rect 1176 3680 1182 3692
rect 2501 3689 2513 3692
rect 2547 3689 2559 3723
rect 2501 3683 2559 3689
rect 62942 3680 62948 3732
rect 63000 3720 63006 3732
rect 64690 3720 64696 3732
rect 63000 3692 64696 3720
rect 63000 3680 63006 3692
rect 64690 3680 64696 3692
rect 64748 3680 64754 3732
rect 1394 3612 1400 3664
rect 1452 3652 1458 3664
rect 2777 3655 2835 3661
rect 2777 3652 2789 3655
rect 1452 3624 2789 3652
rect 1452 3612 1458 3624
rect 2777 3621 2789 3624
rect 2823 3621 2835 3655
rect 2777 3615 2835 3621
rect 28442 3612 28448 3664
rect 28500 3652 28506 3664
rect 30466 3652 30472 3664
rect 28500 3624 30472 3652
rect 28500 3612 28506 3624
rect 30466 3612 30472 3624
rect 30524 3612 30530 3664
rect 1670 3544 1676 3596
rect 1728 3584 1734 3596
rect 3053 3587 3111 3593
rect 3053 3584 3065 3587
rect 1728 3556 3065 3584
rect 1728 3544 1734 3556
rect 3053 3553 3065 3556
rect 3099 3553 3111 3587
rect 3053 3547 3111 3553
rect 25406 3544 25412 3596
rect 25464 3584 25470 3596
rect 27430 3584 27436 3596
rect 25464 3556 27436 3584
rect 25464 3544 25470 3556
rect 27430 3544 27436 3556
rect 27488 3544 27494 3596
rect 28166 3544 28172 3596
rect 28224 3584 28230 3596
rect 30190 3584 30196 3596
rect 28224 3556 30196 3584
rect 28224 3544 28230 3556
rect 30190 3544 30196 3556
rect 30248 3544 30254 3596
rect 65702 3544 65708 3596
rect 65760 3584 65766 3596
rect 67450 3584 67456 3596
rect 65760 3556 67456 3584
rect 65760 3544 65766 3556
rect 67450 3544 67456 3556
rect 67508 3544 67514 3596
rect 1946 3476 1952 3528
rect 2004 3516 2010 3528
rect 3329 3519 3387 3525
rect 3329 3516 3341 3519
rect 2004 3488 3341 3516
rect 2004 3476 2010 3488
rect 3329 3485 3341 3488
rect 3375 3485 3387 3519
rect 3329 3479 3387 3485
rect 24578 3476 24584 3528
rect 24636 3516 24642 3528
rect 26326 3516 26332 3528
rect 24636 3488 26332 3516
rect 24636 3476 24642 3488
rect 26326 3476 26332 3488
rect 26384 3476 26390 3528
rect 27890 3476 27896 3528
rect 27948 3516 27954 3528
rect 29914 3516 29920 3528
rect 27948 3488 29920 3516
rect 27948 3476 27954 3488
rect 29914 3476 29920 3488
rect 29972 3476 29978 3528
rect 64598 3476 64604 3528
rect 64656 3516 64662 3528
rect 66346 3516 66352 3528
rect 64656 3488 66352 3516
rect 64656 3476 64662 3488
rect 66346 3476 66352 3488
rect 66404 3476 66410 3528
rect 14918 3408 14924 3460
rect 14976 3448 14982 3460
rect 16114 3448 16120 3460
rect 14976 3420 16120 3448
rect 14976 3408 14982 3420
rect 16114 3408 16120 3420
rect 16172 3408 16178 3460
rect 17678 3408 17684 3460
rect 17736 3448 17742 3460
rect 19150 3448 19156 3460
rect 17736 3420 19156 3448
rect 17736 3408 17742 3420
rect 19150 3408 19156 3420
rect 19208 3408 19214 3460
rect 21542 3408 21548 3460
rect 21600 3448 21606 3460
rect 23290 3448 23296 3460
rect 21600 3420 23296 3448
rect 21600 3408 21606 3420
rect 23290 3408 23296 3420
rect 23348 3408 23354 3460
rect 23474 3408 23480 3460
rect 23532 3448 23538 3460
rect 25222 3448 25228 3460
rect 23532 3420 25228 3448
rect 23532 3408 23538 3420
rect 25222 3408 25228 3420
rect 25280 3408 25286 3460
rect 28994 3408 29000 3460
rect 29052 3448 29058 3460
rect 31018 3448 31024 3460
rect 29052 3420 31024 3448
rect 29052 3408 29058 3420
rect 31018 3408 31024 3420
rect 31076 3408 31082 3460
rect 56318 3408 56324 3460
rect 56376 3448 56382 3460
rect 57330 3448 57336 3460
rect 56376 3420 57336 3448
rect 56376 3408 56382 3420
rect 57330 3408 57336 3420
rect 57388 3408 57394 3460
rect 59906 3408 59912 3460
rect 59964 3448 59970 3460
rect 61378 3448 61384 3460
rect 59964 3420 61384 3448
rect 59964 3408 59970 3420
rect 61378 3408 61384 3420
rect 61436 3408 61442 3460
rect 61562 3408 61568 3460
rect 61620 3448 61626 3460
rect 62942 3448 62948 3460
rect 61620 3420 62948 3448
rect 61620 3408 61626 3420
rect 62942 3408 62948 3420
rect 63000 3408 63006 3460
rect 65978 3408 65984 3460
rect 66036 3448 66042 3460
rect 67726 3448 67732 3460
rect 66036 3420 67732 3448
rect 66036 3408 66042 3420
rect 67726 3408 67732 3420
rect 67784 3408 67790 3460
rect 14642 3340 14648 3392
rect 14700 3380 14706 3392
rect 15838 3380 15844 3392
rect 14700 3352 15844 3380
rect 14700 3340 14706 3352
rect 15838 3340 15844 3352
rect 15896 3340 15902 3392
rect 17954 3340 17960 3392
rect 18012 3380 18018 3392
rect 19426 3380 19432 3392
rect 18012 3352 19432 3380
rect 18012 3340 18018 3352
rect 19426 3340 19432 3352
rect 19484 3340 19490 3392
rect 20162 3340 20168 3392
rect 20220 3380 20226 3392
rect 21634 3380 21640 3392
rect 20220 3352 21640 3380
rect 20220 3340 20226 3352
rect 21634 3340 21640 3352
rect 21692 3340 21698 3392
rect 21818 3340 21824 3392
rect 21876 3380 21882 3392
rect 23566 3380 23572 3392
rect 21876 3352 23572 3380
rect 21876 3340 21882 3352
rect 23566 3340 23572 3352
rect 23624 3340 23630 3392
rect 24302 3340 24308 3392
rect 24360 3380 24366 3392
rect 26050 3380 26056 3392
rect 24360 3352 26056 3380
rect 24360 3340 24366 3352
rect 26050 3340 26056 3352
rect 26108 3340 26114 3392
rect 26234 3340 26240 3392
rect 26292 3380 26298 3392
rect 28258 3380 28264 3392
rect 26292 3352 28264 3380
rect 26292 3340 26298 3352
rect 28258 3340 28264 3352
rect 28316 3340 28322 3392
rect 28718 3340 28724 3392
rect 28776 3380 28782 3392
rect 30742 3380 30748 3392
rect 28776 3352 30748 3380
rect 28776 3340 28782 3352
rect 30742 3340 30748 3352
rect 30800 3340 30806 3392
rect 61286 3340 61292 3392
rect 61344 3380 61350 3392
rect 62758 3380 62764 3392
rect 61344 3352 62764 3380
rect 61344 3340 61350 3352
rect 62758 3340 62764 3352
rect 62816 3340 62822 3392
rect 65426 3340 65432 3392
rect 65484 3380 65490 3392
rect 67174 3380 67180 3392
rect 65484 3352 67180 3380
rect 65484 3340 65490 3352
rect 67174 3340 67180 3352
rect 67232 3340 67238 3392
rect 1104 3290 72864 3312
rect 1104 3238 3078 3290
rect 3130 3238 15078 3290
rect 15130 3238 27078 3290
rect 27130 3238 39078 3290
rect 39130 3238 51078 3290
rect 51130 3238 63078 3290
rect 63130 3238 72864 3290
rect 1104 3216 72864 3238
rect 11882 3136 11888 3188
rect 11940 3176 11946 3188
rect 13078 3176 13084 3188
rect 11940 3148 13084 3176
rect 11940 3136 11946 3148
rect 13078 3136 13084 3148
rect 13136 3136 13142 3188
rect 14366 3136 14372 3188
rect 14424 3176 14430 3188
rect 14424 3148 15608 3176
rect 14424 3136 14430 3148
rect 4154 3068 4160 3120
rect 4212 3108 4218 3120
rect 4212 3080 5028 3108
rect 4212 3068 4218 3080
rect 2222 3040 2228 3052
rect 2183 3012 2228 3040
rect 2222 3000 2228 3012
rect 2280 3000 2286 3052
rect 2498 3040 2504 3052
rect 2459 3012 2504 3040
rect 2498 3000 2504 3012
rect 2556 3000 2562 3052
rect 2774 3040 2780 3052
rect 2735 3012 2780 3040
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 3602 3000 3608 3052
rect 3660 3040 3666 3052
rect 5000 3049 5028 3080
rect 5258 3068 5264 3120
rect 5316 3108 5322 3120
rect 5316 3080 6132 3108
rect 5316 3068 5322 3080
rect 4433 3043 4491 3049
rect 4433 3040 4445 3043
rect 3660 3012 4445 3040
rect 3660 3000 3666 3012
rect 4433 3009 4445 3012
rect 4479 3009 4491 3043
rect 4433 3003 4491 3009
rect 4985 3043 5043 3049
rect 4985 3009 4997 3043
rect 5031 3009 5043 3043
rect 4985 3003 5043 3009
rect 5074 3000 5080 3052
rect 5132 3040 5138 3052
rect 6104 3049 6132 3080
rect 6362 3068 6368 3120
rect 6420 3108 6426 3120
rect 6420 3080 7328 3108
rect 6420 3068 6426 3080
rect 5813 3043 5871 3049
rect 5813 3040 5825 3043
rect 5132 3012 5825 3040
rect 5132 3000 5138 3012
rect 5813 3009 5825 3012
rect 5859 3009 5871 3043
rect 5813 3003 5871 3009
rect 6089 3043 6147 3049
rect 6089 3009 6101 3043
rect 6135 3009 6147 3043
rect 6089 3003 6147 3009
rect 6178 3000 6184 3052
rect 6236 3040 6242 3052
rect 7300 3049 7328 3080
rect 8294 3068 8300 3120
rect 8352 3108 8358 3120
rect 8352 3080 9260 3108
rect 8352 3068 8358 3080
rect 7009 3043 7067 3049
rect 7009 3040 7021 3043
rect 6236 3012 7021 3040
rect 6236 3000 6242 3012
rect 7009 3009 7021 3012
rect 7055 3009 7067 3043
rect 7009 3003 7067 3009
rect 7285 3043 7343 3049
rect 7285 3009 7297 3043
rect 7331 3009 7343 3043
rect 7285 3003 7343 3009
rect 7466 3000 7472 3052
rect 7524 3040 7530 3052
rect 9232 3049 9260 3080
rect 9398 3068 9404 3120
rect 9456 3108 9462 3120
rect 9456 3080 10364 3108
rect 9456 3068 9462 3080
rect 8389 3043 8447 3049
rect 8389 3040 8401 3043
rect 7524 3012 8401 3040
rect 7524 3000 7530 3012
rect 8389 3009 8401 3012
rect 8435 3009 8447 3043
rect 8389 3003 8447 3009
rect 9217 3043 9275 3049
rect 9217 3009 9229 3043
rect 9263 3009 9275 3043
rect 10042 3040 10048 3052
rect 10003 3012 10048 3040
rect 9217 3003 9275 3009
rect 10042 3000 10048 3012
rect 10100 3000 10106 3052
rect 10336 3049 10364 3080
rect 11330 3068 11336 3120
rect 11388 3108 11394 3120
rect 11388 3080 12572 3108
rect 11388 3068 11394 3080
rect 10321 3043 10379 3049
rect 10321 3009 10333 3043
rect 10367 3009 10379 3043
rect 10321 3003 10379 3009
rect 10502 3000 10508 3052
rect 10560 3040 10566 3052
rect 12544 3049 12572 3080
rect 12710 3068 12716 3120
rect 12768 3108 12774 3120
rect 13170 3108 13176 3120
rect 12768 3080 13176 3108
rect 12768 3068 12774 3080
rect 13170 3068 13176 3080
rect 13228 3068 13234 3120
rect 13262 3068 13268 3120
rect 13320 3108 13326 3120
rect 13320 3080 14504 3108
rect 13320 3068 13326 3080
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 10560 3012 11713 3040
rect 10560 3000 10566 3012
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 12529 3043 12587 3049
rect 12529 3009 12541 3043
rect 12575 3009 12587 3043
rect 12529 3003 12587 3009
rect 12986 3000 12992 3052
rect 13044 3040 13050 3052
rect 14476 3049 14504 3080
rect 15580 3049 15608 3148
rect 16850 3136 16856 3188
rect 16908 3176 16914 3188
rect 16908 3148 18368 3176
rect 16908 3136 16914 3148
rect 16298 3068 16304 3120
rect 16356 3108 16362 3120
rect 16356 3080 17816 3108
rect 16356 3068 16362 3080
rect 14185 3043 14243 3049
rect 14185 3040 14197 3043
rect 13044 3012 14197 3040
rect 13044 3000 13050 3012
rect 14185 3009 14197 3012
rect 14231 3009 14243 3043
rect 14185 3003 14243 3009
rect 14461 3043 14519 3049
rect 14461 3009 14473 3043
rect 14507 3009 14519 3043
rect 14461 3003 14519 3009
rect 15565 3043 15623 3049
rect 15565 3009 15577 3043
rect 15611 3009 15623 3043
rect 15565 3003 15623 3009
rect 15746 3000 15752 3052
rect 15804 3040 15810 3052
rect 17788 3049 17816 3080
rect 18340 3049 18368 3148
rect 19334 3136 19340 3188
rect 19392 3176 19398 3188
rect 19392 3148 20116 3176
rect 19392 3136 19398 3148
rect 18506 3068 18512 3120
rect 18564 3108 18570 3120
rect 18564 3080 20024 3108
rect 18564 3068 18570 3080
rect 17221 3043 17279 3049
rect 17221 3040 17233 3043
rect 15804 3012 17233 3040
rect 15804 3000 15810 3012
rect 17221 3009 17233 3012
rect 17267 3009 17279 3043
rect 17221 3003 17279 3009
rect 17773 3043 17831 3049
rect 17773 3009 17785 3043
rect 17819 3009 17831 3043
rect 17773 3003 17831 3009
rect 18325 3043 18383 3049
rect 18325 3009 18337 3043
rect 18371 3009 18383 3043
rect 19150 3040 19156 3052
rect 19111 3012 19156 3040
rect 18325 3003 18383 3009
rect 19150 3000 19156 3012
rect 19208 3000 19214 3052
rect 19426 3040 19432 3052
rect 19387 3012 19432 3040
rect 19426 3000 19432 3012
rect 19484 3000 19490 3052
rect 19996 3049 20024 3080
rect 19981 3043 20039 3049
rect 19981 3009 19993 3043
rect 20027 3009 20039 3043
rect 20088 3040 20116 3148
rect 20438 3136 20444 3188
rect 20496 3176 20502 3188
rect 20496 3148 22232 3176
rect 20496 3136 20502 3148
rect 20162 3068 20168 3120
rect 20220 3108 20226 3120
rect 20220 3080 21404 3108
rect 20220 3068 20226 3080
rect 21376 3049 21404 3080
rect 20809 3043 20867 3049
rect 20809 3040 20821 3043
rect 20088 3012 20821 3040
rect 19981 3003 20039 3009
rect 20809 3009 20821 3012
rect 20855 3009 20867 3043
rect 20809 3003 20867 3009
rect 21361 3043 21419 3049
rect 21361 3009 21373 3043
rect 21407 3009 21419 3043
rect 21634 3040 21640 3052
rect 21595 3012 21640 3040
rect 21361 3003 21419 3009
rect 21634 3000 21640 3012
rect 21692 3000 21698 3052
rect 22204 3049 22232 3148
rect 22922 3136 22928 3188
rect 22980 3176 22986 3188
rect 22980 3148 24716 3176
rect 22980 3136 22986 3148
rect 22278 3068 22284 3120
rect 22336 3108 22342 3120
rect 22336 3080 23888 3108
rect 22336 3068 22342 3080
rect 22189 3043 22247 3049
rect 22189 3009 22201 3043
rect 22235 3009 22247 3043
rect 22189 3003 22247 3009
rect 22370 3000 22376 3052
rect 22428 3040 22434 3052
rect 23290 3040 23296 3052
rect 22428 3012 23152 3040
rect 23251 3012 23296 3040
rect 22428 3000 22434 3012
rect 2133 2975 2191 2981
rect 2133 2941 2145 2975
rect 2179 2972 2191 2975
rect 2406 2972 2412 2984
rect 2179 2944 2412 2972
rect 2179 2941 2191 2944
rect 2133 2935 2191 2941
rect 2406 2932 2412 2944
rect 2464 2932 2470 2984
rect 3326 2932 3332 2984
rect 3384 2932 3390 2984
rect 3878 2932 3884 2984
rect 3936 2972 3942 2984
rect 4709 2975 4767 2981
rect 4709 2972 4721 2975
rect 3936 2944 4721 2972
rect 3936 2932 3942 2944
rect 4709 2941 4721 2944
rect 4755 2941 4767 2975
rect 4709 2935 4767 2941
rect 5534 2932 5540 2984
rect 5592 2972 5598 2984
rect 6457 2975 6515 2981
rect 6457 2972 6469 2975
rect 5592 2944 6469 2972
rect 5592 2932 5598 2944
rect 6457 2941 6469 2944
rect 6503 2941 6515 2975
rect 6457 2935 6515 2941
rect 6638 2932 6644 2984
rect 6696 2972 6702 2984
rect 7561 2975 7619 2981
rect 7561 2972 7573 2975
rect 6696 2944 7573 2972
rect 6696 2932 6702 2944
rect 7561 2941 7573 2944
rect 7607 2941 7619 2975
rect 7561 2935 7619 2941
rect 7742 2932 7748 2984
rect 7800 2972 7806 2984
rect 8665 2975 8723 2981
rect 8665 2972 8677 2975
rect 7800 2944 8677 2972
rect 7800 2932 7806 2944
rect 8665 2941 8677 2944
rect 8711 2941 8723 2975
rect 8665 2935 8723 2941
rect 8846 2932 8852 2984
rect 8904 2972 8910 2984
rect 9769 2975 9827 2981
rect 9769 2972 9781 2975
rect 8904 2944 9781 2972
rect 8904 2932 8910 2944
rect 9769 2941 9781 2944
rect 9815 2941 9827 2975
rect 9769 2935 9827 2941
rect 9950 2932 9956 2984
rect 10008 2972 10014 2984
rect 10873 2975 10931 2981
rect 10873 2972 10885 2975
rect 10008 2944 10885 2972
rect 10008 2932 10014 2944
rect 10873 2941 10885 2944
rect 10919 2941 10931 2975
rect 10873 2935 10931 2941
rect 11054 2932 11060 2984
rect 11112 2972 11118 2984
rect 12253 2975 12311 2981
rect 12253 2972 12265 2975
rect 11112 2944 12265 2972
rect 11112 2932 11118 2944
rect 12253 2941 12265 2944
rect 12299 2941 12311 2975
rect 12253 2935 12311 2941
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 13633 2975 13691 2981
rect 13633 2972 13645 2975
rect 12492 2944 13645 2972
rect 12492 2932 12498 2944
rect 13633 2941 13645 2944
rect 13679 2941 13691 2975
rect 13633 2935 13691 2941
rect 13814 2932 13820 2984
rect 13872 2972 13878 2984
rect 15013 2975 15071 2981
rect 15013 2972 15025 2975
rect 13872 2944 15025 2972
rect 13872 2932 13878 2944
rect 15013 2941 15025 2944
rect 15059 2941 15071 2975
rect 15013 2935 15071 2941
rect 15470 2932 15476 2984
rect 15528 2972 15534 2984
rect 16945 2975 17003 2981
rect 16945 2972 16957 2975
rect 15528 2944 16957 2972
rect 15528 2932 15534 2944
rect 16945 2941 16957 2944
rect 16991 2941 17003 2975
rect 16945 2935 17003 2941
rect 17126 2932 17132 2984
rect 17184 2972 17190 2984
rect 18601 2975 18659 2981
rect 18601 2972 18613 2975
rect 17184 2944 18613 2972
rect 17184 2932 17190 2944
rect 18601 2941 18613 2944
rect 18647 2941 18659 2975
rect 18601 2935 18659 2941
rect 18782 2932 18788 2984
rect 18840 2972 18846 2984
rect 20257 2975 20315 2981
rect 20257 2972 20269 2975
rect 18840 2944 20269 2972
rect 18840 2932 18846 2944
rect 20257 2941 20269 2944
rect 20303 2941 20315 2975
rect 20257 2935 20315 2941
rect 21266 2932 21272 2984
rect 21324 2972 21330 2984
rect 21913 2975 21971 2981
rect 21913 2972 21925 2975
rect 21324 2944 21925 2972
rect 21324 2932 21330 2944
rect 21913 2941 21925 2944
rect 21959 2941 21971 2975
rect 22738 2972 22744 2984
rect 22699 2944 22744 2972
rect 21913 2935 21971 2941
rect 22738 2932 22744 2944
rect 22796 2932 22802 2984
rect 23124 2972 23152 3012
rect 23290 3000 23296 3012
rect 23348 3000 23354 3052
rect 23566 3040 23572 3052
rect 23527 3012 23572 3040
rect 23566 3000 23572 3012
rect 23624 3000 23630 3052
rect 23860 3049 23888 3080
rect 23845 3043 23903 3049
rect 23845 3009 23857 3043
rect 23891 3009 23903 3043
rect 23845 3003 23903 3009
rect 23934 3000 23940 3052
rect 23992 3040 23998 3052
rect 24688 3049 24716 3148
rect 29270 3136 29276 3188
rect 29328 3176 29334 3188
rect 31294 3176 31300 3188
rect 29328 3148 31300 3176
rect 29328 3136 29334 3148
rect 31294 3136 31300 3148
rect 31352 3136 31358 3188
rect 54386 3136 54392 3188
rect 54444 3176 54450 3188
rect 54444 3148 55628 3176
rect 54444 3136 54450 3148
rect 24854 3068 24860 3120
rect 24912 3108 24918 3120
rect 24912 3080 26648 3108
rect 24912 3068 24918 3080
rect 24673 3043 24731 3049
rect 23992 3012 24624 3040
rect 23992 3000 23998 3012
rect 24121 2975 24179 2981
rect 24121 2972 24133 2975
rect 23124 2944 24133 2972
rect 24121 2941 24133 2944
rect 24167 2941 24179 2975
rect 24121 2935 24179 2941
rect 24210 2932 24216 2984
rect 24268 2972 24274 2984
rect 24596 2972 24624 3012
rect 24673 3009 24685 3043
rect 24719 3009 24731 3043
rect 25222 3040 25228 3052
rect 25183 3012 25228 3040
rect 24673 3003 24731 3009
rect 25222 3000 25228 3012
rect 25280 3000 25286 3052
rect 26050 3040 26056 3052
rect 26011 3012 26056 3040
rect 26050 3000 26056 3012
rect 26108 3000 26114 3052
rect 26326 3040 26332 3052
rect 26287 3012 26332 3040
rect 26326 3000 26332 3012
rect 26384 3000 26390 3052
rect 26620 3049 26648 3080
rect 26786 3068 26792 3120
rect 26844 3108 26850 3120
rect 26844 3080 28856 3108
rect 26844 3068 26850 3080
rect 26605 3043 26663 3049
rect 26605 3009 26617 3043
rect 26651 3009 26663 3043
rect 26878 3040 26884 3052
rect 26839 3012 26884 3040
rect 26605 3003 26663 3009
rect 26878 3000 26884 3012
rect 26936 3000 26942 3052
rect 27430 3040 27436 3052
rect 27391 3012 27436 3040
rect 27430 3000 27436 3012
rect 27488 3000 27494 3052
rect 27522 3000 27528 3052
rect 27580 3040 27586 3052
rect 28258 3040 28264 3052
rect 27580 3012 28120 3040
rect 28219 3012 28264 3040
rect 27580 3000 27586 3012
rect 25501 2975 25559 2981
rect 25501 2972 25513 2975
rect 24268 2944 24532 2972
rect 24596 2944 25513 2972
rect 24268 2932 24274 2944
rect 566 2864 572 2916
rect 624 2904 630 2916
rect 3053 2907 3111 2913
rect 3053 2904 3065 2907
rect 624 2876 3065 2904
rect 624 2864 630 2876
rect 3053 2873 3065 2876
rect 3099 2873 3111 2907
rect 3344 2904 3372 2932
rect 4157 2907 4215 2913
rect 4157 2904 4169 2907
rect 3344 2876 4169 2904
rect 3053 2867 3111 2873
rect 4157 2873 4169 2876
rect 4203 2873 4215 2907
rect 4157 2867 4215 2873
rect 4430 2864 4436 2916
rect 4488 2904 4494 2916
rect 5261 2907 5319 2913
rect 5261 2904 5273 2907
rect 4488 2876 5273 2904
rect 4488 2864 4494 2876
rect 5261 2873 5273 2876
rect 5307 2873 5319 2907
rect 5261 2867 5319 2873
rect 5810 2864 5816 2916
rect 5868 2904 5874 2916
rect 6733 2907 6791 2913
rect 6733 2904 6745 2907
rect 5868 2876 6745 2904
rect 5868 2864 5874 2876
rect 6733 2873 6745 2876
rect 6779 2873 6791 2907
rect 6733 2867 6791 2873
rect 6914 2864 6920 2916
rect 6972 2904 6978 2916
rect 7650 2904 7656 2916
rect 6972 2876 7656 2904
rect 6972 2864 6978 2876
rect 7650 2864 7656 2876
rect 7708 2864 7714 2916
rect 8113 2907 8171 2913
rect 8113 2904 8125 2907
rect 7760 2876 8125 2904
rect 842 2796 848 2848
rect 900 2836 906 2848
rect 3329 2839 3387 2845
rect 3329 2836 3341 2839
rect 900 2808 3341 2836
rect 900 2796 906 2808
rect 3329 2805 3341 2808
rect 3375 2805 3387 2839
rect 3329 2799 3387 2805
rect 3510 2796 3516 2848
rect 3568 2836 3574 2848
rect 3605 2839 3663 2845
rect 3605 2836 3617 2839
rect 3568 2808 3617 2836
rect 3568 2796 3574 2808
rect 3605 2805 3617 2808
rect 3651 2805 3663 2839
rect 3605 2799 3663 2805
rect 3786 2796 3792 2848
rect 3844 2836 3850 2848
rect 3881 2839 3939 2845
rect 3881 2836 3893 2839
rect 3844 2808 3893 2836
rect 3844 2796 3850 2808
rect 3881 2805 3893 2808
rect 3927 2805 3939 2839
rect 3881 2799 3939 2805
rect 4706 2796 4712 2848
rect 4764 2836 4770 2848
rect 5537 2839 5595 2845
rect 5537 2836 5549 2839
rect 4764 2808 5549 2836
rect 4764 2796 4770 2808
rect 5537 2805 5549 2808
rect 5583 2805 5595 2839
rect 5537 2799 5595 2805
rect 7190 2796 7196 2848
rect 7248 2836 7254 2848
rect 7760 2836 7788 2876
rect 8113 2873 8125 2876
rect 8159 2873 8171 2907
rect 8113 2867 8171 2873
rect 8570 2864 8576 2916
rect 8628 2904 8634 2916
rect 9493 2907 9551 2913
rect 9493 2904 9505 2907
rect 8628 2876 9505 2904
rect 8628 2864 8634 2876
rect 9493 2873 9505 2876
rect 9539 2873 9551 2907
rect 9493 2867 9551 2873
rect 9674 2864 9680 2916
rect 9732 2904 9738 2916
rect 10597 2907 10655 2913
rect 10597 2904 10609 2907
rect 9732 2876 10609 2904
rect 9732 2864 9738 2876
rect 10597 2873 10609 2876
rect 10643 2873 10655 2907
rect 10597 2867 10655 2873
rect 10778 2864 10784 2916
rect 10836 2904 10842 2916
rect 11977 2907 12035 2913
rect 11977 2904 11989 2907
rect 10836 2876 11989 2904
rect 10836 2864 10842 2876
rect 11977 2873 11989 2876
rect 12023 2873 12035 2907
rect 11977 2867 12035 2873
rect 12158 2864 12164 2916
rect 12216 2904 12222 2916
rect 13357 2907 13415 2913
rect 13357 2904 13369 2907
rect 12216 2876 13369 2904
rect 12216 2864 12222 2876
rect 13357 2873 13369 2876
rect 13403 2873 13415 2907
rect 13357 2867 13415 2873
rect 13538 2864 13544 2916
rect 13596 2904 13602 2916
rect 14737 2907 14795 2913
rect 14737 2904 14749 2907
rect 13596 2876 14749 2904
rect 13596 2864 13602 2876
rect 14737 2873 14749 2876
rect 14783 2873 14795 2907
rect 14737 2867 14795 2873
rect 15194 2864 15200 2916
rect 15252 2904 15258 2916
rect 16393 2907 16451 2913
rect 16393 2904 16405 2907
rect 15252 2876 16405 2904
rect 15252 2864 15258 2876
rect 16393 2873 16405 2876
rect 16439 2873 16451 2907
rect 16393 2867 16451 2873
rect 16574 2864 16580 2916
rect 16632 2904 16638 2916
rect 18049 2907 18107 2913
rect 18049 2904 18061 2907
rect 16632 2876 18061 2904
rect 16632 2864 16638 2876
rect 18049 2873 18061 2876
rect 18095 2873 18107 2907
rect 18877 2907 18935 2913
rect 18877 2904 18889 2907
rect 18049 2867 18107 2873
rect 18156 2876 18889 2904
rect 7248 2808 7788 2836
rect 7248 2796 7254 2808
rect 7834 2796 7840 2848
rect 7892 2836 7898 2848
rect 7892 2808 7937 2836
rect 7892 2796 7898 2808
rect 8018 2796 8024 2848
rect 8076 2836 8082 2848
rect 8941 2839 8999 2845
rect 8941 2836 8953 2839
rect 8076 2808 8953 2836
rect 8076 2796 8082 2808
rect 8941 2805 8953 2808
rect 8987 2805 8999 2839
rect 8941 2799 8999 2805
rect 10226 2796 10232 2848
rect 10284 2836 10290 2848
rect 11149 2839 11207 2845
rect 11149 2836 11161 2839
rect 10284 2808 11161 2836
rect 10284 2796 10290 2808
rect 11149 2805 11161 2808
rect 11195 2805 11207 2839
rect 11149 2799 11207 2805
rect 11606 2796 11612 2848
rect 11664 2836 11670 2848
rect 12805 2839 12863 2845
rect 12805 2836 12817 2839
rect 11664 2808 12817 2836
rect 11664 2796 11670 2808
rect 12805 2805 12817 2808
rect 12851 2805 12863 2839
rect 13078 2836 13084 2848
rect 13039 2808 13084 2836
rect 12805 2799 12863 2805
rect 13078 2796 13084 2808
rect 13136 2796 13142 2848
rect 13170 2796 13176 2848
rect 13228 2836 13234 2848
rect 13909 2839 13967 2845
rect 13909 2836 13921 2839
rect 13228 2808 13921 2836
rect 13228 2796 13234 2808
rect 13909 2805 13921 2808
rect 13955 2805 13967 2839
rect 13909 2799 13967 2805
rect 14090 2796 14096 2848
rect 14148 2836 14154 2848
rect 15289 2839 15347 2845
rect 15289 2836 15301 2839
rect 14148 2808 15301 2836
rect 14148 2796 14154 2808
rect 15289 2805 15301 2808
rect 15335 2805 15347 2839
rect 15838 2836 15844 2848
rect 15799 2808 15844 2836
rect 15289 2799 15347 2805
rect 15838 2796 15844 2808
rect 15896 2796 15902 2848
rect 16114 2836 16120 2848
rect 16075 2808 16120 2836
rect 16114 2796 16120 2808
rect 16172 2796 16178 2848
rect 17494 2836 17500 2848
rect 17455 2808 17500 2836
rect 17494 2796 17500 2808
rect 17552 2796 17558 2848
rect 17586 2796 17592 2848
rect 17644 2836 17650 2848
rect 18156 2836 18184 2876
rect 18877 2873 18889 2876
rect 18923 2873 18935 2907
rect 18877 2867 18935 2873
rect 19058 2864 19064 2916
rect 19116 2904 19122 2916
rect 20533 2907 20591 2913
rect 20533 2904 20545 2907
rect 19116 2876 20545 2904
rect 19116 2864 19122 2876
rect 20533 2873 20545 2876
rect 20579 2873 20591 2907
rect 20533 2867 20591 2873
rect 20714 2864 20720 2916
rect 20772 2904 20778 2916
rect 22465 2907 22523 2913
rect 22465 2904 22477 2907
rect 20772 2876 22477 2904
rect 20772 2864 20778 2876
rect 22465 2873 22477 2876
rect 22511 2873 22523 2907
rect 22465 2867 22523 2873
rect 22646 2864 22652 2916
rect 22704 2904 22710 2916
rect 24397 2907 24455 2913
rect 24397 2904 24409 2907
rect 22704 2876 24409 2904
rect 22704 2864 22710 2876
rect 24397 2873 24409 2876
rect 24443 2873 24455 2907
rect 24504 2904 24532 2944
rect 25501 2941 25513 2944
rect 25547 2941 25559 2975
rect 25501 2935 25559 2941
rect 25958 2932 25964 2984
rect 26016 2972 26022 2984
rect 27985 2975 28043 2981
rect 27985 2972 27997 2975
rect 26016 2944 27997 2972
rect 26016 2932 26022 2944
rect 27985 2941 27997 2944
rect 28031 2941 28043 2975
rect 28092 2972 28120 3012
rect 28258 3000 28264 3012
rect 28316 3000 28322 3052
rect 28828 3049 28856 3080
rect 29822 3068 29828 3120
rect 29880 3108 29886 3120
rect 29880 3080 32352 3108
rect 29880 3068 29886 3080
rect 28813 3043 28871 3049
rect 28813 3009 28825 3043
rect 28859 3009 28871 3043
rect 29086 3040 29092 3052
rect 29047 3012 29092 3040
rect 28813 3003 28871 3009
rect 29086 3000 29092 3012
rect 29144 3000 29150 3052
rect 29914 3040 29920 3052
rect 29875 3012 29920 3040
rect 29914 3000 29920 3012
rect 29972 3000 29978 3052
rect 30190 3040 30196 3052
rect 30151 3012 30196 3040
rect 30190 3000 30196 3012
rect 30248 3000 30254 3052
rect 30374 3000 30380 3052
rect 30432 3040 30438 3052
rect 32324 3049 32352 3080
rect 48314 3068 48320 3120
rect 48372 3108 48378 3120
rect 48372 3080 49280 3108
rect 48372 3068 48378 3080
rect 32033 3043 32091 3049
rect 32033 3040 32045 3043
rect 30432 3012 32045 3040
rect 30432 3000 30438 3012
rect 32033 3009 32045 3012
rect 32079 3009 32091 3043
rect 32033 3003 32091 3009
rect 32309 3043 32367 3049
rect 32309 3009 32321 3043
rect 32355 3009 32367 3043
rect 32309 3003 32367 3009
rect 36170 3000 36176 3052
rect 36228 3040 36234 3052
rect 36265 3043 36323 3049
rect 36265 3040 36277 3043
rect 36228 3012 36277 3040
rect 36228 3000 36234 3012
rect 36265 3009 36277 3012
rect 36311 3009 36323 3043
rect 36265 3003 36323 3009
rect 36446 3000 36452 3052
rect 36504 3040 36510 3052
rect 36541 3043 36599 3049
rect 36541 3040 36553 3043
rect 36504 3012 36553 3040
rect 36504 3000 36510 3012
rect 36541 3009 36553 3012
rect 36587 3009 36599 3043
rect 36541 3003 36599 3009
rect 36998 3000 37004 3052
rect 37056 3040 37062 3052
rect 37093 3043 37151 3049
rect 37093 3040 37105 3043
rect 37056 3012 37105 3040
rect 37056 3000 37062 3012
rect 37093 3009 37105 3012
rect 37139 3009 37151 3043
rect 37093 3003 37151 3009
rect 37274 3000 37280 3052
rect 37332 3040 37338 3052
rect 37369 3043 37427 3049
rect 37369 3040 37381 3043
rect 37332 3012 37381 3040
rect 37332 3000 37338 3012
rect 37369 3009 37381 3012
rect 37415 3009 37427 3043
rect 37369 3003 37427 3009
rect 37550 3000 37556 3052
rect 37608 3040 37614 3052
rect 37921 3043 37979 3049
rect 37921 3040 37933 3043
rect 37608 3012 37933 3040
rect 37608 3000 37614 3012
rect 37921 3009 37933 3012
rect 37967 3009 37979 3043
rect 37921 3003 37979 3009
rect 38102 3000 38108 3052
rect 38160 3040 38166 3052
rect 38473 3043 38531 3049
rect 38473 3040 38485 3043
rect 38160 3012 38485 3040
rect 38160 3000 38166 3012
rect 38473 3009 38485 3012
rect 38519 3009 38531 3043
rect 38473 3003 38531 3009
rect 38654 3000 38660 3052
rect 38712 3040 38718 3052
rect 39025 3043 39083 3049
rect 39025 3040 39037 3043
rect 38712 3012 39037 3040
rect 38712 3000 38718 3012
rect 39025 3009 39037 3012
rect 39071 3009 39083 3043
rect 39025 3003 39083 3009
rect 39206 3000 39212 3052
rect 39264 3040 39270 3052
rect 39577 3043 39635 3049
rect 39577 3040 39589 3043
rect 39264 3012 39589 3040
rect 39264 3000 39270 3012
rect 39577 3009 39589 3012
rect 39623 3009 39635 3043
rect 39577 3003 39635 3009
rect 39758 3000 39764 3052
rect 39816 3040 39822 3052
rect 40129 3043 40187 3049
rect 40129 3040 40141 3043
rect 39816 3012 40141 3040
rect 39816 3000 39822 3012
rect 40129 3009 40141 3012
rect 40175 3009 40187 3043
rect 40129 3003 40187 3009
rect 40310 3000 40316 3052
rect 40368 3040 40374 3052
rect 40681 3043 40739 3049
rect 40681 3040 40693 3043
rect 40368 3012 40693 3040
rect 40368 3000 40374 3012
rect 40681 3009 40693 3012
rect 40727 3009 40739 3043
rect 40681 3003 40739 3009
rect 40862 3000 40868 3052
rect 40920 3040 40926 3052
rect 41233 3043 41291 3049
rect 41233 3040 41245 3043
rect 40920 3012 41245 3040
rect 40920 3000 40926 3012
rect 41233 3009 41245 3012
rect 41279 3009 41291 3043
rect 41233 3003 41291 3009
rect 41414 3000 41420 3052
rect 41472 3040 41478 3052
rect 41785 3043 41843 3049
rect 41785 3040 41797 3043
rect 41472 3012 41797 3040
rect 41472 3000 41478 3012
rect 41785 3009 41797 3012
rect 41831 3009 41843 3043
rect 41785 3003 41843 3009
rect 41966 3000 41972 3052
rect 42024 3040 42030 3052
rect 42337 3043 42395 3049
rect 42337 3040 42349 3043
rect 42024 3012 42349 3040
rect 42024 3000 42030 3012
rect 42337 3009 42349 3012
rect 42383 3009 42395 3043
rect 42337 3003 42395 3009
rect 42518 3000 42524 3052
rect 42576 3040 42582 3052
rect 43165 3043 43223 3049
rect 43165 3040 43177 3043
rect 42576 3012 43177 3040
rect 42576 3000 42582 3012
rect 43165 3009 43177 3012
rect 43211 3009 43223 3043
rect 43165 3003 43223 3009
rect 43346 3000 43352 3052
rect 43404 3040 43410 3052
rect 43993 3043 44051 3049
rect 43993 3040 44005 3043
rect 43404 3012 44005 3040
rect 43404 3000 43410 3012
rect 43993 3009 44005 3012
rect 44039 3009 44051 3043
rect 43993 3003 44051 3009
rect 44174 3000 44180 3052
rect 44232 3040 44238 3052
rect 44821 3043 44879 3049
rect 44821 3040 44833 3043
rect 44232 3012 44833 3040
rect 44232 3000 44238 3012
rect 44821 3009 44833 3012
rect 44867 3009 44879 3043
rect 45646 3040 45652 3052
rect 45607 3012 45652 3040
rect 44821 3003 44879 3009
rect 45646 3000 45652 3012
rect 45704 3000 45710 3052
rect 45830 3000 45836 3052
rect 45888 3040 45894 3052
rect 46477 3043 46535 3049
rect 46477 3040 46489 3043
rect 45888 3012 46489 3040
rect 45888 3000 45894 3012
rect 46477 3009 46489 3012
rect 46523 3009 46535 3043
rect 46477 3003 46535 3009
rect 46658 3000 46664 3052
rect 46716 3040 46722 3052
rect 47305 3043 47363 3049
rect 47305 3040 47317 3043
rect 46716 3012 47317 3040
rect 46716 3000 46722 3012
rect 47305 3009 47317 3012
rect 47351 3009 47363 3043
rect 47305 3003 47363 3009
rect 48038 3000 48044 3052
rect 48096 3040 48102 3052
rect 49252 3049 49280 3080
rect 50246 3068 50252 3120
rect 50304 3108 50310 3120
rect 50304 3080 51212 3108
rect 50304 3068 50310 3080
rect 48961 3043 49019 3049
rect 48961 3040 48973 3043
rect 48096 3012 48973 3040
rect 48096 3000 48102 3012
rect 48961 3009 48973 3012
rect 49007 3009 49019 3043
rect 48961 3003 49019 3009
rect 49237 3043 49295 3049
rect 49237 3009 49249 3043
rect 49283 3009 49295 3043
rect 49237 3003 49295 3009
rect 49418 3000 49424 3052
rect 49476 3040 49482 3052
rect 51184 3049 51212 3080
rect 51626 3068 51632 3120
rect 51684 3108 51690 3120
rect 51684 3080 52592 3108
rect 51684 3068 51690 3080
rect 50341 3043 50399 3049
rect 50341 3040 50353 3043
rect 49476 3012 50353 3040
rect 49476 3000 49482 3012
rect 50341 3009 50353 3012
rect 50387 3009 50399 3043
rect 50341 3003 50399 3009
rect 51169 3043 51227 3049
rect 51169 3009 51181 3043
rect 51215 3009 51227 3043
rect 51994 3040 52000 3052
rect 51955 3012 52000 3040
rect 51169 3003 51227 3009
rect 51994 3000 52000 3012
rect 52052 3000 52058 3052
rect 52564 3049 52592 3080
rect 53282 3068 53288 3120
rect 53340 3108 53346 3120
rect 53340 3080 54524 3108
rect 53340 3068 53346 3080
rect 52549 3043 52607 3049
rect 52549 3009 52561 3043
rect 52595 3009 52607 3043
rect 52549 3003 52607 3009
rect 52730 3000 52736 3052
rect 52788 3040 52794 3052
rect 53929 3043 53987 3049
rect 53929 3040 53941 3043
rect 52788 3012 53941 3040
rect 52788 3000 52794 3012
rect 53929 3009 53941 3012
rect 53975 3009 53987 3043
rect 53929 3003 53987 3009
rect 54110 3000 54116 3052
rect 54168 3040 54174 3052
rect 54496 3049 54524 3080
rect 54481 3043 54539 3049
rect 54168 3012 54432 3040
rect 54168 3000 54174 3012
rect 29365 2975 29423 2981
rect 29365 2972 29377 2975
rect 28092 2944 29377 2972
rect 27985 2935 28043 2941
rect 29365 2941 29377 2944
rect 29411 2941 29423 2975
rect 29365 2935 29423 2941
rect 30098 2932 30104 2984
rect 30156 2972 30162 2984
rect 32677 2975 32735 2981
rect 32677 2972 32689 2975
rect 30156 2944 32689 2972
rect 30156 2932 30162 2944
rect 32677 2941 32689 2944
rect 32723 2941 32735 2975
rect 32677 2935 32735 2941
rect 37826 2932 37832 2984
rect 37884 2972 37890 2984
rect 38197 2975 38255 2981
rect 38197 2972 38209 2975
rect 37884 2944 38209 2972
rect 37884 2932 37890 2944
rect 38197 2941 38209 2944
rect 38243 2941 38255 2975
rect 38197 2935 38255 2941
rect 38378 2932 38384 2984
rect 38436 2972 38442 2984
rect 38749 2975 38807 2981
rect 38749 2972 38761 2975
rect 38436 2944 38761 2972
rect 38436 2932 38442 2944
rect 38749 2941 38761 2944
rect 38795 2941 38807 2975
rect 38749 2935 38807 2941
rect 38930 2932 38936 2984
rect 38988 2972 38994 2984
rect 39301 2975 39359 2981
rect 39301 2972 39313 2975
rect 38988 2944 39313 2972
rect 38988 2932 38994 2944
rect 39301 2941 39313 2944
rect 39347 2941 39359 2975
rect 39301 2935 39359 2941
rect 39482 2932 39488 2984
rect 39540 2972 39546 2984
rect 39853 2975 39911 2981
rect 39853 2972 39865 2975
rect 39540 2944 39865 2972
rect 39540 2932 39546 2944
rect 39853 2941 39865 2944
rect 39899 2941 39911 2975
rect 39853 2935 39911 2941
rect 40034 2932 40040 2984
rect 40092 2972 40098 2984
rect 40405 2975 40463 2981
rect 40405 2972 40417 2975
rect 40092 2944 40417 2972
rect 40092 2932 40098 2944
rect 40405 2941 40417 2944
rect 40451 2941 40463 2975
rect 40405 2935 40463 2941
rect 40586 2932 40592 2984
rect 40644 2972 40650 2984
rect 40957 2975 41015 2981
rect 40957 2972 40969 2975
rect 40644 2944 40969 2972
rect 40644 2932 40650 2944
rect 40957 2941 40969 2944
rect 41003 2941 41015 2975
rect 40957 2935 41015 2941
rect 41138 2932 41144 2984
rect 41196 2972 41202 2984
rect 41509 2975 41567 2981
rect 41509 2972 41521 2975
rect 41196 2944 41521 2972
rect 41196 2932 41202 2944
rect 41509 2941 41521 2944
rect 41555 2941 41567 2975
rect 41509 2935 41567 2941
rect 41690 2932 41696 2984
rect 41748 2972 41754 2984
rect 42061 2975 42119 2981
rect 42061 2972 42073 2975
rect 41748 2944 42073 2972
rect 41748 2932 41754 2944
rect 42061 2941 42073 2944
rect 42107 2941 42119 2975
rect 42061 2935 42119 2941
rect 42242 2932 42248 2984
rect 42300 2972 42306 2984
rect 42613 2975 42671 2981
rect 42613 2972 42625 2975
rect 42300 2944 42625 2972
rect 42300 2932 42306 2944
rect 42613 2941 42625 2944
rect 42659 2941 42671 2975
rect 42613 2935 42671 2941
rect 42794 2932 42800 2984
rect 42852 2972 42858 2984
rect 43441 2975 43499 2981
rect 43441 2972 43453 2975
rect 42852 2944 43453 2972
rect 42852 2932 42858 2944
rect 43441 2941 43453 2944
rect 43487 2941 43499 2975
rect 43441 2935 43499 2941
rect 43622 2932 43628 2984
rect 43680 2972 43686 2984
rect 44269 2975 44327 2981
rect 44269 2972 44281 2975
rect 43680 2944 44281 2972
rect 43680 2932 43686 2944
rect 44269 2941 44281 2944
rect 44315 2941 44327 2975
rect 44269 2935 44327 2941
rect 44450 2932 44456 2984
rect 44508 2972 44514 2984
rect 45097 2975 45155 2981
rect 45097 2972 45109 2975
rect 44508 2944 45109 2972
rect 44508 2932 44514 2944
rect 45097 2941 45109 2944
rect 45143 2941 45155 2975
rect 45097 2935 45155 2941
rect 45278 2932 45284 2984
rect 45336 2972 45342 2984
rect 45925 2975 45983 2981
rect 45925 2972 45937 2975
rect 45336 2944 45937 2972
rect 45336 2932 45342 2944
rect 45925 2941 45937 2944
rect 45971 2941 45983 2975
rect 45925 2935 45983 2941
rect 46106 2932 46112 2984
rect 46164 2972 46170 2984
rect 46753 2975 46811 2981
rect 46753 2972 46765 2975
rect 46164 2944 46765 2972
rect 46164 2932 46170 2944
rect 46753 2941 46765 2944
rect 46799 2941 46811 2975
rect 46753 2935 46811 2941
rect 46934 2932 46940 2984
rect 46992 2972 46998 2984
rect 47581 2975 47639 2981
rect 47581 2972 47593 2975
rect 46992 2944 47593 2972
rect 46992 2932 46998 2944
rect 47581 2941 47593 2944
rect 47627 2941 47639 2975
rect 47581 2935 47639 2941
rect 47762 2932 47768 2984
rect 47820 2972 47826 2984
rect 47820 2944 48176 2972
rect 47820 2932 47826 2944
rect 25777 2907 25835 2913
rect 25777 2904 25789 2907
rect 24504 2876 25789 2904
rect 24397 2867 24455 2873
rect 25777 2873 25789 2876
rect 25823 2873 25835 2907
rect 27706 2904 27712 2916
rect 27667 2876 27712 2904
rect 25777 2867 25835 2873
rect 27706 2864 27712 2876
rect 27764 2864 27770 2916
rect 27798 2864 27804 2916
rect 27856 2904 27862 2916
rect 27856 2876 29454 2904
rect 27856 2864 27862 2876
rect 17644 2808 18184 2836
rect 17644 2796 17650 2808
rect 18230 2796 18236 2848
rect 18288 2836 18294 2848
rect 19705 2839 19763 2845
rect 19705 2836 19717 2839
rect 18288 2808 19717 2836
rect 18288 2796 18294 2808
rect 19705 2805 19717 2808
rect 19751 2805 19763 2839
rect 19705 2799 19763 2805
rect 19794 2796 19800 2848
rect 19852 2836 19858 2848
rect 21085 2839 21143 2845
rect 21085 2836 21097 2839
rect 19852 2808 21097 2836
rect 19852 2796 19858 2808
rect 21085 2805 21097 2808
rect 21131 2805 21143 2839
rect 21085 2799 21143 2805
rect 21913 2839 21971 2845
rect 21913 2805 21925 2839
rect 21959 2836 21971 2839
rect 23017 2839 23075 2845
rect 23017 2836 23029 2839
rect 21959 2808 23029 2836
rect 21959 2805 21971 2808
rect 21913 2799 21971 2805
rect 23017 2805 23029 2808
rect 23063 2805 23075 2839
rect 23017 2799 23075 2805
rect 23198 2796 23204 2848
rect 23256 2836 23262 2848
rect 24949 2839 25007 2845
rect 24949 2836 24961 2839
rect 23256 2808 24961 2836
rect 23256 2796 23262 2808
rect 24949 2805 24961 2808
rect 24995 2805 25007 2839
rect 24949 2799 25007 2805
rect 25682 2796 25688 2848
rect 25740 2836 25746 2848
rect 27614 2836 27620 2848
rect 25740 2808 27620 2836
rect 25740 2796 25746 2808
rect 27614 2796 27620 2808
rect 27672 2796 27678 2848
rect 28534 2836 28540 2848
rect 28495 2808 28540 2836
rect 28534 2796 28540 2808
rect 28592 2796 28598 2848
rect 29426 2836 29454 2876
rect 29546 2864 29552 2916
rect 29604 2904 29610 2916
rect 31573 2907 31631 2913
rect 31573 2904 31585 2907
rect 29604 2876 31585 2904
rect 29604 2864 29610 2876
rect 31573 2873 31585 2876
rect 31619 2873 31631 2907
rect 31573 2867 31631 2873
rect 36722 2864 36728 2916
rect 36780 2904 36786 2916
rect 36817 2907 36875 2913
rect 36817 2904 36829 2907
rect 36780 2876 36829 2904
rect 36780 2864 36786 2876
rect 36817 2873 36829 2876
rect 36863 2873 36875 2907
rect 36817 2867 36875 2873
rect 43070 2864 43076 2916
rect 43128 2904 43134 2916
rect 43717 2907 43775 2913
rect 43717 2904 43729 2907
rect 43128 2876 43729 2904
rect 43128 2864 43134 2876
rect 43717 2873 43729 2876
rect 43763 2873 43775 2907
rect 43717 2867 43775 2873
rect 43898 2864 43904 2916
rect 43956 2904 43962 2916
rect 44545 2907 44603 2913
rect 44545 2904 44557 2907
rect 43956 2876 44557 2904
rect 43956 2864 43962 2876
rect 44545 2873 44557 2876
rect 44591 2873 44603 2907
rect 44545 2867 44603 2873
rect 44726 2864 44732 2916
rect 44784 2904 44790 2916
rect 45373 2907 45431 2913
rect 45373 2904 45385 2907
rect 44784 2876 45385 2904
rect 44784 2864 44790 2876
rect 45373 2873 45385 2876
rect 45419 2873 45431 2907
rect 45373 2867 45431 2873
rect 45554 2864 45560 2916
rect 45612 2904 45618 2916
rect 46201 2907 46259 2913
rect 46201 2904 46213 2907
rect 45612 2876 46213 2904
rect 45612 2864 45618 2876
rect 46201 2873 46213 2876
rect 46247 2873 46259 2907
rect 46201 2867 46259 2873
rect 46382 2864 46388 2916
rect 46440 2904 46446 2916
rect 47029 2907 47087 2913
rect 47029 2904 47041 2907
rect 46440 2876 47041 2904
rect 46440 2864 46446 2876
rect 47029 2873 47041 2876
rect 47075 2873 47087 2907
rect 47029 2867 47087 2873
rect 47210 2864 47216 2916
rect 47268 2904 47274 2916
rect 47857 2907 47915 2913
rect 47857 2904 47869 2907
rect 47268 2876 47869 2904
rect 47268 2864 47274 2876
rect 47857 2873 47869 2876
rect 47903 2873 47915 2907
rect 48148 2904 48176 2944
rect 48590 2932 48596 2984
rect 48648 2972 48654 2984
rect 49513 2975 49571 2981
rect 49513 2972 49525 2975
rect 48648 2944 49525 2972
rect 48648 2932 48654 2944
rect 49513 2941 49525 2944
rect 49559 2941 49571 2975
rect 49513 2935 49571 2941
rect 49694 2932 49700 2984
rect 49752 2972 49758 2984
rect 50617 2975 50675 2981
rect 50617 2972 50629 2975
rect 49752 2944 50629 2972
rect 49752 2932 49758 2944
rect 50617 2941 50629 2944
rect 50663 2941 50675 2975
rect 50617 2935 50675 2941
rect 50798 2932 50804 2984
rect 50856 2972 50862 2984
rect 51721 2975 51779 2981
rect 51721 2972 51733 2975
rect 50856 2944 51733 2972
rect 50856 2932 50862 2944
rect 51721 2941 51733 2944
rect 51767 2941 51779 2975
rect 51721 2935 51779 2941
rect 51902 2932 51908 2984
rect 51960 2972 51966 2984
rect 52825 2975 52883 2981
rect 52825 2972 52837 2975
rect 51960 2944 52837 2972
rect 51960 2932 51966 2944
rect 52825 2941 52837 2944
rect 52871 2941 52883 2975
rect 52825 2935 52883 2941
rect 53006 2932 53012 2984
rect 53064 2972 53070 2984
rect 54205 2975 54263 2981
rect 54205 2972 54217 2975
rect 53064 2944 54217 2972
rect 53064 2932 53070 2944
rect 54205 2941 54217 2944
rect 54251 2941 54263 2975
rect 54404 2972 54432 3012
rect 54481 3009 54493 3043
rect 54527 3009 54539 3043
rect 54481 3003 54539 3009
rect 54662 3000 54668 3052
rect 54720 3040 54726 3052
rect 55600 3049 55628 3148
rect 56870 3136 56876 3188
rect 56928 3176 56934 3188
rect 56928 3148 58112 3176
rect 56928 3136 56934 3148
rect 55766 3068 55772 3120
rect 55824 3108 55830 3120
rect 55824 3080 57008 3108
rect 55824 3068 55830 3080
rect 55585 3043 55643 3049
rect 54720 3012 55444 3040
rect 54720 3000 54726 3012
rect 55309 2975 55367 2981
rect 55309 2972 55321 2975
rect 54404 2944 55321 2972
rect 54205 2935 54263 2941
rect 55309 2941 55321 2944
rect 55355 2941 55367 2975
rect 55416 2972 55444 3012
rect 55585 3009 55597 3043
rect 55631 3009 55643 3043
rect 55585 3003 55643 3009
rect 55674 3000 55680 3052
rect 55732 3040 55738 3052
rect 56980 3049 57008 3080
rect 58084 3049 58112 3148
rect 58802 3136 58808 3188
rect 58860 3176 58866 3188
rect 58860 3148 60320 3176
rect 58860 3136 58866 3148
rect 58250 3068 58256 3120
rect 58308 3108 58314 3120
rect 58308 3080 59768 3108
rect 58308 3068 58314 3080
rect 56689 3043 56747 3049
rect 56689 3040 56701 3043
rect 55732 3012 56701 3040
rect 55732 3000 55738 3012
rect 56689 3009 56701 3012
rect 56735 3009 56747 3043
rect 56689 3003 56747 3009
rect 56965 3043 57023 3049
rect 56965 3009 56977 3043
rect 57011 3009 57023 3043
rect 56965 3003 57023 3009
rect 58069 3043 58127 3049
rect 58069 3009 58081 3043
rect 58115 3009 58127 3043
rect 58069 3003 58127 3009
rect 58158 3000 58164 3052
rect 58216 3040 58222 3052
rect 59740 3049 59768 3080
rect 59449 3043 59507 3049
rect 59449 3040 59461 3043
rect 58216 3012 59461 3040
rect 58216 3000 58222 3012
rect 59449 3009 59461 3012
rect 59495 3009 59507 3043
rect 59449 3003 59507 3009
rect 59725 3043 59783 3049
rect 59725 3009 59737 3043
rect 59771 3009 59783 3043
rect 59725 3003 59783 3009
rect 59814 3000 59820 3052
rect 59872 3040 59878 3052
rect 60292 3049 60320 3148
rect 61010 3136 61016 3188
rect 61068 3176 61074 3188
rect 61068 3148 62528 3176
rect 61068 3136 61074 3148
rect 60366 3068 60372 3120
rect 60424 3108 60430 3120
rect 60424 3080 61700 3108
rect 60424 3068 60430 3080
rect 60277 3043 60335 3049
rect 59872 3012 60228 3040
rect 59872 3000 59878 3012
rect 55861 2975 55919 2981
rect 55861 2972 55873 2975
rect 55416 2944 55873 2972
rect 55309 2935 55367 2941
rect 55861 2941 55873 2944
rect 55907 2941 55919 2975
rect 55861 2935 55919 2941
rect 56042 2932 56048 2984
rect 56100 2972 56106 2984
rect 56100 2944 56548 2972
rect 56100 2932 56106 2944
rect 48685 2907 48743 2913
rect 48685 2904 48697 2907
rect 48148 2876 48697 2904
rect 47857 2867 47915 2873
rect 48685 2873 48697 2876
rect 48731 2873 48743 2907
rect 48685 2867 48743 2873
rect 48866 2864 48872 2916
rect 48924 2904 48930 2916
rect 49789 2907 49847 2913
rect 49789 2904 49801 2907
rect 48924 2876 49801 2904
rect 48924 2864 48930 2876
rect 49789 2873 49801 2876
rect 49835 2873 49847 2907
rect 49789 2867 49847 2873
rect 49970 2864 49976 2916
rect 50028 2904 50034 2916
rect 50893 2907 50951 2913
rect 50893 2904 50905 2907
rect 50028 2876 50905 2904
rect 50028 2864 50034 2876
rect 50893 2873 50905 2876
rect 50939 2873 50951 2907
rect 50893 2867 50951 2873
rect 51350 2864 51356 2916
rect 51408 2904 51414 2916
rect 52273 2907 52331 2913
rect 52273 2904 52285 2907
rect 51408 2876 52285 2904
rect 51408 2864 51414 2876
rect 52273 2873 52285 2876
rect 52319 2873 52331 2907
rect 52273 2867 52331 2873
rect 52454 2864 52460 2916
rect 52512 2904 52518 2916
rect 53653 2907 53711 2913
rect 53653 2904 53665 2907
rect 52512 2876 53665 2904
rect 52512 2864 52518 2876
rect 53653 2873 53665 2876
rect 53699 2873 53711 2907
rect 53653 2867 53711 2873
rect 53834 2864 53840 2916
rect 53892 2904 53898 2916
rect 55033 2907 55091 2913
rect 55033 2904 55045 2907
rect 53892 2876 55045 2904
rect 53892 2864 53898 2876
rect 55033 2873 55045 2876
rect 55079 2873 55091 2907
rect 55033 2867 55091 2873
rect 55214 2864 55220 2916
rect 55272 2904 55278 2916
rect 56413 2907 56471 2913
rect 56413 2904 56425 2907
rect 55272 2876 56425 2904
rect 55272 2864 55278 2876
rect 56413 2873 56425 2876
rect 56459 2873 56471 2907
rect 56413 2867 56471 2873
rect 29641 2839 29699 2845
rect 29641 2836 29653 2839
rect 29426 2808 29653 2836
rect 29641 2805 29653 2808
rect 29687 2805 29699 2839
rect 30466 2836 30472 2848
rect 30427 2808 30472 2836
rect 29641 2799 29699 2805
rect 30466 2796 30472 2808
rect 30524 2796 30530 2848
rect 30742 2836 30748 2848
rect 30703 2808 30748 2836
rect 30742 2796 30748 2808
rect 30800 2796 30806 2848
rect 31018 2836 31024 2848
rect 30979 2808 31024 2836
rect 31018 2796 31024 2808
rect 31076 2796 31082 2848
rect 31294 2836 31300 2848
rect 31255 2808 31300 2836
rect 31294 2796 31300 2808
rect 31352 2796 31358 2848
rect 47486 2796 47492 2848
rect 47544 2836 47550 2848
rect 48409 2839 48467 2845
rect 48409 2836 48421 2839
rect 47544 2808 48421 2836
rect 47544 2796 47550 2808
rect 48409 2805 48421 2808
rect 48455 2805 48467 2839
rect 48409 2799 48467 2805
rect 49142 2796 49148 2848
rect 49200 2836 49206 2848
rect 50065 2839 50123 2845
rect 50065 2836 50077 2839
rect 49200 2808 50077 2836
rect 49200 2796 49206 2808
rect 50065 2805 50077 2808
rect 50111 2805 50123 2839
rect 50065 2799 50123 2805
rect 50522 2796 50528 2848
rect 50580 2836 50586 2848
rect 51445 2839 51503 2845
rect 51445 2836 51457 2839
rect 50580 2808 51457 2836
rect 50580 2796 50586 2808
rect 51445 2805 51457 2808
rect 51491 2805 51503 2839
rect 51445 2799 51503 2805
rect 52178 2796 52184 2848
rect 52236 2836 52242 2848
rect 53101 2839 53159 2845
rect 53101 2836 53113 2839
rect 52236 2808 53113 2836
rect 52236 2796 52242 2808
rect 53101 2805 53113 2808
rect 53147 2805 53159 2839
rect 53101 2799 53159 2805
rect 53558 2796 53564 2848
rect 53616 2836 53622 2848
rect 54757 2839 54815 2845
rect 54757 2836 54769 2839
rect 53616 2808 54769 2836
rect 53616 2796 53622 2808
rect 54757 2805 54769 2808
rect 54803 2805 54815 2839
rect 54757 2799 54815 2805
rect 54938 2796 54944 2848
rect 54996 2836 55002 2848
rect 56137 2839 56195 2845
rect 56137 2836 56149 2839
rect 54996 2808 56149 2836
rect 54996 2796 55002 2808
rect 56137 2805 56149 2808
rect 56183 2805 56195 2839
rect 56520 2836 56548 2944
rect 57238 2932 57244 2984
rect 57296 2972 57302 2984
rect 58345 2975 58403 2981
rect 58345 2972 58357 2975
rect 57296 2944 58357 2972
rect 57296 2932 57302 2944
rect 58345 2941 58357 2944
rect 58391 2941 58403 2975
rect 58345 2935 58403 2941
rect 58526 2932 58532 2984
rect 58584 2972 58590 2984
rect 60001 2975 60059 2981
rect 60001 2972 60013 2975
rect 58584 2944 60013 2972
rect 58584 2932 58590 2944
rect 60001 2941 60013 2944
rect 60047 2941 60059 2975
rect 60200 2972 60228 3012
rect 60277 3009 60289 3043
rect 60323 3009 60335 3043
rect 60277 3003 60335 3009
rect 60458 3000 60464 3052
rect 60516 3040 60522 3052
rect 61378 3040 61384 3052
rect 60516 3012 61240 3040
rect 61339 3012 61384 3040
rect 60516 3000 60522 3012
rect 61105 2975 61163 2981
rect 61105 2972 61117 2975
rect 60200 2944 61117 2972
rect 60001 2935 60059 2941
rect 61105 2941 61117 2944
rect 61151 2941 61163 2975
rect 61212 2972 61240 3012
rect 61378 3000 61384 3012
rect 61436 3000 61442 3052
rect 61672 3049 61700 3080
rect 62500 3049 62528 3148
rect 64046 3136 64052 3188
rect 64104 3176 64110 3188
rect 64104 3148 65840 3176
rect 64104 3136 64110 3148
rect 63310 3068 63316 3120
rect 63368 3108 63374 3120
rect 63368 3080 65012 3108
rect 63368 3068 63374 3080
rect 61657 3043 61715 3049
rect 61657 3009 61669 3043
rect 61703 3009 61715 3043
rect 61657 3003 61715 3009
rect 62485 3043 62543 3049
rect 62485 3009 62497 3043
rect 62531 3009 62543 3043
rect 62758 3040 62764 3052
rect 62719 3012 62764 3040
rect 62485 3003 62543 3009
rect 62758 3000 62764 3012
rect 62816 3000 62822 3052
rect 62942 3000 62948 3052
rect 63000 3040 63006 3052
rect 63037 3043 63095 3049
rect 63037 3040 63049 3043
rect 63000 3012 63049 3040
rect 63000 3000 63006 3012
rect 63037 3009 63049 3012
rect 63083 3009 63095 3043
rect 63037 3003 63095 3009
rect 63770 3000 63776 3052
rect 63828 3040 63834 3052
rect 64690 3040 64696 3052
rect 63828 3012 64552 3040
rect 64651 3012 64696 3040
rect 63828 3000 63834 3012
rect 61933 2975 61991 2981
rect 61933 2972 61945 2975
rect 61212 2944 61945 2972
rect 61105 2935 61163 2941
rect 61933 2941 61945 2944
rect 61979 2941 61991 2975
rect 61933 2935 61991 2941
rect 62390 2932 62396 2984
rect 62448 2972 62454 2984
rect 64141 2975 64199 2981
rect 64141 2972 64153 2975
rect 62448 2944 64153 2972
rect 62448 2932 62454 2944
rect 64141 2941 64153 2944
rect 64187 2941 64199 2975
rect 64524 2972 64552 3012
rect 64690 3000 64696 3012
rect 64748 3000 64754 3052
rect 64984 3049 65012 3080
rect 64969 3043 65027 3049
rect 64969 3009 64981 3043
rect 65015 3009 65027 3043
rect 64969 3003 65027 3009
rect 65058 3000 65064 3052
rect 65116 3040 65122 3052
rect 65812 3049 65840 3148
rect 66254 3136 66260 3188
rect 66312 3176 66318 3188
rect 68002 3176 68008 3188
rect 66312 3148 68008 3176
rect 66312 3136 66318 3148
rect 68002 3136 68008 3148
rect 68060 3136 68066 3188
rect 66806 3068 66812 3120
rect 66864 3108 66870 3120
rect 66864 3080 69060 3108
rect 66864 3068 66870 3080
rect 65797 3043 65855 3049
rect 65116 3012 65748 3040
rect 65116 3000 65122 3012
rect 65521 2975 65579 2981
rect 65521 2972 65533 2975
rect 64524 2944 65533 2972
rect 64141 2935 64199 2941
rect 65521 2941 65533 2944
rect 65567 2941 65579 2975
rect 65720 2972 65748 3012
rect 65797 3009 65809 3043
rect 65843 3009 65855 3043
rect 66346 3040 66352 3052
rect 66307 3012 66352 3040
rect 65797 3003 65855 3009
rect 66346 3000 66352 3012
rect 66404 3000 66410 3052
rect 67174 3040 67180 3052
rect 67135 3012 67180 3040
rect 67174 3000 67180 3012
rect 67232 3000 67238 3052
rect 67358 3000 67364 3052
rect 67416 3040 67422 3052
rect 69032 3049 69060 3080
rect 68741 3043 68799 3049
rect 68741 3040 68753 3043
rect 67416 3012 68753 3040
rect 67416 3000 67422 3012
rect 68741 3009 68753 3012
rect 68787 3009 68799 3043
rect 68741 3003 68799 3009
rect 69017 3043 69075 3049
rect 69017 3009 69029 3043
rect 69063 3009 69075 3043
rect 69017 3003 69075 3009
rect 66625 2975 66683 2981
rect 66625 2972 66637 2975
rect 65720 2944 66637 2972
rect 65521 2935 65579 2941
rect 66625 2941 66637 2944
rect 66671 2941 66683 2975
rect 66625 2935 66683 2941
rect 67082 2932 67088 2984
rect 67140 2972 67146 2984
rect 69385 2975 69443 2981
rect 69385 2972 69397 2975
rect 67140 2944 69397 2972
rect 67140 2932 67146 2944
rect 69385 2941 69397 2944
rect 69431 2941 69443 2975
rect 69385 2935 69443 2941
rect 56594 2864 56600 2916
rect 56652 2904 56658 2916
rect 57793 2907 57851 2913
rect 57793 2904 57805 2907
rect 56652 2876 57805 2904
rect 56652 2864 56658 2876
rect 57793 2873 57805 2876
rect 57839 2873 57851 2907
rect 57793 2867 57851 2873
rect 58066 2864 58072 2916
rect 58124 2904 58130 2916
rect 58124 2876 59032 2904
rect 58124 2864 58130 2876
rect 57241 2839 57299 2845
rect 57241 2836 57253 2839
rect 56520 2808 57253 2836
rect 56137 2799 56195 2805
rect 57241 2805 57253 2808
rect 57287 2805 57299 2839
rect 57241 2799 57299 2805
rect 57330 2796 57336 2848
rect 57388 2836 57394 2848
rect 57517 2839 57575 2845
rect 57517 2836 57529 2839
rect 57388 2808 57529 2836
rect 57388 2796 57394 2808
rect 57517 2805 57529 2808
rect 57563 2805 57575 2839
rect 57517 2799 57575 2805
rect 57606 2796 57612 2848
rect 57664 2836 57670 2848
rect 58897 2839 58955 2845
rect 58897 2836 58909 2839
rect 57664 2808 58909 2836
rect 57664 2796 57670 2808
rect 58897 2805 58909 2808
rect 58943 2805 58955 2839
rect 59004 2836 59032 2876
rect 59078 2864 59084 2916
rect 59136 2904 59142 2916
rect 59136 2876 59308 2904
rect 59136 2864 59142 2876
rect 59173 2839 59231 2845
rect 59173 2836 59185 2839
rect 59004 2808 59185 2836
rect 58897 2799 58955 2805
rect 59173 2805 59185 2808
rect 59219 2805 59231 2839
rect 59280 2836 59308 2876
rect 59354 2864 59360 2916
rect 59412 2904 59418 2916
rect 60829 2907 60887 2913
rect 60829 2904 60841 2907
rect 59412 2876 60841 2904
rect 59412 2864 59418 2876
rect 60829 2873 60841 2876
rect 60875 2873 60887 2907
rect 60829 2867 60887 2873
rect 61838 2864 61844 2916
rect 61896 2904 61902 2916
rect 63313 2907 63371 2913
rect 63313 2904 63325 2907
rect 61896 2876 63325 2904
rect 61896 2864 61902 2876
rect 63313 2873 63325 2876
rect 63359 2873 63371 2907
rect 63313 2867 63371 2873
rect 63494 2864 63500 2916
rect 63552 2904 63558 2916
rect 65058 2904 65064 2916
rect 63552 2876 65064 2904
rect 63552 2864 63558 2876
rect 65058 2864 65064 2876
rect 65116 2864 65122 2916
rect 66073 2907 66131 2913
rect 66073 2904 66085 2907
rect 65168 2876 66085 2904
rect 60553 2839 60611 2845
rect 60553 2836 60565 2839
rect 59280 2808 60565 2836
rect 59173 2799 59231 2805
rect 60553 2805 60565 2808
rect 60599 2805 60611 2839
rect 60553 2799 60611 2805
rect 60734 2796 60740 2848
rect 60792 2836 60798 2848
rect 62209 2839 62267 2845
rect 62209 2836 62221 2839
rect 60792 2808 62221 2836
rect 60792 2796 60798 2808
rect 62209 2805 62221 2808
rect 62255 2805 62267 2839
rect 62209 2799 62267 2805
rect 62298 2796 62304 2848
rect 62356 2836 62362 2848
rect 63589 2839 63647 2845
rect 63589 2836 63601 2839
rect 62356 2808 63601 2836
rect 62356 2796 62362 2808
rect 63589 2805 63601 2808
rect 63635 2805 63647 2839
rect 64414 2836 64420 2848
rect 64375 2808 64420 2836
rect 63589 2799 63647 2805
rect 64414 2796 64420 2808
rect 64472 2796 64478 2848
rect 64506 2796 64512 2848
rect 64564 2836 64570 2848
rect 65168 2836 65196 2876
rect 66073 2873 66085 2876
rect 66119 2873 66131 2907
rect 66073 2867 66131 2873
rect 66530 2864 66536 2916
rect 66588 2904 66594 2916
rect 67450 2904 67456 2916
rect 66588 2876 67312 2904
rect 67411 2876 67456 2904
rect 66588 2864 66594 2876
rect 64564 2808 65196 2836
rect 64564 2796 64570 2808
rect 65242 2796 65248 2848
rect 65300 2836 65306 2848
rect 65300 2808 65345 2836
rect 65300 2796 65306 2808
rect 65426 2796 65432 2848
rect 65484 2836 65490 2848
rect 66901 2839 66959 2845
rect 66901 2836 66913 2839
rect 65484 2808 66913 2836
rect 65484 2796 65490 2808
rect 66901 2805 66913 2808
rect 66947 2805 66959 2839
rect 67284 2836 67312 2876
rect 67450 2864 67456 2876
rect 67508 2864 67514 2916
rect 67726 2904 67732 2916
rect 67687 2876 67732 2904
rect 67726 2864 67732 2876
rect 67784 2864 67790 2916
rect 68002 2904 68008 2916
rect 67963 2876 68008 2904
rect 68002 2864 68008 2876
rect 68060 2864 68066 2916
rect 68281 2839 68339 2845
rect 68281 2836 68293 2839
rect 67284 2808 68293 2836
rect 66901 2799 66959 2805
rect 68281 2805 68293 2808
rect 68327 2805 68339 2839
rect 68281 2799 68339 2805
rect 1104 2746 72864 2768
rect 1104 2694 9078 2746
rect 9130 2694 21078 2746
rect 21130 2694 33078 2746
rect 33130 2694 45078 2746
rect 45130 2694 57078 2746
rect 57130 2694 69078 2746
rect 69130 2694 72864 2746
rect 1104 2672 72864 2694
rect 2958 2592 2964 2644
rect 3016 2632 3022 2644
rect 3053 2635 3111 2641
rect 3053 2632 3065 2635
rect 3016 2604 3065 2632
rect 3016 2592 3022 2604
rect 3053 2601 3065 2604
rect 3099 2601 3111 2635
rect 3053 2595 3111 2601
rect 16022 2524 16028 2576
rect 16080 2564 16086 2576
rect 17494 2564 17500 2576
rect 16080 2536 17500 2564
rect 16080 2524 16086 2536
rect 17494 2524 17500 2536
rect 17552 2524 17558 2576
rect 62666 2524 62672 2576
rect 62724 2564 62730 2576
rect 64414 2564 64420 2576
rect 62724 2536 64420 2564
rect 62724 2524 62730 2536
rect 64414 2524 64420 2536
rect 64472 2524 64478 2576
rect 2774 2496 2780 2508
rect 2735 2468 2780 2496
rect 2774 2456 2780 2468
rect 2832 2456 2838 2508
rect 2498 2428 2504 2440
rect 2459 2400 2504 2428
rect 2498 2388 2504 2400
rect 2556 2388 2562 2440
rect 1104 2202 72864 2224
rect 1104 2150 3078 2202
rect 3130 2150 15078 2202
rect 15130 2150 27078 2202
rect 27130 2150 39078 2202
rect 39130 2150 51078 2202
rect 51130 2150 63078 2202
rect 63130 2150 72864 2202
rect 1104 2128 72864 2150
rect 1394 1844 1400 1896
rect 1452 1884 1458 1896
rect 3145 1887 3203 1893
rect 3145 1884 3157 1887
rect 1452 1856 3157 1884
rect 1452 1844 1458 1856
rect 3145 1853 3157 1856
rect 3191 1853 3203 1887
rect 3145 1847 3203 1853
rect 30098 1776 30104 1828
rect 30156 1816 30162 1828
rect 31021 1819 31079 1825
rect 31021 1816 31033 1819
rect 30156 1788 31033 1816
rect 30156 1776 30162 1788
rect 31021 1785 31033 1788
rect 31067 1785 31079 1819
rect 31021 1779 31079 1785
rect 2222 1748 2228 1760
rect 2183 1720 2228 1748
rect 2222 1708 2228 1720
rect 2280 1708 2286 1760
rect 2314 1708 2320 1760
rect 2372 1748 2378 1760
rect 2501 1751 2559 1757
rect 2501 1748 2513 1751
rect 2372 1720 2513 1748
rect 2372 1708 2378 1720
rect 2501 1717 2513 1720
rect 2547 1717 2559 1751
rect 2501 1711 2559 1717
rect 2774 1708 2780 1760
rect 2832 1748 2838 1760
rect 2869 1751 2927 1757
rect 2869 1748 2881 1751
rect 2832 1720 2881 1748
rect 2832 1708 2838 1720
rect 2869 1717 2881 1720
rect 2915 1717 2927 1751
rect 2869 1711 2927 1717
rect 2958 1708 2964 1760
rect 3016 1748 3022 1760
rect 3421 1751 3479 1757
rect 3421 1748 3433 1751
rect 3016 1720 3433 1748
rect 3016 1708 3022 1720
rect 3421 1717 3433 1720
rect 3467 1717 3479 1751
rect 3421 1711 3479 1717
rect 3878 1708 3884 1760
rect 3936 1748 3942 1760
rect 4065 1751 4123 1757
rect 4065 1748 4077 1751
rect 3936 1720 4077 1748
rect 3936 1708 3942 1720
rect 4065 1717 4077 1720
rect 4111 1717 4123 1751
rect 4065 1711 4123 1717
rect 6638 1708 6644 1760
rect 6696 1748 6702 1760
rect 7009 1751 7067 1757
rect 7009 1748 7021 1751
rect 6696 1720 7021 1748
rect 6696 1708 6702 1720
rect 7009 1717 7021 1720
rect 7055 1717 7067 1751
rect 7009 1711 7067 1717
rect 8570 1708 8576 1760
rect 8628 1748 8634 1760
rect 8941 1751 8999 1757
rect 8941 1748 8953 1751
rect 8628 1720 8953 1748
rect 8628 1708 8634 1720
rect 8941 1717 8953 1720
rect 8987 1717 8999 1751
rect 8941 1711 8999 1717
rect 9398 1708 9404 1760
rect 9456 1748 9462 1760
rect 9861 1751 9919 1757
rect 9861 1748 9873 1751
rect 9456 1720 9873 1748
rect 9456 1708 9462 1720
rect 9861 1717 9873 1720
rect 9907 1717 9919 1751
rect 9861 1711 9919 1717
rect 11606 1708 11612 1760
rect 11664 1748 11670 1760
rect 11885 1751 11943 1757
rect 11885 1748 11897 1751
rect 11664 1720 11897 1748
rect 11664 1708 11670 1720
rect 11885 1717 11897 1720
rect 11931 1717 11943 1751
rect 11885 1711 11943 1717
rect 12986 1708 12992 1760
rect 13044 1748 13050 1760
rect 13265 1751 13323 1757
rect 13265 1748 13277 1751
rect 13044 1720 13277 1748
rect 13044 1708 13050 1720
rect 13265 1717 13277 1720
rect 13311 1717 13323 1751
rect 13265 1711 13323 1717
rect 14918 1708 14924 1760
rect 14976 1748 14982 1760
rect 15197 1751 15255 1757
rect 15197 1748 15209 1751
rect 14976 1720 15209 1748
rect 14976 1708 14982 1720
rect 15197 1717 15209 1720
rect 15243 1717 15255 1751
rect 15197 1711 15255 1717
rect 15746 1708 15752 1760
rect 15804 1748 15810 1760
rect 16117 1751 16175 1757
rect 16117 1748 16129 1751
rect 15804 1720 16129 1748
rect 15804 1708 15810 1720
rect 16117 1717 16129 1720
rect 16163 1717 16175 1751
rect 16117 1711 16175 1717
rect 19886 1708 19892 1760
rect 19944 1748 19950 1760
rect 20349 1751 20407 1757
rect 20349 1748 20361 1751
rect 19944 1720 20361 1748
rect 19944 1708 19950 1720
rect 20349 1717 20361 1720
rect 20395 1717 20407 1751
rect 20349 1711 20407 1717
rect 25958 1708 25964 1760
rect 26016 1748 26022 1760
rect 26697 1751 26755 1757
rect 26697 1748 26709 1751
rect 26016 1720 26709 1748
rect 26016 1708 26022 1720
rect 26697 1717 26709 1720
rect 26743 1717 26755 1751
rect 26697 1711 26755 1717
rect 29822 1708 29828 1760
rect 29880 1748 29886 1760
rect 30745 1751 30803 1757
rect 30745 1748 30757 1751
rect 29880 1720 30757 1748
rect 29880 1708 29886 1720
rect 30745 1717 30757 1720
rect 30791 1717 30803 1751
rect 30745 1711 30803 1717
rect 31478 1708 31484 1760
rect 31536 1748 31542 1760
rect 32677 1751 32735 1757
rect 32677 1748 32689 1751
rect 31536 1720 32689 1748
rect 31536 1708 31542 1720
rect 32677 1717 32689 1720
rect 32723 1717 32735 1751
rect 32677 1711 32735 1717
rect 38565 1751 38623 1757
rect 38565 1717 38577 1751
rect 38611 1748 38623 1751
rect 38930 1748 38936 1760
rect 38611 1720 38936 1748
rect 38611 1717 38623 1720
rect 38565 1711 38623 1717
rect 38930 1708 38936 1720
rect 38988 1708 38994 1760
rect 43993 1751 44051 1757
rect 43993 1717 44005 1751
rect 44039 1748 44051 1751
rect 44174 1748 44180 1760
rect 44039 1720 44180 1748
rect 44039 1717 44051 1720
rect 43993 1711 44051 1717
rect 44174 1708 44180 1720
rect 44232 1708 44238 1760
rect 46845 1751 46903 1757
rect 46845 1717 46857 1751
rect 46891 1748 46903 1751
rect 46934 1748 46940 1760
rect 46891 1720 46940 1748
rect 46891 1717 46903 1720
rect 46845 1711 46903 1717
rect 46934 1708 46940 1720
rect 46992 1708 46998 1760
rect 50522 1748 50528 1760
rect 50483 1720 50528 1748
rect 50522 1708 50528 1720
rect 50580 1708 50586 1760
rect 52454 1708 52460 1760
rect 52512 1748 52518 1760
rect 52549 1751 52607 1757
rect 52549 1748 52561 1751
rect 52512 1720 52561 1748
rect 52512 1708 52518 1720
rect 52549 1717 52561 1720
rect 52595 1717 52607 1751
rect 54386 1748 54392 1760
rect 54347 1720 54392 1748
rect 52549 1711 52607 1717
rect 54386 1708 54392 1720
rect 54444 1708 54450 1760
rect 57422 1708 57428 1760
rect 57480 1748 57486 1760
rect 57517 1751 57575 1757
rect 57517 1748 57529 1751
rect 57480 1720 57529 1748
rect 57480 1708 57486 1720
rect 57517 1717 57529 1720
rect 57563 1717 57575 1751
rect 57517 1711 57575 1717
rect 63494 1708 63500 1760
rect 63552 1748 63558 1760
rect 64141 1751 64199 1757
rect 64141 1748 64153 1751
rect 63552 1720 64153 1748
rect 63552 1708 63558 1720
rect 64141 1717 64153 1720
rect 64187 1717 64199 1751
rect 64141 1711 64199 1717
rect 67634 1708 67640 1760
rect 67692 1748 67698 1760
rect 68189 1751 68247 1757
rect 68189 1748 68201 1751
rect 67692 1720 68201 1748
rect 67692 1708 67698 1720
rect 68189 1717 68201 1720
rect 68235 1717 68247 1751
rect 68189 1711 68247 1717
rect 69198 1708 69204 1760
rect 69256 1748 69262 1760
rect 69569 1751 69627 1757
rect 69569 1748 69581 1751
rect 69256 1720 69581 1748
rect 69256 1708 69262 1720
rect 69569 1717 69581 1720
rect 69615 1717 69627 1751
rect 69569 1711 69627 1717
rect 1104 1658 72864 1680
rect 1104 1606 9078 1658
rect 9130 1606 21078 1658
rect 21130 1606 33078 1658
rect 33130 1606 45078 1658
rect 45130 1606 57078 1658
rect 57130 1606 69078 1658
rect 69130 1606 72864 1658
rect 1104 1584 72864 1606
rect 1118 1504 1124 1556
rect 1176 1544 1182 1556
rect 2777 1547 2835 1553
rect 2777 1544 2789 1547
rect 1176 1516 2789 1544
rect 1176 1504 1182 1516
rect 2777 1513 2789 1516
rect 2823 1513 2835 1547
rect 2777 1507 2835 1513
rect 24026 1504 24032 1556
rect 24084 1544 24090 1556
rect 24857 1547 24915 1553
rect 24857 1544 24869 1547
rect 24084 1516 24869 1544
rect 24084 1504 24090 1516
rect 24857 1513 24869 1516
rect 24903 1513 24915 1547
rect 24857 1507 24915 1513
rect 25406 1504 25412 1556
rect 25464 1544 25470 1556
rect 26329 1547 26387 1553
rect 26329 1544 26341 1547
rect 25464 1516 26341 1544
rect 25464 1504 25470 1516
rect 26329 1513 26341 1516
rect 26375 1513 26387 1547
rect 26329 1507 26387 1513
rect 27430 1504 27436 1556
rect 27488 1544 27494 1556
rect 28721 1547 28779 1553
rect 28721 1544 28733 1547
rect 27488 1516 28733 1544
rect 27488 1504 27494 1516
rect 28721 1513 28733 1516
rect 28767 1513 28779 1547
rect 28721 1507 28779 1513
rect 29546 1504 29552 1556
rect 29604 1544 29610 1556
rect 30837 1547 30895 1553
rect 30837 1544 30849 1547
rect 29604 1516 30849 1544
rect 29604 1504 29610 1516
rect 30837 1513 30849 1516
rect 30883 1513 30895 1547
rect 30837 1507 30895 1513
rect 31202 1504 31208 1556
rect 31260 1544 31266 1556
rect 32125 1547 32183 1553
rect 32125 1544 32137 1547
rect 31260 1516 32137 1544
rect 31260 1504 31266 1516
rect 32125 1513 32137 1516
rect 32171 1513 32183 1547
rect 32125 1507 32183 1513
rect 2133 1479 2191 1485
rect 2133 1445 2145 1479
rect 2179 1476 2191 1479
rect 2498 1476 2504 1488
rect 2179 1448 2504 1476
rect 2179 1445 2191 1448
rect 2133 1439 2191 1445
rect 2498 1436 2504 1448
rect 2556 1436 2562 1488
rect 3326 1436 3332 1488
rect 3384 1476 3390 1488
rect 4157 1479 4215 1485
rect 4157 1476 4169 1479
rect 3384 1448 4169 1476
rect 3384 1436 3390 1448
rect 4157 1445 4169 1448
rect 4203 1445 4215 1479
rect 4157 1439 4215 1445
rect 4430 1436 4436 1488
rect 4488 1476 4494 1488
rect 4709 1479 4767 1485
rect 4709 1476 4721 1479
rect 4488 1448 4721 1476
rect 4488 1436 4494 1448
rect 4709 1445 4721 1448
rect 4755 1445 4767 1479
rect 4709 1439 4767 1445
rect 4982 1436 4988 1488
rect 5040 1476 5046 1488
rect 5353 1479 5411 1485
rect 5353 1476 5365 1479
rect 5040 1448 5365 1476
rect 5040 1436 5046 1448
rect 5353 1445 5365 1448
rect 5399 1445 5411 1479
rect 5353 1439 5411 1445
rect 7742 1436 7748 1488
rect 7800 1476 7806 1488
rect 8113 1479 8171 1485
rect 8113 1476 8125 1479
rect 7800 1448 8125 1476
rect 7800 1436 7806 1448
rect 8113 1445 8125 1448
rect 8159 1445 8171 1479
rect 8113 1439 8171 1445
rect 9306 1436 9312 1488
rect 9364 1476 9370 1488
rect 9585 1479 9643 1485
rect 9585 1476 9597 1479
rect 9364 1448 9597 1476
rect 9364 1436 9370 1448
rect 9585 1445 9597 1448
rect 9631 1445 9643 1479
rect 9585 1439 9643 1445
rect 9950 1436 9956 1488
rect 10008 1476 10014 1488
rect 10321 1479 10379 1485
rect 10321 1476 10333 1479
rect 10008 1448 10333 1476
rect 10008 1436 10014 1448
rect 10321 1445 10333 1448
rect 10367 1445 10379 1479
rect 10321 1439 10379 1445
rect 11882 1436 11888 1488
rect 11940 1476 11946 1488
rect 12253 1479 12311 1485
rect 12253 1476 12265 1479
rect 11940 1448 12265 1476
rect 11940 1436 11946 1448
rect 12253 1445 12265 1448
rect 12299 1445 12311 1479
rect 12253 1439 12311 1445
rect 12710 1436 12716 1488
rect 12768 1476 12774 1488
rect 12989 1479 13047 1485
rect 12989 1476 13001 1479
rect 12768 1448 13001 1476
rect 12768 1436 12774 1448
rect 12989 1445 13001 1448
rect 13035 1445 13047 1479
rect 12989 1439 13047 1445
rect 13538 1436 13544 1488
rect 13596 1476 13602 1488
rect 13817 1479 13875 1485
rect 13817 1476 13829 1479
rect 13596 1448 13829 1476
rect 13596 1436 13602 1448
rect 13817 1445 13829 1448
rect 13863 1445 13875 1479
rect 13817 1439 13875 1445
rect 14090 1436 14096 1488
rect 14148 1476 14154 1488
rect 14553 1479 14611 1485
rect 14553 1476 14565 1479
rect 14148 1448 14565 1476
rect 14148 1436 14154 1448
rect 14553 1445 14565 1448
rect 14599 1445 14611 1479
rect 14553 1439 14611 1445
rect 15194 1436 15200 1488
rect 15252 1476 15258 1488
rect 15565 1479 15623 1485
rect 15565 1476 15577 1479
rect 15252 1448 15577 1476
rect 15252 1436 15258 1448
rect 15565 1445 15577 1448
rect 15611 1445 15623 1479
rect 15565 1439 15623 1445
rect 16298 1436 16304 1488
rect 16356 1476 16362 1488
rect 16577 1479 16635 1485
rect 16577 1476 16589 1479
rect 16356 1448 16589 1476
rect 16356 1436 16362 1448
rect 16577 1445 16589 1448
rect 16623 1445 16635 1479
rect 16577 1439 16635 1445
rect 17126 1436 17132 1488
rect 17184 1476 17190 1488
rect 17497 1479 17555 1485
rect 17497 1476 17509 1479
rect 17184 1448 17509 1476
rect 17184 1436 17190 1448
rect 17497 1445 17509 1448
rect 17543 1445 17555 1479
rect 17497 1439 17555 1445
rect 17954 1436 17960 1488
rect 18012 1476 18018 1488
rect 18325 1479 18383 1485
rect 18325 1476 18337 1479
rect 18012 1448 18337 1476
rect 18012 1436 18018 1448
rect 18325 1445 18337 1448
rect 18371 1445 18383 1479
rect 18325 1439 18383 1445
rect 18782 1436 18788 1488
rect 18840 1476 18846 1488
rect 19153 1479 19211 1485
rect 19153 1476 19165 1479
rect 18840 1448 19165 1476
rect 18840 1436 18846 1448
rect 19153 1445 19165 1448
rect 19199 1445 19211 1479
rect 19153 1439 19211 1445
rect 20162 1436 20168 1488
rect 20220 1476 20226 1488
rect 20625 1479 20683 1485
rect 20625 1476 20637 1479
rect 20220 1448 20637 1476
rect 20220 1436 20226 1448
rect 20625 1445 20637 1448
rect 20671 1445 20683 1479
rect 20625 1439 20683 1445
rect 21266 1436 21272 1488
rect 21324 1476 21330 1488
rect 21453 1479 21511 1485
rect 21453 1476 21465 1479
rect 21324 1448 21465 1476
rect 21324 1436 21330 1448
rect 21453 1445 21465 1448
rect 21499 1445 21511 1479
rect 21453 1439 21511 1445
rect 22646 1436 22652 1488
rect 22704 1476 22710 1488
rect 23385 1479 23443 1485
rect 23385 1476 23397 1479
rect 22704 1448 23397 1476
rect 22704 1436 22710 1448
rect 23385 1445 23397 1448
rect 23431 1445 23443 1479
rect 23385 1439 23443 1445
rect 23474 1436 23480 1488
rect 23532 1476 23538 1488
rect 24305 1479 24363 1485
rect 24305 1476 24317 1479
rect 23532 1448 24317 1476
rect 23532 1436 23538 1448
rect 24305 1445 24317 1448
rect 24351 1445 24363 1479
rect 24305 1439 24363 1445
rect 24578 1436 24584 1488
rect 24636 1476 24642 1488
rect 25501 1479 25559 1485
rect 25501 1476 25513 1479
rect 24636 1448 25513 1476
rect 24636 1436 24642 1448
rect 25501 1445 25513 1448
rect 25547 1445 25559 1479
rect 25501 1439 25559 1445
rect 26510 1436 26516 1488
rect 26568 1476 26574 1488
rect 27341 1479 27399 1485
rect 27341 1476 27353 1479
rect 26568 1448 27353 1476
rect 26568 1436 26574 1448
rect 27341 1445 27353 1448
rect 27387 1445 27399 1479
rect 27341 1439 27399 1445
rect 27890 1436 27896 1488
rect 27948 1476 27954 1488
rect 28997 1479 29055 1485
rect 28997 1476 29009 1479
rect 27948 1448 29009 1476
rect 27948 1436 27954 1448
rect 28997 1445 29009 1448
rect 29043 1445 29055 1479
rect 28997 1439 29055 1445
rect 29270 1436 29276 1488
rect 29328 1476 29334 1488
rect 30561 1479 30619 1485
rect 30561 1476 30573 1479
rect 29328 1448 30573 1476
rect 29328 1436 29334 1448
rect 30561 1445 30573 1448
rect 30607 1445 30619 1479
rect 30561 1439 30619 1445
rect 30650 1436 30656 1488
rect 30708 1476 30714 1488
rect 31573 1479 31631 1485
rect 31573 1476 31585 1479
rect 30708 1448 31585 1476
rect 30708 1436 30714 1448
rect 31573 1445 31585 1448
rect 31619 1445 31631 1479
rect 31573 1439 31631 1445
rect 32030 1436 32036 1488
rect 32088 1476 32094 1488
rect 32861 1479 32919 1485
rect 32861 1476 32873 1479
rect 32088 1448 32873 1476
rect 32088 1436 32094 1448
rect 32861 1445 32873 1448
rect 32907 1445 32919 1479
rect 32861 1439 32919 1445
rect 37829 1479 37887 1485
rect 37829 1445 37841 1479
rect 37875 1476 37887 1479
rect 38102 1476 38108 1488
rect 37875 1448 38108 1476
rect 37875 1445 37887 1448
rect 37829 1439 37887 1445
rect 38102 1436 38108 1448
rect 38160 1436 38166 1488
rect 39117 1479 39175 1485
rect 39117 1445 39129 1479
rect 39163 1476 39175 1479
rect 39482 1476 39488 1488
rect 39163 1448 39488 1476
rect 39163 1445 39175 1448
rect 39117 1439 39175 1445
rect 39482 1436 39488 1448
rect 39540 1436 39546 1488
rect 40221 1479 40279 1485
rect 40221 1445 40233 1479
rect 40267 1476 40279 1479
rect 40586 1476 40592 1488
rect 40267 1448 40592 1476
rect 40267 1445 40279 1448
rect 40221 1439 40279 1445
rect 40586 1436 40592 1448
rect 40644 1436 40650 1488
rect 41417 1479 41475 1485
rect 41417 1445 41429 1479
rect 41463 1476 41475 1479
rect 41690 1476 41696 1488
rect 41463 1448 41696 1476
rect 41463 1445 41475 1448
rect 41417 1439 41475 1445
rect 41690 1436 41696 1448
rect 41748 1436 41754 1488
rect 41969 1479 42027 1485
rect 41969 1445 41981 1479
rect 42015 1476 42027 1479
rect 42242 1476 42248 1488
rect 42015 1448 42248 1476
rect 42015 1445 42027 1448
rect 41969 1439 42027 1445
rect 42242 1436 42248 1448
rect 42300 1436 42306 1488
rect 42521 1479 42579 1485
rect 42521 1445 42533 1479
rect 42567 1476 42579 1479
rect 42794 1476 42800 1488
rect 42567 1448 42800 1476
rect 42567 1445 42579 1448
rect 42521 1439 42579 1445
rect 42794 1436 42800 1448
rect 42852 1436 42858 1488
rect 43073 1479 43131 1485
rect 43073 1445 43085 1479
rect 43119 1476 43131 1479
rect 43346 1476 43352 1488
rect 43119 1448 43352 1476
rect 43119 1445 43131 1448
rect 43073 1439 43131 1445
rect 43346 1436 43352 1448
rect 43404 1436 43410 1488
rect 59906 1436 59912 1488
rect 59964 1476 59970 1488
rect 60185 1479 60243 1485
rect 60185 1476 60197 1479
rect 59964 1448 60197 1476
rect 59964 1436 59970 1448
rect 60185 1445 60197 1448
rect 60231 1445 60243 1479
rect 60185 1439 60243 1445
rect 60734 1436 60740 1488
rect 60792 1476 60798 1488
rect 61013 1479 61071 1485
rect 61013 1476 61025 1479
rect 60792 1448 61025 1476
rect 60792 1436 60798 1448
rect 61013 1445 61025 1448
rect 61059 1445 61071 1479
rect 61013 1439 61071 1445
rect 61286 1436 61292 1488
rect 61344 1476 61350 1488
rect 61565 1479 61623 1485
rect 61565 1476 61577 1479
rect 61344 1448 61577 1476
rect 61344 1436 61350 1448
rect 61565 1445 61577 1448
rect 61611 1445 61623 1479
rect 61565 1439 61623 1445
rect 61838 1436 61844 1488
rect 61896 1476 61902 1488
rect 62117 1479 62175 1485
rect 62117 1476 62129 1479
rect 61896 1448 62129 1476
rect 61896 1436 61902 1448
rect 62117 1445 62129 1448
rect 62163 1445 62175 1479
rect 62117 1439 62175 1445
rect 64598 1436 64604 1488
rect 64656 1476 64662 1488
rect 65245 1479 65303 1485
rect 65245 1476 65257 1479
rect 64656 1448 65257 1476
rect 64656 1436 64662 1448
rect 65245 1445 65257 1448
rect 65291 1445 65303 1479
rect 65245 1439 65303 1445
rect 65702 1436 65708 1488
rect 65760 1476 65766 1488
rect 66441 1479 66499 1485
rect 66441 1476 66453 1479
rect 65760 1448 66453 1476
rect 65760 1436 65766 1448
rect 66441 1445 66453 1448
rect 66487 1445 66499 1479
rect 66441 1439 66499 1445
rect 66530 1436 66536 1488
rect 66588 1476 66594 1488
rect 67269 1479 67327 1485
rect 67269 1476 67281 1479
rect 66588 1448 67281 1476
rect 66588 1436 66594 1448
rect 67269 1445 67281 1448
rect 67315 1445 67327 1479
rect 67269 1439 67327 1445
rect 67910 1436 67916 1488
rect 67968 1476 67974 1488
rect 68465 1479 68523 1485
rect 68465 1476 68477 1479
rect 67968 1448 68477 1476
rect 67968 1436 67974 1448
rect 68465 1445 68477 1448
rect 68511 1445 68523 1479
rect 68465 1439 68523 1445
rect 68738 1436 68744 1488
rect 68796 1476 68802 1488
rect 69293 1479 69351 1485
rect 69293 1476 69305 1479
rect 68796 1448 69305 1476
rect 68796 1436 68802 1448
rect 69293 1445 69305 1448
rect 69339 1445 69351 1479
rect 69293 1439 69351 1445
rect 69566 1436 69572 1488
rect 69624 1476 69630 1488
rect 70029 1479 70087 1485
rect 70029 1476 70041 1479
rect 69624 1448 70041 1476
rect 69624 1436 69630 1448
rect 70029 1445 70041 1448
rect 70075 1445 70087 1479
rect 70029 1439 70087 1445
rect 1670 1408 1676 1420
rect 1631 1380 1676 1408
rect 1670 1368 1676 1380
rect 1728 1368 1734 1420
rect 1762 1368 1768 1420
rect 1820 1408 1826 1420
rect 3053 1411 3111 1417
rect 3053 1408 3065 1411
rect 1820 1380 3065 1408
rect 1820 1368 1826 1380
rect 3053 1377 3065 1380
rect 3099 1377 3111 1411
rect 3053 1371 3111 1377
rect 5258 1368 5264 1420
rect 5316 1408 5322 1420
rect 5629 1411 5687 1417
rect 5629 1408 5641 1411
rect 5316 1380 5641 1408
rect 5316 1368 5322 1380
rect 5629 1377 5641 1380
rect 5675 1377 5687 1411
rect 5629 1371 5687 1377
rect 5810 1368 5816 1420
rect 5868 1408 5874 1420
rect 6181 1411 6239 1417
rect 6181 1408 6193 1411
rect 5868 1380 6193 1408
rect 5868 1368 5874 1380
rect 6181 1377 6193 1380
rect 6227 1377 6239 1411
rect 6181 1371 6239 1377
rect 6362 1368 6368 1420
rect 6420 1408 6426 1420
rect 6825 1411 6883 1417
rect 6825 1408 6837 1411
rect 6420 1380 6837 1408
rect 6420 1368 6426 1380
rect 6825 1377 6837 1380
rect 6871 1377 6883 1411
rect 6825 1371 6883 1377
rect 7190 1368 7196 1420
rect 7248 1408 7254 1420
rect 7561 1411 7619 1417
rect 7561 1408 7573 1411
rect 7248 1380 7573 1408
rect 7248 1368 7254 1380
rect 7561 1377 7573 1380
rect 7607 1377 7619 1411
rect 7561 1371 7619 1377
rect 8018 1368 8024 1420
rect 8076 1408 8082 1420
rect 8389 1411 8447 1417
rect 8389 1408 8401 1411
rect 8076 1380 8401 1408
rect 8076 1368 8082 1380
rect 8389 1377 8401 1380
rect 8435 1377 8447 1411
rect 8389 1371 8447 1377
rect 10226 1368 10232 1420
rect 10284 1408 10290 1420
rect 10597 1411 10655 1417
rect 10597 1408 10609 1411
rect 10284 1380 10609 1408
rect 10284 1368 10290 1380
rect 10597 1377 10609 1380
rect 10643 1377 10655 1411
rect 10597 1371 10655 1377
rect 10778 1368 10784 1420
rect 10836 1408 10842 1420
rect 11241 1411 11299 1417
rect 11241 1408 11253 1411
rect 10836 1380 11253 1408
rect 10836 1368 10842 1380
rect 11241 1377 11253 1380
rect 11287 1377 11299 1411
rect 11241 1371 11299 1377
rect 12158 1368 12164 1420
rect 12216 1408 12222 1420
rect 13265 1411 13323 1417
rect 13265 1408 13277 1411
rect 12216 1380 13277 1408
rect 12216 1368 12222 1380
rect 13265 1377 13277 1380
rect 13311 1377 13323 1411
rect 13265 1371 13323 1377
rect 15470 1368 15476 1420
rect 15528 1408 15534 1420
rect 15841 1411 15899 1417
rect 15841 1408 15853 1411
rect 15528 1380 15853 1408
rect 15528 1368 15534 1380
rect 15841 1377 15853 1380
rect 15887 1377 15899 1411
rect 15841 1371 15899 1377
rect 17402 1368 17408 1420
rect 17460 1408 17466 1420
rect 17773 1411 17831 1417
rect 17773 1408 17785 1411
rect 17460 1380 17785 1408
rect 17460 1368 17466 1380
rect 17773 1377 17785 1380
rect 17819 1377 17831 1411
rect 17773 1371 17831 1377
rect 18230 1368 18236 1420
rect 18288 1408 18294 1420
rect 18601 1411 18659 1417
rect 18601 1408 18613 1411
rect 18288 1380 18613 1408
rect 18288 1368 18294 1380
rect 18601 1377 18613 1380
rect 18647 1377 18659 1411
rect 18601 1371 18659 1377
rect 19058 1368 19064 1420
rect 19116 1408 19122 1420
rect 19429 1411 19487 1417
rect 19429 1408 19441 1411
rect 19116 1380 19441 1408
rect 19116 1368 19122 1380
rect 19429 1377 19441 1380
rect 19475 1377 19487 1411
rect 19429 1371 19487 1377
rect 20714 1368 20720 1420
rect 20772 1408 20778 1420
rect 21177 1411 21235 1417
rect 21177 1408 21189 1411
rect 20772 1380 21189 1408
rect 20772 1368 20778 1380
rect 21177 1377 21189 1380
rect 21223 1377 21235 1411
rect 21177 1371 21235 1377
rect 21542 1368 21548 1420
rect 21600 1408 21606 1420
rect 22097 1411 22155 1417
rect 22097 1408 22109 1411
rect 21600 1380 22109 1408
rect 21600 1368 21606 1380
rect 22097 1377 22109 1380
rect 22143 1377 22155 1411
rect 22097 1371 22155 1377
rect 22370 1368 22376 1420
rect 22428 1408 22434 1420
rect 23109 1411 23167 1417
rect 23109 1408 23121 1411
rect 22428 1380 23121 1408
rect 22428 1368 22434 1380
rect 23109 1377 23121 1380
rect 23155 1377 23167 1411
rect 23109 1371 23167 1377
rect 23198 1368 23204 1420
rect 23256 1408 23262 1420
rect 23753 1411 23811 1417
rect 23753 1408 23765 1411
rect 23256 1380 23765 1408
rect 23256 1368 23262 1380
rect 23753 1377 23765 1380
rect 23799 1377 23811 1411
rect 25225 1411 25283 1417
rect 25225 1408 25237 1411
rect 23753 1371 23811 1377
rect 24320 1380 25237 1408
rect 24320 1352 24348 1380
rect 25225 1377 25237 1380
rect 25271 1377 25283 1411
rect 25777 1411 25835 1417
rect 25777 1408 25789 1411
rect 25225 1371 25283 1377
rect 25424 1380 25789 1408
rect 566 1300 572 1352
rect 624 1340 630 1352
rect 2225 1343 2283 1349
rect 2225 1340 2237 1343
rect 624 1312 2237 1340
rect 624 1300 630 1312
rect 2225 1309 2237 1312
rect 2271 1309 2283 1343
rect 2225 1303 2283 1309
rect 2501 1343 2559 1349
rect 2501 1309 2513 1343
rect 2547 1309 2559 1343
rect 2501 1303 2559 1309
rect 3329 1343 3387 1349
rect 3329 1309 3341 1343
rect 3375 1309 3387 1343
rect 3329 1303 3387 1309
rect 842 1232 848 1284
rect 900 1272 906 1284
rect 2516 1272 2544 1303
rect 900 1244 2544 1272
rect 900 1232 906 1244
rect 1946 1164 1952 1216
rect 2004 1204 2010 1216
rect 3344 1204 3372 1303
rect 3602 1300 3608 1352
rect 3660 1340 3666 1352
rect 3881 1343 3939 1349
rect 3881 1340 3893 1343
rect 3660 1312 3893 1340
rect 3660 1300 3666 1312
rect 3881 1309 3893 1312
rect 3927 1309 3939 1343
rect 3881 1303 3939 1309
rect 4246 1300 4252 1352
rect 4304 1340 4310 1352
rect 4433 1343 4491 1349
rect 4433 1340 4445 1343
rect 4304 1312 4445 1340
rect 4304 1300 4310 1312
rect 4433 1309 4445 1312
rect 4479 1309 4491 1343
rect 4433 1303 4491 1309
rect 4706 1300 4712 1352
rect 4764 1340 4770 1352
rect 5077 1343 5135 1349
rect 5077 1340 5089 1343
rect 4764 1312 5089 1340
rect 4764 1300 4770 1312
rect 5077 1309 5089 1312
rect 5123 1309 5135 1343
rect 5077 1303 5135 1309
rect 5534 1300 5540 1352
rect 5592 1340 5598 1352
rect 5905 1343 5963 1349
rect 5905 1340 5917 1343
rect 5592 1312 5917 1340
rect 5592 1300 5598 1312
rect 5905 1309 5917 1312
rect 5951 1309 5963 1343
rect 5905 1303 5963 1309
rect 6086 1300 6092 1352
rect 6144 1340 6150 1352
rect 6549 1343 6607 1349
rect 6549 1340 6561 1343
rect 6144 1312 6561 1340
rect 6144 1300 6150 1312
rect 6549 1309 6561 1312
rect 6595 1309 6607 1343
rect 6549 1303 6607 1309
rect 6914 1300 6920 1352
rect 6972 1340 6978 1352
rect 7285 1343 7343 1349
rect 7285 1340 7297 1343
rect 6972 1312 7297 1340
rect 6972 1300 6978 1312
rect 7285 1309 7297 1312
rect 7331 1309 7343 1343
rect 7285 1303 7343 1309
rect 7466 1300 7472 1352
rect 7524 1340 7530 1352
rect 7837 1343 7895 1349
rect 7837 1340 7849 1343
rect 7524 1312 7849 1340
rect 7524 1300 7530 1312
rect 7837 1309 7849 1312
rect 7883 1309 7895 1343
rect 7837 1303 7895 1309
rect 8294 1300 8300 1352
rect 8352 1340 8358 1352
rect 8757 1343 8815 1349
rect 8757 1340 8769 1343
rect 8352 1312 8769 1340
rect 8352 1300 8358 1312
rect 8757 1309 8769 1312
rect 8803 1309 8815 1343
rect 8757 1303 8815 1309
rect 8846 1300 8852 1352
rect 8904 1340 8910 1352
rect 9309 1343 9367 1349
rect 9309 1340 9321 1343
rect 8904 1312 9321 1340
rect 8904 1300 8910 1312
rect 9309 1309 9321 1312
rect 9355 1309 9367 1343
rect 9309 1303 9367 1309
rect 9674 1300 9680 1352
rect 9732 1340 9738 1352
rect 10045 1343 10103 1349
rect 10045 1340 10057 1343
rect 9732 1312 10057 1340
rect 9732 1300 9738 1312
rect 10045 1309 10057 1312
rect 10091 1309 10103 1343
rect 10045 1303 10103 1309
rect 10502 1300 10508 1352
rect 10560 1340 10566 1352
rect 10965 1343 11023 1349
rect 10965 1340 10977 1343
rect 10560 1312 10977 1340
rect 10560 1300 10566 1312
rect 10965 1309 10977 1312
rect 11011 1309 11023 1343
rect 10965 1303 11023 1309
rect 11054 1300 11060 1352
rect 11112 1340 11118 1352
rect 11517 1343 11575 1349
rect 11517 1340 11529 1343
rect 11112 1312 11529 1340
rect 11112 1300 11118 1312
rect 11517 1309 11529 1312
rect 11563 1309 11575 1343
rect 11517 1303 11575 1309
rect 11885 1343 11943 1349
rect 11885 1309 11897 1343
rect 11931 1309 11943 1343
rect 11885 1303 11943 1309
rect 11330 1232 11336 1284
rect 11388 1272 11394 1284
rect 11900 1272 11928 1303
rect 12434 1300 12440 1352
rect 12492 1340 12498 1352
rect 12713 1343 12771 1349
rect 12713 1340 12725 1343
rect 12492 1312 12725 1340
rect 12492 1300 12498 1312
rect 12713 1309 12725 1312
rect 12759 1309 12771 1343
rect 12713 1303 12771 1309
rect 13354 1300 13360 1352
rect 13412 1340 13418 1352
rect 13541 1343 13599 1349
rect 13541 1340 13553 1343
rect 13412 1312 13553 1340
rect 13412 1300 13418 1312
rect 13541 1309 13553 1312
rect 13587 1309 13599 1343
rect 13541 1303 13599 1309
rect 13814 1300 13820 1352
rect 13872 1340 13878 1352
rect 14093 1343 14151 1349
rect 14093 1340 14105 1343
rect 13872 1312 14105 1340
rect 13872 1300 13878 1312
rect 14093 1309 14105 1312
rect 14139 1309 14151 1343
rect 14093 1303 14151 1309
rect 14642 1300 14648 1352
rect 14700 1340 14706 1352
rect 14921 1343 14979 1349
rect 14921 1340 14933 1343
rect 14700 1312 14933 1340
rect 14700 1300 14706 1312
rect 14921 1309 14933 1312
rect 14967 1309 14979 1343
rect 14921 1303 14979 1309
rect 15197 1343 15255 1349
rect 15197 1309 15209 1343
rect 15243 1309 15255 1343
rect 15197 1303 15255 1309
rect 11388 1244 11928 1272
rect 11388 1232 11394 1244
rect 14366 1232 14372 1284
rect 14424 1272 14430 1284
rect 15212 1272 15240 1303
rect 16022 1300 16028 1352
rect 16080 1340 16086 1352
rect 16301 1343 16359 1349
rect 16301 1340 16313 1343
rect 16080 1312 16313 1340
rect 16080 1300 16086 1312
rect 16301 1309 16313 1312
rect 16347 1309 16359 1343
rect 16850 1340 16856 1352
rect 16811 1312 16856 1340
rect 16301 1303 16359 1309
rect 16850 1300 16856 1312
rect 16908 1300 16914 1352
rect 17221 1343 17279 1349
rect 17221 1309 17233 1343
rect 17267 1309 17279 1343
rect 17221 1303 17279 1309
rect 14424 1244 15240 1272
rect 14424 1232 14430 1244
rect 16574 1232 16580 1284
rect 16632 1272 16638 1284
rect 17236 1272 17264 1303
rect 17678 1300 17684 1352
rect 17736 1340 17742 1352
rect 18049 1343 18107 1349
rect 18049 1340 18061 1343
rect 17736 1312 18061 1340
rect 17736 1300 17742 1312
rect 18049 1309 18061 1312
rect 18095 1309 18107 1343
rect 18049 1303 18107 1309
rect 18506 1300 18512 1352
rect 18564 1340 18570 1352
rect 18877 1343 18935 1349
rect 18877 1340 18889 1343
rect 18564 1312 18889 1340
rect 18564 1300 18570 1312
rect 18877 1309 18889 1312
rect 18923 1309 18935 1343
rect 18877 1303 18935 1309
rect 19334 1300 19340 1352
rect 19392 1340 19398 1352
rect 19889 1343 19947 1349
rect 19889 1340 19901 1343
rect 19392 1312 19901 1340
rect 19392 1300 19398 1312
rect 19889 1309 19901 1312
rect 19935 1309 19947 1343
rect 19889 1303 19947 1309
rect 20165 1343 20223 1349
rect 20165 1309 20177 1343
rect 20211 1309 20223 1343
rect 20165 1303 20223 1309
rect 20901 1343 20959 1349
rect 20901 1309 20913 1343
rect 20947 1309 20959 1343
rect 20901 1303 20959 1309
rect 16632 1244 17264 1272
rect 16632 1232 16638 1244
rect 19610 1232 19616 1284
rect 19668 1272 19674 1284
rect 20180 1272 20208 1303
rect 19668 1244 20208 1272
rect 19668 1232 19674 1244
rect 20438 1232 20444 1284
rect 20496 1272 20502 1284
rect 20916 1272 20944 1303
rect 21266 1300 21272 1352
rect 21324 1340 21330 1352
rect 21729 1343 21787 1349
rect 21729 1340 21741 1343
rect 21324 1312 21741 1340
rect 21324 1300 21330 1312
rect 21729 1309 21741 1312
rect 21775 1309 21787 1343
rect 21729 1303 21787 1309
rect 21818 1300 21824 1352
rect 21876 1340 21882 1352
rect 22557 1343 22615 1349
rect 22557 1340 22569 1343
rect 21876 1312 22569 1340
rect 21876 1300 21882 1312
rect 22557 1309 22569 1312
rect 22603 1309 22615 1343
rect 22557 1303 22615 1309
rect 22833 1343 22891 1349
rect 22833 1309 22845 1343
rect 22879 1309 22891 1343
rect 24029 1343 24087 1349
rect 24029 1340 24041 1343
rect 22833 1303 22891 1309
rect 23538 1312 24041 1340
rect 20496 1244 20944 1272
rect 20496 1232 20502 1244
rect 22094 1232 22100 1284
rect 22152 1272 22158 1284
rect 22848 1272 22876 1303
rect 22152 1244 22876 1272
rect 22152 1232 22158 1244
rect 22922 1232 22928 1284
rect 22980 1272 22986 1284
rect 23538 1272 23566 1312
rect 24029 1309 24041 1312
rect 24075 1309 24087 1343
rect 24029 1303 24087 1309
rect 24302 1300 24308 1352
rect 24360 1300 24366 1352
rect 24581 1343 24639 1349
rect 24581 1309 24593 1343
rect 24627 1309 24639 1343
rect 24581 1303 24639 1309
rect 22980 1244 23566 1272
rect 22980 1232 22986 1244
rect 23750 1232 23756 1284
rect 23808 1272 23814 1284
rect 24596 1272 24624 1303
rect 24854 1300 24860 1352
rect 24912 1340 24918 1352
rect 25424 1340 25452 1380
rect 25777 1377 25789 1380
rect 25823 1377 25835 1411
rect 25777 1371 25835 1377
rect 26234 1368 26240 1420
rect 26292 1408 26298 1420
rect 26973 1411 27031 1417
rect 26973 1408 26985 1411
rect 26292 1380 26985 1408
rect 26292 1368 26298 1380
rect 26973 1377 26985 1380
rect 27019 1377 27031 1411
rect 26973 1371 27031 1377
rect 27614 1368 27620 1420
rect 27672 1408 27678 1420
rect 28445 1411 28503 1417
rect 28445 1408 28457 1411
rect 27672 1380 28457 1408
rect 27672 1368 27678 1380
rect 28445 1377 28457 1380
rect 28491 1377 28503 1411
rect 28445 1371 28503 1377
rect 28718 1368 28724 1420
rect 28776 1408 28782 1420
rect 29825 1411 29883 1417
rect 29825 1408 29837 1411
rect 28776 1380 29837 1408
rect 28776 1368 28782 1380
rect 29825 1377 29837 1380
rect 29871 1377 29883 1411
rect 29825 1371 29883 1377
rect 30374 1368 30380 1420
rect 30432 1408 30438 1420
rect 31297 1411 31355 1417
rect 31297 1408 31309 1411
rect 30432 1380 31309 1408
rect 30432 1368 30438 1380
rect 31297 1377 31309 1380
rect 31343 1377 31355 1411
rect 31297 1371 31355 1377
rect 32306 1368 32312 1420
rect 32364 1408 32370 1420
rect 33229 1411 33287 1417
rect 33229 1408 33241 1411
rect 32364 1380 33241 1408
rect 32364 1368 32370 1380
rect 33229 1377 33241 1380
rect 33275 1377 33287 1411
rect 33229 1371 33287 1377
rect 38841 1411 38899 1417
rect 38841 1377 38853 1411
rect 38887 1408 38899 1411
rect 39206 1408 39212 1420
rect 38887 1380 39212 1408
rect 38887 1377 38899 1380
rect 38841 1371 38899 1377
rect 39206 1368 39212 1380
rect 39264 1368 39270 1420
rect 39393 1411 39451 1417
rect 39393 1377 39405 1411
rect 39439 1408 39451 1411
rect 39758 1408 39764 1420
rect 39439 1380 39764 1408
rect 39439 1377 39451 1380
rect 39393 1371 39451 1377
rect 39758 1368 39764 1380
rect 39816 1368 39822 1420
rect 39945 1411 40003 1417
rect 39945 1377 39957 1411
rect 39991 1408 40003 1411
rect 40310 1408 40316 1420
rect 39991 1380 40316 1408
rect 39991 1377 40003 1380
rect 39945 1371 40003 1377
rect 40310 1368 40316 1380
rect 40368 1368 40374 1420
rect 40773 1411 40831 1417
rect 40773 1377 40785 1411
rect 40819 1408 40831 1411
rect 41138 1408 41144 1420
rect 40819 1380 41144 1408
rect 40819 1377 40831 1380
rect 40773 1371 40831 1377
rect 41138 1368 41144 1380
rect 41196 1368 41202 1420
rect 49142 1368 49148 1420
rect 49200 1408 49206 1420
rect 49513 1411 49571 1417
rect 49513 1408 49525 1411
rect 49200 1380 49525 1408
rect 49200 1368 49206 1380
rect 49513 1377 49525 1380
rect 49559 1377 49571 1411
rect 49513 1371 49571 1377
rect 49694 1368 49700 1420
rect 49752 1408 49758 1420
rect 50341 1411 50399 1417
rect 50341 1408 50353 1411
rect 49752 1380 50353 1408
rect 49752 1368 49758 1380
rect 50341 1377 50353 1380
rect 50387 1377 50399 1411
rect 50341 1371 50399 1377
rect 51902 1368 51908 1420
rect 51960 1408 51966 1420
rect 52365 1411 52423 1417
rect 52365 1408 52377 1411
rect 51960 1380 52377 1408
rect 51960 1368 51966 1380
rect 52365 1377 52377 1380
rect 52411 1377 52423 1411
rect 52365 1371 52423 1377
rect 62390 1368 62396 1420
rect 62448 1408 62454 1420
rect 62853 1411 62911 1417
rect 62853 1408 62865 1411
rect 62448 1380 62865 1408
rect 62448 1368 62454 1380
rect 62853 1377 62865 1380
rect 62899 1377 62911 1411
rect 62853 1371 62911 1377
rect 62942 1368 62948 1420
rect 63000 1408 63006 1420
rect 63405 1411 63463 1417
rect 63405 1408 63417 1411
rect 63000 1380 63417 1408
rect 63000 1368 63006 1380
rect 63405 1377 63417 1380
rect 63451 1377 63463 1411
rect 63405 1371 63463 1377
rect 64046 1368 64052 1420
rect 64104 1408 64110 1420
rect 64417 1411 64475 1417
rect 64417 1408 64429 1411
rect 64104 1380 64429 1408
rect 64104 1368 64110 1380
rect 64417 1377 64429 1380
rect 64463 1377 64475 1411
rect 64417 1371 64475 1377
rect 65426 1368 65432 1420
rect 65484 1408 65490 1420
rect 66165 1411 66223 1417
rect 66165 1408 66177 1411
rect 65484 1380 66177 1408
rect 65484 1368 65490 1380
rect 66165 1377 66177 1380
rect 66211 1377 66223 1411
rect 66165 1371 66223 1377
rect 66254 1368 66260 1420
rect 66312 1408 66318 1420
rect 66993 1411 67051 1417
rect 66993 1408 67005 1411
rect 66312 1380 67005 1408
rect 66312 1368 66318 1380
rect 66993 1377 67005 1380
rect 67039 1377 67051 1411
rect 66993 1371 67051 1377
rect 67358 1368 67364 1420
rect 67416 1408 67422 1420
rect 68189 1411 68247 1417
rect 68189 1408 68201 1411
rect 67416 1380 68201 1408
rect 67416 1368 67422 1380
rect 68189 1377 68201 1380
rect 68235 1377 68247 1411
rect 68189 1371 68247 1377
rect 69842 1368 69848 1420
rect 69900 1408 69906 1420
rect 70581 1411 70639 1417
rect 70581 1408 70593 1411
rect 69900 1380 70593 1408
rect 69900 1368 69906 1380
rect 70581 1377 70593 1380
rect 70627 1377 70639 1411
rect 70581 1371 70639 1377
rect 24912 1312 25452 1340
rect 26053 1343 26111 1349
rect 24912 1300 24918 1312
rect 26053 1309 26065 1343
rect 26099 1309 26111 1343
rect 26053 1303 26111 1309
rect 26605 1343 26663 1349
rect 26605 1309 26617 1343
rect 26651 1309 26663 1343
rect 26605 1303 26663 1309
rect 23808 1244 24624 1272
rect 23808 1232 23814 1244
rect 25130 1232 25136 1284
rect 25188 1272 25194 1284
rect 26068 1272 26096 1303
rect 25188 1244 26096 1272
rect 25188 1232 25194 1244
rect 2004 1176 3372 1204
rect 2004 1164 2010 1176
rect 25682 1164 25688 1216
rect 25740 1204 25746 1216
rect 26620 1204 26648 1303
rect 26786 1300 26792 1352
rect 26844 1340 26850 1352
rect 27893 1343 27951 1349
rect 27893 1340 27905 1343
rect 26844 1312 27905 1340
rect 26844 1300 26850 1312
rect 27893 1309 27905 1312
rect 27939 1309 27951 1343
rect 27893 1303 27951 1309
rect 28169 1343 28227 1349
rect 28169 1309 28181 1343
rect 28215 1309 28227 1343
rect 28169 1303 28227 1309
rect 27246 1232 27252 1284
rect 27304 1272 27310 1284
rect 28184 1272 28212 1303
rect 28258 1300 28264 1352
rect 28316 1340 28322 1352
rect 29273 1343 29331 1349
rect 29273 1340 29285 1343
rect 28316 1312 29285 1340
rect 28316 1300 28322 1312
rect 29273 1309 29285 1312
rect 29319 1309 29331 1343
rect 29273 1303 29331 1309
rect 29549 1343 29607 1349
rect 29549 1309 29561 1343
rect 29595 1309 29607 1343
rect 29549 1303 29607 1309
rect 30101 1343 30159 1349
rect 30101 1309 30113 1343
rect 30147 1309 30159 1343
rect 30101 1303 30159 1309
rect 29564 1272 29592 1303
rect 27304 1244 28212 1272
rect 28460 1244 29592 1272
rect 27304 1232 27310 1244
rect 28460 1216 28488 1244
rect 25740 1176 26648 1204
rect 25740 1164 25746 1176
rect 28442 1164 28448 1216
rect 28500 1164 28506 1216
rect 28994 1164 29000 1216
rect 29052 1204 29058 1216
rect 30116 1204 30144 1303
rect 30926 1300 30932 1352
rect 30984 1340 30990 1352
rect 31849 1343 31907 1349
rect 31849 1340 31861 1343
rect 30984 1312 31861 1340
rect 30984 1300 30990 1312
rect 31849 1309 31861 1312
rect 31895 1309 31907 1343
rect 31849 1303 31907 1309
rect 32585 1343 32643 1349
rect 32585 1309 32597 1343
rect 32631 1309 32643 1343
rect 32585 1303 32643 1309
rect 38105 1343 38163 1349
rect 38105 1309 38117 1343
rect 38151 1340 38163 1343
rect 38286 1340 38292 1352
rect 38151 1312 38292 1340
rect 38151 1309 38163 1312
rect 38105 1303 38163 1309
rect 31754 1232 31760 1284
rect 31812 1272 31818 1284
rect 32600 1272 32628 1303
rect 38286 1300 38292 1312
rect 38344 1300 38350 1352
rect 38381 1343 38439 1349
rect 38381 1309 38393 1343
rect 38427 1340 38439 1343
rect 38654 1340 38660 1352
rect 38427 1312 38660 1340
rect 38427 1309 38439 1312
rect 38381 1303 38439 1309
rect 38654 1300 38660 1312
rect 38712 1300 38718 1352
rect 39669 1343 39727 1349
rect 39669 1309 39681 1343
rect 39715 1340 39727 1343
rect 40034 1340 40040 1352
rect 39715 1312 40040 1340
rect 39715 1309 39727 1312
rect 39669 1303 39727 1309
rect 40034 1300 40040 1312
rect 40092 1300 40098 1352
rect 40497 1343 40555 1349
rect 40497 1309 40509 1343
rect 40543 1340 40555 1343
rect 40862 1340 40868 1352
rect 40543 1312 40868 1340
rect 40543 1309 40555 1312
rect 40497 1303 40555 1309
rect 40862 1300 40868 1312
rect 40920 1300 40926 1352
rect 41049 1343 41107 1349
rect 41049 1309 41061 1343
rect 41095 1340 41107 1343
rect 41322 1340 41328 1352
rect 41095 1312 41328 1340
rect 41095 1309 41107 1312
rect 41049 1303 41107 1309
rect 41322 1300 41328 1312
rect 41380 1300 41386 1352
rect 41693 1343 41751 1349
rect 41693 1309 41705 1343
rect 41739 1340 41751 1343
rect 41966 1340 41972 1352
rect 41739 1312 41972 1340
rect 41739 1309 41751 1312
rect 41693 1303 41751 1309
rect 41966 1300 41972 1312
rect 42024 1300 42030 1352
rect 42245 1343 42303 1349
rect 42245 1309 42257 1343
rect 42291 1340 42303 1343
rect 42518 1340 42524 1352
rect 42291 1312 42524 1340
rect 42291 1309 42303 1312
rect 42245 1303 42303 1309
rect 42518 1300 42524 1312
rect 42576 1300 42582 1352
rect 42797 1343 42855 1349
rect 42797 1309 42809 1343
rect 42843 1340 42855 1343
rect 43070 1340 43076 1352
rect 42843 1312 43076 1340
rect 42843 1309 42855 1312
rect 42797 1303 42855 1309
rect 43070 1300 43076 1312
rect 43128 1300 43134 1352
rect 43349 1343 43407 1349
rect 43349 1309 43361 1343
rect 43395 1340 43407 1343
rect 43622 1340 43628 1352
rect 43395 1312 43628 1340
rect 43395 1309 43407 1312
rect 43349 1303 43407 1309
rect 43622 1300 43628 1312
rect 43680 1300 43686 1352
rect 43717 1343 43775 1349
rect 43717 1309 43729 1343
rect 43763 1340 43775 1343
rect 43898 1340 43904 1352
rect 43763 1312 43904 1340
rect 43763 1309 43775 1312
rect 43717 1303 43775 1309
rect 43898 1300 43904 1312
rect 43956 1300 43962 1352
rect 44269 1343 44327 1349
rect 44269 1309 44281 1343
rect 44315 1340 44327 1343
rect 44450 1340 44456 1352
rect 44315 1312 44456 1340
rect 44315 1309 44327 1312
rect 44269 1303 44327 1309
rect 44450 1300 44456 1312
rect 44508 1300 44514 1352
rect 44545 1343 44603 1349
rect 44545 1309 44557 1343
rect 44591 1340 44603 1343
rect 44726 1340 44732 1352
rect 44591 1312 44732 1340
rect 44591 1309 44603 1312
rect 44545 1303 44603 1309
rect 44726 1300 44732 1312
rect 44784 1300 44790 1352
rect 44821 1343 44879 1349
rect 44821 1309 44833 1343
rect 44867 1340 44879 1343
rect 44910 1340 44916 1352
rect 44867 1312 44916 1340
rect 44867 1309 44879 1312
rect 44821 1303 44879 1309
rect 44910 1300 44916 1312
rect 44968 1300 44974 1352
rect 45097 1343 45155 1349
rect 45097 1309 45109 1343
rect 45143 1340 45155 1343
rect 45278 1340 45284 1352
rect 45143 1312 45284 1340
rect 45143 1309 45155 1312
rect 45097 1303 45155 1309
rect 45278 1300 45284 1312
rect 45336 1300 45342 1352
rect 45373 1343 45431 1349
rect 45373 1309 45385 1343
rect 45419 1340 45431 1343
rect 45554 1340 45560 1352
rect 45419 1312 45560 1340
rect 45419 1309 45431 1312
rect 45373 1303 45431 1309
rect 45554 1300 45560 1312
rect 45612 1300 45618 1352
rect 45649 1343 45707 1349
rect 45649 1309 45661 1343
rect 45695 1340 45707 1343
rect 45830 1340 45836 1352
rect 45695 1312 45836 1340
rect 45695 1309 45707 1312
rect 45649 1303 45707 1309
rect 45830 1300 45836 1312
rect 45888 1300 45894 1352
rect 45925 1343 45983 1349
rect 45925 1309 45937 1343
rect 45971 1340 45983 1343
rect 46106 1340 46112 1352
rect 45971 1312 46112 1340
rect 45971 1309 45983 1312
rect 45925 1303 45983 1309
rect 46106 1300 46112 1312
rect 46164 1300 46170 1352
rect 46293 1343 46351 1349
rect 46293 1309 46305 1343
rect 46339 1340 46351 1343
rect 46382 1340 46388 1352
rect 46339 1312 46388 1340
rect 46339 1309 46351 1312
rect 46293 1303 46351 1309
rect 46382 1300 46388 1312
rect 46440 1300 46446 1352
rect 46658 1300 46664 1352
rect 46716 1340 46722 1352
rect 46753 1343 46811 1349
rect 46753 1340 46765 1343
rect 46716 1312 46765 1340
rect 46716 1300 46722 1312
rect 46753 1309 46765 1312
rect 46799 1309 46811 1343
rect 46753 1303 46811 1309
rect 47121 1343 47179 1349
rect 47121 1309 47133 1343
rect 47167 1340 47179 1343
rect 47210 1340 47216 1352
rect 47167 1312 47216 1340
rect 47167 1309 47179 1312
rect 47121 1303 47179 1309
rect 47210 1300 47216 1312
rect 47268 1300 47274 1352
rect 47397 1343 47455 1349
rect 47397 1309 47409 1343
rect 47443 1340 47455 1343
rect 47486 1340 47492 1352
rect 47443 1312 47492 1340
rect 47443 1309 47455 1312
rect 47397 1303 47455 1309
rect 47486 1300 47492 1312
rect 47544 1300 47550 1352
rect 47673 1343 47731 1349
rect 47673 1309 47685 1343
rect 47719 1340 47731 1343
rect 47762 1340 47768 1352
rect 47719 1312 47768 1340
rect 47719 1309 47731 1312
rect 47673 1303 47731 1309
rect 47762 1300 47768 1312
rect 47820 1300 47826 1352
rect 47949 1343 48007 1349
rect 47949 1309 47961 1343
rect 47995 1340 48007 1343
rect 48038 1340 48044 1352
rect 47995 1312 48044 1340
rect 47995 1309 48007 1312
rect 47949 1303 48007 1309
rect 48038 1300 48044 1312
rect 48096 1300 48102 1352
rect 48225 1343 48283 1349
rect 48225 1309 48237 1343
rect 48271 1340 48283 1343
rect 48314 1340 48320 1352
rect 48271 1312 48320 1340
rect 48271 1309 48283 1312
rect 48225 1303 48283 1309
rect 48314 1300 48320 1312
rect 48372 1300 48378 1352
rect 48590 1340 48596 1352
rect 48551 1312 48596 1340
rect 48590 1300 48596 1312
rect 48648 1300 48654 1352
rect 48866 1340 48872 1352
rect 48827 1312 48872 1340
rect 48866 1300 48872 1312
rect 48924 1300 48930 1352
rect 49418 1340 49424 1352
rect 49379 1312 49424 1340
rect 49418 1300 49424 1312
rect 49476 1300 49482 1352
rect 49970 1340 49976 1352
rect 49931 1312 49976 1340
rect 49970 1300 49976 1312
rect 50028 1300 50034 1352
rect 50246 1340 50252 1352
rect 50207 1312 50252 1340
rect 50246 1300 50252 1312
rect 50304 1300 50310 1352
rect 50798 1300 50804 1352
rect 50856 1340 50862 1352
rect 50893 1343 50951 1349
rect 50893 1340 50905 1343
rect 50856 1312 50905 1340
rect 50856 1300 50862 1312
rect 50893 1309 50905 1312
rect 50939 1309 50951 1343
rect 50893 1303 50951 1309
rect 51169 1343 51227 1349
rect 51169 1309 51181 1343
rect 51215 1340 51227 1343
rect 51258 1340 51264 1352
rect 51215 1312 51264 1340
rect 51215 1309 51227 1312
rect 51169 1303 51227 1309
rect 51258 1300 51264 1312
rect 51316 1300 51322 1352
rect 51350 1300 51356 1352
rect 51408 1340 51414 1352
rect 51445 1343 51503 1349
rect 51445 1340 51457 1343
rect 51408 1312 51457 1340
rect 51408 1300 51414 1312
rect 51445 1309 51457 1312
rect 51491 1309 51503 1343
rect 51445 1303 51503 1309
rect 51626 1300 51632 1352
rect 51684 1340 51690 1352
rect 51721 1343 51779 1349
rect 51721 1340 51733 1343
rect 51684 1312 51733 1340
rect 51684 1300 51690 1312
rect 51721 1309 51733 1312
rect 51767 1309 51779 1343
rect 51721 1303 51779 1309
rect 52178 1300 52184 1352
rect 52236 1340 52242 1352
rect 52273 1343 52331 1349
rect 52273 1340 52285 1343
rect 52236 1312 52285 1340
rect 52236 1300 52242 1312
rect 52273 1309 52285 1312
rect 52319 1309 52331 1343
rect 52273 1303 52331 1309
rect 52730 1300 52736 1352
rect 52788 1340 52794 1352
rect 52825 1343 52883 1349
rect 52825 1340 52837 1343
rect 52788 1312 52837 1340
rect 52788 1300 52794 1312
rect 52825 1309 52837 1312
rect 52871 1309 52883 1343
rect 52825 1303 52883 1309
rect 53006 1300 53012 1352
rect 53064 1340 53070 1352
rect 53282 1340 53288 1352
rect 53064 1312 53109 1340
rect 53243 1312 53288 1340
rect 53064 1300 53070 1312
rect 53282 1300 53288 1312
rect 53340 1300 53346 1352
rect 53558 1340 53564 1352
rect 53519 1312 53564 1340
rect 53558 1300 53564 1312
rect 53616 1300 53622 1352
rect 53834 1340 53840 1352
rect 53795 1312 53840 1340
rect 53834 1300 53840 1312
rect 53892 1300 53898 1352
rect 54110 1340 54116 1352
rect 54071 1312 54116 1340
rect 54110 1300 54116 1312
rect 54168 1300 54174 1352
rect 54662 1340 54668 1352
rect 54623 1312 54668 1340
rect 54662 1300 54668 1312
rect 54720 1300 54726 1352
rect 54938 1340 54944 1352
rect 54899 1312 54944 1340
rect 54938 1300 54944 1312
rect 54996 1300 55002 1352
rect 55214 1340 55220 1352
rect 55175 1312 55220 1340
rect 55214 1300 55220 1312
rect 55272 1300 55278 1352
rect 55490 1300 55496 1352
rect 55548 1340 55554 1352
rect 55585 1343 55643 1349
rect 55585 1340 55597 1343
rect 55548 1312 55597 1340
rect 55548 1300 55554 1312
rect 55585 1309 55597 1312
rect 55631 1309 55643 1343
rect 55585 1303 55643 1309
rect 55766 1300 55772 1352
rect 55824 1340 55830 1352
rect 55861 1343 55919 1349
rect 55861 1340 55873 1343
rect 55824 1312 55873 1340
rect 55824 1300 55830 1312
rect 55861 1309 55873 1312
rect 55907 1309 55919 1343
rect 55861 1303 55919 1309
rect 56042 1300 56048 1352
rect 56100 1340 56106 1352
rect 56137 1343 56195 1349
rect 56137 1340 56149 1343
rect 56100 1312 56149 1340
rect 56100 1300 56106 1312
rect 56137 1309 56149 1312
rect 56183 1309 56195 1343
rect 56137 1303 56195 1309
rect 56318 1300 56324 1352
rect 56376 1340 56382 1352
rect 56413 1343 56471 1349
rect 56413 1340 56425 1343
rect 56376 1312 56425 1340
rect 56376 1300 56382 1312
rect 56413 1309 56425 1312
rect 56459 1309 56471 1343
rect 56413 1303 56471 1309
rect 56594 1300 56600 1352
rect 56652 1340 56658 1352
rect 56689 1343 56747 1349
rect 56689 1340 56701 1343
rect 56652 1312 56701 1340
rect 56652 1300 56658 1312
rect 56689 1309 56701 1312
rect 56735 1309 56747 1343
rect 56689 1303 56747 1309
rect 56870 1300 56876 1352
rect 56928 1340 56934 1352
rect 57241 1343 57299 1349
rect 57241 1340 57253 1343
rect 56928 1312 57253 1340
rect 56928 1300 56934 1312
rect 57241 1309 57253 1312
rect 57287 1309 57299 1343
rect 57241 1303 57299 1309
rect 57330 1300 57336 1352
rect 57388 1340 57394 1352
rect 57517 1343 57575 1349
rect 57517 1340 57529 1343
rect 57388 1312 57529 1340
rect 57388 1300 57394 1312
rect 57517 1309 57529 1312
rect 57563 1309 57575 1343
rect 57517 1303 57575 1309
rect 57698 1300 57704 1352
rect 57756 1340 57762 1352
rect 57793 1343 57851 1349
rect 57793 1340 57805 1343
rect 57756 1312 57805 1340
rect 57756 1300 57762 1312
rect 57793 1309 57805 1312
rect 57839 1309 57851 1343
rect 57793 1303 57851 1309
rect 57974 1300 57980 1352
rect 58032 1340 58038 1352
rect 58069 1343 58127 1349
rect 58069 1340 58081 1343
rect 58032 1312 58081 1340
rect 58032 1300 58038 1312
rect 58069 1309 58081 1312
rect 58115 1309 58127 1343
rect 58069 1303 58127 1309
rect 58250 1300 58256 1352
rect 58308 1340 58314 1352
rect 58437 1343 58495 1349
rect 58437 1340 58449 1343
rect 58308 1312 58449 1340
rect 58308 1300 58314 1312
rect 58437 1309 58449 1312
rect 58483 1309 58495 1343
rect 58437 1303 58495 1309
rect 58526 1300 58532 1352
rect 58584 1340 58590 1352
rect 58713 1343 58771 1349
rect 58713 1340 58725 1343
rect 58584 1312 58725 1340
rect 58584 1300 58590 1312
rect 58713 1309 58725 1312
rect 58759 1309 58771 1343
rect 58713 1303 58771 1309
rect 58802 1300 58808 1352
rect 58860 1340 58866 1352
rect 58989 1343 59047 1349
rect 58989 1340 59001 1343
rect 58860 1312 59001 1340
rect 58860 1300 58866 1312
rect 58989 1309 59001 1312
rect 59035 1309 59047 1343
rect 58989 1303 59047 1309
rect 59078 1300 59084 1352
rect 59136 1340 59142 1352
rect 59265 1343 59323 1349
rect 59265 1340 59277 1343
rect 59136 1312 59277 1340
rect 59136 1300 59142 1312
rect 59265 1309 59277 1312
rect 59311 1309 59323 1343
rect 59265 1303 59323 1309
rect 59354 1300 59360 1352
rect 59412 1340 59418 1352
rect 59541 1343 59599 1349
rect 59541 1340 59553 1343
rect 59412 1312 59553 1340
rect 59412 1300 59418 1312
rect 59541 1309 59553 1312
rect 59587 1309 59599 1343
rect 59541 1303 59599 1309
rect 59630 1300 59636 1352
rect 59688 1340 59694 1352
rect 59909 1343 59967 1349
rect 59909 1340 59921 1343
rect 59688 1312 59921 1340
rect 59688 1300 59694 1312
rect 59909 1309 59921 1312
rect 59955 1309 59967 1343
rect 59909 1303 59967 1309
rect 60274 1300 60280 1352
rect 60332 1340 60338 1352
rect 60461 1343 60519 1349
rect 60461 1340 60473 1343
rect 60332 1312 60473 1340
rect 60332 1300 60338 1312
rect 60461 1309 60473 1312
rect 60507 1309 60519 1343
rect 60461 1303 60519 1309
rect 60550 1300 60556 1352
rect 60608 1340 60614 1352
rect 60737 1343 60795 1349
rect 60737 1340 60749 1343
rect 60608 1312 60749 1340
rect 60608 1300 60614 1312
rect 60737 1309 60749 1312
rect 60783 1309 60795 1343
rect 60737 1303 60795 1309
rect 61010 1300 61016 1352
rect 61068 1340 61074 1352
rect 61289 1343 61347 1349
rect 61289 1340 61301 1343
rect 61068 1312 61301 1340
rect 61068 1300 61074 1312
rect 61289 1309 61301 1312
rect 61335 1309 61347 1343
rect 61289 1303 61347 1309
rect 61562 1300 61568 1352
rect 61620 1340 61626 1352
rect 61841 1343 61899 1349
rect 61841 1340 61853 1343
rect 61620 1312 61853 1340
rect 61620 1300 61626 1312
rect 61841 1309 61853 1312
rect 61887 1309 61899 1343
rect 61841 1303 61899 1309
rect 62114 1300 62120 1352
rect 62172 1340 62178 1352
rect 62577 1343 62635 1349
rect 62577 1340 62589 1343
rect 62172 1312 62589 1340
rect 62172 1300 62178 1312
rect 62577 1309 62589 1312
rect 62623 1309 62635 1343
rect 62577 1303 62635 1309
rect 62666 1300 62672 1352
rect 62724 1340 62730 1352
rect 63129 1343 63187 1349
rect 63129 1340 63141 1343
rect 62724 1312 63141 1340
rect 62724 1300 62730 1312
rect 63129 1309 63141 1312
rect 63175 1309 63187 1343
rect 63129 1303 63187 1309
rect 63218 1300 63224 1352
rect 63276 1340 63282 1352
rect 63681 1343 63739 1349
rect 63276 1300 63310 1340
rect 63681 1309 63693 1343
rect 63727 1309 63739 1343
rect 63681 1303 63739 1309
rect 31812 1244 32628 1272
rect 63282 1272 63310 1300
rect 63696 1272 63724 1303
rect 63770 1300 63776 1352
rect 63828 1340 63834 1352
rect 64141 1343 64199 1349
rect 64141 1340 64153 1343
rect 63828 1312 64153 1340
rect 63828 1300 63834 1312
rect 64141 1309 64153 1312
rect 64187 1309 64199 1343
rect 64141 1303 64199 1309
rect 64322 1300 64328 1352
rect 64380 1340 64386 1352
rect 64693 1343 64751 1349
rect 64693 1340 64705 1343
rect 64380 1312 64705 1340
rect 64380 1300 64386 1312
rect 64693 1309 64705 1312
rect 64739 1309 64751 1343
rect 64693 1303 64751 1309
rect 65150 1300 65156 1352
rect 65208 1340 65214 1352
rect 65613 1343 65671 1349
rect 65613 1340 65625 1343
rect 65208 1312 65625 1340
rect 65208 1300 65214 1312
rect 65613 1309 65625 1312
rect 65659 1309 65671 1343
rect 65613 1303 65671 1309
rect 65889 1343 65947 1349
rect 65889 1309 65901 1343
rect 65935 1309 65947 1343
rect 65889 1303 65947 1309
rect 63282 1244 63724 1272
rect 31812 1232 31818 1244
rect 64874 1232 64880 1284
rect 64932 1272 64938 1284
rect 65904 1272 65932 1303
rect 65978 1300 65984 1352
rect 66036 1340 66042 1352
rect 66717 1343 66775 1349
rect 66717 1340 66729 1343
rect 66036 1312 66729 1340
rect 66036 1300 66042 1312
rect 66717 1309 66729 1312
rect 66763 1309 66775 1343
rect 66717 1303 66775 1309
rect 66806 1300 66812 1352
rect 66864 1340 66870 1352
rect 67545 1343 67603 1349
rect 67545 1340 67557 1343
rect 66864 1312 67557 1340
rect 66864 1300 66870 1312
rect 67545 1309 67557 1312
rect 67591 1309 67603 1343
rect 67545 1303 67603 1309
rect 67913 1343 67971 1349
rect 67913 1309 67925 1343
rect 67959 1309 67971 1343
rect 67913 1303 67971 1309
rect 64932 1244 65932 1272
rect 64932 1232 64938 1244
rect 67082 1232 67088 1284
rect 67140 1272 67146 1284
rect 67928 1272 67956 1303
rect 68278 1300 68284 1352
rect 68336 1340 68342 1352
rect 68741 1343 68799 1349
rect 68741 1340 68753 1343
rect 68336 1312 68753 1340
rect 68336 1300 68342 1312
rect 68741 1309 68753 1312
rect 68787 1309 68799 1343
rect 68741 1303 68799 1309
rect 69017 1343 69075 1349
rect 69017 1309 69029 1343
rect 69063 1309 69075 1343
rect 69017 1303 69075 1309
rect 67140 1244 67956 1272
rect 67140 1232 67146 1244
rect 68462 1232 68468 1284
rect 68520 1272 68526 1284
rect 69032 1272 69060 1303
rect 69382 1300 69388 1352
rect 69440 1340 69446 1352
rect 69753 1343 69811 1349
rect 69753 1340 69765 1343
rect 69440 1312 69765 1340
rect 69440 1300 69446 1312
rect 69753 1309 69765 1312
rect 69799 1309 69811 1343
rect 69753 1303 69811 1309
rect 68520 1244 69060 1272
rect 68520 1232 68526 1244
rect 29052 1176 30144 1204
rect 29052 1164 29058 1176
rect 1104 1114 72864 1136
rect 1104 1062 3078 1114
rect 3130 1062 15078 1114
rect 15130 1062 27078 1114
rect 27130 1062 39078 1114
rect 39130 1062 51078 1114
rect 51130 1062 63078 1114
rect 63130 1062 72864 1114
rect 1104 1040 72864 1062
<< via1 >>
rect 3056 3952 3108 4004
rect 3792 3952 3844 4004
rect 9128 3952 9180 4004
rect 10048 3952 10100 4004
rect 20996 3952 21048 4004
rect 22744 3952 22796 4004
rect 27068 3952 27120 4004
rect 29092 3952 29144 4004
rect 45008 3952 45060 4004
rect 45652 3952 45704 4004
rect 51080 3952 51132 4004
rect 52000 3952 52052 4004
rect 57152 3952 57204 4004
rect 57336 3952 57388 4004
rect 2780 3884 2832 3936
rect 3516 3884 3568 3936
rect 9078 3782 9130 3834
rect 21078 3782 21130 3834
rect 33078 3782 33130 3834
rect 45078 3782 45130 3834
rect 57078 3782 57130 3834
rect 69078 3782 69130 3834
rect 1124 3680 1176 3732
rect 62948 3680 63000 3732
rect 64696 3680 64748 3732
rect 1400 3612 1452 3664
rect 28448 3612 28500 3664
rect 30472 3612 30524 3664
rect 1676 3544 1728 3596
rect 25412 3544 25464 3596
rect 27436 3544 27488 3596
rect 28172 3544 28224 3596
rect 30196 3544 30248 3596
rect 65708 3544 65760 3596
rect 67456 3544 67508 3596
rect 1952 3476 2004 3528
rect 24584 3476 24636 3528
rect 26332 3476 26384 3528
rect 27896 3476 27948 3528
rect 29920 3476 29972 3528
rect 64604 3476 64656 3528
rect 66352 3476 66404 3528
rect 14924 3408 14976 3460
rect 16120 3408 16172 3460
rect 17684 3408 17736 3460
rect 19156 3408 19208 3460
rect 21548 3408 21600 3460
rect 23296 3408 23348 3460
rect 23480 3408 23532 3460
rect 25228 3408 25280 3460
rect 29000 3408 29052 3460
rect 31024 3408 31076 3460
rect 56324 3408 56376 3460
rect 57336 3408 57388 3460
rect 59912 3408 59964 3460
rect 61384 3408 61436 3460
rect 61568 3408 61620 3460
rect 62948 3408 63000 3460
rect 65984 3408 66036 3460
rect 67732 3408 67784 3460
rect 14648 3340 14700 3392
rect 15844 3340 15896 3392
rect 17960 3340 18012 3392
rect 19432 3340 19484 3392
rect 20168 3340 20220 3392
rect 21640 3340 21692 3392
rect 21824 3340 21876 3392
rect 23572 3340 23624 3392
rect 24308 3340 24360 3392
rect 26056 3340 26108 3392
rect 26240 3340 26292 3392
rect 28264 3340 28316 3392
rect 28724 3340 28776 3392
rect 30748 3340 30800 3392
rect 61292 3340 61344 3392
rect 62764 3340 62816 3392
rect 65432 3340 65484 3392
rect 67180 3340 67232 3392
rect 3078 3238 3130 3290
rect 15078 3238 15130 3290
rect 27078 3238 27130 3290
rect 39078 3238 39130 3290
rect 51078 3238 51130 3290
rect 63078 3238 63130 3290
rect 11888 3136 11940 3188
rect 13084 3136 13136 3188
rect 14372 3136 14424 3188
rect 4160 3068 4212 3120
rect 2228 3043 2280 3052
rect 2228 3009 2237 3043
rect 2237 3009 2271 3043
rect 2271 3009 2280 3043
rect 2228 3000 2280 3009
rect 2504 3043 2556 3052
rect 2504 3009 2513 3043
rect 2513 3009 2547 3043
rect 2547 3009 2556 3043
rect 2504 3000 2556 3009
rect 2780 3043 2832 3052
rect 2780 3009 2789 3043
rect 2789 3009 2823 3043
rect 2823 3009 2832 3043
rect 2780 3000 2832 3009
rect 3608 3000 3660 3052
rect 5264 3068 5316 3120
rect 5080 3000 5132 3052
rect 6368 3068 6420 3120
rect 6184 3000 6236 3052
rect 8300 3068 8352 3120
rect 7472 3000 7524 3052
rect 9404 3068 9456 3120
rect 10048 3043 10100 3052
rect 10048 3009 10057 3043
rect 10057 3009 10091 3043
rect 10091 3009 10100 3043
rect 10048 3000 10100 3009
rect 11336 3068 11388 3120
rect 10508 3000 10560 3052
rect 12716 3068 12768 3120
rect 13176 3068 13228 3120
rect 13268 3068 13320 3120
rect 12992 3000 13044 3052
rect 16856 3136 16908 3188
rect 16304 3068 16356 3120
rect 15752 3000 15804 3052
rect 19340 3136 19392 3188
rect 18512 3068 18564 3120
rect 19156 3043 19208 3052
rect 19156 3009 19165 3043
rect 19165 3009 19199 3043
rect 19199 3009 19208 3043
rect 19156 3000 19208 3009
rect 19432 3043 19484 3052
rect 19432 3009 19441 3043
rect 19441 3009 19475 3043
rect 19475 3009 19484 3043
rect 19432 3000 19484 3009
rect 20444 3136 20496 3188
rect 20168 3068 20220 3120
rect 21640 3043 21692 3052
rect 21640 3009 21649 3043
rect 21649 3009 21683 3043
rect 21683 3009 21692 3043
rect 21640 3000 21692 3009
rect 22928 3136 22980 3188
rect 22284 3068 22336 3120
rect 22376 3000 22428 3052
rect 23296 3043 23348 3052
rect 2412 2932 2464 2984
rect 3332 2932 3384 2984
rect 3884 2932 3936 2984
rect 5540 2932 5592 2984
rect 6644 2932 6696 2984
rect 7748 2932 7800 2984
rect 8852 2932 8904 2984
rect 9956 2932 10008 2984
rect 11060 2932 11112 2984
rect 12440 2932 12492 2984
rect 13820 2932 13872 2984
rect 15476 2932 15528 2984
rect 17132 2932 17184 2984
rect 18788 2932 18840 2984
rect 21272 2932 21324 2984
rect 22744 2975 22796 2984
rect 22744 2941 22753 2975
rect 22753 2941 22787 2975
rect 22787 2941 22796 2975
rect 22744 2932 22796 2941
rect 23296 3009 23305 3043
rect 23305 3009 23339 3043
rect 23339 3009 23348 3043
rect 23296 3000 23348 3009
rect 23572 3043 23624 3052
rect 23572 3009 23581 3043
rect 23581 3009 23615 3043
rect 23615 3009 23624 3043
rect 23572 3000 23624 3009
rect 23940 3000 23992 3052
rect 29276 3136 29328 3188
rect 31300 3136 31352 3188
rect 54392 3136 54444 3188
rect 24860 3068 24912 3120
rect 24216 2932 24268 2984
rect 25228 3043 25280 3052
rect 25228 3009 25237 3043
rect 25237 3009 25271 3043
rect 25271 3009 25280 3043
rect 25228 3000 25280 3009
rect 26056 3043 26108 3052
rect 26056 3009 26065 3043
rect 26065 3009 26099 3043
rect 26099 3009 26108 3043
rect 26056 3000 26108 3009
rect 26332 3043 26384 3052
rect 26332 3009 26341 3043
rect 26341 3009 26375 3043
rect 26375 3009 26384 3043
rect 26332 3000 26384 3009
rect 26792 3068 26844 3120
rect 26884 3043 26936 3052
rect 26884 3009 26893 3043
rect 26893 3009 26927 3043
rect 26927 3009 26936 3043
rect 26884 3000 26936 3009
rect 27436 3043 27488 3052
rect 27436 3009 27445 3043
rect 27445 3009 27479 3043
rect 27479 3009 27488 3043
rect 27436 3000 27488 3009
rect 27528 3000 27580 3052
rect 28264 3043 28316 3052
rect 572 2864 624 2916
rect 4436 2864 4488 2916
rect 5816 2864 5868 2916
rect 6920 2864 6972 2916
rect 7656 2864 7708 2916
rect 848 2796 900 2848
rect 3516 2796 3568 2848
rect 3792 2796 3844 2848
rect 4712 2796 4764 2848
rect 7196 2796 7248 2848
rect 8576 2864 8628 2916
rect 9680 2864 9732 2916
rect 10784 2864 10836 2916
rect 12164 2864 12216 2916
rect 13544 2864 13596 2916
rect 15200 2864 15252 2916
rect 16580 2864 16632 2916
rect 7840 2839 7892 2848
rect 7840 2805 7849 2839
rect 7849 2805 7883 2839
rect 7883 2805 7892 2839
rect 7840 2796 7892 2805
rect 8024 2796 8076 2848
rect 10232 2796 10284 2848
rect 11612 2796 11664 2848
rect 13084 2839 13136 2848
rect 13084 2805 13093 2839
rect 13093 2805 13127 2839
rect 13127 2805 13136 2839
rect 13084 2796 13136 2805
rect 13176 2796 13228 2848
rect 14096 2796 14148 2848
rect 15844 2839 15896 2848
rect 15844 2805 15853 2839
rect 15853 2805 15887 2839
rect 15887 2805 15896 2839
rect 15844 2796 15896 2805
rect 16120 2839 16172 2848
rect 16120 2805 16129 2839
rect 16129 2805 16163 2839
rect 16163 2805 16172 2839
rect 16120 2796 16172 2805
rect 17500 2839 17552 2848
rect 17500 2805 17509 2839
rect 17509 2805 17543 2839
rect 17543 2805 17552 2839
rect 17500 2796 17552 2805
rect 17592 2796 17644 2848
rect 19064 2864 19116 2916
rect 20720 2864 20772 2916
rect 22652 2864 22704 2916
rect 25964 2932 26016 2984
rect 28264 3009 28273 3043
rect 28273 3009 28307 3043
rect 28307 3009 28316 3043
rect 28264 3000 28316 3009
rect 29828 3068 29880 3120
rect 29092 3043 29144 3052
rect 29092 3009 29101 3043
rect 29101 3009 29135 3043
rect 29135 3009 29144 3043
rect 29092 3000 29144 3009
rect 29920 3043 29972 3052
rect 29920 3009 29929 3043
rect 29929 3009 29963 3043
rect 29963 3009 29972 3043
rect 29920 3000 29972 3009
rect 30196 3043 30248 3052
rect 30196 3009 30205 3043
rect 30205 3009 30239 3043
rect 30239 3009 30248 3043
rect 30196 3000 30248 3009
rect 30380 3000 30432 3052
rect 48320 3068 48372 3120
rect 36176 3000 36228 3052
rect 36452 3000 36504 3052
rect 37004 3000 37056 3052
rect 37280 3000 37332 3052
rect 37556 3000 37608 3052
rect 38108 3000 38160 3052
rect 38660 3000 38712 3052
rect 39212 3000 39264 3052
rect 39764 3000 39816 3052
rect 40316 3000 40368 3052
rect 40868 3000 40920 3052
rect 41420 3000 41472 3052
rect 41972 3000 42024 3052
rect 42524 3000 42576 3052
rect 43352 3000 43404 3052
rect 44180 3000 44232 3052
rect 45652 3043 45704 3052
rect 45652 3009 45661 3043
rect 45661 3009 45695 3043
rect 45695 3009 45704 3043
rect 45652 3000 45704 3009
rect 45836 3000 45888 3052
rect 46664 3000 46716 3052
rect 48044 3000 48096 3052
rect 50252 3068 50304 3120
rect 49424 3000 49476 3052
rect 51632 3068 51684 3120
rect 52000 3043 52052 3052
rect 52000 3009 52009 3043
rect 52009 3009 52043 3043
rect 52043 3009 52052 3043
rect 52000 3000 52052 3009
rect 53288 3068 53340 3120
rect 52736 3000 52788 3052
rect 54116 3000 54168 3052
rect 30104 2932 30156 2984
rect 37832 2932 37884 2984
rect 38384 2932 38436 2984
rect 38936 2932 38988 2984
rect 39488 2932 39540 2984
rect 40040 2932 40092 2984
rect 40592 2932 40644 2984
rect 41144 2932 41196 2984
rect 41696 2932 41748 2984
rect 42248 2932 42300 2984
rect 42800 2932 42852 2984
rect 43628 2932 43680 2984
rect 44456 2932 44508 2984
rect 45284 2932 45336 2984
rect 46112 2932 46164 2984
rect 46940 2932 46992 2984
rect 47768 2932 47820 2984
rect 27712 2907 27764 2916
rect 27712 2873 27721 2907
rect 27721 2873 27755 2907
rect 27755 2873 27764 2907
rect 27712 2864 27764 2873
rect 27804 2864 27856 2916
rect 18236 2796 18288 2848
rect 19800 2796 19852 2848
rect 23204 2796 23256 2848
rect 25688 2796 25740 2848
rect 27620 2796 27672 2848
rect 28540 2839 28592 2848
rect 28540 2805 28549 2839
rect 28549 2805 28583 2839
rect 28583 2805 28592 2839
rect 28540 2796 28592 2805
rect 29552 2864 29604 2916
rect 36728 2864 36780 2916
rect 43076 2864 43128 2916
rect 43904 2864 43956 2916
rect 44732 2864 44784 2916
rect 45560 2864 45612 2916
rect 46388 2864 46440 2916
rect 47216 2864 47268 2916
rect 48596 2932 48648 2984
rect 49700 2932 49752 2984
rect 50804 2932 50856 2984
rect 51908 2932 51960 2984
rect 53012 2932 53064 2984
rect 54668 3000 54720 3052
rect 56876 3136 56928 3188
rect 55772 3068 55824 3120
rect 55680 3000 55732 3052
rect 58808 3136 58860 3188
rect 58256 3068 58308 3120
rect 58164 3000 58216 3052
rect 59820 3000 59872 3052
rect 61016 3136 61068 3188
rect 60372 3068 60424 3120
rect 56048 2932 56100 2984
rect 48872 2864 48924 2916
rect 49976 2864 50028 2916
rect 51356 2864 51408 2916
rect 52460 2864 52512 2916
rect 53840 2864 53892 2916
rect 55220 2864 55272 2916
rect 30472 2839 30524 2848
rect 30472 2805 30481 2839
rect 30481 2805 30515 2839
rect 30515 2805 30524 2839
rect 30472 2796 30524 2805
rect 30748 2839 30800 2848
rect 30748 2805 30757 2839
rect 30757 2805 30791 2839
rect 30791 2805 30800 2839
rect 30748 2796 30800 2805
rect 31024 2839 31076 2848
rect 31024 2805 31033 2839
rect 31033 2805 31067 2839
rect 31067 2805 31076 2839
rect 31024 2796 31076 2805
rect 31300 2839 31352 2848
rect 31300 2805 31309 2839
rect 31309 2805 31343 2839
rect 31343 2805 31352 2839
rect 31300 2796 31352 2805
rect 47492 2796 47544 2848
rect 49148 2796 49200 2848
rect 50528 2796 50580 2848
rect 52184 2796 52236 2848
rect 53564 2796 53616 2848
rect 54944 2796 54996 2848
rect 57244 2932 57296 2984
rect 58532 2932 58584 2984
rect 60464 3000 60516 3052
rect 61384 3043 61436 3052
rect 61384 3009 61393 3043
rect 61393 3009 61427 3043
rect 61427 3009 61436 3043
rect 61384 3000 61436 3009
rect 64052 3136 64104 3188
rect 63316 3068 63368 3120
rect 62764 3043 62816 3052
rect 62764 3009 62773 3043
rect 62773 3009 62807 3043
rect 62807 3009 62816 3043
rect 62764 3000 62816 3009
rect 62948 3000 63000 3052
rect 63776 3000 63828 3052
rect 64696 3043 64748 3052
rect 62396 2932 62448 2984
rect 64696 3009 64705 3043
rect 64705 3009 64739 3043
rect 64739 3009 64748 3043
rect 64696 3000 64748 3009
rect 65064 3000 65116 3052
rect 66260 3136 66312 3188
rect 68008 3136 68060 3188
rect 66812 3068 66864 3120
rect 66352 3043 66404 3052
rect 66352 3009 66361 3043
rect 66361 3009 66395 3043
rect 66395 3009 66404 3043
rect 66352 3000 66404 3009
rect 67180 3043 67232 3052
rect 67180 3009 67189 3043
rect 67189 3009 67223 3043
rect 67223 3009 67232 3043
rect 67180 3000 67232 3009
rect 67364 3000 67416 3052
rect 67088 2932 67140 2984
rect 56600 2864 56652 2916
rect 58072 2864 58124 2916
rect 57336 2796 57388 2848
rect 57612 2796 57664 2848
rect 59084 2864 59136 2916
rect 59360 2864 59412 2916
rect 61844 2864 61896 2916
rect 63500 2864 63552 2916
rect 65064 2864 65116 2916
rect 60740 2796 60792 2848
rect 62304 2796 62356 2848
rect 64420 2839 64472 2848
rect 64420 2805 64429 2839
rect 64429 2805 64463 2839
rect 64463 2805 64472 2839
rect 64420 2796 64472 2805
rect 64512 2796 64564 2848
rect 66536 2864 66588 2916
rect 67456 2907 67508 2916
rect 65248 2839 65300 2848
rect 65248 2805 65257 2839
rect 65257 2805 65291 2839
rect 65291 2805 65300 2839
rect 65248 2796 65300 2805
rect 65432 2796 65484 2848
rect 67456 2873 67465 2907
rect 67465 2873 67499 2907
rect 67499 2873 67508 2907
rect 67456 2864 67508 2873
rect 67732 2907 67784 2916
rect 67732 2873 67741 2907
rect 67741 2873 67775 2907
rect 67775 2873 67784 2907
rect 67732 2864 67784 2873
rect 68008 2907 68060 2916
rect 68008 2873 68017 2907
rect 68017 2873 68051 2907
rect 68051 2873 68060 2907
rect 68008 2864 68060 2873
rect 9078 2694 9130 2746
rect 21078 2694 21130 2746
rect 33078 2694 33130 2746
rect 45078 2694 45130 2746
rect 57078 2694 57130 2746
rect 69078 2694 69130 2746
rect 2964 2592 3016 2644
rect 16028 2524 16080 2576
rect 17500 2524 17552 2576
rect 62672 2524 62724 2576
rect 64420 2524 64472 2576
rect 2780 2499 2832 2508
rect 2780 2465 2789 2499
rect 2789 2465 2823 2499
rect 2823 2465 2832 2499
rect 2780 2456 2832 2465
rect 2504 2431 2556 2440
rect 2504 2397 2513 2431
rect 2513 2397 2547 2431
rect 2547 2397 2556 2431
rect 2504 2388 2556 2397
rect 3078 2150 3130 2202
rect 15078 2150 15130 2202
rect 27078 2150 27130 2202
rect 39078 2150 39130 2202
rect 51078 2150 51130 2202
rect 63078 2150 63130 2202
rect 1400 1844 1452 1896
rect 30104 1776 30156 1828
rect 2228 1751 2280 1760
rect 2228 1717 2237 1751
rect 2237 1717 2271 1751
rect 2271 1717 2280 1751
rect 2228 1708 2280 1717
rect 2320 1708 2372 1760
rect 2780 1708 2832 1760
rect 2964 1708 3016 1760
rect 3884 1708 3936 1760
rect 6644 1708 6696 1760
rect 8576 1708 8628 1760
rect 9404 1708 9456 1760
rect 11612 1708 11664 1760
rect 12992 1708 13044 1760
rect 14924 1708 14976 1760
rect 15752 1708 15804 1760
rect 19892 1708 19944 1760
rect 25964 1708 26016 1760
rect 29828 1708 29880 1760
rect 31484 1708 31536 1760
rect 38936 1708 38988 1760
rect 44180 1708 44232 1760
rect 46940 1708 46992 1760
rect 50528 1751 50580 1760
rect 50528 1717 50537 1751
rect 50537 1717 50571 1751
rect 50571 1717 50580 1751
rect 50528 1708 50580 1717
rect 52460 1708 52512 1760
rect 54392 1751 54444 1760
rect 54392 1717 54401 1751
rect 54401 1717 54435 1751
rect 54435 1717 54444 1751
rect 54392 1708 54444 1717
rect 57428 1708 57480 1760
rect 63500 1708 63552 1760
rect 67640 1708 67692 1760
rect 69204 1708 69256 1760
rect 9078 1606 9130 1658
rect 21078 1606 21130 1658
rect 33078 1606 33130 1658
rect 45078 1606 45130 1658
rect 57078 1606 57130 1658
rect 69078 1606 69130 1658
rect 1124 1504 1176 1556
rect 24032 1504 24084 1556
rect 25412 1504 25464 1556
rect 27436 1504 27488 1556
rect 29552 1504 29604 1556
rect 31208 1504 31260 1556
rect 2504 1436 2556 1488
rect 3332 1436 3384 1488
rect 4436 1436 4488 1488
rect 4988 1436 5040 1488
rect 7748 1436 7800 1488
rect 9312 1436 9364 1488
rect 9956 1436 10008 1488
rect 11888 1436 11940 1488
rect 12716 1436 12768 1488
rect 13544 1436 13596 1488
rect 14096 1436 14148 1488
rect 15200 1436 15252 1488
rect 16304 1436 16356 1488
rect 17132 1436 17184 1488
rect 17960 1436 18012 1488
rect 18788 1436 18840 1488
rect 20168 1436 20220 1488
rect 21272 1436 21324 1488
rect 22652 1436 22704 1488
rect 23480 1436 23532 1488
rect 24584 1436 24636 1488
rect 26516 1436 26568 1488
rect 27896 1436 27948 1488
rect 29276 1436 29328 1488
rect 30656 1436 30708 1488
rect 32036 1436 32088 1488
rect 38108 1436 38160 1488
rect 39488 1436 39540 1488
rect 40592 1436 40644 1488
rect 41696 1436 41748 1488
rect 42248 1436 42300 1488
rect 42800 1436 42852 1488
rect 43352 1436 43404 1488
rect 59912 1436 59964 1488
rect 60740 1436 60792 1488
rect 61292 1436 61344 1488
rect 61844 1436 61896 1488
rect 64604 1436 64656 1488
rect 65708 1436 65760 1488
rect 66536 1436 66588 1488
rect 67916 1436 67968 1488
rect 68744 1436 68796 1488
rect 69572 1436 69624 1488
rect 1676 1411 1728 1420
rect 1676 1377 1685 1411
rect 1685 1377 1719 1411
rect 1719 1377 1728 1411
rect 1676 1368 1728 1377
rect 1768 1368 1820 1420
rect 5264 1368 5316 1420
rect 5816 1368 5868 1420
rect 6368 1368 6420 1420
rect 7196 1368 7248 1420
rect 8024 1368 8076 1420
rect 10232 1368 10284 1420
rect 10784 1368 10836 1420
rect 12164 1368 12216 1420
rect 15476 1368 15528 1420
rect 17408 1368 17460 1420
rect 18236 1368 18288 1420
rect 19064 1368 19116 1420
rect 20720 1368 20772 1420
rect 21548 1368 21600 1420
rect 22376 1368 22428 1420
rect 23204 1368 23256 1420
rect 572 1300 624 1352
rect 848 1232 900 1284
rect 1952 1164 2004 1216
rect 3608 1300 3660 1352
rect 4252 1300 4304 1352
rect 4712 1300 4764 1352
rect 5540 1300 5592 1352
rect 6092 1300 6144 1352
rect 6920 1300 6972 1352
rect 7472 1300 7524 1352
rect 8300 1300 8352 1352
rect 8852 1300 8904 1352
rect 9680 1300 9732 1352
rect 10508 1300 10560 1352
rect 11060 1300 11112 1352
rect 11336 1232 11388 1284
rect 12440 1300 12492 1352
rect 13360 1300 13412 1352
rect 13820 1300 13872 1352
rect 14648 1300 14700 1352
rect 14372 1232 14424 1284
rect 16028 1300 16080 1352
rect 16856 1343 16908 1352
rect 16856 1309 16865 1343
rect 16865 1309 16899 1343
rect 16899 1309 16908 1343
rect 16856 1300 16908 1309
rect 16580 1232 16632 1284
rect 17684 1300 17736 1352
rect 18512 1300 18564 1352
rect 19340 1300 19392 1352
rect 19616 1232 19668 1284
rect 20444 1232 20496 1284
rect 21272 1300 21324 1352
rect 21824 1300 21876 1352
rect 22100 1232 22152 1284
rect 22928 1232 22980 1284
rect 24308 1300 24360 1352
rect 23756 1232 23808 1284
rect 24860 1300 24912 1352
rect 26240 1368 26292 1420
rect 27620 1368 27672 1420
rect 28724 1368 28776 1420
rect 30380 1368 30432 1420
rect 32312 1368 32364 1420
rect 39212 1368 39264 1420
rect 39764 1368 39816 1420
rect 40316 1368 40368 1420
rect 41144 1368 41196 1420
rect 49148 1368 49200 1420
rect 49700 1368 49752 1420
rect 51908 1368 51960 1420
rect 62396 1368 62448 1420
rect 62948 1368 63000 1420
rect 64052 1368 64104 1420
rect 65432 1368 65484 1420
rect 66260 1368 66312 1420
rect 67364 1368 67416 1420
rect 69848 1368 69900 1420
rect 25136 1232 25188 1284
rect 25688 1164 25740 1216
rect 26792 1300 26844 1352
rect 27252 1232 27304 1284
rect 28264 1300 28316 1352
rect 28448 1164 28500 1216
rect 29000 1164 29052 1216
rect 30932 1300 30984 1352
rect 31760 1232 31812 1284
rect 38292 1300 38344 1352
rect 38660 1300 38712 1352
rect 40040 1300 40092 1352
rect 40868 1300 40920 1352
rect 41328 1300 41380 1352
rect 41972 1300 42024 1352
rect 42524 1300 42576 1352
rect 43076 1300 43128 1352
rect 43628 1300 43680 1352
rect 43904 1300 43956 1352
rect 44456 1300 44508 1352
rect 44732 1300 44784 1352
rect 44916 1300 44968 1352
rect 45284 1300 45336 1352
rect 45560 1300 45612 1352
rect 45836 1300 45888 1352
rect 46112 1300 46164 1352
rect 46388 1300 46440 1352
rect 46664 1300 46716 1352
rect 47216 1300 47268 1352
rect 47492 1300 47544 1352
rect 47768 1300 47820 1352
rect 48044 1300 48096 1352
rect 48320 1300 48372 1352
rect 48596 1343 48648 1352
rect 48596 1309 48605 1343
rect 48605 1309 48639 1343
rect 48639 1309 48648 1343
rect 48596 1300 48648 1309
rect 48872 1343 48924 1352
rect 48872 1309 48881 1343
rect 48881 1309 48915 1343
rect 48915 1309 48924 1343
rect 48872 1300 48924 1309
rect 49424 1343 49476 1352
rect 49424 1309 49433 1343
rect 49433 1309 49467 1343
rect 49467 1309 49476 1343
rect 49424 1300 49476 1309
rect 49976 1343 50028 1352
rect 49976 1309 49985 1343
rect 49985 1309 50019 1343
rect 50019 1309 50028 1343
rect 49976 1300 50028 1309
rect 50252 1343 50304 1352
rect 50252 1309 50261 1343
rect 50261 1309 50295 1343
rect 50295 1309 50304 1343
rect 50252 1300 50304 1309
rect 50804 1300 50856 1352
rect 51264 1300 51316 1352
rect 51356 1300 51408 1352
rect 51632 1300 51684 1352
rect 52184 1300 52236 1352
rect 52736 1300 52788 1352
rect 53012 1343 53064 1352
rect 53012 1309 53021 1343
rect 53021 1309 53055 1343
rect 53055 1309 53064 1343
rect 53288 1343 53340 1352
rect 53012 1300 53064 1309
rect 53288 1309 53297 1343
rect 53297 1309 53331 1343
rect 53331 1309 53340 1343
rect 53288 1300 53340 1309
rect 53564 1343 53616 1352
rect 53564 1309 53573 1343
rect 53573 1309 53607 1343
rect 53607 1309 53616 1343
rect 53564 1300 53616 1309
rect 53840 1343 53892 1352
rect 53840 1309 53849 1343
rect 53849 1309 53883 1343
rect 53883 1309 53892 1343
rect 53840 1300 53892 1309
rect 54116 1343 54168 1352
rect 54116 1309 54125 1343
rect 54125 1309 54159 1343
rect 54159 1309 54168 1343
rect 54116 1300 54168 1309
rect 54668 1343 54720 1352
rect 54668 1309 54677 1343
rect 54677 1309 54711 1343
rect 54711 1309 54720 1343
rect 54668 1300 54720 1309
rect 54944 1343 54996 1352
rect 54944 1309 54953 1343
rect 54953 1309 54987 1343
rect 54987 1309 54996 1343
rect 54944 1300 54996 1309
rect 55220 1343 55272 1352
rect 55220 1309 55229 1343
rect 55229 1309 55263 1343
rect 55263 1309 55272 1343
rect 55220 1300 55272 1309
rect 55496 1300 55548 1352
rect 55772 1300 55824 1352
rect 56048 1300 56100 1352
rect 56324 1300 56376 1352
rect 56600 1300 56652 1352
rect 56876 1300 56928 1352
rect 57336 1300 57388 1352
rect 57704 1300 57756 1352
rect 57980 1300 58032 1352
rect 58256 1300 58308 1352
rect 58532 1300 58584 1352
rect 58808 1300 58860 1352
rect 59084 1300 59136 1352
rect 59360 1300 59412 1352
rect 59636 1300 59688 1352
rect 60280 1300 60332 1352
rect 60556 1300 60608 1352
rect 61016 1300 61068 1352
rect 61568 1300 61620 1352
rect 62120 1300 62172 1352
rect 62672 1300 62724 1352
rect 63224 1300 63276 1352
rect 63776 1300 63828 1352
rect 64328 1300 64380 1352
rect 65156 1300 65208 1352
rect 64880 1232 64932 1284
rect 65984 1300 66036 1352
rect 66812 1300 66864 1352
rect 67088 1232 67140 1284
rect 68284 1300 68336 1352
rect 68468 1232 68520 1284
rect 69388 1300 69440 1352
rect 3078 1062 3130 1114
rect 15078 1062 15130 1114
rect 27078 1062 27130 1114
rect 39078 1062 39130 1114
rect 51078 1062 51130 1114
rect 63078 1062 63130 1114
<< metal2 >>
rect 570 4000 626 5000
rect 846 4000 902 5000
rect 1122 4000 1178 5000
rect 1398 4000 1454 5000
rect 1674 4000 1730 5000
rect 1950 4000 2006 5000
rect 2226 4000 2282 5000
rect 2502 4000 2558 5000
rect 2778 4000 2834 5000
rect 3054 4004 3110 5000
rect 3054 4000 3056 4004
rect 584 2922 612 4000
rect 572 2916 624 2922
rect 572 2858 624 2864
rect 860 2854 888 4000
rect 1136 3738 1164 4000
rect 1124 3732 1176 3738
rect 1124 3674 1176 3680
rect 1412 3670 1440 4000
rect 1400 3664 1452 3670
rect 1400 3606 1452 3612
rect 1688 3602 1716 4000
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1964 3534 1992 4000
rect 1952 3528 2004 3534
rect 1952 3470 2004 3476
rect 2240 3058 2268 4000
rect 2516 3346 2544 4000
rect 2792 3942 2820 4000
rect 3108 4000 3110 4004
rect 3330 4000 3386 5000
rect 3606 4000 3662 5000
rect 3792 4004 3844 4010
rect 3056 3946 3108 3952
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2778 3768 2834 3777
rect 2778 3703 2834 3712
rect 2424 3318 2544 3346
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 2424 2990 2452 3318
rect 2502 3224 2558 3233
rect 2502 3159 2558 3168
rect 2516 3058 2544 3159
rect 2792 3058 2820 3703
rect 3054 3428 3154 3856
rect 3054 3372 3076 3428
rect 3132 3372 3154 3428
rect 3054 3290 3154 3372
rect 3054 3238 3078 3290
rect 3130 3238 3154 3290
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2412 2984 2464 2990
rect 2412 2926 2464 2932
rect 2962 2952 3018 2961
rect 2962 2887 3018 2896
rect 848 2848 900 2854
rect 848 2790 900 2796
rect 2976 2650 3004 2887
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 2778 2544 2834 2553
rect 2778 2479 2780 2488
rect 2832 2479 2834 2488
rect 2780 2450 2832 2456
rect 2504 2440 2556 2446
rect 2504 2382 2556 2388
rect 2516 2145 2544 2382
rect 3054 2202 3154 3238
rect 3344 2990 3372 4000
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 3528 2854 3556 3878
rect 3620 3058 3648 4000
rect 3882 4000 3938 5000
rect 4158 4000 4214 5000
rect 4434 4000 4490 5000
rect 4710 4000 4766 5000
rect 4986 4000 5042 5000
rect 5262 4000 5318 5000
rect 5538 4000 5594 5000
rect 5814 4000 5870 5000
rect 6090 4000 6146 5000
rect 6366 4000 6422 5000
rect 6642 4000 6698 5000
rect 6918 4000 6974 5000
rect 7194 4000 7250 5000
rect 7470 4000 7526 5000
rect 7746 4000 7802 5000
rect 8022 4000 8078 5000
rect 8298 4000 8354 5000
rect 8574 4000 8630 5000
rect 8850 4000 8906 5000
rect 9126 4004 9182 5000
rect 9126 4000 9128 4004
rect 3792 3946 3844 3952
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3804 2854 3832 3946
rect 3896 2990 3924 4000
rect 4172 3126 4200 4000
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 4448 2922 4476 4000
rect 4436 2916 4488 2922
rect 4436 2858 4488 2864
rect 4724 2854 4752 4000
rect 5000 3074 5028 4000
rect 5276 3126 5304 4000
rect 5264 3120 5316 3126
rect 5000 3058 5120 3074
rect 5264 3062 5316 3068
rect 5000 3052 5132 3058
rect 5000 3046 5080 3052
rect 5080 2994 5132 3000
rect 5552 2990 5580 4000
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 5828 2922 5856 4000
rect 6104 3074 6132 4000
rect 6380 3126 6408 4000
rect 6368 3120 6420 3126
rect 6104 3058 6224 3074
rect 6368 3062 6420 3068
rect 6104 3052 6236 3058
rect 6104 3046 6184 3052
rect 6184 2994 6236 3000
rect 6656 2990 6684 4000
rect 6644 2984 6696 2990
rect 6644 2926 6696 2932
rect 6932 2922 6960 4000
rect 5816 2916 5868 2922
rect 5816 2858 5868 2864
rect 6920 2916 6972 2922
rect 6920 2858 6972 2864
rect 7208 2854 7236 4000
rect 7484 3058 7512 4000
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7760 2990 7788 4000
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7656 2916 7708 2922
rect 7656 2858 7708 2864
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3792 2848 3844 2854
rect 3792 2790 3844 2796
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 7668 2802 7696 2858
rect 8036 2854 8064 4000
rect 8312 3126 8340 4000
rect 8300 3120 8352 3126
rect 8300 3062 8352 3068
rect 8588 2922 8616 4000
rect 8864 2990 8892 4000
rect 9180 4000 9182 4004
rect 9402 4000 9458 5000
rect 9678 4000 9734 5000
rect 9954 4000 10010 5000
rect 10048 4004 10100 4010
rect 9128 3946 9180 3952
rect 9054 3834 9154 3856
rect 9054 3782 9078 3834
rect 9130 3782 9154 3834
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8576 2916 8628 2922
rect 8576 2858 8628 2864
rect 7840 2848 7892 2854
rect 7668 2796 7840 2802
rect 7668 2790 7892 2796
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 7668 2774 7880 2790
rect 3054 2150 3078 2202
rect 3130 2150 3154 2202
rect 2502 2136 2558 2145
rect 2502 2071 2558 2080
rect 1400 1896 1452 1902
rect 1400 1838 1452 1844
rect 1124 1556 1176 1562
rect 1124 1498 1176 1504
rect 572 1352 624 1358
rect 572 1294 624 1300
rect 584 1000 612 1294
rect 848 1284 900 1290
rect 848 1226 900 1232
rect 860 1000 888 1226
rect 1136 1000 1164 1498
rect 1412 1000 1440 1838
rect 2228 1760 2280 1766
rect 2226 1728 2228 1737
rect 2320 1760 2372 1766
rect 2280 1728 2282 1737
rect 2320 1702 2372 1708
rect 2780 1760 2832 1766
rect 2780 1702 2832 1708
rect 2964 1760 3016 1766
rect 2964 1702 3016 1708
rect 2226 1663 2282 1672
rect 1674 1456 1730 1465
rect 1674 1391 1676 1400
rect 1728 1391 1730 1400
rect 1768 1420 1820 1426
rect 1676 1362 1728 1368
rect 1768 1362 1820 1368
rect 1780 1170 1808 1362
rect 1688 1142 1808 1170
rect 1952 1216 2004 1222
rect 2332 1170 2360 1702
rect 2504 1488 2556 1494
rect 2504 1430 2556 1436
rect 1952 1158 2004 1164
rect 1688 1000 1716 1142
rect 1964 1000 1992 1158
rect 2240 1142 2360 1170
rect 2240 1000 2268 1142
rect 2516 1000 2544 1430
rect 2792 1000 2820 1702
rect 570 0 626 1000
rect 846 0 902 1000
rect 1122 0 1178 1000
rect 1398 0 1454 1000
rect 1674 0 1730 1000
rect 1950 0 2006 1000
rect 2226 0 2282 1000
rect 2502 0 2558 1000
rect 2778 0 2834 1000
rect 2976 898 3004 1702
rect 3054 1268 3154 2150
rect 9054 2746 9154 3782
rect 9416 3126 9444 4000
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 9692 2922 9720 4000
rect 9968 2990 9996 4000
rect 10230 4000 10286 5000
rect 10506 4000 10562 5000
rect 10782 4000 10838 5000
rect 11058 4000 11114 5000
rect 11334 4000 11390 5000
rect 11610 4000 11666 5000
rect 11886 4000 11942 5000
rect 12162 4000 12218 5000
rect 12438 4000 12494 5000
rect 12714 4000 12770 5000
rect 12990 4000 13046 5000
rect 13266 4000 13322 5000
rect 13542 4000 13598 5000
rect 13818 4000 13874 5000
rect 14094 4000 14150 5000
rect 14370 4000 14426 5000
rect 14646 4000 14702 5000
rect 14922 4000 14978 5000
rect 15198 4000 15254 5000
rect 15474 4000 15530 5000
rect 15750 4000 15806 5000
rect 16026 4000 16082 5000
rect 16302 4000 16358 5000
rect 16578 4000 16634 5000
rect 16854 4000 16910 5000
rect 17130 4000 17186 5000
rect 17406 4000 17462 5000
rect 17682 4000 17738 5000
rect 17958 4000 18014 5000
rect 18234 4000 18290 5000
rect 18510 4000 18566 5000
rect 18786 4000 18842 5000
rect 19062 4000 19118 5000
rect 19338 4000 19394 5000
rect 19614 4000 19670 5000
rect 19890 4000 19946 5000
rect 20166 4000 20222 5000
rect 20442 4000 20498 5000
rect 20718 4000 20774 5000
rect 20994 4004 21050 5000
rect 20994 4000 20996 4004
rect 10048 3946 10100 3952
rect 10060 3058 10088 3946
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 10244 2854 10272 4000
rect 10520 3058 10548 4000
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10796 2922 10824 4000
rect 11072 2990 11100 4000
rect 11348 3126 11376 4000
rect 11336 3120 11388 3126
rect 11336 3062 11388 3068
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 10784 2916 10836 2922
rect 10784 2858 10836 2864
rect 11624 2854 11652 4000
rect 11900 3194 11928 4000
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 12176 2922 12204 4000
rect 12452 2990 12480 4000
rect 12728 3126 12756 4000
rect 12716 3120 12768 3126
rect 12716 3062 12768 3068
rect 13004 3058 13032 4000
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12164 2916 12216 2922
rect 12164 2858 12216 2864
rect 13096 2854 13124 3130
rect 13280 3126 13308 4000
rect 13176 3120 13228 3126
rect 13176 3062 13228 3068
rect 13268 3120 13320 3126
rect 13268 3062 13320 3068
rect 13188 2854 13216 3062
rect 13556 2922 13584 4000
rect 13832 2990 13860 4000
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13544 2916 13596 2922
rect 13544 2858 13596 2864
rect 14108 2854 14136 4000
rect 14384 3194 14412 4000
rect 14660 3398 14688 4000
rect 14936 3466 14964 4000
rect 14924 3460 14976 3466
rect 14924 3402 14976 3408
rect 15054 3428 15154 3856
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 15054 3372 15076 3428
rect 15132 3372 15154 3428
rect 15054 3290 15154 3372
rect 15054 3238 15078 3290
rect 15130 3238 15154 3290
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 13084 2848 13136 2854
rect 13084 2790 13136 2796
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 14096 2848 14148 2854
rect 14096 2790 14148 2796
rect 9054 2694 9078 2746
rect 9130 2694 9154 2746
rect 9054 2348 9154 2694
rect 9054 2292 9076 2348
rect 9132 2292 9154 2348
rect 3884 1760 3936 1766
rect 3884 1702 3936 1708
rect 6644 1760 6696 1766
rect 6644 1702 6696 1708
rect 8576 1760 8628 1766
rect 8576 1702 8628 1708
rect 3332 1488 3384 1494
rect 3332 1430 3384 1436
rect 3054 1212 3076 1268
rect 3132 1212 3154 1268
rect 3054 1114 3154 1212
rect 3054 1062 3078 1114
rect 3130 1062 3154 1114
rect 3054 1040 3154 1062
rect 3344 1000 3372 1430
rect 3608 1352 3660 1358
rect 3608 1294 3660 1300
rect 3620 1000 3648 1294
rect 3896 1000 3924 1702
rect 4436 1488 4488 1494
rect 4436 1430 4488 1436
rect 4988 1488 5040 1494
rect 4988 1430 5040 1436
rect 4252 1352 4304 1358
rect 4172 1312 4252 1340
rect 4172 1000 4200 1312
rect 4252 1294 4304 1300
rect 4448 1000 4476 1430
rect 4712 1352 4764 1358
rect 4712 1294 4764 1300
rect 4724 1000 4752 1294
rect 5000 1000 5028 1430
rect 5264 1420 5316 1426
rect 5264 1362 5316 1368
rect 5816 1420 5868 1426
rect 5816 1362 5868 1368
rect 6368 1420 6420 1426
rect 6368 1362 6420 1368
rect 5276 1000 5304 1362
rect 5540 1352 5592 1358
rect 5540 1294 5592 1300
rect 5552 1000 5580 1294
rect 5828 1000 5856 1362
rect 6092 1352 6144 1358
rect 6092 1294 6144 1300
rect 6104 1000 6132 1294
rect 6380 1000 6408 1362
rect 6656 1000 6684 1702
rect 7748 1488 7800 1494
rect 7748 1430 7800 1436
rect 7196 1420 7248 1426
rect 7196 1362 7248 1368
rect 6920 1352 6972 1358
rect 6920 1294 6972 1300
rect 6932 1000 6960 1294
rect 7208 1000 7236 1362
rect 7472 1352 7524 1358
rect 7472 1294 7524 1300
rect 7484 1000 7512 1294
rect 7760 1000 7788 1430
rect 8024 1420 8076 1426
rect 8024 1362 8076 1368
rect 8036 1000 8064 1362
rect 8300 1352 8352 1358
rect 8300 1294 8352 1300
rect 8312 1000 8340 1294
rect 8588 1000 8616 1702
rect 9054 1658 9154 2292
rect 15054 2202 15154 3238
rect 15212 2922 15240 4000
rect 15488 2990 15516 4000
rect 15764 3058 15792 4000
rect 15844 3392 15896 3398
rect 15844 3334 15896 3340
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 15200 2916 15252 2922
rect 15200 2858 15252 2864
rect 15856 2854 15884 3334
rect 15844 2848 15896 2854
rect 15844 2790 15896 2796
rect 16040 2582 16068 4000
rect 16120 3460 16172 3466
rect 16120 3402 16172 3408
rect 16132 2854 16160 3402
rect 16316 3126 16344 4000
rect 16304 3120 16356 3126
rect 16304 3062 16356 3068
rect 16592 2922 16620 4000
rect 16868 3194 16896 4000
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 17144 2990 17172 4000
rect 17420 3074 17448 4000
rect 17696 3466 17724 4000
rect 17684 3460 17736 3466
rect 17684 3402 17736 3408
rect 17972 3398 18000 4000
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 17420 3046 17632 3074
rect 17132 2984 17184 2990
rect 17132 2926 17184 2932
rect 16580 2916 16632 2922
rect 16580 2858 16632 2864
rect 17604 2854 17632 3046
rect 18248 2854 18276 4000
rect 18524 3126 18552 4000
rect 18512 3120 18564 3126
rect 18512 3062 18564 3068
rect 18800 2990 18828 4000
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 19076 2922 19104 4000
rect 19156 3460 19208 3466
rect 19156 3402 19208 3408
rect 19168 3058 19196 3402
rect 19352 3194 19380 4000
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19444 3058 19472 3334
rect 19156 3052 19208 3058
rect 19156 2994 19208 3000
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19064 2916 19116 2922
rect 19064 2858 19116 2864
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17592 2848 17644 2854
rect 17592 2790 17644 2796
rect 18236 2848 18288 2854
rect 19628 2836 19656 4000
rect 19904 3108 19932 4000
rect 20180 3398 20208 4000
rect 20168 3392 20220 3398
rect 20168 3334 20220 3340
rect 20456 3194 20484 4000
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 20168 3120 20220 3126
rect 19904 3080 20168 3108
rect 20168 3062 20220 3068
rect 20732 2922 20760 4000
rect 21048 4000 21050 4004
rect 21270 4000 21326 5000
rect 21546 4000 21602 5000
rect 21822 4000 21878 5000
rect 22098 4000 22154 5000
rect 22374 4000 22430 5000
rect 22650 4000 22706 5000
rect 22744 4004 22796 4010
rect 20996 3946 21048 3952
rect 21054 3834 21154 3856
rect 21054 3782 21078 3834
rect 21130 3782 21154 3834
rect 20720 2916 20772 2922
rect 20720 2858 20772 2864
rect 19800 2848 19852 2854
rect 19628 2808 19800 2836
rect 18236 2790 18288 2796
rect 19800 2790 19852 2796
rect 17512 2582 17540 2790
rect 21054 2746 21154 3782
rect 21284 2990 21312 4000
rect 21560 3466 21588 4000
rect 21548 3460 21600 3466
rect 21548 3402 21600 3408
rect 21836 3398 21864 4000
rect 21640 3392 21692 3398
rect 21640 3334 21692 3340
rect 21824 3392 21876 3398
rect 21824 3334 21876 3340
rect 21652 3058 21680 3334
rect 22112 3108 22140 4000
rect 22284 3120 22336 3126
rect 22112 3080 22284 3108
rect 22284 3062 22336 3068
rect 22388 3058 22416 4000
rect 21640 3052 21692 3058
rect 21640 2994 21692 3000
rect 22376 3052 22428 3058
rect 22376 2994 22428 3000
rect 21272 2984 21324 2990
rect 21272 2926 21324 2932
rect 22664 2922 22692 4000
rect 22926 4000 22982 5000
rect 23202 4000 23258 5000
rect 23478 4000 23534 5000
rect 23754 4000 23810 5000
rect 24030 4000 24086 5000
rect 24306 4000 24362 5000
rect 24582 4000 24638 5000
rect 24858 4000 24914 5000
rect 25134 4000 25190 5000
rect 25410 4000 25466 5000
rect 25686 4000 25742 5000
rect 25962 4000 26018 5000
rect 26238 4000 26294 5000
rect 26514 4000 26570 5000
rect 26790 4000 26846 5000
rect 27066 4004 27122 5000
rect 27066 4000 27068 4004
rect 22744 3946 22796 3952
rect 22756 2990 22784 3946
rect 22940 3194 22968 4000
rect 22928 3188 22980 3194
rect 22928 3130 22980 3136
rect 22744 2984 22796 2990
rect 22744 2926 22796 2932
rect 22652 2916 22704 2922
rect 22652 2858 22704 2864
rect 23216 2854 23244 4000
rect 23492 3466 23520 4000
rect 23296 3460 23348 3466
rect 23296 3402 23348 3408
rect 23480 3460 23532 3466
rect 23480 3402 23532 3408
rect 23308 3058 23336 3402
rect 23572 3392 23624 3398
rect 23572 3334 23624 3340
rect 23584 3058 23612 3334
rect 23768 3074 23796 4000
rect 24044 3210 24072 4000
rect 24320 3398 24348 4000
rect 24596 3534 24624 4000
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24308 3392 24360 3398
rect 24308 3334 24360 3340
rect 24044 3182 24256 3210
rect 23768 3058 23980 3074
rect 23296 3052 23348 3058
rect 23296 2994 23348 3000
rect 23572 3052 23624 3058
rect 23768 3052 23992 3058
rect 23768 3046 23940 3052
rect 23572 2994 23624 3000
rect 23940 2994 23992 3000
rect 24228 2990 24256 3182
rect 24872 3126 24900 4000
rect 24860 3120 24912 3126
rect 25148 3097 25176 4000
rect 25424 3602 25452 4000
rect 25412 3596 25464 3602
rect 25412 3538 25464 3544
rect 25228 3460 25280 3466
rect 25228 3402 25280 3408
rect 24860 3062 24912 3068
rect 25134 3088 25190 3097
rect 25240 3058 25268 3402
rect 25134 3023 25190 3032
rect 25228 3052 25280 3058
rect 25228 2994 25280 3000
rect 24216 2984 24268 2990
rect 24216 2926 24268 2932
rect 25700 2854 25728 4000
rect 25976 2990 26004 4000
rect 26252 3398 26280 4000
rect 26332 3528 26384 3534
rect 26332 3470 26384 3476
rect 26056 3392 26108 3398
rect 26056 3334 26108 3340
rect 26240 3392 26292 3398
rect 26240 3334 26292 3340
rect 26068 3058 26096 3334
rect 26344 3058 26372 3470
rect 26056 3052 26108 3058
rect 26056 2994 26108 3000
rect 26332 3052 26384 3058
rect 26332 2994 26384 3000
rect 25964 2984 26016 2990
rect 26528 2961 26556 4000
rect 26804 3126 26832 4000
rect 27120 4000 27122 4004
rect 27342 4000 27398 5000
rect 27618 4000 27674 5000
rect 27894 4000 27950 5000
rect 28170 4000 28226 5000
rect 28446 4000 28502 5000
rect 28722 4000 28778 5000
rect 28998 4000 29054 5000
rect 29092 4004 29144 4010
rect 27068 3946 27120 3952
rect 27054 3428 27154 3856
rect 27356 3754 27384 4000
rect 27356 3726 27568 3754
rect 27436 3596 27488 3602
rect 27436 3538 27488 3544
rect 27054 3372 27076 3428
rect 27132 3372 27154 3428
rect 27054 3290 27154 3372
rect 27054 3238 27078 3290
rect 27130 3238 27154 3290
rect 26792 3120 26844 3126
rect 26792 3062 26844 3068
rect 26882 3088 26938 3097
rect 26882 3023 26884 3032
rect 26936 3023 26938 3032
rect 26884 2994 26936 3000
rect 25964 2926 26016 2932
rect 26514 2952 26570 2961
rect 26514 2887 26570 2896
rect 23204 2848 23256 2854
rect 23204 2790 23256 2796
rect 25688 2848 25740 2854
rect 25688 2790 25740 2796
rect 21054 2694 21078 2746
rect 21130 2694 21154 2746
rect 16028 2576 16080 2582
rect 16028 2518 16080 2524
rect 17500 2576 17552 2582
rect 17500 2518 17552 2524
rect 15054 2150 15078 2202
rect 15130 2150 15154 2202
rect 9404 1760 9456 1766
rect 9404 1702 9456 1708
rect 11612 1760 11664 1766
rect 11612 1702 11664 1708
rect 12992 1760 13044 1766
rect 12992 1702 13044 1708
rect 14924 1760 14976 1766
rect 14924 1702 14976 1708
rect 9054 1606 9078 1658
rect 9130 1606 9154 1658
rect 8852 1352 8904 1358
rect 8852 1294 8904 1300
rect 8864 1000 8892 1294
rect 9054 1040 9154 1606
rect 9312 1488 9364 1494
rect 9312 1430 9364 1436
rect 3054 898 3110 1000
rect 2976 870 3110 898
rect 3054 0 3110 870
rect 3330 0 3386 1000
rect 3606 0 3662 1000
rect 3882 0 3938 1000
rect 4158 0 4214 1000
rect 4434 0 4490 1000
rect 4710 0 4766 1000
rect 4986 0 5042 1000
rect 5262 0 5318 1000
rect 5538 0 5594 1000
rect 5814 0 5870 1000
rect 6090 0 6146 1000
rect 6366 0 6422 1000
rect 6642 0 6698 1000
rect 6918 0 6974 1000
rect 7194 0 7250 1000
rect 7470 0 7526 1000
rect 7746 0 7802 1000
rect 8022 0 8078 1000
rect 8298 0 8354 1000
rect 8574 0 8630 1000
rect 8850 0 8906 1000
rect 9126 898 9182 1000
rect 9324 898 9352 1430
rect 9416 1000 9444 1702
rect 9956 1488 10008 1494
rect 9956 1430 10008 1436
rect 9680 1352 9732 1358
rect 9680 1294 9732 1300
rect 9692 1000 9720 1294
rect 9968 1000 9996 1430
rect 10232 1420 10284 1426
rect 10232 1362 10284 1368
rect 10784 1420 10836 1426
rect 10784 1362 10836 1368
rect 10244 1000 10272 1362
rect 10508 1352 10560 1358
rect 10508 1294 10560 1300
rect 10520 1000 10548 1294
rect 10796 1000 10824 1362
rect 11060 1352 11112 1358
rect 11060 1294 11112 1300
rect 11072 1000 11100 1294
rect 11336 1284 11388 1290
rect 11336 1226 11388 1232
rect 11348 1000 11376 1226
rect 11624 1000 11652 1702
rect 11888 1488 11940 1494
rect 11888 1430 11940 1436
rect 12716 1488 12768 1494
rect 12716 1430 12768 1436
rect 11900 1000 11928 1430
rect 12164 1420 12216 1426
rect 12164 1362 12216 1368
rect 12176 1000 12204 1362
rect 12440 1352 12492 1358
rect 12440 1294 12492 1300
rect 12452 1000 12480 1294
rect 12728 1000 12756 1430
rect 13004 1000 13032 1702
rect 13544 1488 13596 1494
rect 13544 1430 13596 1436
rect 14096 1488 14148 1494
rect 14096 1430 14148 1436
rect 13360 1352 13412 1358
rect 13280 1312 13360 1340
rect 13280 1000 13308 1312
rect 13360 1294 13412 1300
rect 13556 1000 13584 1430
rect 13820 1352 13872 1358
rect 13820 1294 13872 1300
rect 13832 1000 13860 1294
rect 14108 1000 14136 1430
rect 14648 1352 14700 1358
rect 14648 1294 14700 1300
rect 14372 1284 14424 1290
rect 14372 1226 14424 1232
rect 14384 1000 14412 1226
rect 14660 1000 14688 1294
rect 14936 1000 14964 1702
rect 15054 1268 15154 2150
rect 21054 2348 21154 2694
rect 21054 2292 21076 2348
rect 21132 2292 21154 2348
rect 15752 1760 15804 1766
rect 15752 1702 15804 1708
rect 19892 1760 19944 1766
rect 19892 1702 19944 1708
rect 15200 1488 15252 1494
rect 15200 1430 15252 1436
rect 15054 1212 15076 1268
rect 15132 1212 15154 1268
rect 15054 1114 15154 1212
rect 15054 1062 15078 1114
rect 15130 1062 15154 1114
rect 15054 1040 15154 1062
rect 15212 1000 15240 1430
rect 15476 1420 15528 1426
rect 15476 1362 15528 1368
rect 15488 1000 15516 1362
rect 15764 1000 15792 1702
rect 16304 1488 16356 1494
rect 16304 1430 16356 1436
rect 17132 1488 17184 1494
rect 17132 1430 17184 1436
rect 17960 1488 18012 1494
rect 17960 1430 18012 1436
rect 18788 1488 18840 1494
rect 18788 1430 18840 1436
rect 16028 1352 16080 1358
rect 16028 1294 16080 1300
rect 16040 1000 16068 1294
rect 16316 1000 16344 1430
rect 16856 1352 16908 1358
rect 16856 1294 16908 1300
rect 16580 1284 16632 1290
rect 16580 1226 16632 1232
rect 16592 1000 16620 1226
rect 16868 1000 16896 1294
rect 17144 1000 17172 1430
rect 17408 1420 17460 1426
rect 17408 1362 17460 1368
rect 17420 1000 17448 1362
rect 17684 1352 17736 1358
rect 17684 1294 17736 1300
rect 17696 1000 17724 1294
rect 17972 1000 18000 1430
rect 18236 1420 18288 1426
rect 18236 1362 18288 1368
rect 18248 1000 18276 1362
rect 18512 1352 18564 1358
rect 18512 1294 18564 1300
rect 18524 1000 18552 1294
rect 18800 1000 18828 1430
rect 19064 1420 19116 1426
rect 19064 1362 19116 1368
rect 19076 1000 19104 1362
rect 19340 1352 19392 1358
rect 19340 1294 19392 1300
rect 19352 1000 19380 1294
rect 19616 1284 19668 1290
rect 19616 1226 19668 1232
rect 19628 1000 19656 1226
rect 19904 1000 19932 1702
rect 21054 1658 21154 2292
rect 27054 2202 27154 3238
rect 27448 3058 27476 3538
rect 27540 3058 27568 3726
rect 27632 3074 27660 4000
rect 27908 3534 27936 4000
rect 28184 3602 28212 4000
rect 28460 3670 28488 4000
rect 28448 3664 28500 3670
rect 28448 3606 28500 3612
rect 28172 3596 28224 3602
rect 28172 3538 28224 3544
rect 27896 3528 27948 3534
rect 27896 3470 27948 3476
rect 28736 3398 28764 4000
rect 29012 3466 29040 4000
rect 29274 4000 29330 5000
rect 29550 4000 29606 5000
rect 29826 4000 29882 5000
rect 30102 4000 30158 5000
rect 30378 4000 30434 5000
rect 36174 4000 36230 5000
rect 36450 4000 36506 5000
rect 36726 4000 36782 5000
rect 37002 4000 37058 5000
rect 37278 4000 37334 5000
rect 37554 4000 37610 5000
rect 37830 4000 37886 5000
rect 38106 4000 38162 5000
rect 38382 4000 38438 5000
rect 38658 4000 38714 5000
rect 38934 4000 38990 5000
rect 39210 4000 39266 5000
rect 39486 4000 39542 5000
rect 39762 4000 39818 5000
rect 40038 4000 40094 5000
rect 40314 4000 40370 5000
rect 40590 4000 40646 5000
rect 40866 4000 40922 5000
rect 41142 4000 41198 5000
rect 41418 4000 41474 5000
rect 41694 4000 41750 5000
rect 41970 4000 42026 5000
rect 42246 4000 42302 5000
rect 42522 4000 42578 5000
rect 42798 4000 42854 5000
rect 43074 4000 43130 5000
rect 43350 4000 43406 5000
rect 43626 4000 43682 5000
rect 43902 4000 43958 5000
rect 44178 4000 44234 5000
rect 44454 4000 44510 5000
rect 44730 4000 44786 5000
rect 45006 4004 45062 5000
rect 45006 4000 45008 4004
rect 29092 3946 29144 3952
rect 29000 3460 29052 3466
rect 29000 3402 29052 3408
rect 28264 3392 28316 3398
rect 28264 3334 28316 3340
rect 28724 3392 28776 3398
rect 28724 3334 28776 3340
rect 27436 3052 27488 3058
rect 27436 2994 27488 3000
rect 27528 3052 27580 3058
rect 27632 3046 27844 3074
rect 28276 3058 28304 3334
rect 29104 3058 29132 3946
rect 29288 3194 29316 4000
rect 29276 3188 29328 3194
rect 29276 3130 29328 3136
rect 27528 2994 27580 3000
rect 27816 2922 27844 3046
rect 28264 3052 28316 3058
rect 28264 2994 28316 3000
rect 29092 3052 29144 3058
rect 29092 2994 29144 3000
rect 28538 2952 28594 2961
rect 27712 2916 27764 2922
rect 27712 2858 27764 2864
rect 27804 2916 27856 2922
rect 29564 2922 29592 4000
rect 29840 3126 29868 4000
rect 29920 3528 29972 3534
rect 29920 3470 29972 3476
rect 29828 3120 29880 3126
rect 29828 3062 29880 3068
rect 29932 3058 29960 3470
rect 29920 3052 29972 3058
rect 29920 2994 29972 3000
rect 30116 2990 30144 4000
rect 30196 3596 30248 3602
rect 30196 3538 30248 3544
rect 30208 3058 30236 3538
rect 30392 3058 30420 4000
rect 33054 3834 33154 3856
rect 33054 3782 33078 3834
rect 33130 3782 33154 3834
rect 30472 3664 30524 3670
rect 30472 3606 30524 3612
rect 30196 3052 30248 3058
rect 30196 2994 30248 3000
rect 30380 3052 30432 3058
rect 30380 2994 30432 3000
rect 30104 2984 30156 2990
rect 30104 2926 30156 2932
rect 28538 2887 28594 2896
rect 29552 2916 29604 2922
rect 27804 2858 27856 2864
rect 27620 2848 27672 2854
rect 27724 2802 27752 2858
rect 28552 2854 28580 2887
rect 29552 2858 29604 2864
rect 30484 2854 30512 3606
rect 31024 3460 31076 3466
rect 31024 3402 31076 3408
rect 30748 3392 30800 3398
rect 30748 3334 30800 3340
rect 30760 2854 30788 3334
rect 31036 2854 31064 3402
rect 31300 3188 31352 3194
rect 31300 3130 31352 3136
rect 31312 2854 31340 3130
rect 27672 2796 27752 2802
rect 27620 2790 27752 2796
rect 28540 2848 28592 2854
rect 28540 2790 28592 2796
rect 30472 2848 30524 2854
rect 30472 2790 30524 2796
rect 30748 2848 30800 2854
rect 30748 2790 30800 2796
rect 31024 2848 31076 2854
rect 31024 2790 31076 2796
rect 31300 2848 31352 2854
rect 31300 2790 31352 2796
rect 27632 2774 27752 2790
rect 27054 2150 27078 2202
rect 27130 2150 27154 2202
rect 25964 1760 26016 1766
rect 25964 1702 26016 1708
rect 21054 1606 21078 1658
rect 21130 1606 21154 1658
rect 20168 1488 20220 1494
rect 20168 1430 20220 1436
rect 20180 1000 20208 1430
rect 20720 1420 20772 1426
rect 20720 1362 20772 1368
rect 20444 1284 20496 1290
rect 20444 1226 20496 1232
rect 20456 1000 20484 1226
rect 20732 1000 20760 1362
rect 21054 1040 21154 1606
rect 24032 1556 24084 1562
rect 24032 1498 24084 1504
rect 25412 1556 25464 1562
rect 25412 1498 25464 1504
rect 21272 1488 21324 1494
rect 21192 1448 21272 1476
rect 9126 870 9352 898
rect 9126 0 9182 870
rect 9402 0 9458 1000
rect 9678 0 9734 1000
rect 9954 0 10010 1000
rect 10230 0 10286 1000
rect 10506 0 10562 1000
rect 10782 0 10838 1000
rect 11058 0 11114 1000
rect 11334 0 11390 1000
rect 11610 0 11666 1000
rect 11886 0 11942 1000
rect 12162 0 12218 1000
rect 12438 0 12494 1000
rect 12714 0 12770 1000
rect 12990 0 13046 1000
rect 13266 0 13322 1000
rect 13542 0 13598 1000
rect 13818 0 13874 1000
rect 14094 0 14150 1000
rect 14370 0 14426 1000
rect 14646 0 14702 1000
rect 14922 0 14978 1000
rect 15198 0 15254 1000
rect 15474 0 15530 1000
rect 15750 0 15806 1000
rect 16026 0 16082 1000
rect 16302 0 16358 1000
rect 16578 0 16634 1000
rect 16854 0 16910 1000
rect 17130 0 17186 1000
rect 17406 0 17462 1000
rect 17682 0 17738 1000
rect 17958 0 18014 1000
rect 18234 0 18290 1000
rect 18510 0 18566 1000
rect 18786 0 18842 1000
rect 19062 0 19118 1000
rect 19338 0 19394 1000
rect 19614 0 19670 1000
rect 19890 0 19946 1000
rect 20166 0 20222 1000
rect 20442 0 20498 1000
rect 20718 0 20774 1000
rect 20994 898 21050 1000
rect 21192 898 21220 1448
rect 21272 1430 21324 1436
rect 22652 1488 22704 1494
rect 22652 1430 22704 1436
rect 23480 1488 23532 1494
rect 23480 1430 23532 1436
rect 21548 1420 21600 1426
rect 21548 1362 21600 1368
rect 22376 1420 22428 1426
rect 22376 1362 22428 1368
rect 21272 1352 21324 1358
rect 21272 1294 21324 1300
rect 21284 1000 21312 1294
rect 21560 1000 21588 1362
rect 21824 1352 21876 1358
rect 21824 1294 21876 1300
rect 21836 1000 21864 1294
rect 22100 1284 22152 1290
rect 22100 1226 22152 1232
rect 22112 1000 22140 1226
rect 22388 1000 22416 1362
rect 22664 1000 22692 1430
rect 23204 1420 23256 1426
rect 23204 1362 23256 1368
rect 22928 1284 22980 1290
rect 22928 1226 22980 1232
rect 22940 1000 22968 1226
rect 23216 1000 23244 1362
rect 23492 1000 23520 1430
rect 23756 1284 23808 1290
rect 23756 1226 23808 1232
rect 23768 1000 23796 1226
rect 24044 1000 24072 1498
rect 24584 1488 24636 1494
rect 24584 1430 24636 1436
rect 24308 1352 24360 1358
rect 24308 1294 24360 1300
rect 24320 1000 24348 1294
rect 24596 1000 24624 1430
rect 24860 1352 24912 1358
rect 24860 1294 24912 1300
rect 24872 1000 24900 1294
rect 25136 1284 25188 1290
rect 25136 1226 25188 1232
rect 25148 1000 25176 1226
rect 25424 1000 25452 1498
rect 25688 1216 25740 1222
rect 25688 1158 25740 1164
rect 25700 1000 25728 1158
rect 25976 1000 26004 1702
rect 26516 1488 26568 1494
rect 26516 1430 26568 1436
rect 26240 1420 26292 1426
rect 26240 1362 26292 1368
rect 26252 1000 26280 1362
rect 26528 1000 26556 1430
rect 26792 1352 26844 1358
rect 26792 1294 26844 1300
rect 26804 1000 26832 1294
rect 27054 1268 27154 2150
rect 33054 2746 33154 3782
rect 36188 3058 36216 4000
rect 36464 3058 36492 4000
rect 36176 3052 36228 3058
rect 36176 2994 36228 3000
rect 36452 3052 36504 3058
rect 36452 2994 36504 3000
rect 36740 2922 36768 4000
rect 37016 3058 37044 4000
rect 37292 3058 37320 4000
rect 37568 3058 37596 4000
rect 37004 3052 37056 3058
rect 37004 2994 37056 3000
rect 37280 3052 37332 3058
rect 37280 2994 37332 3000
rect 37556 3052 37608 3058
rect 37556 2994 37608 3000
rect 37844 2990 37872 4000
rect 38120 3058 38148 4000
rect 38108 3052 38160 3058
rect 38108 2994 38160 3000
rect 38396 2990 38424 4000
rect 38672 3058 38700 4000
rect 38660 3052 38712 3058
rect 38660 2994 38712 3000
rect 38948 2990 38976 4000
rect 39054 3428 39154 3856
rect 39054 3372 39076 3428
rect 39132 3372 39154 3428
rect 39054 3290 39154 3372
rect 39054 3238 39078 3290
rect 39130 3238 39154 3290
rect 37832 2984 37884 2990
rect 37832 2926 37884 2932
rect 38384 2984 38436 2990
rect 38384 2926 38436 2932
rect 38936 2984 38988 2990
rect 38936 2926 38988 2932
rect 36728 2916 36780 2922
rect 36728 2858 36780 2864
rect 33054 2694 33078 2746
rect 33130 2694 33154 2746
rect 33054 2348 33154 2694
rect 33054 2292 33076 2348
rect 33132 2292 33154 2348
rect 30104 1828 30156 1834
rect 30104 1770 30156 1776
rect 29828 1760 29880 1766
rect 29828 1702 29880 1708
rect 27436 1556 27488 1562
rect 27356 1516 27436 1544
rect 27054 1212 27076 1268
rect 27132 1212 27154 1268
rect 27252 1284 27304 1290
rect 27252 1226 27304 1232
rect 27054 1114 27154 1212
rect 27054 1062 27078 1114
rect 27130 1062 27154 1114
rect 27054 1040 27154 1062
rect 20994 870 21220 898
rect 20994 0 21050 870
rect 21270 0 21326 1000
rect 21546 0 21602 1000
rect 21822 0 21878 1000
rect 22098 0 22154 1000
rect 22374 0 22430 1000
rect 22650 0 22706 1000
rect 22926 0 22982 1000
rect 23202 0 23258 1000
rect 23478 0 23534 1000
rect 23754 0 23810 1000
rect 24030 0 24086 1000
rect 24306 0 24362 1000
rect 24582 0 24638 1000
rect 24858 0 24914 1000
rect 25134 0 25190 1000
rect 25410 0 25466 1000
rect 25686 0 25742 1000
rect 25962 0 26018 1000
rect 26238 0 26294 1000
rect 26514 0 26570 1000
rect 26790 0 26846 1000
rect 27066 898 27122 1000
rect 27264 898 27292 1226
rect 27356 1000 27384 1516
rect 27436 1498 27488 1504
rect 29552 1556 29604 1562
rect 29552 1498 29604 1504
rect 27896 1488 27948 1494
rect 27896 1430 27948 1436
rect 29276 1488 29328 1494
rect 29276 1430 29328 1436
rect 27620 1420 27672 1426
rect 27620 1362 27672 1368
rect 27632 1000 27660 1362
rect 27908 1000 27936 1430
rect 28724 1420 28776 1426
rect 28724 1362 28776 1368
rect 28264 1352 28316 1358
rect 28184 1312 28264 1340
rect 28184 1000 28212 1312
rect 28264 1294 28316 1300
rect 28448 1216 28500 1222
rect 28448 1158 28500 1164
rect 28460 1000 28488 1158
rect 28736 1000 28764 1362
rect 29000 1216 29052 1222
rect 29000 1158 29052 1164
rect 29012 1000 29040 1158
rect 29288 1000 29316 1430
rect 29564 1000 29592 1498
rect 29840 1000 29868 1702
rect 30116 1000 30144 1770
rect 31484 1760 31536 1766
rect 31484 1702 31536 1708
rect 31208 1556 31260 1562
rect 31208 1498 31260 1504
rect 30656 1488 30708 1494
rect 30656 1430 30708 1436
rect 30380 1420 30432 1426
rect 30380 1362 30432 1368
rect 30392 1000 30420 1362
rect 30668 1000 30696 1430
rect 30932 1352 30984 1358
rect 30932 1294 30984 1300
rect 30944 1000 30972 1294
rect 31220 1000 31248 1498
rect 31496 1000 31524 1702
rect 33054 1658 33154 2292
rect 39054 2202 39154 3238
rect 39224 3058 39252 4000
rect 39212 3052 39264 3058
rect 39212 2994 39264 3000
rect 39500 2990 39528 4000
rect 39776 3058 39804 4000
rect 39764 3052 39816 3058
rect 39764 2994 39816 3000
rect 40052 2990 40080 4000
rect 40328 3058 40356 4000
rect 40316 3052 40368 3058
rect 40316 2994 40368 3000
rect 40604 2990 40632 4000
rect 40880 3058 40908 4000
rect 40868 3052 40920 3058
rect 40868 2994 40920 3000
rect 41156 2990 41184 4000
rect 41432 3058 41460 4000
rect 41420 3052 41472 3058
rect 41420 2994 41472 3000
rect 41708 2990 41736 4000
rect 41984 3058 42012 4000
rect 41972 3052 42024 3058
rect 41972 2994 42024 3000
rect 42260 2990 42288 4000
rect 42536 3058 42564 4000
rect 42524 3052 42576 3058
rect 42524 2994 42576 3000
rect 42812 2990 42840 4000
rect 39488 2984 39540 2990
rect 39488 2926 39540 2932
rect 40040 2984 40092 2990
rect 40040 2926 40092 2932
rect 40592 2984 40644 2990
rect 40592 2926 40644 2932
rect 41144 2984 41196 2990
rect 41144 2926 41196 2932
rect 41696 2984 41748 2990
rect 41696 2926 41748 2932
rect 42248 2984 42300 2990
rect 42248 2926 42300 2932
rect 42800 2984 42852 2990
rect 42800 2926 42852 2932
rect 43088 2922 43116 4000
rect 43364 3058 43392 4000
rect 43352 3052 43404 3058
rect 43352 2994 43404 3000
rect 43640 2990 43668 4000
rect 43628 2984 43680 2990
rect 43628 2926 43680 2932
rect 43916 2922 43944 4000
rect 44192 3058 44220 4000
rect 44180 3052 44232 3058
rect 44180 2994 44232 3000
rect 44468 2990 44496 4000
rect 44456 2984 44508 2990
rect 44456 2926 44508 2932
rect 44744 2922 44772 4000
rect 45060 4000 45062 4004
rect 45282 4000 45338 5000
rect 45558 4000 45614 5000
rect 45652 4004 45704 4010
rect 45008 3946 45060 3952
rect 45054 3834 45154 3856
rect 45054 3782 45078 3834
rect 45130 3782 45154 3834
rect 43076 2916 43128 2922
rect 43076 2858 43128 2864
rect 43904 2916 43956 2922
rect 43904 2858 43956 2864
rect 44732 2916 44784 2922
rect 44732 2858 44784 2864
rect 39054 2150 39078 2202
rect 39130 2150 39154 2202
rect 38936 1760 38988 1766
rect 38936 1702 38988 1708
rect 33054 1606 33078 1658
rect 33130 1606 33154 1658
rect 32036 1488 32088 1494
rect 32036 1430 32088 1436
rect 31760 1284 31812 1290
rect 31760 1226 31812 1232
rect 31772 1000 31800 1226
rect 32048 1000 32076 1430
rect 32312 1420 32364 1426
rect 32312 1362 32364 1368
rect 32324 1000 32352 1362
rect 33054 1040 33154 1606
rect 38108 1488 38160 1494
rect 38108 1430 38160 1436
rect 38120 1000 38148 1430
rect 38292 1352 38344 1358
rect 38660 1352 38712 1358
rect 38344 1312 38424 1340
rect 38292 1294 38344 1300
rect 38396 1000 38424 1312
rect 38660 1294 38712 1300
rect 38672 1000 38700 1294
rect 38948 1000 38976 1702
rect 39054 1268 39154 2150
rect 45054 2746 45154 3782
rect 45296 2990 45324 4000
rect 45284 2984 45336 2990
rect 45284 2926 45336 2932
rect 45572 2922 45600 4000
rect 45834 4000 45890 5000
rect 46110 4000 46166 5000
rect 46386 4000 46442 5000
rect 46662 4000 46718 5000
rect 46938 4000 46994 5000
rect 47214 4000 47270 5000
rect 47490 4000 47546 5000
rect 47766 4000 47822 5000
rect 48042 4000 48098 5000
rect 48318 4000 48374 5000
rect 48594 4000 48650 5000
rect 48870 4000 48926 5000
rect 49146 4000 49202 5000
rect 49422 4000 49478 5000
rect 49698 4000 49754 5000
rect 49974 4000 50030 5000
rect 50250 4000 50306 5000
rect 50526 4000 50582 5000
rect 50802 4000 50858 5000
rect 51078 4004 51134 5000
rect 51078 4000 51080 4004
rect 45652 3946 45704 3952
rect 45664 3058 45692 3946
rect 45848 3058 45876 4000
rect 45652 3052 45704 3058
rect 45652 2994 45704 3000
rect 45836 3052 45888 3058
rect 45836 2994 45888 3000
rect 46124 2990 46152 4000
rect 46112 2984 46164 2990
rect 46112 2926 46164 2932
rect 46400 2922 46428 4000
rect 46676 3058 46704 4000
rect 46664 3052 46716 3058
rect 46664 2994 46716 3000
rect 46952 2990 46980 4000
rect 46940 2984 46992 2990
rect 46940 2926 46992 2932
rect 47228 2922 47256 4000
rect 45560 2916 45612 2922
rect 45560 2858 45612 2864
rect 46388 2916 46440 2922
rect 46388 2858 46440 2864
rect 47216 2916 47268 2922
rect 47216 2858 47268 2864
rect 47504 2854 47532 4000
rect 47780 2990 47808 4000
rect 48056 3058 48084 4000
rect 48332 3126 48360 4000
rect 48320 3120 48372 3126
rect 48320 3062 48372 3068
rect 48044 3052 48096 3058
rect 48044 2994 48096 3000
rect 48608 2990 48636 4000
rect 47768 2984 47820 2990
rect 47768 2926 47820 2932
rect 48596 2984 48648 2990
rect 48596 2926 48648 2932
rect 48884 2922 48912 4000
rect 48872 2916 48924 2922
rect 48872 2858 48924 2864
rect 49160 2854 49188 4000
rect 49436 3058 49464 4000
rect 49424 3052 49476 3058
rect 49424 2994 49476 3000
rect 49712 2990 49740 4000
rect 49700 2984 49752 2990
rect 49700 2926 49752 2932
rect 49988 2922 50016 4000
rect 50264 3126 50292 4000
rect 50252 3120 50304 3126
rect 50252 3062 50304 3068
rect 49976 2916 50028 2922
rect 49976 2858 50028 2864
rect 50540 2854 50568 4000
rect 50816 2990 50844 4000
rect 51132 4000 51134 4004
rect 51354 4000 51410 5000
rect 51630 4000 51686 5000
rect 51906 4000 51962 5000
rect 52000 4004 52052 4010
rect 51080 3946 51132 3952
rect 51054 3428 51154 3856
rect 51054 3372 51076 3428
rect 51132 3372 51154 3428
rect 51054 3290 51154 3372
rect 51054 3238 51078 3290
rect 51130 3238 51154 3290
rect 50804 2984 50856 2990
rect 50804 2926 50856 2932
rect 47492 2848 47544 2854
rect 47492 2790 47544 2796
rect 49148 2848 49200 2854
rect 49148 2790 49200 2796
rect 50528 2848 50580 2854
rect 50528 2790 50580 2796
rect 45054 2694 45078 2746
rect 45130 2694 45154 2746
rect 45054 2348 45154 2694
rect 45054 2292 45076 2348
rect 45132 2292 45154 2348
rect 44180 1760 44232 1766
rect 44180 1702 44232 1708
rect 39488 1488 39540 1494
rect 39488 1430 39540 1436
rect 40592 1488 40644 1494
rect 40592 1430 40644 1436
rect 41696 1488 41748 1494
rect 41696 1430 41748 1436
rect 42248 1488 42300 1494
rect 42248 1430 42300 1436
rect 42800 1488 42852 1494
rect 42800 1430 42852 1436
rect 43352 1488 43404 1494
rect 43352 1430 43404 1436
rect 39212 1420 39264 1426
rect 39212 1362 39264 1368
rect 39054 1212 39076 1268
rect 39132 1212 39154 1268
rect 39054 1114 39154 1212
rect 39054 1062 39078 1114
rect 39130 1062 39154 1114
rect 39054 1040 39154 1062
rect 39224 1000 39252 1362
rect 39500 1000 39528 1430
rect 39764 1420 39816 1426
rect 39764 1362 39816 1368
rect 40316 1420 40368 1426
rect 40316 1362 40368 1368
rect 39776 1000 39804 1362
rect 40040 1352 40092 1358
rect 40040 1294 40092 1300
rect 40052 1000 40080 1294
rect 40328 1000 40356 1362
rect 40604 1000 40632 1430
rect 41144 1420 41196 1426
rect 41144 1362 41196 1368
rect 40868 1352 40920 1358
rect 40868 1294 40920 1300
rect 40880 1000 40908 1294
rect 41156 1000 41184 1362
rect 41328 1352 41380 1358
rect 41380 1312 41460 1340
rect 41328 1294 41380 1300
rect 41432 1000 41460 1312
rect 41708 1000 41736 1430
rect 41972 1352 42024 1358
rect 41972 1294 42024 1300
rect 41984 1000 42012 1294
rect 42260 1000 42288 1430
rect 42524 1352 42576 1358
rect 42524 1294 42576 1300
rect 42536 1000 42564 1294
rect 42812 1000 42840 1430
rect 43076 1352 43128 1358
rect 43076 1294 43128 1300
rect 43088 1000 43116 1294
rect 43364 1000 43392 1430
rect 43628 1352 43680 1358
rect 43628 1294 43680 1300
rect 43904 1352 43956 1358
rect 43904 1294 43956 1300
rect 43640 1000 43668 1294
rect 43916 1000 43944 1294
rect 44192 1000 44220 1702
rect 45054 1658 45154 2292
rect 51054 2202 51154 3238
rect 51368 2922 51396 4000
rect 51644 3126 51672 4000
rect 51632 3120 51684 3126
rect 51632 3062 51684 3068
rect 51920 2990 51948 4000
rect 52182 4000 52238 5000
rect 52458 4000 52514 5000
rect 52734 4000 52790 5000
rect 53010 4000 53066 5000
rect 53286 4000 53342 5000
rect 53562 4000 53618 5000
rect 53838 4000 53894 5000
rect 54114 4000 54170 5000
rect 54390 4000 54446 5000
rect 54666 4000 54722 5000
rect 54942 4000 54998 5000
rect 55218 4000 55274 5000
rect 55494 4000 55550 5000
rect 55770 4000 55826 5000
rect 56046 4000 56102 5000
rect 56322 4000 56378 5000
rect 56598 4000 56654 5000
rect 56874 4000 56930 5000
rect 57150 4004 57206 5000
rect 57150 4000 57152 4004
rect 52000 3946 52052 3952
rect 52012 3058 52040 3946
rect 52000 3052 52052 3058
rect 52000 2994 52052 3000
rect 51908 2984 51960 2990
rect 51908 2926 51960 2932
rect 51356 2916 51408 2922
rect 51356 2858 51408 2864
rect 52196 2854 52224 4000
rect 52472 2922 52500 4000
rect 52748 3058 52776 4000
rect 52736 3052 52788 3058
rect 52736 2994 52788 3000
rect 53024 2990 53052 4000
rect 53300 3126 53328 4000
rect 53288 3120 53340 3126
rect 53288 3062 53340 3068
rect 53012 2984 53064 2990
rect 53012 2926 53064 2932
rect 52460 2916 52512 2922
rect 52460 2858 52512 2864
rect 53576 2854 53604 4000
rect 53852 2922 53880 4000
rect 54128 3058 54156 4000
rect 54404 3194 54432 4000
rect 54392 3188 54444 3194
rect 54392 3130 54444 3136
rect 54680 3058 54708 4000
rect 54116 3052 54168 3058
rect 54116 2994 54168 3000
rect 54668 3052 54720 3058
rect 54668 2994 54720 3000
rect 53840 2916 53892 2922
rect 53840 2858 53892 2864
rect 54956 2854 54984 4000
rect 55232 2922 55260 4000
rect 55508 3074 55536 4000
rect 55784 3126 55812 4000
rect 55772 3120 55824 3126
rect 55508 3058 55720 3074
rect 55772 3062 55824 3068
rect 55508 3052 55732 3058
rect 55508 3046 55680 3052
rect 55680 2994 55732 3000
rect 56060 2990 56088 4000
rect 56336 3466 56364 4000
rect 56324 3460 56376 3466
rect 56324 3402 56376 3408
rect 56048 2984 56100 2990
rect 56048 2926 56100 2932
rect 56612 2922 56640 4000
rect 56888 3194 56916 4000
rect 57204 4000 57206 4004
rect 57336 4004 57388 4010
rect 57152 3946 57204 3952
rect 57426 4000 57482 5000
rect 57702 4000 57758 5000
rect 57978 4000 58034 5000
rect 58254 4000 58310 5000
rect 58530 4000 58586 5000
rect 58806 4000 58862 5000
rect 59082 4000 59138 5000
rect 59358 4000 59414 5000
rect 59634 4000 59690 5000
rect 59910 4000 59966 5000
rect 60186 4000 60242 5000
rect 60462 4000 60518 5000
rect 60738 4000 60794 5000
rect 61014 4000 61070 5000
rect 61290 4000 61346 5000
rect 61566 4000 61622 5000
rect 61842 4000 61898 5000
rect 62118 4000 62174 5000
rect 62394 4000 62450 5000
rect 62670 4000 62726 5000
rect 62946 4000 63002 5000
rect 63222 4000 63278 5000
rect 63498 4000 63554 5000
rect 63774 4000 63830 5000
rect 64050 4000 64106 5000
rect 64326 4000 64382 5000
rect 64602 4000 64658 5000
rect 64878 4000 64934 5000
rect 65154 4000 65210 5000
rect 65430 4000 65486 5000
rect 65706 4000 65762 5000
rect 65982 4000 66038 5000
rect 66258 4000 66314 5000
rect 66534 4000 66590 5000
rect 66810 4000 66866 5000
rect 67086 4000 67142 5000
rect 67362 4000 67418 5000
rect 57336 3946 57388 3952
rect 57054 3834 57154 3856
rect 57054 3782 57078 3834
rect 57130 3782 57154 3834
rect 56876 3188 56928 3194
rect 56876 3130 56928 3136
rect 55220 2916 55272 2922
rect 55220 2858 55272 2864
rect 56600 2916 56652 2922
rect 56600 2858 56652 2864
rect 52184 2848 52236 2854
rect 52184 2790 52236 2796
rect 53564 2848 53616 2854
rect 53564 2790 53616 2796
rect 54944 2848 54996 2854
rect 54944 2790 54996 2796
rect 51054 2150 51078 2202
rect 51130 2150 51154 2202
rect 46940 1760 46992 1766
rect 46940 1702 46992 1708
rect 50528 1760 50580 1766
rect 50528 1702 50580 1708
rect 45054 1606 45078 1658
rect 45130 1606 45154 1658
rect 44456 1352 44508 1358
rect 44456 1294 44508 1300
rect 44732 1352 44784 1358
rect 44732 1294 44784 1300
rect 44916 1352 44968 1358
rect 44916 1294 44968 1300
rect 44468 1000 44496 1294
rect 44744 1000 44772 1294
rect 27066 870 27292 898
rect 27066 0 27122 870
rect 27342 0 27398 1000
rect 27618 0 27674 1000
rect 27894 0 27950 1000
rect 28170 0 28226 1000
rect 28446 0 28502 1000
rect 28722 0 28778 1000
rect 28998 0 29054 1000
rect 29274 0 29330 1000
rect 29550 0 29606 1000
rect 29826 0 29882 1000
rect 30102 0 30158 1000
rect 30378 0 30434 1000
rect 30654 0 30710 1000
rect 30930 0 30986 1000
rect 31206 0 31262 1000
rect 31482 0 31538 1000
rect 31758 0 31814 1000
rect 32034 0 32090 1000
rect 32310 0 32366 1000
rect 38106 0 38162 1000
rect 38382 0 38438 1000
rect 38658 0 38714 1000
rect 38934 0 38990 1000
rect 39210 0 39266 1000
rect 39486 0 39542 1000
rect 39762 0 39818 1000
rect 40038 0 40094 1000
rect 40314 0 40370 1000
rect 40590 0 40646 1000
rect 40866 0 40922 1000
rect 41142 0 41198 1000
rect 41418 0 41474 1000
rect 41694 0 41750 1000
rect 41970 0 42026 1000
rect 42246 0 42302 1000
rect 42522 0 42578 1000
rect 42798 0 42854 1000
rect 43074 0 43130 1000
rect 43350 0 43406 1000
rect 43626 0 43682 1000
rect 43902 0 43958 1000
rect 44178 0 44234 1000
rect 44454 0 44510 1000
rect 44730 0 44786 1000
rect 44928 898 44956 1294
rect 45054 1040 45154 1606
rect 45284 1352 45336 1358
rect 45284 1294 45336 1300
rect 45560 1352 45612 1358
rect 45560 1294 45612 1300
rect 45836 1352 45888 1358
rect 45836 1294 45888 1300
rect 46112 1352 46164 1358
rect 46112 1294 46164 1300
rect 46388 1352 46440 1358
rect 46388 1294 46440 1300
rect 46664 1352 46716 1358
rect 46664 1294 46716 1300
rect 45296 1000 45324 1294
rect 45572 1000 45600 1294
rect 45848 1000 45876 1294
rect 46124 1000 46152 1294
rect 46400 1000 46428 1294
rect 46676 1000 46704 1294
rect 46952 1000 46980 1702
rect 49148 1420 49200 1426
rect 49148 1362 49200 1368
rect 49700 1420 49752 1426
rect 49700 1362 49752 1368
rect 47216 1352 47268 1358
rect 47216 1294 47268 1300
rect 47492 1352 47544 1358
rect 47492 1294 47544 1300
rect 47768 1352 47820 1358
rect 47768 1294 47820 1300
rect 48044 1352 48096 1358
rect 48044 1294 48096 1300
rect 48320 1352 48372 1358
rect 48320 1294 48372 1300
rect 48596 1352 48648 1358
rect 48596 1294 48648 1300
rect 48872 1352 48924 1358
rect 48872 1294 48924 1300
rect 47228 1000 47256 1294
rect 47504 1000 47532 1294
rect 47780 1000 47808 1294
rect 48056 1000 48084 1294
rect 48332 1000 48360 1294
rect 48608 1000 48636 1294
rect 48884 1000 48912 1294
rect 49160 1000 49188 1362
rect 49424 1352 49476 1358
rect 49424 1294 49476 1300
rect 49436 1000 49464 1294
rect 49712 1000 49740 1362
rect 49976 1352 50028 1358
rect 49976 1294 50028 1300
rect 50252 1352 50304 1358
rect 50252 1294 50304 1300
rect 49988 1000 50016 1294
rect 50264 1000 50292 1294
rect 50540 1000 50568 1702
rect 50804 1352 50856 1358
rect 50804 1294 50856 1300
rect 50816 1000 50844 1294
rect 51054 1268 51154 2150
rect 57054 2746 57154 3782
rect 57348 3618 57376 3946
rect 57256 3590 57376 3618
rect 57256 2990 57284 3590
rect 57336 3460 57388 3466
rect 57336 3402 57388 3408
rect 57244 2984 57296 2990
rect 57244 2926 57296 2932
rect 57348 2854 57376 3402
rect 57440 2958 57468 4000
rect 57716 2958 57744 4000
rect 57992 3040 58020 4000
rect 58268 3126 58296 4000
rect 58256 3120 58308 3126
rect 58256 3062 58308 3068
rect 58164 3052 58216 3058
rect 57992 3012 58164 3040
rect 58164 2994 58216 3000
rect 58544 2990 58572 4000
rect 58820 3194 58848 4000
rect 58808 3188 58860 3194
rect 58808 3130 58860 3136
rect 58532 2984 58584 2990
rect 57440 2930 57652 2958
rect 57716 2930 57836 2958
rect 57624 2854 57652 2930
rect 57336 2848 57388 2854
rect 57336 2790 57388 2796
rect 57612 2848 57664 2854
rect 57612 2790 57664 2796
rect 57808 2802 57836 2930
rect 58532 2926 58584 2932
rect 59096 2922 59124 4000
rect 59372 2922 59400 4000
rect 59648 3040 59676 4000
rect 59924 3466 59952 4000
rect 59912 3460 59964 3466
rect 59912 3402 59964 3408
rect 60200 3108 60228 4000
rect 60372 3120 60424 3126
rect 60200 3080 60372 3108
rect 60372 3062 60424 3068
rect 60476 3058 60504 4000
rect 59820 3052 59872 3058
rect 59648 3012 59820 3040
rect 59820 2994 59872 3000
rect 60464 3052 60516 3058
rect 60464 2994 60516 3000
rect 58072 2916 58124 2922
rect 58072 2858 58124 2864
rect 59084 2916 59136 2922
rect 59084 2858 59136 2864
rect 59360 2916 59412 2922
rect 59360 2858 59412 2864
rect 58084 2802 58112 2858
rect 60752 2854 60780 4000
rect 61028 3194 61056 4000
rect 61304 3398 61332 4000
rect 61580 3466 61608 4000
rect 61384 3460 61436 3466
rect 61384 3402 61436 3408
rect 61568 3460 61620 3466
rect 61568 3402 61620 3408
rect 61292 3392 61344 3398
rect 61292 3334 61344 3340
rect 61016 3188 61068 3194
rect 61016 3130 61068 3136
rect 61396 3058 61424 3402
rect 61384 3052 61436 3058
rect 61384 2994 61436 3000
rect 61856 2922 61884 4000
rect 62132 2938 62160 4000
rect 62408 2990 62436 4000
rect 62396 2984 62448 2990
rect 61844 2916 61896 2922
rect 62132 2910 62344 2938
rect 62396 2926 62448 2932
rect 61844 2858 61896 2864
rect 62316 2854 62344 2910
rect 57808 2774 58112 2802
rect 60740 2848 60792 2854
rect 60740 2790 60792 2796
rect 62304 2848 62356 2854
rect 62304 2790 62356 2796
rect 57054 2694 57078 2746
rect 57130 2694 57154 2746
rect 57054 2348 57154 2694
rect 62684 2582 62712 4000
rect 62960 3738 62988 4000
rect 63236 3924 63264 4000
rect 63236 3896 63356 3924
rect 62948 3732 63000 3738
rect 62948 3674 63000 3680
rect 62948 3460 63000 3466
rect 62948 3402 63000 3408
rect 63054 3428 63154 3856
rect 62764 3392 62816 3398
rect 62764 3334 62816 3340
rect 62776 3058 62804 3334
rect 62960 3058 62988 3402
rect 63054 3372 63076 3428
rect 63132 3372 63154 3428
rect 63054 3290 63154 3372
rect 63054 3238 63078 3290
rect 63130 3238 63154 3290
rect 62764 3052 62816 3058
rect 62764 2994 62816 3000
rect 62948 3052 63000 3058
rect 62948 2994 63000 3000
rect 62672 2576 62724 2582
rect 62672 2518 62724 2524
rect 57054 2292 57076 2348
rect 57132 2292 57154 2348
rect 52460 1760 52512 1766
rect 52460 1702 52512 1708
rect 54392 1760 54444 1766
rect 54392 1702 54444 1708
rect 51908 1420 51960 1426
rect 51908 1362 51960 1368
rect 51264 1352 51316 1358
rect 51264 1294 51316 1300
rect 51356 1352 51408 1358
rect 51356 1294 51408 1300
rect 51632 1352 51684 1358
rect 51632 1294 51684 1300
rect 51054 1212 51076 1268
rect 51132 1212 51154 1268
rect 51054 1114 51154 1212
rect 51054 1062 51078 1114
rect 51130 1062 51154 1114
rect 51054 1040 51154 1062
rect 45006 898 45062 1000
rect 44928 870 45062 898
rect 45006 0 45062 870
rect 45282 0 45338 1000
rect 45558 0 45614 1000
rect 45834 0 45890 1000
rect 46110 0 46166 1000
rect 46386 0 46442 1000
rect 46662 0 46718 1000
rect 46938 0 46994 1000
rect 47214 0 47270 1000
rect 47490 0 47546 1000
rect 47766 0 47822 1000
rect 48042 0 48098 1000
rect 48318 0 48374 1000
rect 48594 0 48650 1000
rect 48870 0 48926 1000
rect 49146 0 49202 1000
rect 49422 0 49478 1000
rect 49698 0 49754 1000
rect 49974 0 50030 1000
rect 50250 0 50306 1000
rect 50526 0 50582 1000
rect 50802 0 50858 1000
rect 51078 898 51134 1000
rect 51276 898 51304 1294
rect 51368 1000 51396 1294
rect 51644 1000 51672 1294
rect 51920 1000 51948 1362
rect 52184 1352 52236 1358
rect 52184 1294 52236 1300
rect 52196 1000 52224 1294
rect 52472 1000 52500 1702
rect 52736 1352 52788 1358
rect 52736 1294 52788 1300
rect 53012 1352 53064 1358
rect 53012 1294 53064 1300
rect 53288 1352 53340 1358
rect 53288 1294 53340 1300
rect 53564 1352 53616 1358
rect 53564 1294 53616 1300
rect 53840 1352 53892 1358
rect 53840 1294 53892 1300
rect 54116 1352 54168 1358
rect 54116 1294 54168 1300
rect 52748 1000 52776 1294
rect 53024 1000 53052 1294
rect 53300 1000 53328 1294
rect 53576 1000 53604 1294
rect 53852 1000 53880 1294
rect 54128 1000 54156 1294
rect 54404 1000 54432 1702
rect 57054 1658 57154 2292
rect 63054 2202 63154 3238
rect 63328 3126 63356 3896
rect 63316 3120 63368 3126
rect 63316 3062 63368 3068
rect 63512 2922 63540 4000
rect 63788 3058 63816 4000
rect 64064 3194 64092 4000
rect 64052 3188 64104 3194
rect 64052 3130 64104 3136
rect 63776 3052 63828 3058
rect 63776 2994 63828 3000
rect 64340 2938 64368 4000
rect 64616 3534 64644 4000
rect 64696 3732 64748 3738
rect 64696 3674 64748 3680
rect 64604 3528 64656 3534
rect 64604 3470 64656 3476
rect 64708 3058 64736 3674
rect 64892 3074 64920 4000
rect 64892 3058 65104 3074
rect 64696 3052 64748 3058
rect 64892 3052 65116 3058
rect 64892 3046 65064 3052
rect 64696 2994 64748 3000
rect 65064 2994 65116 3000
rect 65168 2958 65196 4000
rect 65444 3398 65472 4000
rect 65720 3602 65748 4000
rect 65708 3596 65760 3602
rect 65708 3538 65760 3544
rect 65996 3466 66024 4000
rect 65984 3460 66036 3466
rect 65984 3402 66036 3408
rect 65432 3392 65484 3398
rect 65432 3334 65484 3340
rect 66272 3194 66300 4000
rect 66352 3528 66404 3534
rect 66352 3470 66404 3476
rect 66260 3188 66312 3194
rect 66260 3130 66312 3136
rect 66364 3058 66392 3470
rect 66352 3052 66404 3058
rect 66352 2994 66404 3000
rect 63500 2916 63552 2922
rect 64340 2910 64552 2938
rect 65168 2930 65472 2958
rect 63500 2858 63552 2864
rect 64524 2854 64552 2910
rect 65064 2916 65116 2922
rect 65064 2858 65116 2864
rect 64420 2848 64472 2854
rect 64420 2790 64472 2796
rect 64512 2848 64564 2854
rect 64512 2790 64564 2796
rect 65076 2802 65104 2858
rect 65444 2854 65472 2930
rect 66548 2922 66576 4000
rect 66824 3126 66852 4000
rect 66812 3120 66864 3126
rect 66812 3062 66864 3068
rect 67100 2990 67128 4000
rect 67180 3392 67232 3398
rect 67180 3334 67232 3340
rect 67192 3058 67220 3334
rect 67376 3058 67404 4000
rect 69054 3834 69154 3856
rect 69054 3782 69078 3834
rect 69130 3782 69154 3834
rect 67456 3596 67508 3602
rect 67456 3538 67508 3544
rect 67180 3052 67232 3058
rect 67180 2994 67232 3000
rect 67364 3052 67416 3058
rect 67364 2994 67416 3000
rect 67088 2984 67140 2990
rect 67088 2926 67140 2932
rect 67468 2922 67496 3538
rect 67732 3460 67784 3466
rect 67732 3402 67784 3408
rect 67744 2922 67772 3402
rect 68008 3188 68060 3194
rect 68008 3130 68060 3136
rect 68020 2922 68048 3130
rect 66536 2916 66588 2922
rect 66536 2858 66588 2864
rect 67456 2916 67508 2922
rect 67456 2858 67508 2864
rect 67732 2916 67784 2922
rect 67732 2858 67784 2864
rect 68008 2916 68060 2922
rect 68008 2858 68060 2864
rect 65248 2848 65300 2854
rect 65076 2796 65248 2802
rect 65076 2790 65300 2796
rect 65432 2848 65484 2854
rect 65432 2790 65484 2796
rect 64432 2582 64460 2790
rect 65076 2774 65288 2790
rect 69054 2746 69154 3782
rect 69054 2694 69078 2746
rect 69130 2694 69154 2746
rect 64420 2576 64472 2582
rect 64420 2518 64472 2524
rect 63054 2150 63078 2202
rect 63130 2150 63154 2202
rect 57428 1760 57480 1766
rect 57428 1702 57480 1708
rect 57054 1606 57078 1658
rect 57130 1606 57154 1658
rect 54668 1352 54720 1358
rect 54668 1294 54720 1300
rect 54944 1352 54996 1358
rect 54944 1294 54996 1300
rect 55220 1352 55272 1358
rect 55220 1294 55272 1300
rect 55496 1352 55548 1358
rect 55496 1294 55548 1300
rect 55772 1352 55824 1358
rect 55772 1294 55824 1300
rect 56048 1352 56100 1358
rect 56048 1294 56100 1300
rect 56324 1352 56376 1358
rect 56324 1294 56376 1300
rect 56600 1352 56652 1358
rect 56600 1294 56652 1300
rect 56876 1352 56928 1358
rect 56876 1294 56928 1300
rect 54680 1000 54708 1294
rect 54956 1000 54984 1294
rect 55232 1000 55260 1294
rect 55508 1000 55536 1294
rect 55784 1000 55812 1294
rect 56060 1000 56088 1294
rect 56336 1000 56364 1294
rect 56612 1000 56640 1294
rect 56888 1000 56916 1294
rect 57054 1040 57154 1606
rect 57336 1352 57388 1358
rect 57336 1294 57388 1300
rect 51078 870 51304 898
rect 51078 0 51134 870
rect 51354 0 51410 1000
rect 51630 0 51686 1000
rect 51906 0 51962 1000
rect 52182 0 52238 1000
rect 52458 0 52514 1000
rect 52734 0 52790 1000
rect 53010 0 53066 1000
rect 53286 0 53342 1000
rect 53562 0 53618 1000
rect 53838 0 53894 1000
rect 54114 0 54170 1000
rect 54390 0 54446 1000
rect 54666 0 54722 1000
rect 54942 0 54998 1000
rect 55218 0 55274 1000
rect 55494 0 55550 1000
rect 55770 0 55826 1000
rect 56046 0 56102 1000
rect 56322 0 56378 1000
rect 56598 0 56654 1000
rect 56874 0 56930 1000
rect 57150 898 57206 1000
rect 57348 898 57376 1294
rect 57440 1000 57468 1702
rect 59912 1488 59964 1494
rect 59912 1430 59964 1436
rect 60740 1488 60792 1494
rect 60740 1430 60792 1436
rect 61292 1488 61344 1494
rect 61292 1430 61344 1436
rect 61844 1488 61896 1494
rect 61844 1430 61896 1436
rect 57704 1352 57756 1358
rect 57704 1294 57756 1300
rect 57980 1352 58032 1358
rect 57980 1294 58032 1300
rect 58256 1352 58308 1358
rect 58256 1294 58308 1300
rect 58532 1352 58584 1358
rect 58532 1294 58584 1300
rect 58808 1352 58860 1358
rect 58808 1294 58860 1300
rect 59084 1352 59136 1358
rect 59084 1294 59136 1300
rect 59360 1352 59412 1358
rect 59360 1294 59412 1300
rect 59636 1352 59688 1358
rect 59636 1294 59688 1300
rect 57716 1000 57744 1294
rect 57992 1000 58020 1294
rect 58268 1000 58296 1294
rect 58544 1000 58572 1294
rect 58820 1000 58848 1294
rect 59096 1000 59124 1294
rect 59372 1000 59400 1294
rect 59648 1000 59676 1294
rect 59924 1000 59952 1430
rect 60280 1352 60332 1358
rect 60200 1312 60280 1340
rect 60200 1000 60228 1312
rect 60556 1352 60608 1358
rect 60280 1294 60332 1300
rect 60476 1312 60556 1340
rect 60476 1000 60504 1312
rect 60556 1294 60608 1300
rect 60752 1000 60780 1430
rect 61016 1352 61068 1358
rect 61016 1294 61068 1300
rect 61028 1000 61056 1294
rect 61304 1000 61332 1430
rect 61568 1352 61620 1358
rect 61568 1294 61620 1300
rect 61580 1000 61608 1294
rect 61856 1000 61884 1430
rect 62396 1420 62448 1426
rect 62396 1362 62448 1368
rect 62948 1420 63000 1426
rect 62948 1362 63000 1368
rect 62120 1352 62172 1358
rect 62120 1294 62172 1300
rect 62132 1000 62160 1294
rect 62408 1000 62436 1362
rect 62672 1352 62724 1358
rect 62672 1294 62724 1300
rect 62684 1000 62712 1294
rect 62960 1000 62988 1362
rect 63054 1268 63154 2150
rect 69054 2348 69154 2694
rect 69054 2292 69076 2348
rect 69132 2292 69154 2348
rect 63500 1760 63552 1766
rect 63500 1702 63552 1708
rect 67640 1760 67692 1766
rect 67640 1702 67692 1708
rect 63224 1352 63276 1358
rect 63224 1294 63276 1300
rect 63054 1212 63076 1268
rect 63132 1212 63154 1268
rect 63054 1114 63154 1212
rect 63054 1062 63078 1114
rect 63130 1062 63154 1114
rect 63054 1040 63154 1062
rect 63236 1000 63264 1294
rect 63512 1000 63540 1702
rect 64604 1488 64656 1494
rect 64604 1430 64656 1436
rect 65708 1488 65760 1494
rect 65708 1430 65760 1436
rect 66536 1488 66588 1494
rect 66536 1430 66588 1436
rect 64052 1420 64104 1426
rect 64052 1362 64104 1368
rect 63776 1352 63828 1358
rect 63776 1294 63828 1300
rect 63788 1000 63816 1294
rect 64064 1000 64092 1362
rect 64328 1352 64380 1358
rect 64328 1294 64380 1300
rect 64340 1000 64368 1294
rect 64616 1000 64644 1430
rect 65432 1420 65484 1426
rect 65432 1362 65484 1368
rect 65156 1352 65208 1358
rect 65156 1294 65208 1300
rect 64880 1284 64932 1290
rect 64880 1226 64932 1232
rect 64892 1000 64920 1226
rect 65168 1000 65196 1294
rect 65444 1000 65472 1362
rect 65720 1000 65748 1430
rect 66260 1420 66312 1426
rect 66260 1362 66312 1368
rect 65984 1352 66036 1358
rect 65984 1294 66036 1300
rect 65996 1000 66024 1294
rect 66272 1000 66300 1362
rect 66548 1000 66576 1430
rect 67364 1420 67416 1426
rect 67364 1362 67416 1368
rect 66812 1352 66864 1358
rect 66812 1294 66864 1300
rect 66824 1000 66852 1294
rect 67088 1284 67140 1290
rect 67088 1226 67140 1232
rect 67100 1000 67128 1226
rect 67376 1000 67404 1362
rect 67652 1000 67680 1702
rect 69054 1658 69154 2292
rect 69204 1760 69256 1766
rect 69204 1702 69256 1708
rect 69054 1606 69078 1658
rect 69130 1606 69154 1658
rect 67916 1488 67968 1494
rect 67916 1430 67968 1436
rect 68744 1488 68796 1494
rect 68744 1430 68796 1436
rect 67928 1000 67956 1430
rect 68284 1352 68336 1358
rect 68204 1312 68284 1340
rect 68204 1000 68232 1312
rect 68284 1294 68336 1300
rect 68468 1284 68520 1290
rect 68468 1226 68520 1232
rect 68480 1000 68508 1226
rect 68756 1000 68784 1430
rect 69054 1040 69154 1606
rect 57150 870 57376 898
rect 57150 0 57206 870
rect 57426 0 57482 1000
rect 57702 0 57758 1000
rect 57978 0 58034 1000
rect 58254 0 58310 1000
rect 58530 0 58586 1000
rect 58806 0 58862 1000
rect 59082 0 59138 1000
rect 59358 0 59414 1000
rect 59634 0 59690 1000
rect 59910 0 59966 1000
rect 60186 0 60242 1000
rect 60462 0 60518 1000
rect 60738 0 60794 1000
rect 61014 0 61070 1000
rect 61290 0 61346 1000
rect 61566 0 61622 1000
rect 61842 0 61898 1000
rect 62118 0 62174 1000
rect 62394 0 62450 1000
rect 62670 0 62726 1000
rect 62946 0 63002 1000
rect 63222 0 63278 1000
rect 63498 0 63554 1000
rect 63774 0 63830 1000
rect 64050 0 64106 1000
rect 64326 0 64382 1000
rect 64602 0 64658 1000
rect 64878 0 64934 1000
rect 65154 0 65210 1000
rect 65430 0 65486 1000
rect 65706 0 65762 1000
rect 65982 0 66038 1000
rect 66258 0 66314 1000
rect 66534 0 66590 1000
rect 66810 0 66866 1000
rect 67086 0 67142 1000
rect 67362 0 67418 1000
rect 67638 0 67694 1000
rect 67914 0 67970 1000
rect 68190 0 68246 1000
rect 68466 0 68522 1000
rect 68742 0 68798 1000
rect 69018 898 69074 1000
rect 69216 898 69244 1702
rect 69572 1488 69624 1494
rect 69572 1430 69624 1436
rect 69388 1352 69440 1358
rect 69308 1312 69388 1340
rect 69308 1000 69336 1312
rect 69388 1294 69440 1300
rect 69584 1000 69612 1430
rect 69848 1420 69900 1426
rect 69848 1362 69900 1368
rect 69860 1000 69888 1362
rect 69018 870 69244 898
rect 69018 0 69074 870
rect 69294 0 69350 1000
rect 69570 0 69626 1000
rect 69846 0 69902 1000
<< via2 >>
rect 2778 3712 2834 3768
rect 2502 3168 2558 3224
rect 3076 3372 3132 3428
rect 2962 2896 3018 2952
rect 2778 2508 2834 2544
rect 2778 2488 2780 2508
rect 2780 2488 2832 2508
rect 2832 2488 2834 2508
rect 2502 2080 2558 2136
rect 2226 1708 2228 1728
rect 2228 1708 2280 1728
rect 2280 1708 2282 1728
rect 2226 1672 2282 1708
rect 1674 1420 1730 1456
rect 1674 1400 1676 1420
rect 1676 1400 1728 1420
rect 1728 1400 1730 1420
rect 15076 3372 15132 3428
rect 9076 2292 9132 2348
rect 3076 1212 3132 1268
rect 25134 3032 25190 3088
rect 27076 3372 27132 3428
rect 26882 3052 26938 3088
rect 26882 3032 26884 3052
rect 26884 3032 26936 3052
rect 26936 3032 26938 3052
rect 26514 2896 26570 2952
rect 21076 2292 21132 2348
rect 15076 1212 15132 1268
rect 28538 2896 28594 2952
rect 39076 3372 39132 3428
rect 33076 2292 33132 2348
rect 27076 1212 27132 1268
rect 51076 3372 51132 3428
rect 45076 2292 45132 2348
rect 39076 1212 39132 1268
rect 63076 3372 63132 3428
rect 57076 2292 57132 2348
rect 51076 1212 51132 1268
rect 69076 2292 69132 2348
rect 63076 1212 63132 1268
<< metal3 >>
rect 0 3770 1000 3800
rect 2773 3770 2839 3773
rect 0 3768 2839 3770
rect 0 3712 2778 3768
rect 2834 3712 2839 3768
rect 0 3710 2839 3712
rect 0 3680 1000 3710
rect 2773 3707 2839 3710
rect 1104 3428 72864 3450
rect 0 3362 1000 3392
rect 1104 3372 3076 3428
rect 3132 3372 15076 3428
rect 15132 3372 27076 3428
rect 27132 3372 39076 3428
rect 39132 3372 51076 3428
rect 51132 3372 63076 3428
rect 63132 3372 72864 3428
rect 0 3272 1042 3362
rect 1104 3350 72864 3372
rect 982 3226 1042 3272
rect 2497 3226 2563 3229
rect 982 3224 2563 3226
rect 982 3168 2502 3224
rect 2558 3168 2563 3224
rect 982 3166 2563 3168
rect 2497 3163 2563 3166
rect 25129 3090 25195 3093
rect 26877 3090 26943 3093
rect 25129 3088 26943 3090
rect 25129 3032 25134 3088
rect 25190 3032 26882 3088
rect 26938 3032 26943 3088
rect 25129 3030 26943 3032
rect 25129 3027 25195 3030
rect 26877 3027 26943 3030
rect 0 2954 1000 2984
rect 2957 2954 3023 2957
rect 0 2952 3023 2954
rect 0 2896 2962 2952
rect 3018 2896 3023 2952
rect 0 2894 3023 2896
rect 0 2864 1000 2894
rect 2957 2891 3023 2894
rect 26509 2954 26575 2957
rect 28533 2954 28599 2957
rect 26509 2952 28599 2954
rect 26509 2896 26514 2952
rect 26570 2896 28538 2952
rect 28594 2896 28599 2952
rect 26509 2894 28599 2896
rect 26509 2891 26575 2894
rect 28533 2891 28599 2894
rect 0 2546 1000 2576
rect 2773 2546 2839 2549
rect 0 2544 2839 2546
rect 0 2488 2778 2544
rect 2834 2488 2839 2544
rect 0 2486 2839 2488
rect 0 2456 1000 2486
rect 2773 2483 2839 2486
rect 1104 2348 72864 2370
rect 1104 2292 9076 2348
rect 9132 2292 21076 2348
rect 21132 2292 33076 2348
rect 33132 2292 45076 2348
rect 45132 2292 57076 2348
rect 57132 2292 69076 2348
rect 69132 2292 72864 2348
rect 1104 2270 72864 2292
rect 0 2138 1000 2168
rect 2497 2138 2563 2141
rect 0 2136 2563 2138
rect 0 2080 2502 2136
rect 2558 2080 2563 2136
rect 0 2078 2563 2080
rect 0 2048 1000 2078
rect 2497 2075 2563 2078
rect 0 1730 1000 1760
rect 2221 1730 2287 1733
rect 0 1728 2287 1730
rect 0 1672 2226 1728
rect 2282 1672 2287 1728
rect 0 1670 2287 1672
rect 0 1640 1000 1670
rect 2221 1667 2287 1670
rect 1669 1458 1735 1461
rect 982 1456 1735 1458
rect 982 1400 1674 1456
rect 1730 1400 1735 1456
rect 982 1398 1735 1400
rect 982 1352 1042 1398
rect 1669 1395 1735 1398
rect 0 1262 1042 1352
rect 1104 1268 72864 1290
rect 0 1232 1000 1262
rect 1104 1212 3076 1268
rect 3132 1212 15076 1268
rect 15132 1212 27076 1268
rect 27132 1212 39076 1268
rect 39132 1212 51076 1268
rect 51132 1212 63076 1268
rect 63132 1212 72864 1268
rect 1104 1190 72864 1212
use sky130_fd_sc_hd__conb_1  insts\[174\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 2208 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[183\]
timestamp 1618914159
transform -1 0 2208 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[205\]
timestamp 1618914159
transform 1 0 1656 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[206\]
timestamp 1618914159
transform 1 0 2208 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 1104 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1618914159
transform 1 0 1104 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3
timestamp 1618914159
transform 1 0 1380 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 1380 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 2116 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[103\]
timestamp 1618914159
transform 1 0 2484 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[114\]
timestamp 1618914159
transform 1 0 2760 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[121\]
timestamp 1618914159
transform 1 0 3036 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[158\]
timestamp 1618914159
transform 1 0 3312 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[15\]
timestamp 1618914159
transform 1 0 2484 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[181\]
timestamp 1618914159
transform 1 0 2852 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[196\]
timestamp 1618914159
transform 1 0 3128 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[19\]
timestamp 1618914159
transform 1 0 3404 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_18
timestamp 1618914159
transform 1 0 2760 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[141\]
timestamp 1618914159
transform 1 0 3864 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[163\]
timestamp 1618914159
transform 1 0 4140 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[165\]
timestamp 1618914159
transform 1 0 4416 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[167\]
timestamp 1618914159
transform 1 0 4048 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 3772 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 3588 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 3680 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_35 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[117\]
timestamp 1618914159
transform 1 0 5612 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[132\]
timestamp 1618914159
transform 1 0 5060 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[143\]
timestamp 1618914159
transform 1 0 4692 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[176\]
timestamp 1618914159
transform 1 0 5336 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42
timestamp 1618914159
transform 1 0 4968 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_47
timestamp 1618914159
transform 1 0 5428 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[110\]
timestamp 1618914159
transform 1 0 6164 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[139\]
timestamp 1618914159
transform 1 0 6808 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[172\]
timestamp 1618914159
transform 1 0 6532 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[187\]
timestamp 1618914159
transform 1 0 6992 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[192\]
timestamp 1618914159
transform 1 0 5888 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_11
timestamp 1618914159
transform 1 0 6440 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_36
timestamp 1618914159
transform 1 0 6348 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_55
timestamp 1618914159
transform 1 0 6164 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_58 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 6440 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  insts\[125\]
timestamp 1618914159
transform 1 0 7268 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[138\]
timestamp 1618914159
transform 1 0 7544 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[152\]
timestamp 1618914159
transform 1 0 7820 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[17\]
timestamp 1618914159
transform 1 0 8096 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65
timestamp 1618914159
transform 1 0 7084 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_67
timestamp 1618914159
transform 1 0 7268 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82
timestamp 1618914159
transform 1 0 8648 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[14\]
timestamp 1618914159
transform 1 0 8372 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[106\]
timestamp 1618914159
transform 1 0 8740 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88
timestamp 1618914159
transform 1 0 9200 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86
timestamp 1618914159
transform 1 0 9016 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_12
timestamp 1618914159
transform 1 0 9108 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[189\]
timestamp 1618914159
transform 1 0 8924 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[155\]
timestamp 1618914159
transform 1 0 9292 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_88
timestamp 1618914159
transform 1 0 9200 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_79
timestamp 1618914159
transform 1 0 8372 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  insts\[109\]
timestamp 1618914159
transform 1 0 10304 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[157\]
timestamp 1618914159
transform 1 0 9568 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[160\]
timestamp 1618914159
transform 1 0 10028 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[198\]
timestamp 1618914159
transform 1 0 9844 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_95
timestamp 1618914159
transform 1 0 9844 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_94
timestamp 1618914159
transform 1 0 9752 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1618914159
transform 1 0 10120 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[102\]
timestamp 1618914159
transform 1 0 10580 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[133\]
timestamp 1618914159
transform 1 0 11224 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[166\]
timestamp 1618914159
transform 1 0 10948 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[16\]
timestamp 1618914159
transform 1 0 11500 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_37
timestamp 1618914159
transform 1 0 11592 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106
timestamp 1618914159
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_110
timestamp 1618914159
transform 1 0 11224 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_115
timestamp 1618914159
transform 1 0 11684 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[119\]
timestamp 1618914159
transform 1 0 12236 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[122\]
timestamp 1618914159
transform 1 0 11868 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[124\]
timestamp 1618914159
transform 1 0 12696 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[173\]
timestamp 1618914159
transform 1 0 11868 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_13
timestamp 1618914159
transform 1 0 11776 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120
timestamp 1618914159
transform 1 0 12144 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_124
timestamp 1618914159
transform 1 0 12512 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_120
timestamp 1618914159
transform 1 0 12144 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[135\]
timestamp 1618914159
transform 1 0 13800 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[154\]
timestamp 1618914159
transform 1 0 12972 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[170\]
timestamp 1618914159
transform 1 0 13524 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[177\]
timestamp 1618914159
transform 1 0 13248 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[188\]
timestamp 1618914159
transform 1 0 14076 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[202\]
timestamp 1618914159
transform 1 0 13248 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1618914159
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[116\]
timestamp 1618914159
transform 1 0 14904 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[178\]
timestamp 1618914159
transform 1 0 14536 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[191\]
timestamp 1618914159
transform 1 0 15180 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[195\]
timestamp 1618914159
transform 1 0 15180 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_14
timestamp 1618914159
transform 1 0 14444 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_144
timestamp 1618914159
transform 1 0 14352 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149
timestamp 1618914159
transform 1 0 14812 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_147
timestamp 1618914159
transform 1 0 14628 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  insts\[128\]
timestamp 1618914159
transform 1 0 15824 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[151\]
timestamp 1618914159
transform 1 0 15548 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[184\]
timestamp 1618914159
transform 1 0 16284 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[1\]
timestamp 1618914159
transform 1 0 16100 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156
timestamp 1618914159
transform 1 0 15456 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_163
timestamp 1618914159
transform 1 0 16100 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_156
timestamp 1618914159
transform 1 0 15456 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_162
timestamp 1618914159
transform 1 0 16008 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_166
timestamp 1618914159
transform 1 0 16376 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  insts\[147\]
timestamp 1618914159
transform 1 0 17204 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[149\]
timestamp 1618914159
transform 1 0 17480 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[162\]
timestamp 1618914159
transform 1 0 16560 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[169\]
timestamp 1618914159
transform 1 0 16836 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_15
timestamp 1618914159
transform 1 0 17112 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_38
timestamp 1618914159
transform 1 0 16836 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_170
timestamp 1618914159
transform 1 0 16744 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_172
timestamp 1618914159
transform 1 0 16928 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[10\]
timestamp 1618914159
transform 1 0 17756 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[112\]
timestamp 1618914159
transform 1 0 18032 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[118\]
timestamp 1618914159
transform 1 0 18584 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[12\]
timestamp 1618914159
transform 1 0 18308 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1618914159
transform 1 0 18032 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[120\]
timestamp 1618914159
transform 1 0 18860 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[126\]
timestamp 1618914159
transform 1 0 19412 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[129\]
timestamp 1618914159
transform 1 0 19872 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[146\]
timestamp 1618914159
transform 1 0 19136 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_16
timestamp 1618914159
transform 1 0 19780 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_202
timestamp 1618914159
transform 1 0 19688 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1618914159
transform 1 0 19136 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[131\]
timestamp 1618914159
transform 1 0 20148 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[137\]
timestamp 1618914159
transform 1 0 20884 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[142\]
timestamp 1618914159
transform 1 0 21160 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[194\]
timestamp 1618914159
transform 1 0 20608 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[201\]
timestamp 1618914159
transform 1 0 20332 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_210
timestamp 1618914159
transform 1 0 20424 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_208
timestamp 1618914159
transform 1 0 20240 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_212
timestamp 1618914159
transform 1 0 20608 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[100\]
timestamp 1618914159
transform 1 0 21436 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[13\]
timestamp 1618914159
transform 1 0 21712 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[150\]
timestamp 1618914159
transform 1 0 22080 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_39
timestamp 1618914159
transform 1 0 22080 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_227
timestamp 1618914159
transform 1 0 21988 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_231
timestamp 1618914159
transform 1 0 22356 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_224
timestamp 1618914159
transform 1 0 21712 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_229
timestamp 1618914159
transform 1 0 22172 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[153\]
timestamp 1618914159
transform 1 0 22540 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[156\]
timestamp 1618914159
transform 1 0 22816 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[159\]
timestamp 1618914159
transform 1 0 23092 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[161\]
timestamp 1618914159
transform 1 0 23368 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_17
timestamp 1618914159
transform 1 0 22448 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_241
timestamp 1618914159
transform 1 0 23276 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[148\]
timestamp 1618914159
transform 1 0 23736 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[164\]
timestamp 1618914159
transform 1 0 24012 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[171\]
timestamp 1618914159
transform 1 0 24288 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[175\]
timestamp 1618914159
transform 1 0 24564 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_245
timestamp 1618914159
transform 1 0 23644 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_253
timestamp 1618914159
transform 1 0 24380 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[179\]
timestamp 1618914159
transform 1 0 24840 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[182\]
timestamp 1618914159
transform 1 0 25208 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[186\]
timestamp 1618914159
transform 1 0 25484 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[18\]
timestamp 1618914159
transform 1 0 25760 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_18
timestamp 1618914159
transform 1 0 25116 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_265
timestamp 1618914159
transform 1 0 25484 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[104\]
timestamp 1618914159
transform 1 0 26956 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[193\]
timestamp 1618914159
transform 1 0 26036 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[197\]
timestamp 1618914159
transform 1 0 26312 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[200\]
timestamp 1618914159
transform 1 0 26588 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[203\]
timestamp 1618914159
transform 1 0 26680 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_280
timestamp 1618914159
transform 1 0 26864 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_277
timestamp 1618914159
transform 1 0 26588 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1618914159
transform 1 0 26956 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  insts\[108\]
timestamp 1618914159
transform 1 0 27324 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[111\]
timestamp 1618914159
transform 1 0 27876 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[115\]
timestamp 1618914159
transform 1 0 28152 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_19
timestamp 1618914159
transform 1 0 27784 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_40
timestamp 1618914159
transform 1 0 27324 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_284
timestamp 1618914159
transform 1 0 27232 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_288
timestamp 1618914159
transform 1 0 27600 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_286
timestamp 1618914159
transform 1 0 27416 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[113\]
timestamp 1618914159
transform 1 0 28428 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[11\]
timestamp 1618914159
transform 1 0 28704 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[127\]
timestamp 1618914159
transform 1 0 28980 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[130\]
timestamp 1618914159
transform 1 0 29256 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_298
timestamp 1618914159
transform 1 0 28520 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[134\]
timestamp 1618914159
transform 1 0 29532 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[140\]
timestamp 1618914159
transform 1 0 29808 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[144\]
timestamp 1618914159
transform 1 0 30084 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[168\]
timestamp 1618914159
transform 1 0 30544 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_20
timestamp 1618914159
transform 1 0 30452 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_318
timestamp 1618914159
transform 1 0 30360 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_310
timestamp 1618914159
transform 1 0 29624 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[101\]
timestamp 1618914159
transform 1 0 31280 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[123\]
timestamp 1618914159
transform 1 0 31556 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[180\]
timestamp 1618914159
transform 1 0 30820 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[190\]
timestamp 1618914159
transform 1 0 30728 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[199\]
timestamp 1618914159
transform 1 0 31004 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_326
timestamp 1618914159
transform 1 0 31096 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_328
timestamp 1618914159
transform 1 0 31280 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[105\]
timestamp 1618914159
transform 1 0 32844 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[107\]
timestamp 1618914159
transform 1 0 32568 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[136\]
timestamp 1618914159
transform 1 0 31832 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[145\]
timestamp 1618914159
transform 1 0 32108 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[185\]
timestamp 1618914159
transform 1 0 32660 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_41
timestamp 1618914159
transform 1 0 32568 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_340
timestamp 1618914159
transform 1 0 32384 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_340
timestamp 1618914159
transform 1 0 32384 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_346
timestamp 1618914159
transform 1 0 32936 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[0\]
timestamp 1618914159
transform 1 0 33212 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_21
timestamp 1618914159
transform 1 0 33120 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_352
timestamp 1618914159
transform 1 0 33488 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_358
timestamp 1618914159
transform 1 0 34040 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_364
timestamp 1618914159
transform 1 0 34592 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_370
timestamp 1618914159
transform 1 0 35144 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_22
timestamp 1618914159
transform 1 0 35788 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_376
timestamp 1618914159
transform 1 0 35696 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_378
timestamp 1618914159
transform 1 0 35880 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_382
timestamp 1618914159
transform 1 0 36248 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[383\]
timestamp 1618914159
transform -1 0 37904 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_390
timestamp 1618914159
transform 1 0 36984 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_396
timestamp 1618914159
transform 1 0 37536 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_394
timestamp 1618914159
transform 1 0 37352 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_404
timestamp 1618914159
transform 1 0 38272 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_400
timestamp 1618914159
transform 1 0 37904 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_398
timestamp 1618914159
transform 1 0 37720 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_42
timestamp 1618914159
transform 1 0 37812 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[323\]
timestamp 1618914159
transform -1 0 38456 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[312\]
timestamp 1618914159
transform -1 0 38180 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_407
timestamp 1618914159
transform 1 0 38548 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_23
timestamp 1618914159
transform 1 0 38456 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[404\]
timestamp 1618914159
transform -1 0 38640 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[330\]
timestamp 1618914159
transform -1 0 38916 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_408
timestamp 1618914159
transform 1 0 38640 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[367\]
timestamp 1618914159
transform -1 0 39192 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[369\]
timestamp 1618914159
transform -1 0 39468 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[390\]
timestamp 1618914159
transform -1 0 40020 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[392\]
timestamp 1618914159
transform -1 0 39744 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[408\]
timestamp 1618914159
transform -1 0 40296 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_420
timestamp 1618914159
transform 1 0 39744 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[350\]
timestamp 1618914159
transform -1 0 40848 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[372\]
timestamp 1618914159
transform -1 0 40572 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[374\]
timestamp 1618914159
transform -1 0 41492 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[376\]
timestamp 1618914159
transform -1 0 41124 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_24
timestamp 1618914159
transform 1 0 41124 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_432
timestamp 1618914159
transform 1 0 40848 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[326\]
timestamp 1618914159
transform -1 0 42596 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[341\]
timestamp 1618914159
transform -1 0 42044 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[352\]
timestamp 1618914159
transform -1 0 41768 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[385\]
timestamp 1618914159
transform -1 0 42320 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_444
timestamp 1618914159
transform 1 0 41952 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[31\]
timestamp 1618914159
transform -1 0 43148 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[348\]
timestamp 1618914159
transform -1 0 43792 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[381\]
timestamp 1618914159
transform -1 0 43424 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[400\]
timestamp 1618914159
transform -1 0 42872 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_43
timestamp 1618914159
transform 1 0 43056 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_460
timestamp 1618914159
transform 1 0 43424 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_457
timestamp 1618914159
transform 1 0 43148 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  insts\[334\]
timestamp 1618914159
transform -1 0 44344 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[347\]
timestamp 1618914159
transform -1 0 44620 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[361\]
timestamp 1618914159
transform -1 0 44896 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[396\]
timestamp 1618914159
transform -1 0 44068 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_25
timestamp 1618914159
transform 1 0 43792 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_465
timestamp 1618914159
transform 1 0 43884 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_463
timestamp 1618914159
transform 1 0 43700 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_467
timestamp 1618914159
transform 1 0 44068 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[315\]
timestamp 1618914159
transform -1 0 45724 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[359\]
timestamp 1618914159
transform -1 0 45448 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[389\]
timestamp 1618914159
transform -1 0 45172 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[398\]
timestamp 1618914159
transform -1 0 46000 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_479
timestamp 1618914159
transform 1 0 45172 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_491
timestamp 1618914159
transform 1 0 46276 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_492
timestamp 1618914159
transform 1 0 46368 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_488
timestamp 1618914159
transform 1 0 46000 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_26
timestamp 1618914159
transform 1 0 46460 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[366\]
timestamp 1618914159
transform -1 0 46828 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[364\]
timestamp 1618914159
transform -1 0 46368 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_497
timestamp 1618914159
transform 1 0 46828 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[406\]
timestamp 1618914159
transform -1 0 46920 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[36\]
timestamp 1618914159
transform -1 0 47196 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_498
timestamp 1618914159
transform 1 0 46920 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[311\]
timestamp 1618914159
transform -1 0 47748 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[318\]
timestamp 1618914159
transform -1 0 47472 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[342\]
timestamp 1618914159
transform -1 0 48300 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[375\]
timestamp 1618914159
transform -1 0 48024 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_44
timestamp 1618914159
transform 1 0 48300 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_513
timestamp 1618914159
transform 1 0 48300 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_510
timestamp 1618914159
transform 1 0 48024 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[328\]
timestamp 1618914159
transform -1 0 49496 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[331\]
timestamp 1618914159
transform -1 0 48944 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[379\]
timestamp 1618914159
transform -1 0 48668 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[382\]
timestamp 1618914159
transform 1 0 49496 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_27
timestamp 1618914159
transform 1 0 49128 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_520
timestamp 1618914159
transform 1 0 48944 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_514
timestamp 1618914159
transform 1 0 48392 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_526
timestamp 1618914159
transform 1 0 49496 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[333\]
timestamp 1618914159
transform -1 0 50048 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[363\]
timestamp 1618914159
transform -1 0 50324 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[37\]
timestamp 1618914159
transform -1 0 50968 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[386\]
timestamp 1618914159
transform 1 0 50324 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[411\]
timestamp 1618914159
transform -1 0 50600 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_538
timestamp 1618914159
transform 1 0 50600 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_534
timestamp 1618914159
transform 1 0 50232 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_538
timestamp 1618914159
transform 1 0 50600 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[344\]
timestamp 1618914159
transform -1 0 51244 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[387\]
timestamp 1618914159
transform -1 0 51796 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[397\]
timestamp 1618914159
transform -1 0 51520 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_28
timestamp 1618914159
transform 1 0 51796 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_550
timestamp 1618914159
transform 1 0 51704 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  insts\[325\]
timestamp 1618914159
transform -1 0 52348 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[337\]
timestamp 1618914159
transform 1 0 52992 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[360\]
timestamp 1618914159
transform -1 0 52900 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[3\]
timestamp 1618914159
transform 1 0 52348 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[403\]
timestamp 1618914159
transform -1 0 52624 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_552
timestamp 1618914159
transform 1 0 51888 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_563
timestamp 1618914159
transform 1 0 52900 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_556
timestamp 1618914159
transform 1 0 52256 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_560
timestamp 1618914159
transform 1 0 52624 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[356\]
timestamp 1618914159
transform 1 0 54096 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[371\]
timestamp 1618914159
transform 1 0 53820 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[393\]
timestamp 1618914159
transform 1 0 53544 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[409\]
timestamp 1618914159
transform 1 0 53268 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_45
timestamp 1618914159
transform 1 0 53544 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_568
timestamp 1618914159
transform 1 0 53360 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_571
timestamp 1618914159
transform 1 0 53636 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[319\]
timestamp 1618914159
transform 1 0 54924 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[321\]
timestamp 1618914159
transform 1 0 55200 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[358\]
timestamp 1618914159
transform 1 0 54648 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[378\]
timestamp 1618914159
transform 1 0 54372 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_29
timestamp 1618914159
transform 1 0 54464 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_579
timestamp 1618914159
transform 1 0 54372 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_581
timestamp 1618914159
transform 1 0 54556 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_582
timestamp 1618914159
transform 1 0 54648 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[327\]
timestamp 1618914159
transform 1 0 55844 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[32\]
timestamp 1618914159
transform 1 0 56120 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[339\]
timestamp 1618914159
transform 1 0 55568 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[355\]
timestamp 1618914159
transform 1 0 56396 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_591
timestamp 1618914159
transform 1 0 55476 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_594
timestamp 1618914159
transform 1 0 55752 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_607
timestamp 1618914159
transform 1 0 56948 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_30
timestamp 1618914159
transform 1 0 57132 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[335\]
timestamp 1618914159
transform 1 0 56672 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_612
timestamp 1618914159
transform 1 0 57408 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[410\]
timestamp 1618914159
transform 1 0 57500 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[402\]
timestamp 1618914159
transform 1 0 57776 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[340\]
timestamp 1618914159
transform 1 0 57500 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[338\]
timestamp 1618914159
transform 1 0 57224 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_616
timestamp 1618914159
transform 1 0 57776 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_606
timestamp 1618914159
transform 1 0 56856 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  insts\[30\]
timestamp 1618914159
transform 1 0 58696 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[346\]
timestamp 1618914159
transform 1 0 58052 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[349\]
timestamp 1618914159
transform 1 0 58972 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[351\]
timestamp 1618914159
transform 1 0 58420 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46
timestamp 1618914159
transform 1 0 58788 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_622
timestamp 1618914159
transform 1 0 58328 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_624
timestamp 1618914159
transform 1 0 58512 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_628
timestamp 1618914159
transform 1 0 58880 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[35\]
timestamp 1618914159
transform 1 0 59248 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[362\]
timestamp 1618914159
transform 1 0 59524 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[365\]
timestamp 1618914159
transform 1 0 59892 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_31
timestamp 1618914159
transform 1 0 59800 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_640
timestamp 1618914159
transform 1 0 59984 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[357\]
timestamp 1618914159
transform 1 0 60996 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[368\]
timestamp 1618914159
transform 1 0 60168 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[370\]
timestamp 1618914159
transform 1 0 60444 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[373\]
timestamp 1618914159
transform 1 0 60720 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[380\]
timestamp 1618914159
transform 1 0 61272 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_652
timestamp 1618914159
transform 1 0 61088 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[384\]
timestamp 1618914159
transform 1 0 61548 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[388\]
timestamp 1618914159
transform 1 0 61824 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[391\]
timestamp 1618914159
transform 1 0 62100 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_32
timestamp 1618914159
transform 1 0 62468 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_666
timestamp 1618914159
transform 1 0 62376 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_664
timestamp 1618914159
transform 1 0 62192 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[395\]
timestamp 1618914159
transform 1 0 62560 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[399\]
timestamp 1618914159
transform 1 0 62836 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[401\]
timestamp 1618914159
transform 1 0 63112 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[405\]
timestamp 1618914159
transform 1 0 63388 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[40\]
timestamp 1618914159
transform 1 0 63664 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_676
timestamp 1618914159
transform 1 0 63296 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[313\]
timestamp 1618914159
transform 1 0 64124 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[317\]
timestamp 1618914159
transform 1 0 64400 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[320\]
timestamp 1618914159
transform 1 0 64676 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[412\]
timestamp 1618914159
transform 1 0 64124 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1618914159
transform 1 0 64032 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_683
timestamp 1618914159
transform 1 0 63940 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_688
timestamp 1618914159
transform 1 0 64400 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[322\]
timestamp 1618914159
transform 1 0 65596 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[324\]
timestamp 1618914159
transform 1 0 65228 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[329\]
timestamp 1618914159
transform 1 0 65872 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_33
timestamp 1618914159
transform 1 0 65136 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_694
timestamp 1618914159
transform 1 0 64952 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_700
timestamp 1618914159
transform 1 0 65504 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_700
timestamp 1618914159
transform 1 0 65504 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[336\]
timestamp 1618914159
transform 1 0 66148 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[33\]
timestamp 1618914159
transform 1 0 66424 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[343\]
timestamp 1618914159
transform 1 0 66700 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[34\]
timestamp 1618914159
transform 1 0 66976 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_712
timestamp 1618914159
transform 1 0 66608 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[353\]
timestamp 1618914159
transform 1 0 67252 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[377\]
timestamp 1618914159
transform 1 0 67528 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[38\]
timestamp 1618914159
transform 1 0 67896 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[39\]
timestamp 1618914159
transform 1 0 68172 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[407\]
timestamp 1618914159
transform 1 0 68172 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_34
timestamp 1618914159
transform 1 0 67804 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_724
timestamp 1618914159
transform 1 0 67712 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_728
timestamp 1618914159
transform 1 0 68080 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[345\]
timestamp 1618914159
transform 1 0 69000 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[332\]
timestamp 1618914159
transform 1 0 68724 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[310\]
timestamp 1618914159
transform 1 0 68448 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_742
timestamp 1618914159
transform 1 0 69368 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_740
timestamp 1618914159
transform 1 0 69184 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_744
timestamp 1618914159
transform 1 0 69552 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1618914159
transform 1 0 69276 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[394\]
timestamp 1618914159
transform 1 0 69552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[354\]
timestamp 1618914159
transform 1 0 69276 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_732
timestamp 1618914159
transform 1 0 68448 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[309\]
timestamp 1618914159
transform 1 0 70564 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[314\]
timestamp 1618914159
transform 1 0 70012 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[316\]
timestamp 1618914159
transform 1 0 69736 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_35
timestamp 1618914159
transform 1 0 70472 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_752
timestamp 1618914159
transform 1 0 70288 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_747
timestamp 1618914159
transform 1 0 69828 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_758
timestamp 1618914159
transform 1 0 70840 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_770
timestamp 1618914159
transform 1 0 71944 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_759
timestamp 1618914159
transform 1 0 70932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1618914159
transform -1 0 72864 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1618914159
transform -1 0 72864 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_776
timestamp 1618914159
transform 1 0 72496 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_771
timestamp 1618914159
transform 1 0 72036 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1618914159
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1618914159
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[207\]
timestamp 1618914159
transform 1 0 2484 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[208\]
timestamp 1618914159
transform 1 0 2760 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[209\]
timestamp 1618914159
transform 1 0 3036 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1618914159
transform 1 0 3312 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1618914159
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_28
timestamp 1618914159
transform 1 0 3680 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_30
timestamp 1618914159
transform 1 0 3864 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_42
timestamp 1618914159
transform 1 0 4968 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_54
timestamp 1618914159
transform 1 0 6072 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_66
timestamp 1618914159
transform 1 0 7176 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1618914159
transform 1 0 9016 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_78
timestamp 1618914159
transform 1 0 8280 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_87
timestamp 1618914159
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_99
timestamp 1618914159
transform 1 0 10212 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_111
timestamp 1618914159
transform 1 0 11316 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1618914159
transform 1 0 12420 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_135
timestamp 1618914159
transform 1 0 13524 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1618914159
transform 1 0 14260 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_144
timestamp 1618914159
transform 1 0 14352 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_156
timestamp 1618914159
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_168
timestamp 1618914159
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_180
timestamp 1618914159
transform 1 0 17664 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_192
timestamp 1618914159
transform 1 0 18768 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1618914159
transform 1 0 19504 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_201
timestamp 1618914159
transform 1 0 19596 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_213
timestamp 1618914159
transform 1 0 20700 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_225
timestamp 1618914159
transform 1 0 21804 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_237
timestamp 1618914159
transform 1 0 22908 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_249
timestamp 1618914159
transform 1 0 24012 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1618914159
transform 1 0 24748 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_258
timestamp 1618914159
transform 1 0 24840 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_270
timestamp 1618914159
transform 1 0 25944 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_282
timestamp 1618914159
transform 1 0 27048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_294
timestamp 1618914159
transform 1 0 28152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_306
timestamp 1618914159
transform 1 0 29256 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1618914159
transform 1 0 29992 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_315
timestamp 1618914159
transform 1 0 30084 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_327
timestamp 1618914159
transform 1 0 31188 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_339
timestamp 1618914159
transform 1 0 32292 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_351
timestamp 1618914159
transform 1 0 33396 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1618914159
transform 1 0 35236 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_363
timestamp 1618914159
transform 1 0 34500 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_372
timestamp 1618914159
transform 1 0 35328 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_384
timestamp 1618914159
transform 1 0 36432 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_396
timestamp 1618914159
transform 1 0 37536 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_408
timestamp 1618914159
transform 1 0 38640 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_420
timestamp 1618914159
transform 1 0 39744 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1618914159
transform 1 0 40480 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_429
timestamp 1618914159
transform 1 0 40572 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_441
timestamp 1618914159
transform 1 0 41676 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_453
timestamp 1618914159
transform 1 0 42780 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_465
timestamp 1618914159
transform 1 0 43884 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1618914159
transform 1 0 45724 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_477
timestamp 1618914159
transform 1 0 44988 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_486
timestamp 1618914159
transform 1 0 45816 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_498
timestamp 1618914159
transform 1 0 46920 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_510
timestamp 1618914159
transform 1 0 48024 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_522
timestamp 1618914159
transform 1 0 49128 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_534
timestamp 1618914159
transform 1 0 50232 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1618914159
transform 1 0 50968 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_543
timestamp 1618914159
transform 1 0 51060 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_555
timestamp 1618914159
transform 1 0 52164 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_567
timestamp 1618914159
transform 1 0 53268 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_579
timestamp 1618914159
transform 1 0 54372 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1618914159
transform 1 0 56212 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_591
timestamp 1618914159
transform 1 0 55476 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_600
timestamp 1618914159
transform 1 0 56304 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_612
timestamp 1618914159
transform 1 0 57408 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_624
timestamp 1618914159
transform 1 0 58512 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_636
timestamp 1618914159
transform 1 0 59616 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_648
timestamp 1618914159
transform 1 0 60720 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1618914159
transform 1 0 61456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_657
timestamp 1618914159
transform 1 0 61548 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_669
timestamp 1618914159
transform 1 0 62652 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_681
timestamp 1618914159
transform 1 0 63756 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_693
timestamp 1618914159
transform 1 0 64860 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_705
timestamp 1618914159
transform 1 0 65964 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1618914159
transform 1 0 66700 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_714
timestamp 1618914159
transform 1 0 66792 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_726
timestamp 1618914159
transform 1 0 67896 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_738
timestamp 1618914159
transform 1 0 69000 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_750
timestamp 1618914159
transform 1 0 70104 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1618914159
transform 1 0 71944 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_762
timestamp 1618914159
transform 1 0 71208 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1618914159
transform -1 0 72864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_771
timestamp 1618914159
transform 1 0 72036 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  insts\[217\]
timestamp 1618914159
transform 1 0 2208 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[218\]
timestamp 1618914159
transform -1 0 2208 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1618914159
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1618914159
transform 1 0 1380 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  insts\[20\]
timestamp 1618914159
transform 1 0 2484 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[210\]
timestamp 1618914159
transform 1 0 2760 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[211\]
timestamp 1618914159
transform 1 0 3036 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[212\]
timestamp 1618914159
transform 1 0 3312 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[219\]
timestamp 1618914159
transform 1 0 3588 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[21\]
timestamp 1618914159
transform 1 0 3864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[220\]
timestamp 1618914159
transform 1 0 4140 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[221\]
timestamp 1618914159
transform 1 0 4416 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[222\]
timestamp 1618914159
transform 1 0 4692 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[223\]
timestamp 1618914159
transform 1 0 4968 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[224\]
timestamp 1618914159
transform 1 0 5244 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[225\]
timestamp 1618914159
transform 1 0 5520 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[226\]
timestamp 1618914159
transform 1 0 5796 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[227\]
timestamp 1618914159
transform 1 0 6072 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[228\]
timestamp 1618914159
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[229\]
timestamp 1618914159
transform 1 0 6716 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[22\]
timestamp 1618914159
transform 1 0 6992 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1618914159
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[230\]
timestamp 1618914159
transform 1 0 7268 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[231\]
timestamp 1618914159
transform 1 0 7544 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[232\]
timestamp 1618914159
transform 1 0 7820 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[233\]
timestamp 1618914159
transform 1 0 8096 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[234\]
timestamp 1618914159
transform 1 0 8372 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[235\]
timestamp 1618914159
transform 1 0 8648 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[236\]
timestamp 1618914159
transform 1 0 8924 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[237\]
timestamp 1618914159
transform 1 0 9200 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[238\]
timestamp 1618914159
transform 1 0 9476 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[239\]
timestamp 1618914159
transform 1 0 9752 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[23\]
timestamp 1618914159
transform 1 0 10028 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[240\]
timestamp 1618914159
transform 1 0 10304 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[241\]
timestamp 1618914159
transform 1 0 10580 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[242\]
timestamp 1618914159
transform 1 0 10856 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[243\]
timestamp 1618914159
transform 1 0 11132 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[244\]
timestamp 1618914159
transform 1 0 11684 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1618914159
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_112
timestamp 1618914159
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[245\]
timestamp 1618914159
transform 1 0 11960 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[246\]
timestamp 1618914159
transform 1 0 12236 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[247\]
timestamp 1618914159
transform 1 0 12512 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[248\]
timestamp 1618914159
transform 1 0 12788 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[249\]
timestamp 1618914159
transform 1 0 13064 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[24\]
timestamp 1618914159
transform 1 0 13340 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[250\]
timestamp 1618914159
transform 1 0 13616 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[251\]
timestamp 1618914159
transform 1 0 13892 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[252\]
timestamp 1618914159
transform 1 0 14168 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[253\]
timestamp 1618914159
transform 1 0 14444 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[254\]
timestamp 1618914159
transform 1 0 14720 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[255\]
timestamp 1618914159
transform 1 0 14996 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[256\]
timestamp 1618914159
transform 1 0 15272 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[257\]
timestamp 1618914159
transform 1 0 15548 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[258\]
timestamp 1618914159
transform 1 0 15824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[259\]
timestamp 1618914159
transform 1 0 16100 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[25\]
timestamp 1618914159
transform 1 0 16376 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[260\]
timestamp 1618914159
transform 1 0 16928 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[261\]
timestamp 1618914159
transform 1 0 17204 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[262\]
timestamp 1618914159
transform 1 0 17480 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1618914159
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1618914159
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[263\]
timestamp 1618914159
transform 1 0 17756 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[264\]
timestamp 1618914159
transform 1 0 18032 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[265\]
timestamp 1618914159
transform 1 0 18308 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[266\]
timestamp 1618914159
transform 1 0 18584 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[267\]
timestamp 1618914159
transform 1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[268\]
timestamp 1618914159
transform 1 0 19136 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[269\]
timestamp 1618914159
transform 1 0 19412 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[26\]
timestamp 1618914159
transform 1 0 19688 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[270\]
timestamp 1618914159
transform 1 0 19964 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[271\]
timestamp 1618914159
transform 1 0 20240 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[272\]
timestamp 1618914159
transform 1 0 20516 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[273\]
timestamp 1618914159
transform 1 0 20792 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[274\]
timestamp 1618914159
transform 1 0 21068 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[275\]
timestamp 1618914159
transform 1 0 21344 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[276\]
timestamp 1618914159
transform 1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[277\]
timestamp 1618914159
transform 1 0 22172 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1618914159
transform 1 0 22080 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_226
timestamp 1618914159
transform 1 0 21896 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[278\]
timestamp 1618914159
transform 1 0 22448 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[279\]
timestamp 1618914159
transform 1 0 22724 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[27\]
timestamp 1618914159
transform 1 0 23000 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[280\]
timestamp 1618914159
transform 1 0 23276 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[281\]
timestamp 1618914159
transform 1 0 23552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[282\]
timestamp 1618914159
transform 1 0 23828 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[283\]
timestamp 1618914159
transform 1 0 24104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[284\]
timestamp 1618914159
transform 1 0 24380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[285\]
timestamp 1618914159
transform 1 0 24656 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[286\]
timestamp 1618914159
transform 1 0 24932 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[287\]
timestamp 1618914159
transform 1 0 25208 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[288\]
timestamp 1618914159
transform 1 0 25484 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[289\]
timestamp 1618914159
transform 1 0 25760 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[28\]
timestamp 1618914159
transform 1 0 26036 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[290\]
timestamp 1618914159
transform 1 0 26312 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[291\]
timestamp 1618914159
transform 1 0 26588 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[292\]
timestamp 1618914159
transform 1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[293\]
timestamp 1618914159
transform 1 0 27416 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[294\]
timestamp 1618914159
transform 1 0 27692 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[295\]
timestamp 1618914159
transform 1 0 27968 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[296\]
timestamp 1618914159
transform 1 0 28244 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1618914159
transform 1 0 27324 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_283
timestamp 1618914159
transform 1 0 27140 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[297\]
timestamp 1618914159
transform 1 0 28520 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[298\]
timestamp 1618914159
transform 1 0 28796 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[299\]
timestamp 1618914159
transform 1 0 29072 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[29\]
timestamp 1618914159
transform 1 0 29348 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[2\]
timestamp 1618914159
transform 1 0 29624 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[300\]
timestamp 1618914159
transform 1 0 29900 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[301\]
timestamp 1618914159
transform 1 0 30176 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[302\]
timestamp 1618914159
transform 1 0 30452 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[303\]
timestamp 1618914159
transform 1 0 30728 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[304\]
timestamp 1618914159
transform 1 0 31004 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[305\]
timestamp 1618914159
transform 1 0 31280 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[306\]
timestamp 1618914159
transform 1 0 31556 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[204\]
timestamp 1618914159
transform 1 0 32016 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[307\]
timestamp 1618914159
transform 1 0 32292 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[308\]
timestamp 1618914159
transform 1 0 32660 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1618914159
transform 1 0 32568 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1618914159
transform 1 0 31832 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_346
timestamp 1618914159
transform 1 0 32936 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_358
timestamp 1618914159
transform 1 0 34040 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_370
timestamp 1618914159
transform 1 0 35144 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[414\]
timestamp 1618914159
transform 1 0 36248 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[415\]
timestamp 1618914159
transform 1 0 36524 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[416\]
timestamp 1618914159
transform 1 0 36800 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[417\]
timestamp 1618914159
transform 1 0 37076 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[418\]
timestamp 1618914159
transform 1 0 37352 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_397
timestamp 1618914159
transform 1 0 37628 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[419\]
timestamp 1618914159
transform 1 0 37904 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[41\]
timestamp 1618914159
transform 1 0 38180 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[420\]
timestamp 1618914159
transform 1 0 38456 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[421\]
timestamp 1618914159
transform 1 0 38732 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1618914159
transform 1 0 37812 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[422\]
timestamp 1618914159
transform 1 0 39008 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[423\]
timestamp 1618914159
transform 1 0 39284 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[424\]
timestamp 1618914159
transform 1 0 39560 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[425\]
timestamp 1618914159
transform 1 0 39836 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[426\]
timestamp 1618914159
transform 1 0 40112 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[427\]
timestamp 1618914159
transform 1 0 40388 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[428\]
timestamp 1618914159
transform 1 0 40664 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[429\]
timestamp 1618914159
transform 1 0 40940 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[42\]
timestamp 1618914159
transform 1 0 41216 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[430\]
timestamp 1618914159
transform 1 0 41492 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[431\]
timestamp 1618914159
transform 1 0 41768 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[432\]
timestamp 1618914159
transform 1 0 42044 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[433\]
timestamp 1618914159
transform 1 0 42320 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[434\]
timestamp 1618914159
transform 1 0 42596 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[435\]
timestamp 1618914159
transform 1 0 43148 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[436\]
timestamp 1618914159
transform 1 0 43424 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1618914159
transform 1 0 43056 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_454
timestamp 1618914159
transform 1 0 42872 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[437\]
timestamp 1618914159
transform 1 0 43700 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[438\]
timestamp 1618914159
transform 1 0 43976 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[439\]
timestamp 1618914159
transform 1 0 44252 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[43\]
timestamp 1618914159
transform 1 0 44528 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[440\]
timestamp 1618914159
transform 1 0 44804 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[441\]
timestamp 1618914159
transform 1 0 45080 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[442\]
timestamp 1618914159
transform 1 0 45356 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[443\]
timestamp 1618914159
transform 1 0 45632 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[444\]
timestamp 1618914159
transform 1 0 45908 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[445\]
timestamp 1618914159
transform 1 0 46184 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[446\]
timestamp 1618914159
transform 1 0 46460 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[447\]
timestamp 1618914159
transform 1 0 46736 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[448\]
timestamp 1618914159
transform 1 0 47012 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[449\]
timestamp 1618914159
transform 1 0 47288 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[44\]
timestamp 1618914159
transform 1 0 47564 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[450\]
timestamp 1618914159
transform 1 0 47840 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1618914159
transform 1 0 48300 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_511
timestamp 1618914159
transform 1 0 48116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[451\]
timestamp 1618914159
transform 1 0 48392 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[452\]
timestamp 1618914159
transform 1 0 48668 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[453\]
timestamp 1618914159
transform 1 0 48944 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[454\]
timestamp 1618914159
transform 1 0 49220 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[455\]
timestamp 1618914159
transform 1 0 49496 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[456\]
timestamp 1618914159
transform 1 0 49772 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[457\]
timestamp 1618914159
transform 1 0 50048 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[458\]
timestamp 1618914159
transform 1 0 50324 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[459\]
timestamp 1618914159
transform 1 0 50600 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[45\]
timestamp 1618914159
transform 1 0 50876 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[460\]
timestamp 1618914159
transform 1 0 51152 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[461\]
timestamp 1618914159
transform 1 0 51428 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[46\]
timestamp 1618914159
transform 1 0 51704 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[47\]
timestamp 1618914159
transform 1 0 51980 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[48\]
timestamp 1618914159
transform 1 0 52256 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[49\]
timestamp 1618914159
transform 1 0 52532 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[4\]
timestamp 1618914159
transform 1 0 52808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[50\]
timestamp 1618914159
transform 1 0 53084 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[51\]
timestamp 1618914159
transform 1 0 53636 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[52\]
timestamp 1618914159
transform 1 0 53912 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[53\]
timestamp 1618914159
transform 1 0 54188 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1618914159
transform 1 0 53544 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_568
timestamp 1618914159
transform 1 0 53360 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[54\]
timestamp 1618914159
transform 1 0 54464 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[55\]
timestamp 1618914159
transform 1 0 54740 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[56\]
timestamp 1618914159
transform 1 0 55016 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[57\]
timestamp 1618914159
transform 1 0 55292 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[58\]
timestamp 1618914159
transform 1 0 55568 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[59\]
timestamp 1618914159
transform 1 0 55844 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[5\]
timestamp 1618914159
transform 1 0 56120 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[60\]
timestamp 1618914159
transform 1 0 56396 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[61\]
timestamp 1618914159
transform 1 0 56672 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[62\]
timestamp 1618914159
transform 1 0 56948 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[63\]
timestamp 1618914159
transform 1 0 57224 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[64\]
timestamp 1618914159
transform 1 0 57500 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[65\]
timestamp 1618914159
transform 1 0 57776 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[66\]
timestamp 1618914159
transform 1 0 58052 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[67\]
timestamp 1618914159
transform 1 0 58328 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[68\]
timestamp 1618914159
transform 1 0 58880 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1618914159
transform 1 0 58788 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_625
timestamp 1618914159
transform 1 0 58604 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[69\]
timestamp 1618914159
transform 1 0 59156 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[6\]
timestamp 1618914159
transform 1 0 59432 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[70\]
timestamp 1618914159
transform 1 0 59708 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[71\]
timestamp 1618914159
transform 1 0 59984 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[72\]
timestamp 1618914159
transform 1 0 60260 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[73\]
timestamp 1618914159
transform 1 0 60536 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[74\]
timestamp 1618914159
transform 1 0 60812 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[75\]
timestamp 1618914159
transform 1 0 61088 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[76\]
timestamp 1618914159
transform 1 0 61364 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[77\]
timestamp 1618914159
transform 1 0 61640 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[78\]
timestamp 1618914159
transform 1 0 61916 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[79\]
timestamp 1618914159
transform 1 0 62192 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[7\]
timestamp 1618914159
transform 1 0 62468 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[80\]
timestamp 1618914159
transform 1 0 62744 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[81\]
timestamp 1618914159
transform 1 0 63020 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[82\]
timestamp 1618914159
transform 1 0 63296 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[83\]
timestamp 1618914159
transform 1 0 63572 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[84\]
timestamp 1618914159
transform 1 0 64124 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[85\]
timestamp 1618914159
transform 1 0 64400 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[86\]
timestamp 1618914159
transform 1 0 64676 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1618914159
transform 1 0 64032 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_682
timestamp 1618914159
transform 1 0 63848 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[87\]
timestamp 1618914159
transform 1 0 64952 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[88\]
timestamp 1618914159
transform 1 0 65228 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[89\]
timestamp 1618914159
transform 1 0 65504 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[8\]
timestamp 1618914159
transform 1 0 65780 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[90\]
timestamp 1618914159
transform 1 0 66056 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[91\]
timestamp 1618914159
transform 1 0 66332 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[92\]
timestamp 1618914159
transform 1 0 66608 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[93\]
timestamp 1618914159
transform 1 0 66884 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[94\]
timestamp 1618914159
transform 1 0 67160 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[95\]
timestamp 1618914159
transform 1 0 67436 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[96\]
timestamp 1618914159
transform 1 0 67712 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[97\]
timestamp 1618914159
transform 1 0 67988 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[98\]
timestamp 1618914159
transform 1 0 68264 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[413\]
timestamp 1618914159
transform 1 0 68724 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[99\]
timestamp 1618914159
transform 1 0 69000 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[9\]
timestamp 1618914159
transform 1 0 69368 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1618914159
transform 1 0 69276 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_733
timestamp 1618914159
transform 1 0 68540 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_745
timestamp 1618914159
transform 1 0 69644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_757
timestamp 1618914159
transform 1 0 70748 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_769
timestamp 1618914159
transform 1 0 71852 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1618914159
transform -1 0 72864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1618914159
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1618914159
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[213\]
timestamp 1618914159
transform 1 0 2484 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[214\]
timestamp 1618914159
transform 1 0 2760 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[215\]
timestamp 1618914159
transform 1 0 3036 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[216\]
timestamp 1618914159
transform 1 0 3312 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1618914159
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1618914159
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_30
timestamp 1618914159
transform 1 0 3864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_42
timestamp 1618914159
transform 1 0 4968 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1618914159
transform 1 0 6440 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_54
timestamp 1618914159
transform 1 0 6072 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_59
timestamp 1618914159
transform 1 0 6532 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_71
timestamp 1618914159
transform 1 0 7636 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1618914159
transform 1 0 9108 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_83
timestamp 1618914159
transform 1 0 8740 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_88
timestamp 1618914159
transform 1 0 9200 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_100
timestamp 1618914159
transform 1 0 10304 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_112
timestamp 1618914159
transform 1 0 11408 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1618914159
transform 1 0 11776 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1618914159
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1618914159
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1618914159
transform 1 0 14076 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1618914159
transform 1 0 14444 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_146
timestamp 1618914159
transform 1 0 14536 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_158
timestamp 1618914159
transform 1 0 15640 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1618914159
transform 1 0 17112 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_170
timestamp 1618914159
transform 1 0 16744 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_175
timestamp 1618914159
transform 1 0 17204 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_187
timestamp 1618914159
transform 1 0 18308 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1618914159
transform 1 0 19780 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_199
timestamp 1618914159
transform 1 0 19412 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_204
timestamp 1618914159
transform 1 0 19872 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_216
timestamp 1618914159
transform 1 0 20976 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_228
timestamp 1618914159
transform 1 0 22080 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1618914159
transform 1 0 22448 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1618914159
transform 1 0 22540 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_245
timestamp 1618914159
transform 1 0 23644 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1618914159
transform 1 0 25116 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_257
timestamp 1618914159
transform 1 0 24748 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_262
timestamp 1618914159
transform 1 0 25208 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_274
timestamp 1618914159
transform 1 0 26312 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1618914159
transform 1 0 27784 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_286
timestamp 1618914159
transform 1 0 27416 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_291
timestamp 1618914159
transform 1 0 27876 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_303
timestamp 1618914159
transform 1 0 28980 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1618914159
transform 1 0 30452 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_315
timestamp 1618914159
transform 1 0 30084 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_320
timestamp 1618914159
transform 1 0 30544 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_332
timestamp 1618914159
transform 1 0 31648 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_344
timestamp 1618914159
transform 1 0 32752 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1618914159
transform 1 0 33120 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_349
timestamp 1618914159
transform 1 0 33212 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_361
timestamp 1618914159
transform 1 0 34316 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1618914159
transform 1 0 35788 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_373
timestamp 1618914159
transform 1 0 35420 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_378
timestamp 1618914159
transform 1 0 35880 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_390
timestamp 1618914159
transform 1 0 36984 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1618914159
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_402
timestamp 1618914159
transform 1 0 38088 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_407
timestamp 1618914159
transform 1 0 38548 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_419
timestamp 1618914159
transform 1 0 39652 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1618914159
transform 1 0 41124 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_431
timestamp 1618914159
transform 1 0 40756 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_436
timestamp 1618914159
transform 1 0 41216 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_448
timestamp 1618914159
transform 1 0 42320 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_460
timestamp 1618914159
transform 1 0 43424 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1618914159
transform 1 0 43792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_465
timestamp 1618914159
transform 1 0 43884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1618914159
transform 1 0 44988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1618914159
transform 1 0 46460 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_489
timestamp 1618914159
transform 1 0 46092 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_494
timestamp 1618914159
transform 1 0 46552 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_506
timestamp 1618914159
transform 1 0 47656 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1618914159
transform 1 0 49128 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_518
timestamp 1618914159
transform 1 0 48760 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_523
timestamp 1618914159
transform 1 0 49220 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_535
timestamp 1618914159
transform 1 0 50324 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1618914159
transform 1 0 51796 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_547
timestamp 1618914159
transform 1 0 51428 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_552
timestamp 1618914159
transform 1 0 51888 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_564
timestamp 1618914159
transform 1 0 52992 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_576
timestamp 1618914159
transform 1 0 54096 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1618914159
transform 1 0 54464 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_581
timestamp 1618914159
transform 1 0 54556 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_593
timestamp 1618914159
transform 1 0 55660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1618914159
transform 1 0 57132 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_605
timestamp 1618914159
transform 1 0 56764 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_610
timestamp 1618914159
transform 1 0 57224 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_622
timestamp 1618914159
transform 1 0 58328 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1618914159
transform 1 0 59800 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_634
timestamp 1618914159
transform 1 0 59432 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_639
timestamp 1618914159
transform 1 0 59892 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_651
timestamp 1618914159
transform 1 0 60996 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1618914159
transform 1 0 62468 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_663
timestamp 1618914159
transform 1 0 62100 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_668
timestamp 1618914159
transform 1 0 62560 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_680
timestamp 1618914159
transform 1 0 63664 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_692
timestamp 1618914159
transform 1 0 64768 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1618914159
transform 1 0 65136 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_697
timestamp 1618914159
transform 1 0 65228 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_709
timestamp 1618914159
transform 1 0 66332 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1618914159
transform 1 0 67804 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_721
timestamp 1618914159
transform 1 0 67436 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_726
timestamp 1618914159
transform 1 0 67896 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_738
timestamp 1618914159
transform 1 0 69000 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1618914159
transform 1 0 70472 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_750
timestamp 1618914159
transform 1 0 70104 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_755
timestamp 1618914159
transform 1 0 70564 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_767
timestamp 1618914159
transform 1 0 71668 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1618914159
transform -1 0 72864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_775
timestamp 1618914159
transform 1 0 72404 0 -1 3808
box -38 -48 222 592
<< labels >>
rlabel metal2 s 32310 0 32366 1000 6 HI[0]
port 0 nsew signal tristate
rlabel metal2 s 20994 0 21050 1000 6 HI[100]
port 1 nsew signal tristate
rlabel metal2 s 30378 0 30434 1000 6 HI[101]
port 2 nsew signal tristate
rlabel metal2 s 10230 0 10286 1000 6 HI[102]
port 3 nsew signal tristate
rlabel metal2 s 846 0 902 1000 6 HI[103]
port 4 nsew signal tristate
rlabel metal2 s 26238 0 26294 1000 6 HI[104]
port 5 nsew signal tristate
rlabel metal2 s 32034 0 32090 1000 6 HI[105]
port 6 nsew signal tristate
rlabel metal2 s 8298 0 8354 1000 6 HI[106]
port 7 nsew signal tristate
rlabel metal2 s 31758 0 31814 1000 6 HI[107]
port 8 nsew signal tristate
rlabel metal2 s 26514 0 26570 1000 6 HI[108]
port 9 nsew signal tristate
rlabel metal2 s 9954 0 10010 1000 6 HI[109]
port 10 nsew signal tristate
rlabel metal2 s 17406 0 17462 1000 6 HI[10]
port 11 nsew signal tristate
rlabel metal2 s 5814 0 5870 1000 6 HI[110]
port 12 nsew signal tristate
rlabel metal2 s 26790 0 26846 1000 6 HI[111]
port 13 nsew signal tristate
rlabel metal2 s 17682 0 17738 1000 6 HI[112]
port 14 nsew signal tristate
rlabel metal2 s 27618 0 27674 1000 6 HI[113]
port 15 nsew signal tristate
rlabel metal2 s 1122 0 1178 1000 6 HI[114]
port 16 nsew signal tristate
rlabel metal2 s 27066 0 27122 1000 6 HI[115]
port 17 nsew signal tristate
rlabel metal2 s 14646 0 14702 1000 6 HI[116]
port 18 nsew signal tristate
rlabel metal2 s 5262 0 5318 1000 6 HI[117]
port 19 nsew signal tristate
rlabel metal2 s 18234 0 18290 1000 6 HI[118]
port 20 nsew signal tristate
rlabel metal2 s 11886 0 11942 1000 6 HI[119]
port 21 nsew signal tristate
rlabel metal2 s 27342 0 27398 1000 6 HI[11]
port 22 nsew signal tristate
rlabel metal2 s 18510 0 18566 1000 6 HI[120]
port 23 nsew signal tristate
rlabel metal2 s 1674 0 1730 1000 6 HI[121]
port 24 nsew signal tristate
rlabel metal2 s 11334 0 11390 1000 6 HI[122]
port 25 nsew signal tristate
rlabel metal2 s 30654 0 30710 1000 6 HI[123]
port 26 nsew signal tristate
rlabel metal2 s 12438 0 12494 1000 6 HI[124]
port 27 nsew signal tristate
rlabel metal2 s 6918 0 6974 1000 6 HI[125]
port 28 nsew signal tristate
rlabel metal2 s 19062 0 19118 1000 6 HI[126]
port 29 nsew signal tristate
rlabel metal2 s 27894 0 27950 1000 6 HI[127]
port 30 nsew signal tristate
rlabel metal2 s 15474 0 15530 1000 6 HI[128]
port 31 nsew signal tristate
rlabel metal2 s 19338 0 19394 1000 6 HI[129]
port 32 nsew signal tristate
rlabel metal2 s 17958 0 18014 1000 6 HI[12]
port 33 nsew signal tristate
rlabel metal2 s 28170 0 28226 1000 6 HI[130]
port 34 nsew signal tristate
rlabel metal2 s 19614 0 19670 1000 6 HI[131]
port 35 nsew signal tristate
rlabel metal2 s 4710 0 4766 1000 6 HI[132]
port 36 nsew signal tristate
rlabel metal2 s 10782 0 10838 1000 6 HI[133]
port 37 nsew signal tristate
rlabel metal2 s 28446 0 28502 1000 6 HI[134]
port 38 nsew signal tristate
rlabel metal2 s 13542 0 13598 1000 6 HI[135]
port 39 nsew signal tristate
rlabel metal2 s 30930 0 30986 1000 6 HI[136]
port 40 nsew signal tristate
rlabel metal2 s 20442 0 20498 1000 6 HI[137]
port 41 nsew signal tristate
rlabel metal2 s 7194 0 7250 1000 6 HI[138]
port 42 nsew signal tristate
rlabel metal2 s 6366 0 6422 1000 6 HI[139]
port 43 nsew signal tristate
rlabel metal2 s 21270 0 21326 1000 6 HI[13]
port 44 nsew signal tristate
rlabel metal2 s 28722 0 28778 1000 6 HI[140]
port 45 nsew signal tristate
rlabel metal2 s 3606 0 3662 1000 6 HI[141]
port 46 nsew signal tristate
rlabel metal2 s 20718 0 20774 1000 6 HI[142]
port 47 nsew signal tristate
rlabel metal2 s 4434 0 4490 1000 6 HI[143]
port 48 nsew signal tristate
rlabel metal2 s 28998 0 29054 1000 6 HI[144]
port 49 nsew signal tristate
rlabel metal2 s 31206 0 31262 1000 6 HI[145]
port 50 nsew signal tristate
rlabel metal2 s 18786 0 18842 1000 6 HI[146]
port 51 nsew signal tristate
rlabel metal2 s 16578 0 16634 1000 6 HI[147]
port 52 nsew signal tristate
rlabel metal2 s 23202 0 23258 1000 6 HI[148]
port 53 nsew signal tristate
rlabel metal2 s 17130 0 17186 1000 6 HI[149]
port 54 nsew signal tristate
rlabel metal2 s 8022 0 8078 1000 6 HI[14]
port 55 nsew signal tristate
rlabel metal2 s 21546 0 21602 1000 6 HI[150]
port 56 nsew signal tristate
rlabel metal2 s 15198 0 15254 1000 6 HI[151]
port 57 nsew signal tristate
rlabel metal2 s 7470 0 7526 1000 6 HI[152]
port 58 nsew signal tristate
rlabel metal2 s 21822 0 21878 1000 6 HI[153]
port 59 nsew signal tristate
rlabel metal2 s 12714 0 12770 1000 6 HI[154]
port 60 nsew signal tristate
rlabel metal2 s 8850 0 8906 1000 6 HI[155]
port 61 nsew signal tristate
rlabel metal2 s 22098 0 22154 1000 6 HI[156]
port 62 nsew signal tristate
rlabel metal2 s 9126 0 9182 1000 6 HI[157]
port 63 nsew signal tristate
rlabel metal2 s 1950 0 2006 1000 6 HI[158]
port 64 nsew signal tristate
rlabel metal2 s 22374 0 22430 1000 6 HI[159]
port 65 nsew signal tristate
rlabel metal2 s 2226 0 2282 1000 6 HI[15]
port 66 nsew signal tristate
rlabel metal2 s 9678 0 9734 1000 6 HI[160]
port 67 nsew signal tristate
rlabel metal2 s 22650 0 22706 1000 6 HI[161]
port 68 nsew signal tristate
rlabel metal2 s 16302 0 16358 1000 6 HI[162]
port 69 nsew signal tristate
rlabel metal2 s 3330 0 3386 1000 6 HI[163]
port 70 nsew signal tristate
rlabel metal2 s 22926 0 22982 1000 6 HI[164]
port 71 nsew signal tristate
rlabel metal2 s 4158 0 4214 1000 6 HI[165]
port 72 nsew signal tristate
rlabel metal2 s 10506 0 10562 1000 6 HI[166]
port 73 nsew signal tristate
rlabel metal2 s 3882 0 3938 1000 6 HI[167]
port 74 nsew signal tristate
rlabel metal2 s 29274 0 29330 1000 6 HI[168]
port 75 nsew signal tristate
rlabel metal2 s 16854 0 16910 1000 6 HI[169]
port 76 nsew signal tristate
rlabel metal2 s 11058 0 11114 1000 6 HI[16]
port 77 nsew signal tristate
rlabel metal2 s 13266 0 13322 1000 6 HI[170]
port 78 nsew signal tristate
rlabel metal2 s 23478 0 23534 1000 6 HI[171]
port 79 nsew signal tristate
rlabel metal2 s 6090 0 6146 1000 6 HI[172]
port 80 nsew signal tristate
rlabel metal2 s 11610 0 11666 1000 6 HI[173]
port 81 nsew signal tristate
rlabel metal2 s 570 0 626 1000 6 HI[174]
port 82 nsew signal tristate
rlabel metal2 s 23754 0 23810 1000 6 HI[175]
port 83 nsew signal tristate
rlabel metal2 s 4986 0 5042 1000 6 HI[176]
port 84 nsew signal tristate
rlabel metal2 s 12162 0 12218 1000 6 HI[177]
port 85 nsew signal tristate
rlabel metal2 s 14094 0 14150 1000 6 HI[178]
port 86 nsew signal tristate
rlabel metal2 s 24030 0 24086 1000 6 HI[179]
port 87 nsew signal tristate
rlabel metal2 s 7746 0 7802 1000 6 HI[17]
port 88 nsew signal tristate
rlabel metal2 s 29550 0 29606 1000 6 HI[180]
port 89 nsew signal tristate
rlabel metal2 s 2778 0 2834 1000 6 HI[181]
port 90 nsew signal tristate
rlabel metal2 s 24306 0 24362 1000 6 HI[182]
port 91 nsew signal tristate
rlabel metal2 s 2502 0 2558 1000 6 HI[183]
port 92 nsew signal tristate
rlabel metal2 s 16026 0 16082 1000 6 HI[184]
port 93 nsew signal tristate
rlabel metal2 s 31482 0 31538 1000 6 HI[185]
port 94 nsew signal tristate
rlabel metal2 s 24582 0 24638 1000 6 HI[186]
port 95 nsew signal tristate
rlabel metal2 s 6642 0 6698 1000 6 HI[187]
port 96 nsew signal tristate
rlabel metal2 s 13818 0 13874 1000 6 HI[188]
port 97 nsew signal tristate
rlabel metal2 s 8574 0 8630 1000 6 HI[189]
port 98 nsew signal tristate
rlabel metal2 s 24858 0 24914 1000 6 HI[18]
port 99 nsew signal tristate
rlabel metal2 s 29826 0 29882 1000 6 HI[190]
port 100 nsew signal tristate
rlabel metal2 s 14370 0 14426 1000 6 HI[191]
port 101 nsew signal tristate
rlabel metal2 s 5538 0 5594 1000 6 HI[192]
port 102 nsew signal tristate
rlabel metal2 s 25134 0 25190 1000 6 HI[193]
port 103 nsew signal tristate
rlabel metal2 s 20166 0 20222 1000 6 HI[194]
port 104 nsew signal tristate
rlabel metal2 s 14922 0 14978 1000 6 HI[195]
port 105 nsew signal tristate
rlabel metal2 s 1398 0 1454 1000 6 HI[196]
port 106 nsew signal tristate
rlabel metal2 s 25410 0 25466 1000 6 HI[197]
port 107 nsew signal tristate
rlabel metal2 s 9402 0 9458 1000 6 HI[198]
port 108 nsew signal tristate
rlabel metal2 s 30102 0 30158 1000 6 HI[199]
port 109 nsew signal tristate
rlabel metal2 s 3054 0 3110 1000 6 HI[19]
port 110 nsew signal tristate
rlabel metal2 s 15750 0 15806 1000 6 HI[1]
port 111 nsew signal tristate
rlabel metal2 s 25686 0 25742 1000 6 HI[200]
port 112 nsew signal tristate
rlabel metal2 s 19890 0 19946 1000 6 HI[201]
port 113 nsew signal tristate
rlabel metal2 s 12990 0 13046 1000 6 HI[202]
port 114 nsew signal tristate
rlabel metal2 s 25962 0 26018 1000 6 HI[203]
port 115 nsew signal tristate
rlabel metal2 s 30378 4000 30434 5000 6 HI[204]
port 116 nsew signal tristate
rlabel metal3 s 0 1232 1000 1352 6 HI[205]
port 117 nsew signal tristate
rlabel metal3 s 0 1640 1000 1760 6 HI[206]
port 118 nsew signal tristate
rlabel metal3 s 0 2048 1000 2168 6 HI[207]
port 119 nsew signal tristate
rlabel metal3 s 0 2456 1000 2576 6 HI[208]
port 120 nsew signal tristate
rlabel metal3 s 0 2864 1000 2984 6 HI[209]
port 121 nsew signal tristate
rlabel metal3 s 0 3272 1000 3392 6 HI[20]
port 122 nsew signal tristate
rlabel metal3 s 0 3680 1000 3800 6 HI[210]
port 123 nsew signal tristate
rlabel metal2 s 570 4000 626 5000 6 HI[211]
port 124 nsew signal tristate
rlabel metal2 s 846 4000 902 5000 6 HI[212]
port 125 nsew signal tristate
rlabel metal2 s 1122 4000 1178 5000 6 HI[213]
port 126 nsew signal tristate
rlabel metal2 s 1398 4000 1454 5000 6 HI[214]
port 127 nsew signal tristate
rlabel metal2 s 1674 4000 1730 5000 6 HI[215]
port 128 nsew signal tristate
rlabel metal2 s 1950 4000 2006 5000 6 HI[216]
port 129 nsew signal tristate
rlabel metal2 s 2226 4000 2282 5000 6 HI[217]
port 130 nsew signal tristate
rlabel metal2 s 2502 4000 2558 5000 6 HI[218]
port 131 nsew signal tristate
rlabel metal2 s 2778 4000 2834 5000 6 HI[219]
port 132 nsew signal tristate
rlabel metal2 s 3054 4000 3110 5000 6 HI[21]
port 133 nsew signal tristate
rlabel metal2 s 3330 4000 3386 5000 6 HI[220]
port 134 nsew signal tristate
rlabel metal2 s 3606 4000 3662 5000 6 HI[221]
port 135 nsew signal tristate
rlabel metal2 s 3882 4000 3938 5000 6 HI[222]
port 136 nsew signal tristate
rlabel metal2 s 4158 4000 4214 5000 6 HI[223]
port 137 nsew signal tristate
rlabel metal2 s 4434 4000 4490 5000 6 HI[224]
port 138 nsew signal tristate
rlabel metal2 s 4710 4000 4766 5000 6 HI[225]
port 139 nsew signal tristate
rlabel metal2 s 4986 4000 5042 5000 6 HI[226]
port 140 nsew signal tristate
rlabel metal2 s 5262 4000 5318 5000 6 HI[227]
port 141 nsew signal tristate
rlabel metal2 s 5538 4000 5594 5000 6 HI[228]
port 142 nsew signal tristate
rlabel metal2 s 5814 4000 5870 5000 6 HI[229]
port 143 nsew signal tristate
rlabel metal2 s 6090 4000 6146 5000 6 HI[22]
port 144 nsew signal tristate
rlabel metal2 s 6366 4000 6422 5000 6 HI[230]
port 145 nsew signal tristate
rlabel metal2 s 6642 4000 6698 5000 6 HI[231]
port 146 nsew signal tristate
rlabel metal2 s 6918 4000 6974 5000 6 HI[232]
port 147 nsew signal tristate
rlabel metal2 s 7194 4000 7250 5000 6 HI[233]
port 148 nsew signal tristate
rlabel metal2 s 7470 4000 7526 5000 6 HI[234]
port 149 nsew signal tristate
rlabel metal2 s 7746 4000 7802 5000 6 HI[235]
port 150 nsew signal tristate
rlabel metal2 s 8022 4000 8078 5000 6 HI[236]
port 151 nsew signal tristate
rlabel metal2 s 8298 4000 8354 5000 6 HI[237]
port 152 nsew signal tristate
rlabel metal2 s 8574 4000 8630 5000 6 HI[238]
port 153 nsew signal tristate
rlabel metal2 s 8850 4000 8906 5000 6 HI[239]
port 154 nsew signal tristate
rlabel metal2 s 9126 4000 9182 5000 6 HI[23]
port 155 nsew signal tristate
rlabel metal2 s 9402 4000 9458 5000 6 HI[240]
port 156 nsew signal tristate
rlabel metal2 s 9678 4000 9734 5000 6 HI[241]
port 157 nsew signal tristate
rlabel metal2 s 9954 4000 10010 5000 6 HI[242]
port 158 nsew signal tristate
rlabel metal2 s 10230 4000 10286 5000 6 HI[243]
port 159 nsew signal tristate
rlabel metal2 s 10506 4000 10562 5000 6 HI[244]
port 160 nsew signal tristate
rlabel metal2 s 10782 4000 10838 5000 6 HI[245]
port 161 nsew signal tristate
rlabel metal2 s 11058 4000 11114 5000 6 HI[246]
port 162 nsew signal tristate
rlabel metal2 s 11334 4000 11390 5000 6 HI[247]
port 163 nsew signal tristate
rlabel metal2 s 11610 4000 11666 5000 6 HI[248]
port 164 nsew signal tristate
rlabel metal2 s 11886 4000 11942 5000 6 HI[249]
port 165 nsew signal tristate
rlabel metal2 s 12162 4000 12218 5000 6 HI[24]
port 166 nsew signal tristate
rlabel metal2 s 12438 4000 12494 5000 6 HI[250]
port 167 nsew signal tristate
rlabel metal2 s 12714 4000 12770 5000 6 HI[251]
port 168 nsew signal tristate
rlabel metal2 s 12990 4000 13046 5000 6 HI[252]
port 169 nsew signal tristate
rlabel metal2 s 13266 4000 13322 5000 6 HI[253]
port 170 nsew signal tristate
rlabel metal2 s 13542 4000 13598 5000 6 HI[254]
port 171 nsew signal tristate
rlabel metal2 s 13818 4000 13874 5000 6 HI[255]
port 172 nsew signal tristate
rlabel metal2 s 14094 4000 14150 5000 6 HI[256]
port 173 nsew signal tristate
rlabel metal2 s 14370 4000 14426 5000 6 HI[257]
port 174 nsew signal tristate
rlabel metal2 s 14646 4000 14702 5000 6 HI[258]
port 175 nsew signal tristate
rlabel metal2 s 14922 4000 14978 5000 6 HI[259]
port 176 nsew signal tristate
rlabel metal2 s 15198 4000 15254 5000 6 HI[25]
port 177 nsew signal tristate
rlabel metal2 s 15474 4000 15530 5000 6 HI[260]
port 178 nsew signal tristate
rlabel metal2 s 15750 4000 15806 5000 6 HI[261]
port 179 nsew signal tristate
rlabel metal2 s 16026 4000 16082 5000 6 HI[262]
port 180 nsew signal tristate
rlabel metal2 s 16302 4000 16358 5000 6 HI[263]
port 181 nsew signal tristate
rlabel metal2 s 16578 4000 16634 5000 6 HI[264]
port 182 nsew signal tristate
rlabel metal2 s 16854 4000 16910 5000 6 HI[265]
port 183 nsew signal tristate
rlabel metal2 s 17130 4000 17186 5000 6 HI[266]
port 184 nsew signal tristate
rlabel metal2 s 17406 4000 17462 5000 6 HI[267]
port 185 nsew signal tristate
rlabel metal2 s 17682 4000 17738 5000 6 HI[268]
port 186 nsew signal tristate
rlabel metal2 s 17958 4000 18014 5000 6 HI[269]
port 187 nsew signal tristate
rlabel metal2 s 18234 4000 18290 5000 6 HI[26]
port 188 nsew signal tristate
rlabel metal2 s 18510 4000 18566 5000 6 HI[270]
port 189 nsew signal tristate
rlabel metal2 s 18786 4000 18842 5000 6 HI[271]
port 190 nsew signal tristate
rlabel metal2 s 19062 4000 19118 5000 6 HI[272]
port 191 nsew signal tristate
rlabel metal2 s 19338 4000 19394 5000 6 HI[273]
port 192 nsew signal tristate
rlabel metal2 s 19614 4000 19670 5000 6 HI[274]
port 193 nsew signal tristate
rlabel metal2 s 19890 4000 19946 5000 6 HI[275]
port 194 nsew signal tristate
rlabel metal2 s 20166 4000 20222 5000 6 HI[276]
port 195 nsew signal tristate
rlabel metal2 s 20442 4000 20498 5000 6 HI[277]
port 196 nsew signal tristate
rlabel metal2 s 20718 4000 20774 5000 6 HI[278]
port 197 nsew signal tristate
rlabel metal2 s 20994 4000 21050 5000 6 HI[279]
port 198 nsew signal tristate
rlabel metal2 s 21270 4000 21326 5000 6 HI[27]
port 199 nsew signal tristate
rlabel metal2 s 21546 4000 21602 5000 6 HI[280]
port 200 nsew signal tristate
rlabel metal2 s 21822 4000 21878 5000 6 HI[281]
port 201 nsew signal tristate
rlabel metal2 s 22098 4000 22154 5000 6 HI[282]
port 202 nsew signal tristate
rlabel metal2 s 22374 4000 22430 5000 6 HI[283]
port 203 nsew signal tristate
rlabel metal2 s 22650 4000 22706 5000 6 HI[284]
port 204 nsew signal tristate
rlabel metal2 s 22926 4000 22982 5000 6 HI[285]
port 205 nsew signal tristate
rlabel metal2 s 23202 4000 23258 5000 6 HI[286]
port 206 nsew signal tristate
rlabel metal2 s 23478 4000 23534 5000 6 HI[287]
port 207 nsew signal tristate
rlabel metal2 s 23754 4000 23810 5000 6 HI[288]
port 208 nsew signal tristate
rlabel metal2 s 24030 4000 24086 5000 6 HI[289]
port 209 nsew signal tristate
rlabel metal2 s 24306 4000 24362 5000 6 HI[28]
port 210 nsew signal tristate
rlabel metal2 s 24582 4000 24638 5000 6 HI[290]
port 211 nsew signal tristate
rlabel metal2 s 24858 4000 24914 5000 6 HI[291]
port 212 nsew signal tristate
rlabel metal2 s 25134 4000 25190 5000 6 HI[292]
port 213 nsew signal tristate
rlabel metal2 s 25410 4000 25466 5000 6 HI[293]
port 214 nsew signal tristate
rlabel metal2 s 25686 4000 25742 5000 6 HI[294]
port 215 nsew signal tristate
rlabel metal2 s 25962 4000 26018 5000 6 HI[295]
port 216 nsew signal tristate
rlabel metal2 s 26238 4000 26294 5000 6 HI[296]
port 217 nsew signal tristate
rlabel metal2 s 26514 4000 26570 5000 6 HI[297]
port 218 nsew signal tristate
rlabel metal2 s 26790 4000 26846 5000 6 HI[298]
port 219 nsew signal tristate
rlabel metal2 s 27066 4000 27122 5000 6 HI[299]
port 220 nsew signal tristate
rlabel metal2 s 27342 4000 27398 5000 6 HI[29]
port 221 nsew signal tristate
rlabel metal2 s 27618 4000 27674 5000 6 HI[2]
port 222 nsew signal tristate
rlabel metal2 s 27894 4000 27950 5000 6 HI[300]
port 223 nsew signal tristate
rlabel metal2 s 28170 4000 28226 5000 6 HI[301]
port 224 nsew signal tristate
rlabel metal2 s 28446 4000 28502 5000 6 HI[302]
port 225 nsew signal tristate
rlabel metal2 s 28722 4000 28778 5000 6 HI[303]
port 226 nsew signal tristate
rlabel metal2 s 28998 4000 29054 5000 6 HI[304]
port 227 nsew signal tristate
rlabel metal2 s 29274 4000 29330 5000 6 HI[305]
port 228 nsew signal tristate
rlabel metal2 s 29550 4000 29606 5000 6 HI[306]
port 229 nsew signal tristate
rlabel metal2 s 29826 4000 29882 5000 6 HI[307]
port 230 nsew signal tristate
rlabel metal2 s 30102 4000 30158 5000 6 HI[308]
port 231 nsew signal tristate
rlabel metal2 s 69846 0 69902 1000 6 HI[309]
port 232 nsew signal tristate
rlabel metal2 s 58530 0 58586 1000 6 HI[30]
port 233 nsew signal tristate
rlabel metal2 s 67914 0 67970 1000 6 HI[310]
port 234 nsew signal tristate
rlabel metal2 s 47766 0 47822 1000 6 HI[311]
port 235 nsew signal tristate
rlabel metal2 s 38382 0 38438 1000 6 HI[312]
port 236 nsew signal tristate
rlabel metal2 s 63774 0 63830 1000 6 HI[313]
port 237 nsew signal tristate
rlabel metal2 s 69570 0 69626 1000 6 HI[314]
port 238 nsew signal tristate
rlabel metal2 s 45834 0 45890 1000 6 HI[315]
port 239 nsew signal tristate
rlabel metal2 s 69294 0 69350 1000 6 HI[316]
port 240 nsew signal tristate
rlabel metal2 s 64050 0 64106 1000 6 HI[317]
port 241 nsew signal tristate
rlabel metal2 s 47490 0 47546 1000 6 HI[318]
port 242 nsew signal tristate
rlabel metal2 s 54942 0 54998 1000 6 HI[319]
port 243 nsew signal tristate
rlabel metal2 s 43350 0 43406 1000 6 HI[31]
port 244 nsew signal tristate
rlabel metal2 s 64326 0 64382 1000 6 HI[320]
port 245 nsew signal tristate
rlabel metal2 s 55218 0 55274 1000 6 HI[321]
port 246 nsew signal tristate
rlabel metal2 s 65154 0 65210 1000 6 HI[322]
port 247 nsew signal tristate
rlabel metal2 s 38658 0 38714 1000 6 HI[323]
port 248 nsew signal tristate
rlabel metal2 s 64602 0 64658 1000 6 HI[324]
port 249 nsew signal tristate
rlabel metal2 s 52182 0 52238 1000 6 HI[325]
port 250 nsew signal tristate
rlabel metal2 s 42798 0 42854 1000 6 HI[326]
port 251 nsew signal tristate
rlabel metal2 s 55770 0 55826 1000 6 HI[327]
port 252 nsew signal tristate
rlabel metal2 s 49422 0 49478 1000 6 HI[328]
port 253 nsew signal tristate
rlabel metal2 s 64878 0 64934 1000 6 HI[329]
port 254 nsew signal tristate
rlabel metal2 s 56046 0 56102 1000 6 HI[32]
port 255 nsew signal tristate
rlabel metal2 s 39210 0 39266 1000 6 HI[330]
port 256 nsew signal tristate
rlabel metal2 s 48870 0 48926 1000 6 HI[331]
port 257 nsew signal tristate
rlabel metal2 s 68190 0 68246 1000 6 HI[332]
port 258 nsew signal tristate
rlabel metal2 s 49974 0 50030 1000 6 HI[333]
port 259 nsew signal tristate
rlabel metal2 s 44454 0 44510 1000 6 HI[334]
port 260 nsew signal tristate
rlabel metal2 s 56598 0 56654 1000 6 HI[335]
port 261 nsew signal tristate
rlabel metal2 s 65430 0 65486 1000 6 HI[336]
port 262 nsew signal tristate
rlabel metal2 s 53010 0 53066 1000 6 HI[337]
port 263 nsew signal tristate
rlabel metal2 s 56874 0 56930 1000 6 HI[338]
port 264 nsew signal tristate
rlabel metal2 s 55494 0 55550 1000 6 HI[339]
port 265 nsew signal tristate
rlabel metal2 s 65706 0 65762 1000 6 HI[33]
port 266 nsew signal tristate
rlabel metal2 s 57150 0 57206 1000 6 HI[340]
port 267 nsew signal tristate
rlabel metal2 s 42246 0 42302 1000 6 HI[341]
port 268 nsew signal tristate
rlabel metal2 s 48318 0 48374 1000 6 HI[342]
port 269 nsew signal tristate
rlabel metal2 s 65982 0 66038 1000 6 HI[343]
port 270 nsew signal tristate
rlabel metal2 s 51078 0 51134 1000 6 HI[344]
port 271 nsew signal tristate
rlabel metal2 s 68466 0 68522 1000 6 HI[345]
port 272 nsew signal tristate
rlabel metal2 s 57978 0 58034 1000 6 HI[346]
port 273 nsew signal tristate
rlabel metal2 s 44730 0 44786 1000 6 HI[347]
port 274 nsew signal tristate
rlabel metal2 s 43902 0 43958 1000 6 HI[348]
port 275 nsew signal tristate
rlabel metal2 s 58806 0 58862 1000 6 HI[349]
port 276 nsew signal tristate
rlabel metal2 s 66258 0 66314 1000 6 HI[34]
port 277 nsew signal tristate
rlabel metal2 s 41142 0 41198 1000 6 HI[350]
port 278 nsew signal tristate
rlabel metal2 s 58254 0 58310 1000 6 HI[351]
port 279 nsew signal tristate
rlabel metal2 s 41970 0 42026 1000 6 HI[352]
port 280 nsew signal tristate
rlabel metal2 s 66534 0 66590 1000 6 HI[353]
port 281 nsew signal tristate
rlabel metal2 s 68742 0 68798 1000 6 HI[354]
port 282 nsew signal tristate
rlabel metal2 s 56322 0 56378 1000 6 HI[355]
port 283 nsew signal tristate
rlabel metal2 s 54114 0 54170 1000 6 HI[356]
port 284 nsew signal tristate
rlabel metal2 s 60738 0 60794 1000 6 HI[357]
port 285 nsew signal tristate
rlabel metal2 s 54666 0 54722 1000 6 HI[358]
port 286 nsew signal tristate
rlabel metal2 s 45558 0 45614 1000 6 HI[359]
port 287 nsew signal tristate
rlabel metal2 s 59082 0 59138 1000 6 HI[35]
port 288 nsew signal tristate
rlabel metal2 s 52734 0 52790 1000 6 HI[360]
port 289 nsew signal tristate
rlabel metal2 s 45006 0 45062 1000 6 HI[361]
port 290 nsew signal tristate
rlabel metal2 s 59358 0 59414 1000 6 HI[362]
port 291 nsew signal tristate
rlabel metal2 s 50250 0 50306 1000 6 HI[363]
port 292 nsew signal tristate
rlabel metal2 s 46386 0 46442 1000 6 HI[364]
port 293 nsew signal tristate
rlabel metal2 s 59634 0 59690 1000 6 HI[365]
port 294 nsew signal tristate
rlabel metal2 s 46662 0 46718 1000 6 HI[366]
port 295 nsew signal tristate
rlabel metal2 s 39486 0 39542 1000 6 HI[367]
port 296 nsew signal tristate
rlabel metal2 s 59910 0 59966 1000 6 HI[368]
port 297 nsew signal tristate
rlabel metal2 s 39762 0 39818 1000 6 HI[369]
port 298 nsew signal tristate
rlabel metal2 s 47214 0 47270 1000 6 HI[36]
port 299 nsew signal tristate
rlabel metal2 s 60186 0 60242 1000 6 HI[370]
port 300 nsew signal tristate
rlabel metal2 s 53838 0 53894 1000 6 HI[371]
port 301 nsew signal tristate
rlabel metal2 s 40866 0 40922 1000 6 HI[372]
port 302 nsew signal tristate
rlabel metal2 s 60462 0 60518 1000 6 HI[373]
port 303 nsew signal tristate
rlabel metal2 s 41694 0 41750 1000 6 HI[374]
port 304 nsew signal tristate
rlabel metal2 s 48042 0 48098 1000 6 HI[375]
port 305 nsew signal tristate
rlabel metal2 s 41418 0 41474 1000 6 HI[376]
port 306 nsew signal tristate
rlabel metal2 s 66810 0 66866 1000 6 HI[377]
port 307 nsew signal tristate
rlabel metal2 s 54390 0 54446 1000 6 HI[378]
port 308 nsew signal tristate
rlabel metal2 s 48594 0 48650 1000 6 HI[379]
port 309 nsew signal tristate
rlabel metal2 s 50802 0 50858 1000 6 HI[37]
port 310 nsew signal tristate
rlabel metal2 s 61014 0 61070 1000 6 HI[380]
port 311 nsew signal tristate
rlabel metal2 s 43626 0 43682 1000 6 HI[381]
port 312 nsew signal tristate
rlabel metal2 s 49146 0 49202 1000 6 HI[382]
port 313 nsew signal tristate
rlabel metal2 s 38106 0 38162 1000 6 HI[383]
port 314 nsew signal tristate
rlabel metal2 s 61290 0 61346 1000 6 HI[384]
port 315 nsew signal tristate
rlabel metal2 s 42522 0 42578 1000 6 HI[385]
port 316 nsew signal tristate
rlabel metal2 s 49698 0 49754 1000 6 HI[386]
port 317 nsew signal tristate
rlabel metal2 s 51630 0 51686 1000 6 HI[387]
port 318 nsew signal tristate
rlabel metal2 s 61566 0 61622 1000 6 HI[388]
port 319 nsew signal tristate
rlabel metal2 s 45282 0 45338 1000 6 HI[389]
port 320 nsew signal tristate
rlabel metal2 s 67086 0 67142 1000 6 HI[38]
port 321 nsew signal tristate
rlabel metal2 s 40314 0 40370 1000 6 HI[390]
port 322 nsew signal tristate
rlabel metal2 s 61842 0 61898 1000 6 HI[391]
port 323 nsew signal tristate
rlabel metal2 s 40038 0 40094 1000 6 HI[392]
port 324 nsew signal tristate
rlabel metal2 s 53562 0 53618 1000 6 HI[393]
port 325 nsew signal tristate
rlabel metal2 s 69018 0 69074 1000 6 HI[394]
port 326 nsew signal tristate
rlabel metal2 s 62118 0 62174 1000 6 HI[395]
port 327 nsew signal tristate
rlabel metal2 s 44178 0 44234 1000 6 HI[396]
port 328 nsew signal tristate
rlabel metal2 s 51354 0 51410 1000 6 HI[397]
port 329 nsew signal tristate
rlabel metal2 s 46110 0 46166 1000 6 HI[398]
port 330 nsew signal tristate
rlabel metal2 s 62394 0 62450 1000 6 HI[399]
port 331 nsew signal tristate
rlabel metal2 s 67362 0 67418 1000 6 HI[39]
port 332 nsew signal tristate
rlabel metal2 s 51906 0 51962 1000 6 HI[3]
port 333 nsew signal tristate
rlabel metal2 s 43074 0 43130 1000 6 HI[400]
port 334 nsew signal tristate
rlabel metal2 s 62670 0 62726 1000 6 HI[401]
port 335 nsew signal tristate
rlabel metal2 s 57702 0 57758 1000 6 HI[402]
port 336 nsew signal tristate
rlabel metal2 s 52458 0 52514 1000 6 HI[403]
port 337 nsew signal tristate
rlabel metal2 s 38934 0 38990 1000 6 HI[404]
port 338 nsew signal tristate
rlabel metal2 s 62946 0 63002 1000 6 HI[405]
port 339 nsew signal tristate
rlabel metal2 s 46938 0 46994 1000 6 HI[406]
port 340 nsew signal tristate
rlabel metal2 s 67638 0 67694 1000 6 HI[407]
port 341 nsew signal tristate
rlabel metal2 s 40590 0 40646 1000 6 HI[408]
port 342 nsew signal tristate
rlabel metal2 s 53286 0 53342 1000 6 HI[409]
port 343 nsew signal tristate
rlabel metal2 s 63222 0 63278 1000 6 HI[40]
port 344 nsew signal tristate
rlabel metal2 s 57426 0 57482 1000 6 HI[410]
port 345 nsew signal tristate
rlabel metal2 s 50526 0 50582 1000 6 HI[411]
port 346 nsew signal tristate
rlabel metal2 s 63498 0 63554 1000 6 HI[412]
port 347 nsew signal tristate
rlabel metal2 s 67362 4000 67418 5000 6 HI[413]
port 348 nsew signal tristate
rlabel metal2 s 36174 4000 36230 5000 6 HI[414]
port 349 nsew signal tristate
rlabel metal2 s 36450 4000 36506 5000 6 HI[415]
port 350 nsew signal tristate
rlabel metal2 s 36726 4000 36782 5000 6 HI[416]
port 351 nsew signal tristate
rlabel metal2 s 37002 4000 37058 5000 6 HI[417]
port 352 nsew signal tristate
rlabel metal2 s 37278 4000 37334 5000 6 HI[418]
port 353 nsew signal tristate
rlabel metal2 s 37554 4000 37610 5000 6 HI[419]
port 354 nsew signal tristate
rlabel metal2 s 37830 4000 37886 5000 6 HI[41]
port 355 nsew signal tristate
rlabel metal2 s 38106 4000 38162 5000 6 HI[420]
port 356 nsew signal tristate
rlabel metal2 s 38382 4000 38438 5000 6 HI[421]
port 357 nsew signal tristate
rlabel metal2 s 38658 4000 38714 5000 6 HI[422]
port 358 nsew signal tristate
rlabel metal2 s 38934 4000 38990 5000 6 HI[423]
port 359 nsew signal tristate
rlabel metal2 s 39210 4000 39266 5000 6 HI[424]
port 360 nsew signal tristate
rlabel metal2 s 39486 4000 39542 5000 6 HI[425]
port 361 nsew signal tristate
rlabel metal2 s 39762 4000 39818 5000 6 HI[426]
port 362 nsew signal tristate
rlabel metal2 s 40038 4000 40094 5000 6 HI[427]
port 363 nsew signal tristate
rlabel metal2 s 40314 4000 40370 5000 6 HI[428]
port 364 nsew signal tristate
rlabel metal2 s 40590 4000 40646 5000 6 HI[429]
port 365 nsew signal tristate
rlabel metal2 s 40866 4000 40922 5000 6 HI[42]
port 366 nsew signal tristate
rlabel metal2 s 41142 4000 41198 5000 6 HI[430]
port 367 nsew signal tristate
rlabel metal2 s 41418 4000 41474 5000 6 HI[431]
port 368 nsew signal tristate
rlabel metal2 s 41694 4000 41750 5000 6 HI[432]
port 369 nsew signal tristate
rlabel metal2 s 41970 4000 42026 5000 6 HI[433]
port 370 nsew signal tristate
rlabel metal2 s 42246 4000 42302 5000 6 HI[434]
port 371 nsew signal tristate
rlabel metal2 s 42522 4000 42578 5000 6 HI[435]
port 372 nsew signal tristate
rlabel metal2 s 42798 4000 42854 5000 6 HI[436]
port 373 nsew signal tristate
rlabel metal2 s 43074 4000 43130 5000 6 HI[437]
port 374 nsew signal tristate
rlabel metal2 s 43350 4000 43406 5000 6 HI[438]
port 375 nsew signal tristate
rlabel metal2 s 43626 4000 43682 5000 6 HI[439]
port 376 nsew signal tristate
rlabel metal2 s 43902 4000 43958 5000 6 HI[43]
port 377 nsew signal tristate
rlabel metal2 s 44178 4000 44234 5000 6 HI[440]
port 378 nsew signal tristate
rlabel metal2 s 44454 4000 44510 5000 6 HI[441]
port 379 nsew signal tristate
rlabel metal2 s 44730 4000 44786 5000 6 HI[442]
port 380 nsew signal tristate
rlabel metal2 s 45006 4000 45062 5000 6 HI[443]
port 381 nsew signal tristate
rlabel metal2 s 45282 4000 45338 5000 6 HI[444]
port 382 nsew signal tristate
rlabel metal2 s 45558 4000 45614 5000 6 HI[445]
port 383 nsew signal tristate
rlabel metal2 s 45834 4000 45890 5000 6 HI[446]
port 384 nsew signal tristate
rlabel metal2 s 46110 4000 46166 5000 6 HI[447]
port 385 nsew signal tristate
rlabel metal2 s 46386 4000 46442 5000 6 HI[448]
port 386 nsew signal tristate
rlabel metal2 s 46662 4000 46718 5000 6 HI[449]
port 387 nsew signal tristate
rlabel metal2 s 46938 4000 46994 5000 6 HI[44]
port 388 nsew signal tristate
rlabel metal2 s 47214 4000 47270 5000 6 HI[450]
port 389 nsew signal tristate
rlabel metal2 s 47490 4000 47546 5000 6 HI[451]
port 390 nsew signal tristate
rlabel metal2 s 47766 4000 47822 5000 6 HI[452]
port 391 nsew signal tristate
rlabel metal2 s 48042 4000 48098 5000 6 HI[453]
port 392 nsew signal tristate
rlabel metal2 s 48318 4000 48374 5000 6 HI[454]
port 393 nsew signal tristate
rlabel metal2 s 48594 4000 48650 5000 6 HI[455]
port 394 nsew signal tristate
rlabel metal2 s 48870 4000 48926 5000 6 HI[456]
port 395 nsew signal tristate
rlabel metal2 s 49146 4000 49202 5000 6 HI[457]
port 396 nsew signal tristate
rlabel metal2 s 49422 4000 49478 5000 6 HI[458]
port 397 nsew signal tristate
rlabel metal2 s 49698 4000 49754 5000 6 HI[459]
port 398 nsew signal tristate
rlabel metal2 s 49974 4000 50030 5000 6 HI[45]
port 399 nsew signal tristate
rlabel metal2 s 50250 4000 50306 5000 6 HI[460]
port 400 nsew signal tristate
rlabel metal2 s 50526 4000 50582 5000 6 HI[461]
port 401 nsew signal tristate
rlabel metal2 s 50802 4000 50858 5000 6 HI[46]
port 402 nsew signal tristate
rlabel metal2 s 51078 4000 51134 5000 6 HI[47]
port 403 nsew signal tristate
rlabel metal2 s 51354 4000 51410 5000 6 HI[48]
port 404 nsew signal tristate
rlabel metal2 s 51630 4000 51686 5000 6 HI[49]
port 405 nsew signal tristate
rlabel metal2 s 51906 4000 51962 5000 6 HI[4]
port 406 nsew signal tristate
rlabel metal2 s 52182 4000 52238 5000 6 HI[50]
port 407 nsew signal tristate
rlabel metal2 s 52458 4000 52514 5000 6 HI[51]
port 408 nsew signal tristate
rlabel metal2 s 52734 4000 52790 5000 6 HI[52]
port 409 nsew signal tristate
rlabel metal2 s 53010 4000 53066 5000 6 HI[53]
port 410 nsew signal tristate
rlabel metal2 s 53286 4000 53342 5000 6 HI[54]
port 411 nsew signal tristate
rlabel metal2 s 53562 4000 53618 5000 6 HI[55]
port 412 nsew signal tristate
rlabel metal2 s 53838 4000 53894 5000 6 HI[56]
port 413 nsew signal tristate
rlabel metal2 s 54114 4000 54170 5000 6 HI[57]
port 414 nsew signal tristate
rlabel metal2 s 54390 4000 54446 5000 6 HI[58]
port 415 nsew signal tristate
rlabel metal2 s 54666 4000 54722 5000 6 HI[59]
port 416 nsew signal tristate
rlabel metal2 s 54942 4000 54998 5000 6 HI[5]
port 417 nsew signal tristate
rlabel metal2 s 55218 4000 55274 5000 6 HI[60]
port 418 nsew signal tristate
rlabel metal2 s 55494 4000 55550 5000 6 HI[61]
port 419 nsew signal tristate
rlabel metal2 s 55770 4000 55826 5000 6 HI[62]
port 420 nsew signal tristate
rlabel metal2 s 56046 4000 56102 5000 6 HI[63]
port 421 nsew signal tristate
rlabel metal2 s 56322 4000 56378 5000 6 HI[64]
port 422 nsew signal tristate
rlabel metal2 s 56598 4000 56654 5000 6 HI[65]
port 423 nsew signal tristate
rlabel metal2 s 56874 4000 56930 5000 6 HI[66]
port 424 nsew signal tristate
rlabel metal2 s 57150 4000 57206 5000 6 HI[67]
port 425 nsew signal tristate
rlabel metal2 s 57426 4000 57482 5000 6 HI[68]
port 426 nsew signal tristate
rlabel metal2 s 57702 4000 57758 5000 6 HI[69]
port 427 nsew signal tristate
rlabel metal2 s 57978 4000 58034 5000 6 HI[6]
port 428 nsew signal tristate
rlabel metal2 s 58254 4000 58310 5000 6 HI[70]
port 429 nsew signal tristate
rlabel metal2 s 58530 4000 58586 5000 6 HI[71]
port 430 nsew signal tristate
rlabel metal2 s 58806 4000 58862 5000 6 HI[72]
port 431 nsew signal tristate
rlabel metal2 s 59082 4000 59138 5000 6 HI[73]
port 432 nsew signal tristate
rlabel metal2 s 59358 4000 59414 5000 6 HI[74]
port 433 nsew signal tristate
rlabel metal2 s 59634 4000 59690 5000 6 HI[75]
port 434 nsew signal tristate
rlabel metal2 s 59910 4000 59966 5000 6 HI[76]
port 435 nsew signal tristate
rlabel metal2 s 60186 4000 60242 5000 6 HI[77]
port 436 nsew signal tristate
rlabel metal2 s 60462 4000 60518 5000 6 HI[78]
port 437 nsew signal tristate
rlabel metal2 s 60738 4000 60794 5000 6 HI[79]
port 438 nsew signal tristate
rlabel metal2 s 61014 4000 61070 5000 6 HI[7]
port 439 nsew signal tristate
rlabel metal2 s 61290 4000 61346 5000 6 HI[80]
port 440 nsew signal tristate
rlabel metal2 s 61566 4000 61622 5000 6 HI[81]
port 441 nsew signal tristate
rlabel metal2 s 61842 4000 61898 5000 6 HI[82]
port 442 nsew signal tristate
rlabel metal2 s 62118 4000 62174 5000 6 HI[83]
port 443 nsew signal tristate
rlabel metal2 s 62394 4000 62450 5000 6 HI[84]
port 444 nsew signal tristate
rlabel metal2 s 62670 4000 62726 5000 6 HI[85]
port 445 nsew signal tristate
rlabel metal2 s 62946 4000 63002 5000 6 HI[86]
port 446 nsew signal tristate
rlabel metal2 s 63222 4000 63278 5000 6 HI[87]
port 447 nsew signal tristate
rlabel metal2 s 63498 4000 63554 5000 6 HI[88]
port 448 nsew signal tristate
rlabel metal2 s 63774 4000 63830 5000 6 HI[89]
port 449 nsew signal tristate
rlabel metal2 s 64050 4000 64106 5000 6 HI[8]
port 450 nsew signal tristate
rlabel metal2 s 64326 4000 64382 5000 6 HI[90]
port 451 nsew signal tristate
rlabel metal2 s 64602 4000 64658 5000 6 HI[91]
port 452 nsew signal tristate
rlabel metal2 s 64878 4000 64934 5000 6 HI[92]
port 453 nsew signal tristate
rlabel metal2 s 65154 4000 65210 5000 6 HI[93]
port 454 nsew signal tristate
rlabel metal2 s 65430 4000 65486 5000 6 HI[94]
port 455 nsew signal tristate
rlabel metal2 s 65706 4000 65762 5000 6 HI[95]
port 456 nsew signal tristate
rlabel metal2 s 65982 4000 66038 5000 6 HI[96]
port 457 nsew signal tristate
rlabel metal2 s 66258 4000 66314 5000 6 HI[97]
port 458 nsew signal tristate
rlabel metal2 s 66534 4000 66590 5000 6 HI[98]
port 459 nsew signal tristate
rlabel metal2 s 66810 4000 66866 5000 6 HI[99]
port 460 nsew signal tristate
rlabel metal2 s 67086 4000 67142 5000 6 HI[9]
port 461 nsew signal tristate
rlabel metal2 s 63054 1040 63154 3856 6 vccd1
port 462 nsew power bidirectional
rlabel metal2 s 51054 1040 51154 3856 6 vccd1
port 463 nsew power bidirectional
rlabel metal2 s 39054 1040 39154 3856 6 vccd1
port 464 nsew power bidirectional
rlabel metal2 s 27054 1040 27154 3856 6 vccd1
port 465 nsew power bidirectional
rlabel metal2 s 15054 1040 15154 3856 6 vccd1
port 466 nsew power bidirectional
rlabel metal2 s 3054 1040 3154 3856 6 vccd1
port 467 nsew power bidirectional
rlabel metal3 s 1104 3350 72864 3450 6 vccd1
port 468 nsew power bidirectional
rlabel metal3 s 1104 1190 72864 1290 6 vccd1
port 469 nsew power bidirectional
rlabel metal2 s 69054 1040 69154 3856 6 vssd1
port 470 nsew ground bidirectional
rlabel metal2 s 57054 1040 57154 3856 6 vssd1
port 471 nsew ground bidirectional
rlabel metal2 s 45054 1040 45154 3856 6 vssd1
port 472 nsew ground bidirectional
rlabel metal2 s 33054 1040 33154 3856 6 vssd1
port 473 nsew ground bidirectional
rlabel metal2 s 21054 1040 21154 3856 6 vssd1
port 474 nsew ground bidirectional
rlabel metal2 s 9054 1040 9154 3856 6 vssd1
port 475 nsew ground bidirectional
rlabel metal3 s 1104 2270 72864 2370 6 vssd1
port 476 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 74000 5000
<< end >>
