magic
tech sky130A
magscale 1 2
timestamp 1605064556
<< viali >>
rect 2605 6409 2639 6443
rect 1593 6341 1627 6375
rect 2053 6273 2087 6307
rect 2329 6205 2363 6239
rect 4261 6205 4295 6239
rect 4997 6205 5031 6239
rect 3709 5729 3743 5763
rect 4905 5593 4939 5627
rect 5641 5525 5675 5559
rect 2881 5253 2915 5287
rect 5641 5185 5675 5219
rect 3157 5117 3191 5151
rect 1685 4573 1719 4607
rect 2237 4505 2271 4539
rect 1961 4437 1995 4471
rect 3065 4437 3099 4471
rect 3617 4233 3651 4267
rect 4261 4233 4295 4267
rect 1593 4165 1627 4199
rect 5549 4165 5583 4199
rect 2881 4097 2915 4131
rect 3893 4097 3927 4131
rect 4629 4029 4663 4063
rect 2237 3553 2271 3587
rect 1961 3417 1995 3451
rect 1593 3349 1627 3383
rect 1593 3145 1627 3179
rect 2329 3145 2363 3179
rect 5365 3145 5399 3179
rect 1869 2465 1903 2499
rect 4261 2465 4295 2499
rect 5457 2465 5491 2499
<< metal1 >>
rect 3510 7624 3516 7676
rect 3568 7664 3574 7676
rect 5442 7664 5448 7676
rect 3568 7636 5448 7664
rect 3568 7624 3574 7636
rect 5442 7624 5448 7636
rect 5500 7624 5506 7676
rect 1104 7098 5980 7120
rect 1104 7046 2607 7098
rect 2659 7046 2671 7098
rect 2723 7046 2735 7098
rect 2787 7046 2799 7098
rect 2851 7046 4232 7098
rect 4284 7046 4296 7098
rect 4348 7046 4360 7098
rect 4412 7046 4424 7098
rect 4476 7046 5980 7098
rect 1104 7024 5980 7046
rect 1104 6554 5980 6576
rect 1104 6502 1794 6554
rect 1846 6502 1858 6554
rect 1910 6502 1922 6554
rect 1974 6502 1986 6554
rect 2038 6502 3420 6554
rect 3472 6502 3484 6554
rect 3536 6502 3548 6554
rect 3600 6502 3612 6554
rect 3664 6502 5045 6554
rect 5097 6502 5109 6554
rect 5161 6502 5173 6554
rect 5225 6502 5237 6554
rect 5289 6502 5980 6554
rect 1104 6480 5980 6502
rect 2593 6443 2651 6449
rect 2593 6409 2605 6443
rect 2639 6440 2651 6443
rect 4062 6440 4068 6452
rect 2639 6412 4068 6440
rect 2639 6409 2651 6412
rect 2593 6403 2651 6409
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 1581 6375 1639 6381
rect 1581 6341 1593 6375
rect 1627 6372 1639 6375
rect 3142 6372 3148 6384
rect 1627 6344 3148 6372
rect 1627 6341 1639 6344
rect 1581 6335 1639 6341
rect 3142 6332 3148 6344
rect 3200 6332 3206 6384
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6304 2099 6307
rect 4062 6304 4068 6316
rect 2087 6276 4068 6304
rect 2087 6273 2099 6276
rect 2041 6267 2099 6273
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 2314 6236 2320 6248
rect 2275 6208 2320 6236
rect 2314 6196 2320 6208
rect 2372 6196 2378 6248
rect 4249 6239 4307 6245
rect 4249 6205 4261 6239
rect 4295 6236 4307 6239
rect 4522 6236 4528 6248
rect 4295 6208 4528 6236
rect 4295 6205 4307 6208
rect 4249 6199 4307 6205
rect 4522 6196 4528 6208
rect 4580 6196 4586 6248
rect 4985 6239 5043 6245
rect 4985 6205 4997 6239
rect 5031 6236 5043 6239
rect 5718 6236 5724 6248
rect 5031 6208 5724 6236
rect 5031 6205 5043 6208
rect 4985 6199 5043 6205
rect 5718 6196 5724 6208
rect 5776 6196 5782 6248
rect 1104 6010 5980 6032
rect 1104 5958 2607 6010
rect 2659 5958 2671 6010
rect 2723 5958 2735 6010
rect 2787 5958 2799 6010
rect 2851 5958 4232 6010
rect 4284 5958 4296 6010
rect 4348 5958 4360 6010
rect 4412 5958 4424 6010
rect 4476 5958 5980 6010
rect 1104 5936 5980 5958
rect 3697 5763 3755 5769
rect 3697 5729 3709 5763
rect 3743 5760 3755 5763
rect 5902 5760 5908 5772
rect 3743 5732 5908 5760
rect 3743 5729 3755 5732
rect 3697 5723 3755 5729
rect 5902 5720 5908 5732
rect 5960 5720 5966 5772
rect 4893 5627 4951 5633
rect 4893 5593 4905 5627
rect 4939 5624 4951 5627
rect 6454 5624 6460 5636
rect 4939 5596 6460 5624
rect 4939 5593 4951 5596
rect 4893 5587 4951 5593
rect 6454 5584 6460 5596
rect 6512 5584 6518 5636
rect 5626 5556 5632 5568
rect 5587 5528 5632 5556
rect 5626 5516 5632 5528
rect 5684 5516 5690 5568
rect 1104 5466 5980 5488
rect 1104 5414 1794 5466
rect 1846 5414 1858 5466
rect 1910 5414 1922 5466
rect 1974 5414 1986 5466
rect 2038 5414 3420 5466
rect 3472 5414 3484 5466
rect 3536 5414 3548 5466
rect 3600 5414 3612 5466
rect 3664 5414 5045 5466
rect 5097 5414 5109 5466
rect 5161 5414 5173 5466
rect 5225 5414 5237 5466
rect 5289 5414 5980 5466
rect 1104 5392 5980 5414
rect 2498 5312 2504 5364
rect 2556 5352 2562 5364
rect 5626 5352 5632 5364
rect 2556 5324 5632 5352
rect 2556 5312 2562 5324
rect 5626 5312 5632 5324
rect 5684 5312 5690 5364
rect 2869 5287 2927 5293
rect 2869 5253 2881 5287
rect 2915 5284 2927 5287
rect 3970 5284 3976 5296
rect 2915 5256 3976 5284
rect 2915 5253 2927 5256
rect 2869 5247 2927 5253
rect 3970 5244 3976 5256
rect 4028 5244 4034 5296
rect 1302 5176 1308 5228
rect 1360 5216 1366 5228
rect 5629 5219 5687 5225
rect 5629 5216 5641 5219
rect 1360 5188 5641 5216
rect 1360 5176 1366 5188
rect 5629 5185 5641 5188
rect 5675 5185 5687 5219
rect 5629 5179 5687 5185
rect 3145 5151 3203 5157
rect 3145 5117 3157 5151
rect 3191 5148 3203 5151
rect 6362 5148 6368 5160
rect 3191 5120 6368 5148
rect 3191 5117 3203 5120
rect 3145 5111 3203 5117
rect 6362 5108 6368 5120
rect 6420 5108 6426 5160
rect 1104 4922 5980 4944
rect 1104 4870 2607 4922
rect 2659 4870 2671 4922
rect 2723 4870 2735 4922
rect 2787 4870 2799 4922
rect 2851 4870 4232 4922
rect 4284 4870 4296 4922
rect 4348 4870 4360 4922
rect 4412 4870 4424 4922
rect 4476 4870 5980 4922
rect 1104 4848 5980 4870
rect 2130 4700 2136 4752
rect 2188 4740 2194 4752
rect 4798 4740 4804 4752
rect 2188 4712 4804 4740
rect 2188 4700 2194 4712
rect 4798 4700 4804 4712
rect 4856 4700 4862 4752
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4604 1731 4607
rect 4706 4604 4712 4616
rect 1719 4576 4712 4604
rect 1719 4573 1731 4576
rect 1673 4567 1731 4573
rect 4706 4564 4712 4576
rect 4764 4564 4770 4616
rect 2225 4539 2283 4545
rect 2225 4505 2237 4539
rect 2271 4536 2283 4539
rect 4890 4536 4896 4548
rect 2271 4508 4896 4536
rect 2271 4505 2283 4508
rect 2225 4499 2283 4505
rect 4890 4496 4896 4508
rect 4948 4496 4954 4548
rect 1394 4428 1400 4480
rect 1452 4468 1458 4480
rect 1949 4471 2007 4477
rect 1949 4468 1961 4471
rect 1452 4440 1961 4468
rect 1452 4428 1458 4440
rect 1949 4437 1961 4440
rect 1995 4437 2007 4471
rect 3050 4468 3056 4480
rect 3011 4440 3056 4468
rect 1949 4431 2007 4437
rect 3050 4428 3056 4440
rect 3108 4428 3114 4480
rect 1104 4378 5980 4400
rect 1104 4326 1794 4378
rect 1846 4326 1858 4378
rect 1910 4326 1922 4378
rect 1974 4326 1986 4378
rect 2038 4326 3420 4378
rect 3472 4326 3484 4378
rect 3536 4326 3548 4378
rect 3600 4326 3612 4378
rect 3664 4326 5045 4378
rect 5097 4326 5109 4378
rect 5161 4326 5173 4378
rect 5225 4326 5237 4378
rect 5289 4326 5980 4378
rect 1104 4304 5980 4326
rect 3605 4267 3663 4273
rect 3605 4233 3617 4267
rect 3651 4264 3663 4267
rect 3786 4264 3792 4276
rect 3651 4236 3792 4264
rect 3651 4233 3663 4236
rect 3605 4227 3663 4233
rect 3786 4224 3792 4236
rect 3844 4224 3850 4276
rect 3878 4224 3884 4276
rect 3936 4224 3942 4276
rect 4249 4267 4307 4273
rect 4249 4233 4261 4267
rect 4295 4264 4307 4267
rect 4614 4264 4620 4276
rect 4295 4236 4620 4264
rect 4295 4233 4307 4236
rect 4249 4227 4307 4233
rect 4614 4224 4620 4236
rect 4672 4224 4678 4276
rect 1578 4196 1584 4208
rect 1539 4168 1584 4196
rect 1578 4156 1584 4168
rect 1636 4156 1642 4208
rect 3896 4196 3924 4224
rect 5537 4199 5595 4205
rect 5537 4196 5549 4199
rect 3896 4168 5549 4196
rect 5537 4165 5549 4168
rect 5583 4165 5595 4199
rect 5537 4159 5595 4165
rect 1302 4088 1308 4140
rect 1360 4128 1366 4140
rect 2869 4131 2927 4137
rect 2869 4128 2881 4131
rect 1360 4100 2881 4128
rect 1360 4088 1366 4100
rect 2869 4097 2881 4100
rect 2915 4097 2927 4131
rect 2869 4091 2927 4097
rect 3142 4088 3148 4140
rect 3200 4128 3206 4140
rect 3881 4131 3939 4137
rect 3881 4128 3893 4131
rect 3200 4100 3893 4128
rect 3200 4088 3206 4100
rect 3881 4097 3893 4100
rect 3927 4097 3939 4131
rect 3881 4091 3939 4097
rect 2406 4020 2412 4072
rect 2464 4060 2470 4072
rect 4522 4060 4528 4072
rect 2464 4032 4528 4060
rect 2464 4020 2470 4032
rect 4522 4020 4528 4032
rect 4580 4020 4586 4072
rect 4617 4063 4675 4069
rect 4617 4029 4629 4063
rect 4663 4029 4675 4063
rect 4617 4023 4675 4029
rect 1118 3952 1124 4004
rect 1176 3992 1182 4004
rect 3050 3992 3056 4004
rect 1176 3964 3056 3992
rect 1176 3952 1182 3964
rect 3050 3952 3056 3964
rect 3108 3952 3114 4004
rect 566 3884 572 3936
rect 624 3924 630 3936
rect 4632 3924 4660 4023
rect 624 3896 4660 3924
rect 624 3884 630 3896
rect 1104 3834 5980 3856
rect 1104 3782 2607 3834
rect 2659 3782 2671 3834
rect 2723 3782 2735 3834
rect 2787 3782 2799 3834
rect 2851 3782 4232 3834
rect 4284 3782 4296 3834
rect 4348 3782 4360 3834
rect 4412 3782 4424 3834
rect 4476 3782 5980 3834
rect 1104 3760 5980 3782
rect 3234 3720 3240 3732
rect 2240 3692 3240 3720
rect 2240 3593 2268 3692
rect 3234 3680 3240 3692
rect 3292 3680 3298 3732
rect 2225 3587 2283 3593
rect 2225 3553 2237 3587
rect 2271 3553 2283 3587
rect 2225 3547 2283 3553
rect 1949 3451 2007 3457
rect 1949 3417 1961 3451
rect 1995 3448 2007 3451
rect 2958 3448 2964 3460
rect 1995 3420 2964 3448
rect 1995 3417 2007 3420
rect 1949 3411 2007 3417
rect 2958 3408 2964 3420
rect 3016 3408 3022 3460
rect 1581 3383 1639 3389
rect 1581 3349 1593 3383
rect 1627 3380 1639 3383
rect 1670 3380 1676 3392
rect 1627 3352 1676 3380
rect 1627 3349 1639 3352
rect 1581 3343 1639 3349
rect 1670 3340 1676 3352
rect 1728 3340 1734 3392
rect 1104 3290 5980 3312
rect 1104 3238 1794 3290
rect 1846 3238 1858 3290
rect 1910 3238 1922 3290
rect 1974 3238 1986 3290
rect 2038 3238 3420 3290
rect 3472 3238 3484 3290
rect 3536 3238 3548 3290
rect 3600 3238 3612 3290
rect 3664 3238 5045 3290
rect 5097 3238 5109 3290
rect 5161 3238 5173 3290
rect 5225 3238 5237 3290
rect 5289 3238 5980 3290
rect 1104 3216 5980 3238
rect 1486 3136 1492 3188
rect 1544 3176 1550 3188
rect 1581 3179 1639 3185
rect 1581 3176 1593 3179
rect 1544 3148 1593 3176
rect 1544 3136 1550 3148
rect 1581 3145 1593 3148
rect 1627 3145 1639 3179
rect 1581 3139 1639 3145
rect 2317 3179 2375 3185
rect 2317 3145 2329 3179
rect 2363 3176 2375 3179
rect 2866 3176 2872 3188
rect 2363 3148 2872 3176
rect 2363 3145 2375 3148
rect 2317 3139 2375 3145
rect 2866 3136 2872 3148
rect 2924 3136 2930 3188
rect 5350 3176 5356 3188
rect 5311 3148 5356 3176
rect 5350 3136 5356 3148
rect 5408 3136 5414 3188
rect 2314 3000 2320 3052
rect 2372 3040 2378 3052
rect 3786 3040 3792 3052
rect 2372 3012 3792 3040
rect 2372 3000 2378 3012
rect 3786 3000 3792 3012
rect 3844 3000 3850 3052
rect 1104 2746 5980 2768
rect 1104 2694 2607 2746
rect 2659 2694 2671 2746
rect 2723 2694 2735 2746
rect 2787 2694 2799 2746
rect 2851 2694 4232 2746
rect 4284 2694 4296 2746
rect 4348 2694 4360 2746
rect 4412 2694 4424 2746
rect 4476 2694 5980 2746
rect 1104 2672 5980 2694
rect 1857 2499 1915 2505
rect 1857 2465 1869 2499
rect 1903 2496 1915 2499
rect 3050 2496 3056 2508
rect 1903 2468 3056 2496
rect 1903 2465 1915 2468
rect 1857 2459 1915 2465
rect 3050 2456 3056 2468
rect 3108 2456 3114 2508
rect 4249 2499 4307 2505
rect 4249 2465 4261 2499
rect 4295 2496 4307 2499
rect 4798 2496 4804 2508
rect 4295 2468 4804 2496
rect 4295 2465 4307 2468
rect 4249 2459 4307 2465
rect 4798 2456 4804 2468
rect 4856 2456 4862 2508
rect 5442 2496 5448 2508
rect 5403 2468 5448 2496
rect 5442 2456 5448 2468
rect 5500 2456 5506 2508
rect 1104 2202 5980 2224
rect 1104 2150 1794 2202
rect 1846 2150 1858 2202
rect 1910 2150 1922 2202
rect 1974 2150 1986 2202
rect 2038 2150 3420 2202
rect 3472 2150 3484 2202
rect 3536 2150 3548 2202
rect 3600 2150 3612 2202
rect 3664 2150 5045 2202
rect 5097 2150 5109 2202
rect 5161 2150 5173 2202
rect 5225 2150 5237 2202
rect 5289 2150 5980 2202
rect 1104 2128 5980 2150
<< via1 >>
rect 3516 7624 3568 7676
rect 5448 7624 5500 7676
rect 2607 7046 2659 7098
rect 2671 7046 2723 7098
rect 2735 7046 2787 7098
rect 2799 7046 2851 7098
rect 4232 7046 4284 7098
rect 4296 7046 4348 7098
rect 4360 7046 4412 7098
rect 4424 7046 4476 7098
rect 1794 6502 1846 6554
rect 1858 6502 1910 6554
rect 1922 6502 1974 6554
rect 1986 6502 2038 6554
rect 3420 6502 3472 6554
rect 3484 6502 3536 6554
rect 3548 6502 3600 6554
rect 3612 6502 3664 6554
rect 5045 6502 5097 6554
rect 5109 6502 5161 6554
rect 5173 6502 5225 6554
rect 5237 6502 5289 6554
rect 4068 6400 4120 6452
rect 3148 6332 3200 6384
rect 4068 6264 4120 6316
rect 2320 6239 2372 6248
rect 2320 6205 2329 6239
rect 2329 6205 2363 6239
rect 2363 6205 2372 6239
rect 2320 6196 2372 6205
rect 4528 6196 4580 6248
rect 5724 6196 5776 6248
rect 2607 5958 2659 6010
rect 2671 5958 2723 6010
rect 2735 5958 2787 6010
rect 2799 5958 2851 6010
rect 4232 5958 4284 6010
rect 4296 5958 4348 6010
rect 4360 5958 4412 6010
rect 4424 5958 4476 6010
rect 5908 5720 5960 5772
rect 6460 5584 6512 5636
rect 5632 5559 5684 5568
rect 5632 5525 5641 5559
rect 5641 5525 5675 5559
rect 5675 5525 5684 5559
rect 5632 5516 5684 5525
rect 1794 5414 1846 5466
rect 1858 5414 1910 5466
rect 1922 5414 1974 5466
rect 1986 5414 2038 5466
rect 3420 5414 3472 5466
rect 3484 5414 3536 5466
rect 3548 5414 3600 5466
rect 3612 5414 3664 5466
rect 5045 5414 5097 5466
rect 5109 5414 5161 5466
rect 5173 5414 5225 5466
rect 5237 5414 5289 5466
rect 2504 5312 2556 5364
rect 5632 5312 5684 5364
rect 3976 5244 4028 5296
rect 1308 5176 1360 5228
rect 6368 5108 6420 5160
rect 2607 4870 2659 4922
rect 2671 4870 2723 4922
rect 2735 4870 2787 4922
rect 2799 4870 2851 4922
rect 4232 4870 4284 4922
rect 4296 4870 4348 4922
rect 4360 4870 4412 4922
rect 4424 4870 4476 4922
rect 2136 4700 2188 4752
rect 4804 4700 4856 4752
rect 4712 4564 4764 4616
rect 4896 4496 4948 4548
rect 1400 4428 1452 4480
rect 3056 4471 3108 4480
rect 3056 4437 3065 4471
rect 3065 4437 3099 4471
rect 3099 4437 3108 4471
rect 3056 4428 3108 4437
rect 1794 4326 1846 4378
rect 1858 4326 1910 4378
rect 1922 4326 1974 4378
rect 1986 4326 2038 4378
rect 3420 4326 3472 4378
rect 3484 4326 3536 4378
rect 3548 4326 3600 4378
rect 3612 4326 3664 4378
rect 5045 4326 5097 4378
rect 5109 4326 5161 4378
rect 5173 4326 5225 4378
rect 5237 4326 5289 4378
rect 3792 4224 3844 4276
rect 3884 4224 3936 4276
rect 4620 4224 4672 4276
rect 1584 4199 1636 4208
rect 1584 4165 1593 4199
rect 1593 4165 1627 4199
rect 1627 4165 1636 4199
rect 1584 4156 1636 4165
rect 1308 4088 1360 4140
rect 3148 4088 3200 4140
rect 2412 4020 2464 4072
rect 4528 4020 4580 4072
rect 1124 3952 1176 4004
rect 3056 3952 3108 4004
rect 572 3884 624 3936
rect 2607 3782 2659 3834
rect 2671 3782 2723 3834
rect 2735 3782 2787 3834
rect 2799 3782 2851 3834
rect 4232 3782 4284 3834
rect 4296 3782 4348 3834
rect 4360 3782 4412 3834
rect 4424 3782 4476 3834
rect 3240 3680 3292 3732
rect 2964 3408 3016 3460
rect 1676 3340 1728 3392
rect 1794 3238 1846 3290
rect 1858 3238 1910 3290
rect 1922 3238 1974 3290
rect 1986 3238 2038 3290
rect 3420 3238 3472 3290
rect 3484 3238 3536 3290
rect 3548 3238 3600 3290
rect 3612 3238 3664 3290
rect 5045 3238 5097 3290
rect 5109 3238 5161 3290
rect 5173 3238 5225 3290
rect 5237 3238 5289 3290
rect 1492 3136 1544 3188
rect 2872 3136 2924 3188
rect 5356 3179 5408 3188
rect 5356 3145 5365 3179
rect 5365 3145 5399 3179
rect 5399 3145 5408 3179
rect 5356 3136 5408 3145
rect 2320 3000 2372 3052
rect 3792 3000 3844 3052
rect 2607 2694 2659 2746
rect 2671 2694 2723 2746
rect 2735 2694 2787 2746
rect 2799 2694 2851 2746
rect 4232 2694 4284 2746
rect 4296 2694 4348 2746
rect 4360 2694 4412 2746
rect 4424 2694 4476 2746
rect 3056 2456 3108 2508
rect 4804 2456 4856 2508
rect 5448 2499 5500 2508
rect 5448 2465 5457 2499
rect 5457 2465 5491 2499
rect 5491 2465 5500 2499
rect 5448 2456 5500 2465
rect 1794 2150 1846 2202
rect 1858 2150 1910 2202
rect 1922 2150 1974 2202
rect 1986 2150 2038 2202
rect 3420 2150 3472 2202
rect 3484 2150 3536 2202
rect 3548 2150 3600 2202
rect 3612 2150 3664 2202
rect 5045 2150 5097 2202
rect 5109 2150 5161 2202
rect 5173 2150 5225 2202
rect 5237 2150 5289 2202
<< metal2 >>
rect 570 8453 626 9253
rect 1306 8453 1362 9253
rect 1858 8453 1914 9253
rect 2594 8453 2650 9253
rect 3330 8453 3386 9253
rect 3882 8453 3938 9253
rect 4618 8453 4674 9253
rect 5170 8453 5226 9253
rect 5906 8453 5962 9253
rect 6458 8453 6514 9253
rect 1320 5234 1348 8453
rect 1872 6746 1900 8453
rect 2608 7290 2636 8453
rect 2516 7262 2636 7290
rect 1872 6718 2176 6746
rect 1768 6556 2064 6576
rect 1824 6554 1848 6556
rect 1904 6554 1928 6556
rect 1984 6554 2008 6556
rect 1846 6502 1848 6554
rect 1910 6502 1922 6554
rect 1984 6502 1986 6554
rect 1824 6500 1848 6502
rect 1904 6500 1928 6502
rect 1984 6500 2008 6502
rect 1768 6480 2064 6500
rect 1768 5468 2064 5488
rect 1824 5466 1848 5468
rect 1904 5466 1928 5468
rect 1984 5466 2008 5468
rect 1846 5414 1848 5466
rect 1910 5414 1922 5466
rect 1984 5414 1986 5466
rect 1824 5412 1848 5414
rect 1904 5412 1928 5414
rect 1984 5412 2008 5414
rect 1768 5392 2064 5412
rect 1308 5228 1360 5234
rect 1308 5170 1360 5176
rect 2148 4758 2176 6718
rect 2320 6248 2372 6254
rect 2320 6190 2372 6196
rect 2136 4752 2188 4758
rect 1490 4720 1546 4729
rect 2136 4694 2188 4700
rect 1490 4655 1546 4664
rect 1400 4480 1452 4486
rect 1400 4422 1452 4428
rect 1308 4140 1360 4146
rect 1308 4082 1360 4088
rect 1124 4004 1176 4010
rect 1124 3946 1176 3952
rect 572 3936 624 3942
rect 572 3878 624 3884
rect 584 800 612 3878
rect 1136 800 1164 3946
rect 1320 1737 1348 4082
rect 1412 2825 1440 4422
rect 1504 3194 1532 4655
rect 1768 4380 2064 4400
rect 1824 4378 1848 4380
rect 1904 4378 1928 4380
rect 1984 4378 2008 4380
rect 1846 4326 1848 4378
rect 1910 4326 1922 4378
rect 1984 4326 1986 4378
rect 1824 4324 1848 4326
rect 1904 4324 1928 4326
rect 1984 4324 2008 4326
rect 1768 4304 2064 4324
rect 1584 4208 1636 4214
rect 1584 4150 1636 4156
rect 1596 3641 1624 4150
rect 1582 3632 1638 3641
rect 1582 3567 1638 3576
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1492 3188 1544 3194
rect 1492 3130 1544 3136
rect 1398 2816 1454 2825
rect 1398 2751 1454 2760
rect 1306 1728 1362 1737
rect 1306 1663 1362 1672
rect 1688 1442 1716 3334
rect 1768 3292 2064 3312
rect 1824 3290 1848 3292
rect 1904 3290 1928 3292
rect 1984 3290 2008 3292
rect 1846 3238 1848 3290
rect 1910 3238 1922 3290
rect 1984 3238 1986 3290
rect 1824 3236 1848 3238
rect 1904 3236 1928 3238
rect 1984 3236 2008 3238
rect 1768 3216 2064 3236
rect 2332 3058 2360 6190
rect 2516 5370 2544 7262
rect 2581 7100 2877 7120
rect 2637 7098 2661 7100
rect 2717 7098 2741 7100
rect 2797 7098 2821 7100
rect 2659 7046 2661 7098
rect 2723 7046 2735 7098
rect 2797 7046 2799 7098
rect 2637 7044 2661 7046
rect 2717 7044 2741 7046
rect 2797 7044 2821 7046
rect 2581 7024 2877 7044
rect 3344 6882 3372 8453
rect 3514 7712 3570 7721
rect 3514 7647 3516 7656
rect 3568 7647 3570 7656
rect 3516 7618 3568 7624
rect 2976 6854 3372 6882
rect 2581 6012 2877 6032
rect 2637 6010 2661 6012
rect 2717 6010 2741 6012
rect 2797 6010 2821 6012
rect 2659 5958 2661 6010
rect 2723 5958 2735 6010
rect 2797 5958 2799 6010
rect 2637 5956 2661 5958
rect 2717 5956 2741 5958
rect 2797 5956 2821 5958
rect 2581 5936 2877 5956
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2581 4924 2877 4944
rect 2637 4922 2661 4924
rect 2717 4922 2741 4924
rect 2797 4922 2821 4924
rect 2659 4870 2661 4922
rect 2723 4870 2735 4922
rect 2797 4870 2799 4922
rect 2637 4868 2661 4870
rect 2717 4868 2741 4870
rect 2797 4868 2821 4870
rect 2581 4848 2877 4868
rect 2412 4072 2464 4078
rect 2412 4014 2464 4020
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 1768 2204 2064 2224
rect 1824 2202 1848 2204
rect 1904 2202 1928 2204
rect 1984 2202 2008 2204
rect 1846 2150 1848 2202
rect 1910 2150 1922 2202
rect 1984 2150 1986 2202
rect 1824 2148 1848 2150
rect 1904 2148 1928 2150
rect 1984 2148 2008 2150
rect 1768 2128 2064 2148
rect 1688 1414 1900 1442
rect 1872 800 1900 1414
rect 2424 800 2452 4014
rect 2581 3836 2877 3856
rect 2637 3834 2661 3836
rect 2717 3834 2741 3836
rect 2797 3834 2821 3836
rect 2659 3782 2661 3834
rect 2723 3782 2735 3834
rect 2797 3782 2799 3834
rect 2637 3780 2661 3782
rect 2717 3780 2741 3782
rect 2797 3780 2821 3782
rect 2581 3760 2877 3780
rect 2976 3618 3004 6854
rect 3238 6760 3294 6769
rect 3238 6695 3294 6704
rect 3148 6384 3200 6390
rect 3148 6326 3200 6332
rect 3160 4593 3188 6326
rect 3146 4584 3202 4593
rect 3146 4519 3202 4528
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 3068 4010 3096 4422
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3056 4004 3108 4010
rect 3056 3946 3108 3952
rect 2884 3590 3004 3618
rect 3054 3632 3110 3641
rect 2884 3194 2912 3590
rect 3054 3567 3110 3576
rect 2964 3460 3016 3466
rect 2964 3402 3016 3408
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 2581 2748 2877 2768
rect 2637 2746 2661 2748
rect 2717 2746 2741 2748
rect 2797 2746 2821 2748
rect 2659 2694 2661 2746
rect 2723 2694 2735 2746
rect 2797 2694 2799 2746
rect 2637 2692 2661 2694
rect 2717 2692 2741 2694
rect 2797 2692 2821 2694
rect 2581 2672 2877 2692
rect 2976 2553 3004 3402
rect 2962 2544 3018 2553
rect 3068 2514 3096 3567
rect 2962 2479 3018 2488
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 3160 800 3188 4082
rect 3252 3738 3280 6695
rect 3394 6556 3690 6576
rect 3450 6554 3474 6556
rect 3530 6554 3554 6556
rect 3610 6554 3634 6556
rect 3472 6502 3474 6554
rect 3536 6502 3548 6554
rect 3610 6502 3612 6554
rect 3450 6500 3474 6502
rect 3530 6500 3554 6502
rect 3610 6500 3634 6502
rect 3394 6480 3690 6500
rect 3394 5468 3690 5488
rect 3450 5466 3474 5468
rect 3530 5466 3554 5468
rect 3610 5466 3634 5468
rect 3472 5414 3474 5466
rect 3536 5414 3548 5466
rect 3610 5414 3612 5466
rect 3450 5412 3474 5414
rect 3530 5412 3554 5414
rect 3610 5412 3634 5414
rect 3394 5392 3690 5412
rect 3790 5264 3846 5273
rect 3790 5199 3846 5208
rect 3394 4380 3690 4400
rect 3450 4378 3474 4380
rect 3530 4378 3554 4380
rect 3610 4378 3634 4380
rect 3472 4326 3474 4378
rect 3536 4326 3548 4378
rect 3610 4326 3612 4378
rect 3450 4324 3474 4326
rect 3530 4324 3554 4326
rect 3610 4324 3634 4326
rect 3394 4304 3690 4324
rect 3804 4282 3832 5199
rect 3896 4282 3924 8453
rect 4066 7440 4122 7449
rect 4066 7375 4122 7384
rect 4080 6458 4108 7375
rect 4206 7100 4502 7120
rect 4262 7098 4286 7100
rect 4342 7098 4366 7100
rect 4422 7098 4446 7100
rect 4284 7046 4286 7098
rect 4348 7046 4360 7098
rect 4422 7046 4424 7098
rect 4262 7044 4286 7046
rect 4342 7044 4366 7046
rect 4422 7044 4446 7046
rect 4206 7024 4502 7044
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4066 6352 4122 6361
rect 4066 6287 4068 6296
rect 4120 6287 4122 6296
rect 4068 6258 4120 6264
rect 4528 6248 4580 6254
rect 4528 6190 4580 6196
rect 4206 6012 4502 6032
rect 4262 6010 4286 6012
rect 4342 6010 4366 6012
rect 4422 6010 4446 6012
rect 4284 5958 4286 6010
rect 4348 5958 4360 6010
rect 4422 5958 4424 6010
rect 4262 5956 4286 5958
rect 4342 5956 4366 5958
rect 4422 5956 4446 5958
rect 4206 5936 4502 5956
rect 3976 5296 4028 5302
rect 3976 5238 4028 5244
rect 3792 4276 3844 4282
rect 3792 4218 3844 4224
rect 3884 4276 3936 4282
rect 3884 4218 3936 4224
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3394 3292 3690 3312
rect 3450 3290 3474 3292
rect 3530 3290 3554 3292
rect 3610 3290 3634 3292
rect 3472 3238 3474 3290
rect 3536 3238 3548 3290
rect 3610 3238 3612 3290
rect 3450 3236 3474 3238
rect 3530 3236 3554 3238
rect 3610 3236 3634 3238
rect 3394 3216 3690 3236
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 3394 2204 3690 2224
rect 3450 2202 3474 2204
rect 3530 2202 3554 2204
rect 3610 2202 3634 2204
rect 3472 2150 3474 2202
rect 3536 2150 3548 2202
rect 3610 2150 3612 2202
rect 3450 2148 3474 2150
rect 3530 2148 3554 2150
rect 3610 2148 3634 2150
rect 3394 2128 3690 2148
rect 3804 1442 3832 2994
rect 3988 1465 4016 5238
rect 4206 4924 4502 4944
rect 4262 4922 4286 4924
rect 4342 4922 4366 4924
rect 4422 4922 4446 4924
rect 4284 4870 4286 4922
rect 4348 4870 4360 4922
rect 4422 4870 4424 4922
rect 4262 4868 4286 4870
rect 4342 4868 4366 4870
rect 4422 4868 4446 4870
rect 4206 4848 4502 4868
rect 4540 4078 4568 6190
rect 4632 4282 4660 8453
rect 5184 6746 5212 8453
rect 5448 7676 5500 7682
rect 5448 7618 5500 7624
rect 5184 6718 5396 6746
rect 5019 6556 5315 6576
rect 5075 6554 5099 6556
rect 5155 6554 5179 6556
rect 5235 6554 5259 6556
rect 5097 6502 5099 6554
rect 5161 6502 5173 6554
rect 5235 6502 5237 6554
rect 5075 6500 5099 6502
rect 5155 6500 5179 6502
rect 5235 6500 5259 6502
rect 5019 6480 5315 6500
rect 5019 5468 5315 5488
rect 5075 5466 5099 5468
rect 5155 5466 5179 5468
rect 5235 5466 5259 5468
rect 5097 5414 5099 5466
rect 5161 5414 5173 5466
rect 5235 5414 5237 5466
rect 5075 5412 5099 5414
rect 5155 5412 5179 5414
rect 5235 5412 5259 5414
rect 5019 5392 5315 5412
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4206 3836 4502 3856
rect 4262 3834 4286 3836
rect 4342 3834 4366 3836
rect 4422 3834 4446 3836
rect 4284 3782 4286 3834
rect 4348 3782 4360 3834
rect 4422 3782 4424 3834
rect 4262 3780 4286 3782
rect 4342 3780 4366 3782
rect 4422 3780 4446 3782
rect 4206 3760 4502 3780
rect 4206 2748 4502 2768
rect 4262 2746 4286 2748
rect 4342 2746 4366 2748
rect 4422 2746 4446 2748
rect 4284 2694 4286 2746
rect 4348 2694 4360 2746
rect 4422 2694 4424 2746
rect 4262 2692 4286 2694
rect 4342 2692 4366 2694
rect 4422 2692 4446 2694
rect 4206 2672 4502 2692
rect 3712 1414 3832 1442
rect 3974 1456 4030 1465
rect 3712 800 3740 1414
rect 3974 1391 4030 1400
rect 4724 1306 4752 4558
rect 4816 2514 4844 4694
rect 4896 4548 4948 4554
rect 4896 4490 4948 4496
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 4908 1442 4936 4490
rect 5019 4380 5315 4400
rect 5075 4378 5099 4380
rect 5155 4378 5179 4380
rect 5235 4378 5259 4380
rect 5097 4326 5099 4378
rect 5161 4326 5173 4378
rect 5235 4326 5237 4378
rect 5075 4324 5099 4326
rect 5155 4324 5179 4326
rect 5235 4324 5259 4326
rect 5019 4304 5315 4324
rect 5019 3292 5315 3312
rect 5075 3290 5099 3292
rect 5155 3290 5179 3292
rect 5235 3290 5259 3292
rect 5097 3238 5099 3290
rect 5161 3238 5173 3290
rect 5235 3238 5237 3290
rect 5075 3236 5099 3238
rect 5155 3236 5179 3238
rect 5235 3236 5259 3238
rect 5019 3216 5315 3236
rect 5368 3194 5396 6718
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5460 2514 5488 7618
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5644 5370 5672 5510
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5019 2204 5315 2224
rect 5075 2202 5099 2204
rect 5155 2202 5179 2204
rect 5235 2202 5259 2204
rect 5097 2150 5099 2202
rect 5161 2150 5173 2202
rect 5235 2150 5237 2202
rect 5075 2148 5099 2150
rect 5155 2148 5179 2150
rect 5235 2148 5259 2150
rect 5019 2128 5315 2148
rect 4908 1414 5212 1442
rect 4448 1278 4752 1306
rect 4448 800 4476 1278
rect 5184 800 5212 1414
rect 5736 800 5764 6190
rect 5920 5778 5948 8453
rect 6472 5794 6500 8453
rect 5908 5772 5960 5778
rect 5908 5714 5960 5720
rect 6380 5766 6500 5794
rect 6380 5166 6408 5766
rect 6460 5636 6512 5642
rect 6460 5578 6512 5584
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6472 800 6500 5578
rect 570 0 626 800
rect 1122 0 1178 800
rect 1858 0 1914 800
rect 2410 0 2466 800
rect 3146 0 3202 800
rect 3698 0 3754 800
rect 4434 0 4490 800
rect 5170 0 5226 800
rect 5722 0 5778 800
rect 6458 0 6514 800
<< via2 >>
rect 1768 6554 1824 6556
rect 1848 6554 1904 6556
rect 1928 6554 1984 6556
rect 2008 6554 2064 6556
rect 1768 6502 1794 6554
rect 1794 6502 1824 6554
rect 1848 6502 1858 6554
rect 1858 6502 1904 6554
rect 1928 6502 1974 6554
rect 1974 6502 1984 6554
rect 2008 6502 2038 6554
rect 2038 6502 2064 6554
rect 1768 6500 1824 6502
rect 1848 6500 1904 6502
rect 1928 6500 1984 6502
rect 2008 6500 2064 6502
rect 1768 5466 1824 5468
rect 1848 5466 1904 5468
rect 1928 5466 1984 5468
rect 2008 5466 2064 5468
rect 1768 5414 1794 5466
rect 1794 5414 1824 5466
rect 1848 5414 1858 5466
rect 1858 5414 1904 5466
rect 1928 5414 1974 5466
rect 1974 5414 1984 5466
rect 2008 5414 2038 5466
rect 2038 5414 2064 5466
rect 1768 5412 1824 5414
rect 1848 5412 1904 5414
rect 1928 5412 1984 5414
rect 2008 5412 2064 5414
rect 1490 4664 1546 4720
rect 1768 4378 1824 4380
rect 1848 4378 1904 4380
rect 1928 4378 1984 4380
rect 2008 4378 2064 4380
rect 1768 4326 1794 4378
rect 1794 4326 1824 4378
rect 1848 4326 1858 4378
rect 1858 4326 1904 4378
rect 1928 4326 1974 4378
rect 1974 4326 1984 4378
rect 2008 4326 2038 4378
rect 2038 4326 2064 4378
rect 1768 4324 1824 4326
rect 1848 4324 1904 4326
rect 1928 4324 1984 4326
rect 2008 4324 2064 4326
rect 1582 3576 1638 3632
rect 1398 2760 1454 2816
rect 1306 1672 1362 1728
rect 1768 3290 1824 3292
rect 1848 3290 1904 3292
rect 1928 3290 1984 3292
rect 2008 3290 2064 3292
rect 1768 3238 1794 3290
rect 1794 3238 1824 3290
rect 1848 3238 1858 3290
rect 1858 3238 1904 3290
rect 1928 3238 1974 3290
rect 1974 3238 1984 3290
rect 2008 3238 2038 3290
rect 2038 3238 2064 3290
rect 1768 3236 1824 3238
rect 1848 3236 1904 3238
rect 1928 3236 1984 3238
rect 2008 3236 2064 3238
rect 2581 7098 2637 7100
rect 2661 7098 2717 7100
rect 2741 7098 2797 7100
rect 2821 7098 2877 7100
rect 2581 7046 2607 7098
rect 2607 7046 2637 7098
rect 2661 7046 2671 7098
rect 2671 7046 2717 7098
rect 2741 7046 2787 7098
rect 2787 7046 2797 7098
rect 2821 7046 2851 7098
rect 2851 7046 2877 7098
rect 2581 7044 2637 7046
rect 2661 7044 2717 7046
rect 2741 7044 2797 7046
rect 2821 7044 2877 7046
rect 3514 7676 3570 7712
rect 3514 7656 3516 7676
rect 3516 7656 3568 7676
rect 3568 7656 3570 7676
rect 2581 6010 2637 6012
rect 2661 6010 2717 6012
rect 2741 6010 2797 6012
rect 2821 6010 2877 6012
rect 2581 5958 2607 6010
rect 2607 5958 2637 6010
rect 2661 5958 2671 6010
rect 2671 5958 2717 6010
rect 2741 5958 2787 6010
rect 2787 5958 2797 6010
rect 2821 5958 2851 6010
rect 2851 5958 2877 6010
rect 2581 5956 2637 5958
rect 2661 5956 2717 5958
rect 2741 5956 2797 5958
rect 2821 5956 2877 5958
rect 2581 4922 2637 4924
rect 2661 4922 2717 4924
rect 2741 4922 2797 4924
rect 2821 4922 2877 4924
rect 2581 4870 2607 4922
rect 2607 4870 2637 4922
rect 2661 4870 2671 4922
rect 2671 4870 2717 4922
rect 2741 4870 2787 4922
rect 2787 4870 2797 4922
rect 2821 4870 2851 4922
rect 2851 4870 2877 4922
rect 2581 4868 2637 4870
rect 2661 4868 2717 4870
rect 2741 4868 2797 4870
rect 2821 4868 2877 4870
rect 1768 2202 1824 2204
rect 1848 2202 1904 2204
rect 1928 2202 1984 2204
rect 2008 2202 2064 2204
rect 1768 2150 1794 2202
rect 1794 2150 1824 2202
rect 1848 2150 1858 2202
rect 1858 2150 1904 2202
rect 1928 2150 1974 2202
rect 1974 2150 1984 2202
rect 2008 2150 2038 2202
rect 2038 2150 2064 2202
rect 1768 2148 1824 2150
rect 1848 2148 1904 2150
rect 1928 2148 1984 2150
rect 2008 2148 2064 2150
rect 2581 3834 2637 3836
rect 2661 3834 2717 3836
rect 2741 3834 2797 3836
rect 2821 3834 2877 3836
rect 2581 3782 2607 3834
rect 2607 3782 2637 3834
rect 2661 3782 2671 3834
rect 2671 3782 2717 3834
rect 2741 3782 2787 3834
rect 2787 3782 2797 3834
rect 2821 3782 2851 3834
rect 2851 3782 2877 3834
rect 2581 3780 2637 3782
rect 2661 3780 2717 3782
rect 2741 3780 2797 3782
rect 2821 3780 2877 3782
rect 3238 6704 3294 6760
rect 3146 4528 3202 4584
rect 3054 3576 3110 3632
rect 2581 2746 2637 2748
rect 2661 2746 2717 2748
rect 2741 2746 2797 2748
rect 2821 2746 2877 2748
rect 2581 2694 2607 2746
rect 2607 2694 2637 2746
rect 2661 2694 2671 2746
rect 2671 2694 2717 2746
rect 2741 2694 2787 2746
rect 2787 2694 2797 2746
rect 2821 2694 2851 2746
rect 2851 2694 2877 2746
rect 2581 2692 2637 2694
rect 2661 2692 2717 2694
rect 2741 2692 2797 2694
rect 2821 2692 2877 2694
rect 2962 2488 3018 2544
rect 3394 6554 3450 6556
rect 3474 6554 3530 6556
rect 3554 6554 3610 6556
rect 3634 6554 3690 6556
rect 3394 6502 3420 6554
rect 3420 6502 3450 6554
rect 3474 6502 3484 6554
rect 3484 6502 3530 6554
rect 3554 6502 3600 6554
rect 3600 6502 3610 6554
rect 3634 6502 3664 6554
rect 3664 6502 3690 6554
rect 3394 6500 3450 6502
rect 3474 6500 3530 6502
rect 3554 6500 3610 6502
rect 3634 6500 3690 6502
rect 3394 5466 3450 5468
rect 3474 5466 3530 5468
rect 3554 5466 3610 5468
rect 3634 5466 3690 5468
rect 3394 5414 3420 5466
rect 3420 5414 3450 5466
rect 3474 5414 3484 5466
rect 3484 5414 3530 5466
rect 3554 5414 3600 5466
rect 3600 5414 3610 5466
rect 3634 5414 3664 5466
rect 3664 5414 3690 5466
rect 3394 5412 3450 5414
rect 3474 5412 3530 5414
rect 3554 5412 3610 5414
rect 3634 5412 3690 5414
rect 3790 5208 3846 5264
rect 3394 4378 3450 4380
rect 3474 4378 3530 4380
rect 3554 4378 3610 4380
rect 3634 4378 3690 4380
rect 3394 4326 3420 4378
rect 3420 4326 3450 4378
rect 3474 4326 3484 4378
rect 3484 4326 3530 4378
rect 3554 4326 3600 4378
rect 3600 4326 3610 4378
rect 3634 4326 3664 4378
rect 3664 4326 3690 4378
rect 3394 4324 3450 4326
rect 3474 4324 3530 4326
rect 3554 4324 3610 4326
rect 3634 4324 3690 4326
rect 4066 7384 4122 7440
rect 4206 7098 4262 7100
rect 4286 7098 4342 7100
rect 4366 7098 4422 7100
rect 4446 7098 4502 7100
rect 4206 7046 4232 7098
rect 4232 7046 4262 7098
rect 4286 7046 4296 7098
rect 4296 7046 4342 7098
rect 4366 7046 4412 7098
rect 4412 7046 4422 7098
rect 4446 7046 4476 7098
rect 4476 7046 4502 7098
rect 4206 7044 4262 7046
rect 4286 7044 4342 7046
rect 4366 7044 4422 7046
rect 4446 7044 4502 7046
rect 4066 6316 4122 6352
rect 4066 6296 4068 6316
rect 4068 6296 4120 6316
rect 4120 6296 4122 6316
rect 4206 6010 4262 6012
rect 4286 6010 4342 6012
rect 4366 6010 4422 6012
rect 4446 6010 4502 6012
rect 4206 5958 4232 6010
rect 4232 5958 4262 6010
rect 4286 5958 4296 6010
rect 4296 5958 4342 6010
rect 4366 5958 4412 6010
rect 4412 5958 4422 6010
rect 4446 5958 4476 6010
rect 4476 5958 4502 6010
rect 4206 5956 4262 5958
rect 4286 5956 4342 5958
rect 4366 5956 4422 5958
rect 4446 5956 4502 5958
rect 3394 3290 3450 3292
rect 3474 3290 3530 3292
rect 3554 3290 3610 3292
rect 3634 3290 3690 3292
rect 3394 3238 3420 3290
rect 3420 3238 3450 3290
rect 3474 3238 3484 3290
rect 3484 3238 3530 3290
rect 3554 3238 3600 3290
rect 3600 3238 3610 3290
rect 3634 3238 3664 3290
rect 3664 3238 3690 3290
rect 3394 3236 3450 3238
rect 3474 3236 3530 3238
rect 3554 3236 3610 3238
rect 3634 3236 3690 3238
rect 3394 2202 3450 2204
rect 3474 2202 3530 2204
rect 3554 2202 3610 2204
rect 3634 2202 3690 2204
rect 3394 2150 3420 2202
rect 3420 2150 3450 2202
rect 3474 2150 3484 2202
rect 3484 2150 3530 2202
rect 3554 2150 3600 2202
rect 3600 2150 3610 2202
rect 3634 2150 3664 2202
rect 3664 2150 3690 2202
rect 3394 2148 3450 2150
rect 3474 2148 3530 2150
rect 3554 2148 3610 2150
rect 3634 2148 3690 2150
rect 4206 4922 4262 4924
rect 4286 4922 4342 4924
rect 4366 4922 4422 4924
rect 4446 4922 4502 4924
rect 4206 4870 4232 4922
rect 4232 4870 4262 4922
rect 4286 4870 4296 4922
rect 4296 4870 4342 4922
rect 4366 4870 4412 4922
rect 4412 4870 4422 4922
rect 4446 4870 4476 4922
rect 4476 4870 4502 4922
rect 4206 4868 4262 4870
rect 4286 4868 4342 4870
rect 4366 4868 4422 4870
rect 4446 4868 4502 4870
rect 5019 6554 5075 6556
rect 5099 6554 5155 6556
rect 5179 6554 5235 6556
rect 5259 6554 5315 6556
rect 5019 6502 5045 6554
rect 5045 6502 5075 6554
rect 5099 6502 5109 6554
rect 5109 6502 5155 6554
rect 5179 6502 5225 6554
rect 5225 6502 5235 6554
rect 5259 6502 5289 6554
rect 5289 6502 5315 6554
rect 5019 6500 5075 6502
rect 5099 6500 5155 6502
rect 5179 6500 5235 6502
rect 5259 6500 5315 6502
rect 5019 5466 5075 5468
rect 5099 5466 5155 5468
rect 5179 5466 5235 5468
rect 5259 5466 5315 5468
rect 5019 5414 5045 5466
rect 5045 5414 5075 5466
rect 5099 5414 5109 5466
rect 5109 5414 5155 5466
rect 5179 5414 5225 5466
rect 5225 5414 5235 5466
rect 5259 5414 5289 5466
rect 5289 5414 5315 5466
rect 5019 5412 5075 5414
rect 5099 5412 5155 5414
rect 5179 5412 5235 5414
rect 5259 5412 5315 5414
rect 4206 3834 4262 3836
rect 4286 3834 4342 3836
rect 4366 3834 4422 3836
rect 4446 3834 4502 3836
rect 4206 3782 4232 3834
rect 4232 3782 4262 3834
rect 4286 3782 4296 3834
rect 4296 3782 4342 3834
rect 4366 3782 4412 3834
rect 4412 3782 4422 3834
rect 4446 3782 4476 3834
rect 4476 3782 4502 3834
rect 4206 3780 4262 3782
rect 4286 3780 4342 3782
rect 4366 3780 4422 3782
rect 4446 3780 4502 3782
rect 4206 2746 4262 2748
rect 4286 2746 4342 2748
rect 4366 2746 4422 2748
rect 4446 2746 4502 2748
rect 4206 2694 4232 2746
rect 4232 2694 4262 2746
rect 4286 2694 4296 2746
rect 4296 2694 4342 2746
rect 4366 2694 4412 2746
rect 4412 2694 4422 2746
rect 4446 2694 4476 2746
rect 4476 2694 4502 2746
rect 4206 2692 4262 2694
rect 4286 2692 4342 2694
rect 4366 2692 4422 2694
rect 4446 2692 4502 2694
rect 3974 1400 4030 1456
rect 5019 4378 5075 4380
rect 5099 4378 5155 4380
rect 5179 4378 5235 4380
rect 5259 4378 5315 4380
rect 5019 4326 5045 4378
rect 5045 4326 5075 4378
rect 5099 4326 5109 4378
rect 5109 4326 5155 4378
rect 5179 4326 5225 4378
rect 5225 4326 5235 4378
rect 5259 4326 5289 4378
rect 5289 4326 5315 4378
rect 5019 4324 5075 4326
rect 5099 4324 5155 4326
rect 5179 4324 5235 4326
rect 5259 4324 5315 4326
rect 5019 3290 5075 3292
rect 5099 3290 5155 3292
rect 5179 3290 5235 3292
rect 5259 3290 5315 3292
rect 5019 3238 5045 3290
rect 5045 3238 5075 3290
rect 5099 3238 5109 3290
rect 5109 3238 5155 3290
rect 5179 3238 5225 3290
rect 5225 3238 5235 3290
rect 5259 3238 5289 3290
rect 5289 3238 5315 3290
rect 5019 3236 5075 3238
rect 5099 3236 5155 3238
rect 5179 3236 5235 3238
rect 5259 3236 5315 3238
rect 5019 2202 5075 2204
rect 5099 2202 5155 2204
rect 5179 2202 5235 2204
rect 5259 2202 5315 2204
rect 5019 2150 5045 2202
rect 5045 2150 5075 2202
rect 5099 2150 5109 2202
rect 5109 2150 5155 2202
rect 5179 2150 5225 2202
rect 5225 2150 5235 2202
rect 5259 2150 5289 2202
rect 5289 2150 5315 2202
rect 5019 2148 5075 2150
rect 5099 2148 5155 2150
rect 5179 2148 5235 2150
rect 5259 2148 5315 2150
<< metal3 >>
rect 0 7714 800 7744
rect 3509 7714 3575 7717
rect 0 7712 3575 7714
rect 0 7656 3514 7712
rect 3570 7656 3575 7712
rect 0 7654 3575 7656
rect 0 7624 800 7654
rect 3509 7651 3575 7654
rect 4061 7442 4127 7445
rect 6309 7442 7109 7472
rect 4061 7440 7109 7442
rect 4061 7384 4066 7440
rect 4122 7384 7109 7440
rect 4061 7382 7109 7384
rect 4061 7379 4127 7382
rect 6309 7352 7109 7382
rect 2569 7104 2889 7105
rect 2569 7040 2577 7104
rect 2641 7040 2657 7104
rect 2721 7040 2737 7104
rect 2801 7040 2817 7104
rect 2881 7040 2889 7104
rect 2569 7039 2889 7040
rect 4194 7104 4514 7105
rect 4194 7040 4202 7104
rect 4266 7040 4282 7104
rect 4346 7040 4362 7104
rect 4426 7040 4442 7104
rect 4506 7040 4514 7104
rect 4194 7039 4514 7040
rect 3233 6762 3299 6765
rect 1350 6760 3299 6762
rect 1350 6704 3238 6760
rect 3294 6704 3299 6760
rect 1350 6702 3299 6704
rect 0 6626 800 6656
rect 1350 6626 1410 6702
rect 3233 6699 3299 6702
rect 0 6566 1410 6626
rect 0 6536 800 6566
rect 1756 6560 2076 6561
rect 1756 6496 1764 6560
rect 1828 6496 1844 6560
rect 1908 6496 1924 6560
rect 1988 6496 2004 6560
rect 2068 6496 2076 6560
rect 1756 6495 2076 6496
rect 3382 6560 3702 6561
rect 3382 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3702 6560
rect 3382 6495 3702 6496
rect 5007 6560 5327 6561
rect 5007 6496 5015 6560
rect 5079 6496 5095 6560
rect 5159 6496 5175 6560
rect 5239 6496 5255 6560
rect 5319 6496 5327 6560
rect 5007 6495 5327 6496
rect 4061 6354 4127 6357
rect 6309 6354 7109 6384
rect 4061 6352 7109 6354
rect 4061 6296 4066 6352
rect 4122 6296 7109 6352
rect 4061 6294 7109 6296
rect 4061 6291 4127 6294
rect 6309 6264 7109 6294
rect 2569 6016 2889 6017
rect 2569 5952 2577 6016
rect 2641 5952 2657 6016
rect 2721 5952 2737 6016
rect 2801 5952 2817 6016
rect 2881 5952 2889 6016
rect 2569 5951 2889 5952
rect 4194 6016 4514 6017
rect 4194 5952 4202 6016
rect 4266 5952 4282 6016
rect 4346 5952 4362 6016
rect 4426 5952 4442 6016
rect 4506 5952 4514 6016
rect 4194 5951 4514 5952
rect 0 5448 800 5568
rect 6309 5538 7109 5568
rect 5398 5478 7109 5538
rect 1756 5472 2076 5473
rect 1756 5408 1764 5472
rect 1828 5408 1844 5472
rect 1908 5408 1924 5472
rect 1988 5408 2004 5472
rect 2068 5408 2076 5472
rect 1756 5407 2076 5408
rect 3382 5472 3702 5473
rect 3382 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3702 5472
rect 3382 5407 3702 5408
rect 5007 5472 5327 5473
rect 5007 5408 5015 5472
rect 5079 5408 5095 5472
rect 5159 5408 5175 5472
rect 5239 5408 5255 5472
rect 5319 5408 5327 5472
rect 5007 5407 5327 5408
rect 3785 5266 3851 5269
rect 5398 5266 5458 5478
rect 6309 5448 7109 5478
rect 3785 5264 5458 5266
rect 3785 5208 3790 5264
rect 3846 5208 5458 5264
rect 3785 5206 5458 5208
rect 3785 5203 3851 5206
rect 2569 4928 2889 4929
rect 2569 4864 2577 4928
rect 2641 4864 2657 4928
rect 2721 4864 2737 4928
rect 2801 4864 2817 4928
rect 2881 4864 2889 4928
rect 2569 4863 2889 4864
rect 4194 4928 4514 4929
rect 4194 4864 4202 4928
rect 4266 4864 4282 4928
rect 4346 4864 4362 4928
rect 4426 4864 4442 4928
rect 4506 4864 4514 4928
rect 4194 4863 4514 4864
rect 0 4722 800 4752
rect 1485 4722 1551 4725
rect 0 4720 1551 4722
rect 0 4664 1490 4720
rect 1546 4664 1551 4720
rect 0 4662 1551 4664
rect 0 4632 800 4662
rect 1485 4659 1551 4662
rect 3141 4586 3207 4589
rect 3141 4584 5458 4586
rect 3141 4528 3146 4584
rect 3202 4528 5458 4584
rect 3141 4526 5458 4528
rect 3141 4523 3207 4526
rect 5398 4450 5458 4526
rect 6309 4450 7109 4480
rect 5398 4390 7109 4450
rect 1756 4384 2076 4385
rect 1756 4320 1764 4384
rect 1828 4320 1844 4384
rect 1908 4320 1924 4384
rect 1988 4320 2004 4384
rect 2068 4320 2076 4384
rect 1756 4319 2076 4320
rect 3382 4384 3702 4385
rect 3382 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3702 4384
rect 3382 4319 3702 4320
rect 5007 4384 5327 4385
rect 5007 4320 5015 4384
rect 5079 4320 5095 4384
rect 5159 4320 5175 4384
rect 5239 4320 5255 4384
rect 5319 4320 5327 4384
rect 6309 4360 7109 4390
rect 5007 4319 5327 4320
rect 2569 3840 2889 3841
rect 2569 3776 2577 3840
rect 2641 3776 2657 3840
rect 2721 3776 2737 3840
rect 2801 3776 2817 3840
rect 2881 3776 2889 3840
rect 2569 3775 2889 3776
rect 4194 3840 4514 3841
rect 4194 3776 4202 3840
rect 4266 3776 4282 3840
rect 4346 3776 4362 3840
rect 4426 3776 4442 3840
rect 4506 3776 4514 3840
rect 4194 3775 4514 3776
rect 0 3634 800 3664
rect 1577 3634 1643 3637
rect 0 3632 1643 3634
rect 0 3576 1582 3632
rect 1638 3576 1643 3632
rect 0 3574 1643 3576
rect 0 3544 800 3574
rect 1577 3571 1643 3574
rect 3049 3634 3115 3637
rect 6309 3634 7109 3664
rect 3049 3632 7109 3634
rect 3049 3576 3054 3632
rect 3110 3576 7109 3632
rect 3049 3574 7109 3576
rect 3049 3571 3115 3574
rect 6309 3544 7109 3574
rect 1756 3296 2076 3297
rect 1756 3232 1764 3296
rect 1828 3232 1844 3296
rect 1908 3232 1924 3296
rect 1988 3232 2004 3296
rect 2068 3232 2076 3296
rect 1756 3231 2076 3232
rect 3382 3296 3702 3297
rect 3382 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3702 3296
rect 3382 3231 3702 3232
rect 5007 3296 5327 3297
rect 5007 3232 5015 3296
rect 5079 3232 5095 3296
rect 5159 3232 5175 3296
rect 5239 3232 5255 3296
rect 5319 3232 5327 3296
rect 5007 3231 5327 3232
rect 0 2818 800 2848
rect 1393 2818 1459 2821
rect 0 2816 1459 2818
rect 0 2760 1398 2816
rect 1454 2760 1459 2816
rect 0 2758 1459 2760
rect 0 2728 800 2758
rect 1393 2755 1459 2758
rect 2569 2752 2889 2753
rect 2569 2688 2577 2752
rect 2641 2688 2657 2752
rect 2721 2688 2737 2752
rect 2801 2688 2817 2752
rect 2881 2688 2889 2752
rect 2569 2687 2889 2688
rect 4194 2752 4514 2753
rect 4194 2688 4202 2752
rect 4266 2688 4282 2752
rect 4346 2688 4362 2752
rect 4426 2688 4442 2752
rect 4506 2688 4514 2752
rect 4194 2687 4514 2688
rect 2957 2546 3023 2549
rect 6309 2546 7109 2576
rect 2957 2544 7109 2546
rect 2957 2488 2962 2544
rect 3018 2488 7109 2544
rect 2957 2486 7109 2488
rect 2957 2483 3023 2486
rect 6309 2456 7109 2486
rect 1756 2208 2076 2209
rect 1756 2144 1764 2208
rect 1828 2144 1844 2208
rect 1908 2144 1924 2208
rect 1988 2144 2004 2208
rect 2068 2144 2076 2208
rect 1756 2143 2076 2144
rect 3382 2208 3702 2209
rect 3382 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3702 2208
rect 3382 2143 3702 2144
rect 5007 2208 5327 2209
rect 5007 2144 5015 2208
rect 5079 2144 5095 2208
rect 5159 2144 5175 2208
rect 5239 2144 5255 2208
rect 5319 2144 5327 2208
rect 5007 2143 5327 2144
rect 0 1730 800 1760
rect 1301 1730 1367 1733
rect 0 1728 1367 1730
rect 0 1672 1306 1728
rect 1362 1672 1367 1728
rect 0 1670 1367 1672
rect 0 1640 800 1670
rect 1301 1667 1367 1670
rect 3969 1458 4035 1461
rect 6309 1458 7109 1488
rect 3969 1456 7109 1458
rect 3969 1400 3974 1456
rect 4030 1400 7109 1456
rect 3969 1398 7109 1400
rect 3969 1395 4035 1398
rect 6309 1368 7109 1398
<< via3 >>
rect 2577 7100 2641 7104
rect 2577 7044 2581 7100
rect 2581 7044 2637 7100
rect 2637 7044 2641 7100
rect 2577 7040 2641 7044
rect 2657 7100 2721 7104
rect 2657 7044 2661 7100
rect 2661 7044 2717 7100
rect 2717 7044 2721 7100
rect 2657 7040 2721 7044
rect 2737 7100 2801 7104
rect 2737 7044 2741 7100
rect 2741 7044 2797 7100
rect 2797 7044 2801 7100
rect 2737 7040 2801 7044
rect 2817 7100 2881 7104
rect 2817 7044 2821 7100
rect 2821 7044 2877 7100
rect 2877 7044 2881 7100
rect 2817 7040 2881 7044
rect 4202 7100 4266 7104
rect 4202 7044 4206 7100
rect 4206 7044 4262 7100
rect 4262 7044 4266 7100
rect 4202 7040 4266 7044
rect 4282 7100 4346 7104
rect 4282 7044 4286 7100
rect 4286 7044 4342 7100
rect 4342 7044 4346 7100
rect 4282 7040 4346 7044
rect 4362 7100 4426 7104
rect 4362 7044 4366 7100
rect 4366 7044 4422 7100
rect 4422 7044 4426 7100
rect 4362 7040 4426 7044
rect 4442 7100 4506 7104
rect 4442 7044 4446 7100
rect 4446 7044 4502 7100
rect 4502 7044 4506 7100
rect 4442 7040 4506 7044
rect 1764 6556 1828 6560
rect 1764 6500 1768 6556
rect 1768 6500 1824 6556
rect 1824 6500 1828 6556
rect 1764 6496 1828 6500
rect 1844 6556 1908 6560
rect 1844 6500 1848 6556
rect 1848 6500 1904 6556
rect 1904 6500 1908 6556
rect 1844 6496 1908 6500
rect 1924 6556 1988 6560
rect 1924 6500 1928 6556
rect 1928 6500 1984 6556
rect 1984 6500 1988 6556
rect 1924 6496 1988 6500
rect 2004 6556 2068 6560
rect 2004 6500 2008 6556
rect 2008 6500 2064 6556
rect 2064 6500 2068 6556
rect 2004 6496 2068 6500
rect 3390 6556 3454 6560
rect 3390 6500 3394 6556
rect 3394 6500 3450 6556
rect 3450 6500 3454 6556
rect 3390 6496 3454 6500
rect 3470 6556 3534 6560
rect 3470 6500 3474 6556
rect 3474 6500 3530 6556
rect 3530 6500 3534 6556
rect 3470 6496 3534 6500
rect 3550 6556 3614 6560
rect 3550 6500 3554 6556
rect 3554 6500 3610 6556
rect 3610 6500 3614 6556
rect 3550 6496 3614 6500
rect 3630 6556 3694 6560
rect 3630 6500 3634 6556
rect 3634 6500 3690 6556
rect 3690 6500 3694 6556
rect 3630 6496 3694 6500
rect 5015 6556 5079 6560
rect 5015 6500 5019 6556
rect 5019 6500 5075 6556
rect 5075 6500 5079 6556
rect 5015 6496 5079 6500
rect 5095 6556 5159 6560
rect 5095 6500 5099 6556
rect 5099 6500 5155 6556
rect 5155 6500 5159 6556
rect 5095 6496 5159 6500
rect 5175 6556 5239 6560
rect 5175 6500 5179 6556
rect 5179 6500 5235 6556
rect 5235 6500 5239 6556
rect 5175 6496 5239 6500
rect 5255 6556 5319 6560
rect 5255 6500 5259 6556
rect 5259 6500 5315 6556
rect 5315 6500 5319 6556
rect 5255 6496 5319 6500
rect 2577 6012 2641 6016
rect 2577 5956 2581 6012
rect 2581 5956 2637 6012
rect 2637 5956 2641 6012
rect 2577 5952 2641 5956
rect 2657 6012 2721 6016
rect 2657 5956 2661 6012
rect 2661 5956 2717 6012
rect 2717 5956 2721 6012
rect 2657 5952 2721 5956
rect 2737 6012 2801 6016
rect 2737 5956 2741 6012
rect 2741 5956 2797 6012
rect 2797 5956 2801 6012
rect 2737 5952 2801 5956
rect 2817 6012 2881 6016
rect 2817 5956 2821 6012
rect 2821 5956 2877 6012
rect 2877 5956 2881 6012
rect 2817 5952 2881 5956
rect 4202 6012 4266 6016
rect 4202 5956 4206 6012
rect 4206 5956 4262 6012
rect 4262 5956 4266 6012
rect 4202 5952 4266 5956
rect 4282 6012 4346 6016
rect 4282 5956 4286 6012
rect 4286 5956 4342 6012
rect 4342 5956 4346 6012
rect 4282 5952 4346 5956
rect 4362 6012 4426 6016
rect 4362 5956 4366 6012
rect 4366 5956 4422 6012
rect 4422 5956 4426 6012
rect 4362 5952 4426 5956
rect 4442 6012 4506 6016
rect 4442 5956 4446 6012
rect 4446 5956 4502 6012
rect 4502 5956 4506 6012
rect 4442 5952 4506 5956
rect 1764 5468 1828 5472
rect 1764 5412 1768 5468
rect 1768 5412 1824 5468
rect 1824 5412 1828 5468
rect 1764 5408 1828 5412
rect 1844 5468 1908 5472
rect 1844 5412 1848 5468
rect 1848 5412 1904 5468
rect 1904 5412 1908 5468
rect 1844 5408 1908 5412
rect 1924 5468 1988 5472
rect 1924 5412 1928 5468
rect 1928 5412 1984 5468
rect 1984 5412 1988 5468
rect 1924 5408 1988 5412
rect 2004 5468 2068 5472
rect 2004 5412 2008 5468
rect 2008 5412 2064 5468
rect 2064 5412 2068 5468
rect 2004 5408 2068 5412
rect 3390 5468 3454 5472
rect 3390 5412 3394 5468
rect 3394 5412 3450 5468
rect 3450 5412 3454 5468
rect 3390 5408 3454 5412
rect 3470 5468 3534 5472
rect 3470 5412 3474 5468
rect 3474 5412 3530 5468
rect 3530 5412 3534 5468
rect 3470 5408 3534 5412
rect 3550 5468 3614 5472
rect 3550 5412 3554 5468
rect 3554 5412 3610 5468
rect 3610 5412 3614 5468
rect 3550 5408 3614 5412
rect 3630 5468 3694 5472
rect 3630 5412 3634 5468
rect 3634 5412 3690 5468
rect 3690 5412 3694 5468
rect 3630 5408 3694 5412
rect 5015 5468 5079 5472
rect 5015 5412 5019 5468
rect 5019 5412 5075 5468
rect 5075 5412 5079 5468
rect 5015 5408 5079 5412
rect 5095 5468 5159 5472
rect 5095 5412 5099 5468
rect 5099 5412 5155 5468
rect 5155 5412 5159 5468
rect 5095 5408 5159 5412
rect 5175 5468 5239 5472
rect 5175 5412 5179 5468
rect 5179 5412 5235 5468
rect 5235 5412 5239 5468
rect 5175 5408 5239 5412
rect 5255 5468 5319 5472
rect 5255 5412 5259 5468
rect 5259 5412 5315 5468
rect 5315 5412 5319 5468
rect 5255 5408 5319 5412
rect 2577 4924 2641 4928
rect 2577 4868 2581 4924
rect 2581 4868 2637 4924
rect 2637 4868 2641 4924
rect 2577 4864 2641 4868
rect 2657 4924 2721 4928
rect 2657 4868 2661 4924
rect 2661 4868 2717 4924
rect 2717 4868 2721 4924
rect 2657 4864 2721 4868
rect 2737 4924 2801 4928
rect 2737 4868 2741 4924
rect 2741 4868 2797 4924
rect 2797 4868 2801 4924
rect 2737 4864 2801 4868
rect 2817 4924 2881 4928
rect 2817 4868 2821 4924
rect 2821 4868 2877 4924
rect 2877 4868 2881 4924
rect 2817 4864 2881 4868
rect 4202 4924 4266 4928
rect 4202 4868 4206 4924
rect 4206 4868 4262 4924
rect 4262 4868 4266 4924
rect 4202 4864 4266 4868
rect 4282 4924 4346 4928
rect 4282 4868 4286 4924
rect 4286 4868 4342 4924
rect 4342 4868 4346 4924
rect 4282 4864 4346 4868
rect 4362 4924 4426 4928
rect 4362 4868 4366 4924
rect 4366 4868 4422 4924
rect 4422 4868 4426 4924
rect 4362 4864 4426 4868
rect 4442 4924 4506 4928
rect 4442 4868 4446 4924
rect 4446 4868 4502 4924
rect 4502 4868 4506 4924
rect 4442 4864 4506 4868
rect 1764 4380 1828 4384
rect 1764 4324 1768 4380
rect 1768 4324 1824 4380
rect 1824 4324 1828 4380
rect 1764 4320 1828 4324
rect 1844 4380 1908 4384
rect 1844 4324 1848 4380
rect 1848 4324 1904 4380
rect 1904 4324 1908 4380
rect 1844 4320 1908 4324
rect 1924 4380 1988 4384
rect 1924 4324 1928 4380
rect 1928 4324 1984 4380
rect 1984 4324 1988 4380
rect 1924 4320 1988 4324
rect 2004 4380 2068 4384
rect 2004 4324 2008 4380
rect 2008 4324 2064 4380
rect 2064 4324 2068 4380
rect 2004 4320 2068 4324
rect 3390 4380 3454 4384
rect 3390 4324 3394 4380
rect 3394 4324 3450 4380
rect 3450 4324 3454 4380
rect 3390 4320 3454 4324
rect 3470 4380 3534 4384
rect 3470 4324 3474 4380
rect 3474 4324 3530 4380
rect 3530 4324 3534 4380
rect 3470 4320 3534 4324
rect 3550 4380 3614 4384
rect 3550 4324 3554 4380
rect 3554 4324 3610 4380
rect 3610 4324 3614 4380
rect 3550 4320 3614 4324
rect 3630 4380 3694 4384
rect 3630 4324 3634 4380
rect 3634 4324 3690 4380
rect 3690 4324 3694 4380
rect 3630 4320 3694 4324
rect 5015 4380 5079 4384
rect 5015 4324 5019 4380
rect 5019 4324 5075 4380
rect 5075 4324 5079 4380
rect 5015 4320 5079 4324
rect 5095 4380 5159 4384
rect 5095 4324 5099 4380
rect 5099 4324 5155 4380
rect 5155 4324 5159 4380
rect 5095 4320 5159 4324
rect 5175 4380 5239 4384
rect 5175 4324 5179 4380
rect 5179 4324 5235 4380
rect 5235 4324 5239 4380
rect 5175 4320 5239 4324
rect 5255 4380 5319 4384
rect 5255 4324 5259 4380
rect 5259 4324 5315 4380
rect 5315 4324 5319 4380
rect 5255 4320 5319 4324
rect 2577 3836 2641 3840
rect 2577 3780 2581 3836
rect 2581 3780 2637 3836
rect 2637 3780 2641 3836
rect 2577 3776 2641 3780
rect 2657 3836 2721 3840
rect 2657 3780 2661 3836
rect 2661 3780 2717 3836
rect 2717 3780 2721 3836
rect 2657 3776 2721 3780
rect 2737 3836 2801 3840
rect 2737 3780 2741 3836
rect 2741 3780 2797 3836
rect 2797 3780 2801 3836
rect 2737 3776 2801 3780
rect 2817 3836 2881 3840
rect 2817 3780 2821 3836
rect 2821 3780 2877 3836
rect 2877 3780 2881 3836
rect 2817 3776 2881 3780
rect 4202 3836 4266 3840
rect 4202 3780 4206 3836
rect 4206 3780 4262 3836
rect 4262 3780 4266 3836
rect 4202 3776 4266 3780
rect 4282 3836 4346 3840
rect 4282 3780 4286 3836
rect 4286 3780 4342 3836
rect 4342 3780 4346 3836
rect 4282 3776 4346 3780
rect 4362 3836 4426 3840
rect 4362 3780 4366 3836
rect 4366 3780 4422 3836
rect 4422 3780 4426 3836
rect 4362 3776 4426 3780
rect 4442 3836 4506 3840
rect 4442 3780 4446 3836
rect 4446 3780 4502 3836
rect 4502 3780 4506 3836
rect 4442 3776 4506 3780
rect 1764 3292 1828 3296
rect 1764 3236 1768 3292
rect 1768 3236 1824 3292
rect 1824 3236 1828 3292
rect 1764 3232 1828 3236
rect 1844 3292 1908 3296
rect 1844 3236 1848 3292
rect 1848 3236 1904 3292
rect 1904 3236 1908 3292
rect 1844 3232 1908 3236
rect 1924 3292 1988 3296
rect 1924 3236 1928 3292
rect 1928 3236 1984 3292
rect 1984 3236 1988 3292
rect 1924 3232 1988 3236
rect 2004 3292 2068 3296
rect 2004 3236 2008 3292
rect 2008 3236 2064 3292
rect 2064 3236 2068 3292
rect 2004 3232 2068 3236
rect 3390 3292 3454 3296
rect 3390 3236 3394 3292
rect 3394 3236 3450 3292
rect 3450 3236 3454 3292
rect 3390 3232 3454 3236
rect 3470 3292 3534 3296
rect 3470 3236 3474 3292
rect 3474 3236 3530 3292
rect 3530 3236 3534 3292
rect 3470 3232 3534 3236
rect 3550 3292 3614 3296
rect 3550 3236 3554 3292
rect 3554 3236 3610 3292
rect 3610 3236 3614 3292
rect 3550 3232 3614 3236
rect 3630 3292 3694 3296
rect 3630 3236 3634 3292
rect 3634 3236 3690 3292
rect 3690 3236 3694 3292
rect 3630 3232 3694 3236
rect 5015 3292 5079 3296
rect 5015 3236 5019 3292
rect 5019 3236 5075 3292
rect 5075 3236 5079 3292
rect 5015 3232 5079 3236
rect 5095 3292 5159 3296
rect 5095 3236 5099 3292
rect 5099 3236 5155 3292
rect 5155 3236 5159 3292
rect 5095 3232 5159 3236
rect 5175 3292 5239 3296
rect 5175 3236 5179 3292
rect 5179 3236 5235 3292
rect 5235 3236 5239 3292
rect 5175 3232 5239 3236
rect 5255 3292 5319 3296
rect 5255 3236 5259 3292
rect 5259 3236 5315 3292
rect 5315 3236 5319 3292
rect 5255 3232 5319 3236
rect 2577 2748 2641 2752
rect 2577 2692 2581 2748
rect 2581 2692 2637 2748
rect 2637 2692 2641 2748
rect 2577 2688 2641 2692
rect 2657 2748 2721 2752
rect 2657 2692 2661 2748
rect 2661 2692 2717 2748
rect 2717 2692 2721 2748
rect 2657 2688 2721 2692
rect 2737 2748 2801 2752
rect 2737 2692 2741 2748
rect 2741 2692 2797 2748
rect 2797 2692 2801 2748
rect 2737 2688 2801 2692
rect 2817 2748 2881 2752
rect 2817 2692 2821 2748
rect 2821 2692 2877 2748
rect 2877 2692 2881 2748
rect 2817 2688 2881 2692
rect 4202 2748 4266 2752
rect 4202 2692 4206 2748
rect 4206 2692 4262 2748
rect 4262 2692 4266 2748
rect 4202 2688 4266 2692
rect 4282 2748 4346 2752
rect 4282 2692 4286 2748
rect 4286 2692 4342 2748
rect 4342 2692 4346 2748
rect 4282 2688 4346 2692
rect 4362 2748 4426 2752
rect 4362 2692 4366 2748
rect 4366 2692 4422 2748
rect 4422 2692 4426 2748
rect 4362 2688 4426 2692
rect 4442 2748 4506 2752
rect 4442 2692 4446 2748
rect 4446 2692 4502 2748
rect 4502 2692 4506 2748
rect 4442 2688 4506 2692
rect 1764 2204 1828 2208
rect 1764 2148 1768 2204
rect 1768 2148 1824 2204
rect 1824 2148 1828 2204
rect 1764 2144 1828 2148
rect 1844 2204 1908 2208
rect 1844 2148 1848 2204
rect 1848 2148 1904 2204
rect 1904 2148 1908 2204
rect 1844 2144 1908 2148
rect 1924 2204 1988 2208
rect 1924 2148 1928 2204
rect 1928 2148 1984 2204
rect 1984 2148 1988 2204
rect 1924 2144 1988 2148
rect 2004 2204 2068 2208
rect 2004 2148 2008 2204
rect 2008 2148 2064 2204
rect 2064 2148 2068 2204
rect 2004 2144 2068 2148
rect 3390 2204 3454 2208
rect 3390 2148 3394 2204
rect 3394 2148 3450 2204
rect 3450 2148 3454 2204
rect 3390 2144 3454 2148
rect 3470 2204 3534 2208
rect 3470 2148 3474 2204
rect 3474 2148 3530 2204
rect 3530 2148 3534 2204
rect 3470 2144 3534 2148
rect 3550 2204 3614 2208
rect 3550 2148 3554 2204
rect 3554 2148 3610 2204
rect 3610 2148 3614 2204
rect 3550 2144 3614 2148
rect 3630 2204 3694 2208
rect 3630 2148 3634 2204
rect 3634 2148 3690 2204
rect 3690 2148 3694 2204
rect 3630 2144 3694 2148
rect 5015 2204 5079 2208
rect 5015 2148 5019 2204
rect 5019 2148 5075 2204
rect 5075 2148 5079 2204
rect 5015 2144 5079 2148
rect 5095 2204 5159 2208
rect 5095 2148 5099 2204
rect 5099 2148 5155 2204
rect 5155 2148 5159 2204
rect 5095 2144 5159 2148
rect 5175 2204 5239 2208
rect 5175 2148 5179 2204
rect 5179 2148 5235 2204
rect 5235 2148 5239 2204
rect 5175 2144 5239 2148
rect 5255 2204 5319 2208
rect 5255 2148 5259 2204
rect 5259 2148 5315 2204
rect 5315 2148 5319 2204
rect 5255 2144 5319 2148
<< metal4 >>
rect 1756 6560 2076 7120
rect 1756 6496 1764 6560
rect 1828 6496 1844 6560
rect 1908 6496 1924 6560
rect 1988 6496 2004 6560
rect 2068 6496 2076 6560
rect 1756 6326 2076 6496
rect 1756 6090 1798 6326
rect 2034 6090 2076 6326
rect 1756 5472 2076 6090
rect 1756 5408 1764 5472
rect 1828 5408 1844 5472
rect 1908 5408 1924 5472
rect 1988 5408 2004 5472
rect 2068 5408 2076 5472
rect 1756 4694 2076 5408
rect 1756 4458 1798 4694
rect 2034 4458 2076 4694
rect 1756 4384 2076 4458
rect 1756 4320 1764 4384
rect 1828 4320 1844 4384
rect 1908 4320 1924 4384
rect 1988 4320 2004 4384
rect 2068 4320 2076 4384
rect 1756 3296 2076 4320
rect 1756 3232 1764 3296
rect 1828 3232 1844 3296
rect 1908 3232 1924 3296
rect 1988 3232 2004 3296
rect 2068 3232 2076 3296
rect 1756 3062 2076 3232
rect 1756 2826 1798 3062
rect 2034 2826 2076 3062
rect 1756 2208 2076 2826
rect 1756 2144 1764 2208
rect 1828 2144 1844 2208
rect 1908 2144 1924 2208
rect 1988 2144 2004 2208
rect 2068 2144 2076 2208
rect 1756 2128 2076 2144
rect 2569 7104 2889 7120
rect 2569 7040 2577 7104
rect 2641 7040 2657 7104
rect 2721 7040 2737 7104
rect 2801 7040 2817 7104
rect 2881 7040 2889 7104
rect 2569 6016 2889 7040
rect 2569 5952 2577 6016
rect 2641 5952 2657 6016
rect 2721 5952 2737 6016
rect 2801 5952 2817 6016
rect 2881 5952 2889 6016
rect 2569 5510 2889 5952
rect 2569 5274 2611 5510
rect 2847 5274 2889 5510
rect 2569 4928 2889 5274
rect 2569 4864 2577 4928
rect 2641 4864 2657 4928
rect 2721 4864 2737 4928
rect 2801 4864 2817 4928
rect 2881 4864 2889 4928
rect 2569 3878 2889 4864
rect 2569 3840 2611 3878
rect 2847 3840 2889 3878
rect 2569 3776 2577 3840
rect 2881 3776 2889 3840
rect 2569 3642 2611 3776
rect 2847 3642 2889 3776
rect 2569 2752 2889 3642
rect 2569 2688 2577 2752
rect 2641 2688 2657 2752
rect 2721 2688 2737 2752
rect 2801 2688 2817 2752
rect 2881 2688 2889 2752
rect 2569 2128 2889 2688
rect 3382 6560 3702 7120
rect 3382 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3702 6560
rect 3382 6326 3702 6496
rect 3382 6090 3424 6326
rect 3660 6090 3702 6326
rect 3382 5472 3702 6090
rect 3382 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3702 5472
rect 3382 4694 3702 5408
rect 3382 4458 3424 4694
rect 3660 4458 3702 4694
rect 3382 4384 3702 4458
rect 3382 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3702 4384
rect 3382 3296 3702 4320
rect 3382 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3702 3296
rect 3382 3062 3702 3232
rect 3382 2826 3424 3062
rect 3660 2826 3702 3062
rect 3382 2208 3702 2826
rect 3382 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3702 2208
rect 3382 2128 3702 2144
rect 4194 7104 4514 7120
rect 4194 7040 4202 7104
rect 4266 7040 4282 7104
rect 4346 7040 4362 7104
rect 4426 7040 4442 7104
rect 4506 7040 4514 7104
rect 4194 6016 4514 7040
rect 4194 5952 4202 6016
rect 4266 5952 4282 6016
rect 4346 5952 4362 6016
rect 4426 5952 4442 6016
rect 4506 5952 4514 6016
rect 4194 5510 4514 5952
rect 4194 5274 4236 5510
rect 4472 5274 4514 5510
rect 4194 4928 4514 5274
rect 4194 4864 4202 4928
rect 4266 4864 4282 4928
rect 4346 4864 4362 4928
rect 4426 4864 4442 4928
rect 4506 4864 4514 4928
rect 4194 3878 4514 4864
rect 4194 3840 4236 3878
rect 4472 3840 4514 3878
rect 4194 3776 4202 3840
rect 4506 3776 4514 3840
rect 4194 3642 4236 3776
rect 4472 3642 4514 3776
rect 4194 2752 4514 3642
rect 4194 2688 4202 2752
rect 4266 2688 4282 2752
rect 4346 2688 4362 2752
rect 4426 2688 4442 2752
rect 4506 2688 4514 2752
rect 4194 2128 4514 2688
rect 5007 6560 5327 7120
rect 5007 6496 5015 6560
rect 5079 6496 5095 6560
rect 5159 6496 5175 6560
rect 5239 6496 5255 6560
rect 5319 6496 5327 6560
rect 5007 6326 5327 6496
rect 5007 6090 5049 6326
rect 5285 6090 5327 6326
rect 5007 5472 5327 6090
rect 5007 5408 5015 5472
rect 5079 5408 5095 5472
rect 5159 5408 5175 5472
rect 5239 5408 5255 5472
rect 5319 5408 5327 5472
rect 5007 4694 5327 5408
rect 5007 4458 5049 4694
rect 5285 4458 5327 4694
rect 5007 4384 5327 4458
rect 5007 4320 5015 4384
rect 5079 4320 5095 4384
rect 5159 4320 5175 4384
rect 5239 4320 5255 4384
rect 5319 4320 5327 4384
rect 5007 3296 5327 4320
rect 5007 3232 5015 3296
rect 5079 3232 5095 3296
rect 5159 3232 5175 3296
rect 5239 3232 5255 3296
rect 5319 3232 5327 3296
rect 5007 3062 5327 3232
rect 5007 2826 5049 3062
rect 5285 2826 5327 3062
rect 5007 2208 5327 2826
rect 5007 2144 5015 2208
rect 5079 2144 5095 2208
rect 5159 2144 5175 2208
rect 5239 2144 5255 2208
rect 5319 2144 5327 2208
rect 5007 2128 5327 2144
<< via4 >>
rect 1798 6090 2034 6326
rect 1798 4458 2034 4694
rect 1798 2826 2034 3062
rect 2611 5274 2847 5510
rect 2611 3840 2847 3878
rect 2611 3776 2641 3840
rect 2641 3776 2657 3840
rect 2657 3776 2721 3840
rect 2721 3776 2737 3840
rect 2737 3776 2801 3840
rect 2801 3776 2817 3840
rect 2817 3776 2847 3840
rect 2611 3642 2847 3776
rect 3424 6090 3660 6326
rect 3424 4458 3660 4694
rect 3424 2826 3660 3062
rect 4236 5274 4472 5510
rect 4236 3840 4472 3878
rect 4236 3776 4266 3840
rect 4266 3776 4282 3840
rect 4282 3776 4346 3840
rect 4346 3776 4362 3840
rect 4362 3776 4426 3840
rect 4426 3776 4442 3840
rect 4442 3776 4472 3840
rect 4236 3642 4472 3776
rect 5049 6090 5285 6326
rect 5049 4458 5285 4694
rect 5049 2826 5285 3062
<< metal5 >>
rect 1104 6326 5980 6368
rect 1104 6090 1798 6326
rect 2034 6090 3424 6326
rect 3660 6090 5049 6326
rect 5285 6090 5980 6326
rect 1104 6048 5980 6090
rect 1104 5510 5980 5552
rect 1104 5274 2611 5510
rect 2847 5274 4236 5510
rect 4472 5274 5980 5510
rect 1104 5232 5980 5274
rect 1104 4694 5980 4736
rect 1104 4458 1798 4694
rect 2034 4458 3424 4694
rect 3660 4458 5049 4694
rect 5285 4458 5980 4694
rect 1104 4416 5980 4458
rect 1104 3878 5980 3920
rect 1104 3642 2611 3878
rect 2847 3642 4236 3878
rect 4472 3642 5980 3878
rect 1104 3600 5980 3642
rect 1104 3062 5980 3104
rect 1104 2826 1798 3062
rect 2034 2826 3424 3062
rect 3660 2826 5049 3062
rect 5285 2826 5980 3062
rect 1104 2784 5980 2826
use sky130_fd_sc_hd__conb_1  mask_rev_value\[19\] /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 2116 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[20\]
timestamp 1604489732
transform 1 0 1656 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[2\]
timestamp 1604489732
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604489732
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3
timestamp 1604489732
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_9 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_6 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 1656 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_10 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 2024 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 3036 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_14
timestamp 1604489732
transform 1 0 2392 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[17\]
timestamp 1604489732
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_18 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35
timestamp 1604489732
transform 1 0 4324 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_26
timestamp 1604489732
transform 1 0 3496 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_38 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 4600 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[18\]
timestamp 1604489732
transform 1 0 5244 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[26\]
timestamp 1604489732
transform 1 0 5152 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604489732
transform -1 0 5980 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604489732
transform -1 0 5980 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43
timestamp 1604489732
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48
timestamp 1604489732
transform 1 0 5520 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_47
timestamp 1604489732
transform 1 0 5428 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[15\]
timestamp 1604489732
transform 1 0 1748 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[23\]
timestamp 1604489732
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[6\]
timestamp 1604489732
transform 1 0 2024 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604489732
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6
timestamp 1604489732
transform 1 0 1656 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_13
timestamp 1604489732
transform 1 0 2300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_25
timestamp 1604489732
transform 1 0 3404 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_19
timestamp 1604489732
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604489732
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604489732
transform -1 0 5980 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_44
timestamp 1604489732
transform 1 0 5152 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[25\]
timestamp 1604489732
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604489732
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_6
timestamp 1604489732
transform 1 0 1656 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[22\]
timestamp 1604489732
transform 1 0 2668 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[5\]
timestamp 1604489732
transform 1 0 3404 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_14
timestamp 1604489732
transform 1 0 2392 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_20
timestamp 1604489732
transform 1 0 2944 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_24
timestamp 1604489732
transform 1 0 3312 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[0\]
timestamp 1604489732
transform 1 0 4048 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[12\]
timestamp 1604489732
transform 1 0 4416 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[31\]
timestamp 1604489732
transform 1 0 3680 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_31
timestamp 1604489732
transform 1 0 3956 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_35
timestamp 1604489732
transform 1 0 4324 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[7\]
timestamp 1604489732
transform 1 0 5336 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604489732
transform -1 0 5980 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_39
timestamp 1604489732
transform 1 0 4692 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_45
timestamp 1604489732
transform 1 0 5244 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_49
timestamp 1604489732
transform 1 0 5612 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[10\]
timestamp 1604489732
transform 1 0 1472 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[1\]
timestamp 1604489732
transform 1 0 1748 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[8\]
timestamp 1604489732
transform 1 0 2024 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604489732
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1604489732
transform 1 0 1380 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[11\]
timestamp 1604489732
transform 1 0 2852 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_13
timestamp 1604489732
transform 1 0 2300 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_22
timestamp 1604489732
transform 1 0 3128 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_20
timestamp 1604489732
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_30
timestamp 1604489732
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604489732
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604489732
transform -1 0 5980 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_44
timestamp 1604489732
transform 1 0 5152 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604489732
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604489732
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[21\]
timestamp 1604489732
transform 1 0 2668 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[24\]
timestamp 1604489732
transform 1 0 2944 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_15
timestamp 1604489732
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_23
timestamp 1604489732
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_35
timestamp 1604489732
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[27\]
timestamp 1604489732
transform 1 0 5428 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604489732
transform -1 0 5980 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[30\]
timestamp 1604489732
transform 1 0 1840 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[3\]
timestamp 1604489732
transform 1 0 2116 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[4\]
timestamp 1604489732
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604489732
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604489732
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604489732
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_6
timestamp 1604489732
transform 1 0 1656 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[28\]
timestamp 1604489732
transform 1 0 2392 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_15
timestamp 1604489732
transform 1 0 2484 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_23
timestamp 1604489732
transform 1 0 3220 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_17
timestamp 1604489732
transform 1 0 2668 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[13\]
timestamp 1604489732
transform 1 0 3496 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[16\]
timestamp 1604489732
transform 1 0 4048 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_21
timestamp 1604489732
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1604489732
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_32
timestamp 1604489732
transform 1 0 4048 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_38
timestamp 1604489732
transform 1 0 4600 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_29
timestamp 1604489732
transform 1 0 3772 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_35
timestamp 1604489732
transform 1 0 4324 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_39
timestamp 1604489732
transform 1 0 4692 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_42
timestamp 1604489732
transform 1 0 4968 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[29\]
timestamp 1604489732
transform 1 0 4784 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[14\]
timestamp 1604489732
transform 1 0 4692 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_49
timestamp 1604489732
transform 1 0 5612 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_46
timestamp 1604489732
transform 1 0 5336 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604489732
transform -1 0 5980 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604489732
transform -1 0 5980 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[9\]
timestamp 1604489732
transform 1 0 5428 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_43
timestamp 1604489732
transform 1 0 5060 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604489732
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604489732
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604489732
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_22
timestamp 1604489732
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604489732
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604489732
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604489732
transform -1 0 5980 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_44
timestamp 1604489732
transform 1 0 5152 0 -1 7072
box -38 -48 590 592
<< labels >>
rlabel metal2 s 4618 8453 4674 9253 6 mask_rev[0]
port 0 nsew default tristate
rlabel metal2 s 4434 0 4490 800 6 mask_rev[10]
port 1 nsew default tristate
rlabel metal2 s 1122 0 1178 800 6 mask_rev[11]
port 2 nsew default tristate
rlabel metal2 s 570 0 626 800 6 mask_rev[12]
port 3 nsew default tristate
rlabel metal2 s 5906 8453 5962 9253 6 mask_rev[13]
port 4 nsew default tristate
rlabel metal2 s 6458 0 6514 800 6 mask_rev[14]
port 5 nsew default tristate
rlabel metal3 s 6309 2456 7109 2576 6 mask_rev[15]
port 6 nsew default tristate
rlabel metal2 s 2410 0 2466 800 6 mask_rev[16]
port 7 nsew default tristate
rlabel metal2 s 1858 8453 1914 9253 6 mask_rev[17]
port 8 nsew default tristate
rlabel metal3 s 0 7624 800 7744 6 mask_rev[18]
port 9 nsew default tristate
rlabel metal2 s 3330 8453 3386 9253 6 mask_rev[19]
port 10 nsew default tristate
rlabel metal3 s 0 2728 800 2848 6 mask_rev[1]
port 11 nsew default tristate
rlabel metal3 s 6309 3544 7109 3664 6 mask_rev[20]
port 12 nsew default tristate
rlabel metal3 s 6309 1368 7109 1488 6 mask_rev[21]
port 13 nsew default tristate
rlabel metal3 s 0 1640 800 1760 6 mask_rev[22]
port 14 nsew default tristate
rlabel metal2 s 1858 0 1914 800 6 mask_rev[23]
port 15 nsew default tristate
rlabel metal2 s 6458 8453 6514 9253 6 mask_rev[24]
port 16 nsew default tristate
rlabel metal3 s 0 3544 800 3664 6 mask_rev[25]
port 17 nsew default tristate
rlabel metal2 s 5170 8453 5226 9253 6 mask_rev[26]
port 18 nsew default tristate
rlabel metal2 s 1306 8453 1362 9253 6 mask_rev[27]
port 19 nsew default tristate
rlabel metal3 s 6309 7352 7109 7472 6 mask_rev[28]
port 20 nsew default tristate
rlabel metal2 s 5722 0 5778 800 6 mask_rev[29]
port 21 nsew default tristate
rlabel metal3 s 0 4632 800 4752 6 mask_rev[2]
port 22 nsew default tristate
rlabel metal3 s 6309 6264 7109 6384 6 mask_rev[30]
port 23 nsew default tristate
rlabel metal2 s 3146 0 3202 800 6 mask_rev[31]
port 24 nsew default tristate
rlabel metal2 s 3698 0 3754 800 6 mask_rev[3]
port 25 nsew default tristate
rlabel metal3 s 6309 4360 7109 4480 6 mask_rev[4]
port 26 nsew default tristate
rlabel metal3 s 6309 5448 7109 5568 6 mask_rev[5]
port 27 nsew default tristate
rlabel metal3 s 0 6536 800 6656 6 mask_rev[6]
port 28 nsew default tristate
rlabel metal2 s 3882 8453 3938 9253 6 mask_rev[7]
port 29 nsew default tristate
rlabel metal2 s 5170 0 5226 800 6 mask_rev[8]
port 30 nsew default tristate
rlabel metal2 s 2594 8453 2650 9253 6 mask_rev[9]
port 31 nsew default tristate
rlabel metal3 s 0 5448 800 5568 6 vdd1v8
port 32 nsew default bidirectional
rlabel metal2 s 570 8453 626 9253 6 vss
port 33 nsew default bidirectional
rlabel metal5 s 1104 2784 5980 3104 6 VPWR
port 34 nsew default input
rlabel metal5 s 1104 3600 5980 3920 6 VGND
port 35 nsew default input
<< properties >>
string FIXED_BBOX 0 0 7109 9253
<< end >>
