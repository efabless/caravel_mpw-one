VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_core
  CLASS BLOCK ;
  FOREIGN mgmt_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 2150.000 BY 900.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END clock
  PIN core_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 896.000 59.250 900.000 ;
    END
  END core_clk
  PIN core_rstn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 896.000 386.770 900.000 ;
    END
  END core_rstn
  PIN flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END flash_clk
  PIN flash_clk_ieb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END flash_clk_ieb
  PIN flash_clk_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END flash_clk_oeb
  PIN flash_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END flash_csb
  PIN flash_csb_ieb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END flash_csb_ieb
  PIN flash_csb_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END flash_csb_oeb
  PIN flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END flash_io0_di
  PIN flash_io0_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END flash_io0_do
  PIN flash_io0_ieb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END flash_io0_ieb
  PIN flash_io0_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END flash_io0_oeb
  PIN flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END flash_io1_di
  PIN flash_io1_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END flash_io1_do
  PIN flash_io1_ieb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END flash_io1_ieb
  PIN flash_io1_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END flash_io1_oeb
  PIN gpio_in_pad
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END gpio_in_pad
  PIN gpio_inenb_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END gpio_inenb_pad
  PIN gpio_mode0_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END gpio_mode0_pad
  PIN gpio_mode1_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END gpio_mode1_pad
  PIN gpio_out_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END gpio_out_pad
  PIN gpio_outenb_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END gpio_outenb_pad
  PIN jtag_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 337.320 2150.000 337.920 ;
    END
  END jtag_out
  PIN jtag_outenb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 334.600 2150.000 335.200 ;
    END
  END jtag_outenb
  PIN la_input[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 896.000 388.610 900.000 ;
    END
  END la_input[0]
  PIN la_input[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 896.000 384.930 900.000 ;
    END
  END la_input[100]
  PIN la_input[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 896.000 390.450 900.000 ;
    END
  END la_input[101]
  PIN la_input[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 896.000 383.090 900.000 ;
    END
  END la_input[102]
  PIN la_input[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 896.000 392.290 900.000 ;
    END
  END la_input[103]
  PIN la_input[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 896.000 381.250 900.000 ;
    END
  END la_input[104]
  PIN la_input[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 896.000 394.130 900.000 ;
    END
  END la_input[105]
  PIN la_input[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 896.000 379.410 900.000 ;
    END
  END la_input[106]
  PIN la_input[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 896.000 395.970 900.000 ;
    END
  END la_input[107]
  PIN la_input[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 896.000 377.570 900.000 ;
    END
  END la_input[108]
  PIN la_input[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 896.000 397.810 900.000 ;
    END
  END la_input[109]
  PIN la_input[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 896.000 375.730 900.000 ;
    END
  END la_input[10]
  PIN la_input[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 896.000 399.650 900.000 ;
    END
  END la_input[110]
  PIN la_input[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 896.000 373.890 900.000 ;
    END
  END la_input[111]
  PIN la_input[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 896.000 401.490 900.000 ;
    END
  END la_input[112]
  PIN la_input[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 896.000 372.050 900.000 ;
    END
  END la_input[113]
  PIN la_input[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 896.000 403.330 900.000 ;
    END
  END la_input[114]
  PIN la_input[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 896.000 370.210 900.000 ;
    END
  END la_input[115]
  PIN la_input[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 896.000 405.170 900.000 ;
    END
  END la_input[116]
  PIN la_input[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 896.000 368.370 900.000 ;
    END
  END la_input[117]
  PIN la_input[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.730 896.000 407.010 900.000 ;
    END
  END la_input[118]
  PIN la_input[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 896.000 366.530 900.000 ;
    END
  END la_input[119]
  PIN la_input[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 896.000 408.850 900.000 ;
    END
  END la_input[11]
  PIN la_input[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 896.000 364.690 900.000 ;
    END
  END la_input[120]
  PIN la_input[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 896.000 410.690 900.000 ;
    END
  END la_input[121]
  PIN la_input[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 896.000 362.850 900.000 ;
    END
  END la_input[122]
  PIN la_input[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 896.000 412.530 900.000 ;
    END
  END la_input[123]
  PIN la_input[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 896.000 361.010 900.000 ;
    END
  END la_input[124]
  PIN la_input[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 896.000 414.370 900.000 ;
    END
  END la_input[125]
  PIN la_input[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 896.000 359.170 900.000 ;
    END
  END la_input[126]
  PIN la_input[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 896.000 416.210 900.000 ;
    END
  END la_input[127]
  PIN la_input[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 896.000 357.330 900.000 ;
    END
  END la_input[12]
  PIN la_input[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 896.000 418.050 900.000 ;
    END
  END la_input[13]
  PIN la_input[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 896.000 355.490 900.000 ;
    END
  END la_input[14]
  PIN la_input[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.610 896.000 419.890 900.000 ;
    END
  END la_input[15]
  PIN la_input[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 896.000 353.650 900.000 ;
    END
  END la_input[16]
  PIN la_input[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 896.000 421.730 900.000 ;
    END
  END la_input[17]
  PIN la_input[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 896.000 351.810 900.000 ;
    END
  END la_input[18]
  PIN la_input[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 896.000 423.570 900.000 ;
    END
  END la_input[19]
  PIN la_input[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 896.000 349.970 900.000 ;
    END
  END la_input[1]
  PIN la_input[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 896.000 425.410 900.000 ;
    END
  END la_input[20]
  PIN la_input[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 896.000 348.130 900.000 ;
    END
  END la_input[21]
  PIN la_input[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 896.000 427.250 900.000 ;
    END
  END la_input[22]
  PIN la_input[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 896.000 346.290 900.000 ;
    END
  END la_input[23]
  PIN la_input[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 896.000 429.090 900.000 ;
    END
  END la_input[24]
  PIN la_input[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 896.000 344.450 900.000 ;
    END
  END la_input[25]
  PIN la_input[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 896.000 430.930 900.000 ;
    END
  END la_input[26]
  PIN la_input[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 896.000 342.610 900.000 ;
    END
  END la_input[27]
  PIN la_input[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 896.000 432.770 900.000 ;
    END
  END la_input[28]
  PIN la_input[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 896.000 340.770 900.000 ;
    END
  END la_input[29]
  PIN la_input[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 896.000 434.610 900.000 ;
    END
  END la_input[2]
  PIN la_input[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 896.000 338.930 900.000 ;
    END
  END la_input[30]
  PIN la_input[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 896.000 436.450 900.000 ;
    END
  END la_input[31]
  PIN la_input[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 896.000 337.090 900.000 ;
    END
  END la_input[32]
  PIN la_input[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 896.000 438.290 900.000 ;
    END
  END la_input[33]
  PIN la_input[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 896.000 335.250 900.000 ;
    END
  END la_input[34]
  PIN la_input[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 896.000 440.130 900.000 ;
    END
  END la_input[35]
  PIN la_input[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 896.000 333.410 900.000 ;
    END
  END la_input[36]
  PIN la_input[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 896.000 441.970 900.000 ;
    END
  END la_input[37]
  PIN la_input[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 896.000 331.570 900.000 ;
    END
  END la_input[38]
  PIN la_input[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 896.000 443.810 900.000 ;
    END
  END la_input[39]
  PIN la_input[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 896.000 329.730 900.000 ;
    END
  END la_input[3]
  PIN la_input[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 896.000 445.650 900.000 ;
    END
  END la_input[40]
  PIN la_input[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 896.000 327.890 900.000 ;
    END
  END la_input[41]
  PIN la_input[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 896.000 447.490 900.000 ;
    END
  END la_input[42]
  PIN la_input[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 896.000 326.050 900.000 ;
    END
  END la_input[43]
  PIN la_input[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 896.000 449.330 900.000 ;
    END
  END la_input[44]
  PIN la_input[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 896.000 324.210 900.000 ;
    END
  END la_input[45]
  PIN la_input[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 896.000 451.170 900.000 ;
    END
  END la_input[46]
  PIN la_input[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 896.000 322.370 900.000 ;
    END
  END la_input[47]
  PIN la_input[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 896.000 453.010 900.000 ;
    END
  END la_input[48]
  PIN la_input[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 896.000 320.530 900.000 ;
    END
  END la_input[49]
  PIN la_input[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 896.000 454.850 900.000 ;
    END
  END la_input[4]
  PIN la_input[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 896.000 318.690 900.000 ;
    END
  END la_input[50]
  PIN la_input[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 896.000 456.690 900.000 ;
    END
  END la_input[51]
  PIN la_input[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 896.000 316.850 900.000 ;
    END
  END la_input[52]
  PIN la_input[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 896.000 458.530 900.000 ;
    END
  END la_input[53]
  PIN la_input[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 896.000 315.010 900.000 ;
    END
  END la_input[54]
  PIN la_input[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 896.000 460.370 900.000 ;
    END
  END la_input[55]
  PIN la_input[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 896.000 313.170 900.000 ;
    END
  END la_input[56]
  PIN la_input[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.930 896.000 462.210 900.000 ;
    END
  END la_input[57]
  PIN la_input[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 896.000 311.330 900.000 ;
    END
  END la_input[58]
  PIN la_input[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 896.000 464.050 900.000 ;
    END
  END la_input[59]
  PIN la_input[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 896.000 309.490 900.000 ;
    END
  END la_input[5]
  PIN la_input[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 896.000 465.890 900.000 ;
    END
  END la_input[60]
  PIN la_input[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 896.000 307.650 900.000 ;
    END
  END la_input[61]
  PIN la_input[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 896.000 467.730 900.000 ;
    END
  END la_input[62]
  PIN la_input[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 896.000 305.810 900.000 ;
    END
  END la_input[63]
  PIN la_input[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 896.000 469.570 900.000 ;
    END
  END la_input[64]
  PIN la_input[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 896.000 303.970 900.000 ;
    END
  END la_input[65]
  PIN la_input[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 896.000 471.410 900.000 ;
    END
  END la_input[66]
  PIN la_input[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 896.000 302.130 900.000 ;
    END
  END la_input[67]
  PIN la_input[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 896.000 473.250 900.000 ;
    END
  END la_input[68]
  PIN la_input[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 896.000 300.290 900.000 ;
    END
  END la_input[69]
  PIN la_input[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 896.000 475.090 900.000 ;
    END
  END la_input[6]
  PIN la_input[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 896.000 298.450 900.000 ;
    END
  END la_input[70]
  PIN la_input[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 896.000 476.930 900.000 ;
    END
  END la_input[71]
  PIN la_input[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 896.000 296.610 900.000 ;
    END
  END la_input[72]
  PIN la_input[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 896.000 478.770 900.000 ;
    END
  END la_input[73]
  PIN la_input[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 896.000 294.770 900.000 ;
    END
  END la_input[74]
  PIN la_input[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 896.000 480.610 900.000 ;
    END
  END la_input[75]
  PIN la_input[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 896.000 292.930 900.000 ;
    END
  END la_input[76]
  PIN la_input[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 896.000 482.450 900.000 ;
    END
  END la_input[77]
  PIN la_input[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 896.000 291.090 900.000 ;
    END
  END la_input[78]
  PIN la_input[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 896.000 484.290 900.000 ;
    END
  END la_input[79]
  PIN la_input[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 896.000 289.250 900.000 ;
    END
  END la_input[7]
  PIN la_input[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 896.000 486.130 900.000 ;
    END
  END la_input[80]
  PIN la_input[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 896.000 287.410 900.000 ;
    END
  END la_input[81]
  PIN la_input[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 896.000 487.970 900.000 ;
    END
  END la_input[82]
  PIN la_input[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 896.000 285.570 900.000 ;
    END
  END la_input[83]
  PIN la_input[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 896.000 489.810 900.000 ;
    END
  END la_input[84]
  PIN la_input[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 896.000 283.730 900.000 ;
    END
  END la_input[85]
  PIN la_input[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 896.000 491.650 900.000 ;
    END
  END la_input[86]
  PIN la_input[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 896.000 281.890 900.000 ;
    END
  END la_input[87]
  PIN la_input[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 896.000 493.490 900.000 ;
    END
  END la_input[88]
  PIN la_input[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 896.000 280.050 900.000 ;
    END
  END la_input[89]
  PIN la_input[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 896.000 495.330 900.000 ;
    END
  END la_input[8]
  PIN la_input[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 896.000 278.210 900.000 ;
    END
  END la_input[90]
  PIN la_input[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 896.000 497.170 900.000 ;
    END
  END la_input[91]
  PIN la_input[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 896.000 276.370 900.000 ;
    END
  END la_input[92]
  PIN la_input[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 896.000 499.010 900.000 ;
    END
  END la_input[93]
  PIN la_input[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 896.000 274.530 900.000 ;
    END
  END la_input[94]
  PIN la_input[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 896.000 500.850 900.000 ;
    END
  END la_input[95]
  PIN la_input[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 896.000 272.690 900.000 ;
    END
  END la_input[96]
  PIN la_input[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 896.000 502.690 900.000 ;
    END
  END la_input[97]
  PIN la_input[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 896.000 270.850 900.000 ;
    END
  END la_input[98]
  PIN la_input[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 896.000 504.530 900.000 ;
    END
  END la_input[99]
  PIN la_input[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 896.000 269.010 900.000 ;
    END
  END la_input[9]
  PIN la_oen[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 896.000 506.370 900.000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 896.000 267.170 900.000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 896.000 508.210 900.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 896.000 265.330 900.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 896.000 510.050 900.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 896.000 263.490 900.000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.610 896.000 511.890 900.000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 896.000 261.650 900.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 896.000 513.730 900.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 896.000 259.810 900.000 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 896.000 515.570 900.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 896.000 257.970 900.000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 896.000 517.410 900.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 896.000 256.130 900.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 896.000 519.250 900.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 896.000 254.290 900.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 896.000 521.090 900.000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 896.000 252.450 900.000 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 896.000 522.930 900.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 896.000 250.610 900.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 896.000 524.770 900.000 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 896.000 248.770 900.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 896.000 526.610 900.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 896.000 246.930 900.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 896.000 528.450 900.000 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 896.000 245.090 900.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 896.000 530.290 900.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 896.000 243.250 900.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 896.000 532.130 900.000 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 896.000 241.410 900.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 896.000 533.970 900.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 896.000 239.570 900.000 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 896.000 535.810 900.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 896.000 237.730 900.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 896.000 537.650 900.000 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 896.000 235.890 900.000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 896.000 539.490 900.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 896.000 234.050 900.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 896.000 541.330 900.000 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 896.000 232.210 900.000 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 896.000 543.170 900.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 896.000 230.370 900.000 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 896.000 545.010 900.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 896.000 228.530 900.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.570 896.000 546.850 900.000 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 896.000 226.690 900.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.410 896.000 548.690 900.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 896.000 224.850 900.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 896.000 550.530 900.000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 896.000 223.010 900.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 896.000 552.370 900.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 896.000 221.170 900.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 896.000 554.210 900.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 896.000 219.330 900.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 896.000 556.050 900.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 896.000 217.490 900.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 896.000 557.890 900.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 896.000 215.650 900.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 896.000 559.730 900.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 896.000 213.810 900.000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 896.000 561.570 900.000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 896.000 211.970 900.000 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.130 896.000 563.410 900.000 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 896.000 210.130 900.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 896.000 565.250 900.000 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 896.000 208.290 900.000 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 896.000 567.090 900.000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 896.000 206.450 900.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.650 896.000 568.930 900.000 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 896.000 204.610 900.000 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 896.000 570.770 900.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 896.000 202.770 900.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.330 896.000 572.610 900.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 896.000 200.930 900.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 896.000 574.450 900.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 896.000 199.090 900.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 896.000 576.290 900.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 896.000 197.250 900.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 896.000 578.130 900.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 896.000 195.410 900.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 896.000 579.970 900.000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 896.000 193.570 900.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 896.000 581.810 900.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 896.000 191.730 900.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.370 896.000 583.650 900.000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 896.000 189.890 900.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 896.000 585.490 900.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 896.000 188.050 900.000 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 896.000 587.330 900.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 896.000 186.210 900.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 896.000 589.170 900.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 896.000 184.370 900.000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 896.000 591.010 900.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 896.000 182.530 900.000 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 896.000 592.850 900.000 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 896.000 180.690 900.000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 896.000 594.690 900.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 896.000 178.850 900.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 896.000 596.530 900.000 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 896.000 177.010 900.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 896.000 598.370 900.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 896.000 175.170 900.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 896.000 600.210 900.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 896.000 173.330 900.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.770 896.000 602.050 900.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 896.000 171.490 900.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.610 896.000 603.890 900.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 896.000 169.650 900.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 896.000 605.730 900.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 896.000 167.810 900.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.290 896.000 607.570 900.000 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 896.000 165.970 900.000 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 896.000 609.410 900.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 896.000 164.130 900.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 896.000 611.250 900.000 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 896.000 162.290 900.000 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 896.000 613.090 900.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 896.000 160.450 900.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.650 896.000 614.930 900.000 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 896.000 158.610 900.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.490 896.000 616.770 900.000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 896.000 156.770 900.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 896.000 618.610 900.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 896.000 154.930 900.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.170 896.000 620.450 900.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 896.000 153.090 900.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.010 896.000 622.290 900.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 896.000 151.250 900.000 ;
    END
  END la_oen[9]
  PIN la_output[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 896.000 624.130 900.000 ;
    END
  END la_output[0]
  PIN la_output[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 896.000 149.410 900.000 ;
    END
  END la_output[100]
  PIN la_output[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 896.000 625.970 900.000 ;
    END
  END la_output[101]
  PIN la_output[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 896.000 147.570 900.000 ;
    END
  END la_output[102]
  PIN la_output[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 896.000 627.810 900.000 ;
    END
  END la_output[103]
  PIN la_output[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 896.000 145.730 900.000 ;
    END
  END la_output[104]
  PIN la_output[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.370 896.000 629.650 900.000 ;
    END
  END la_output[105]
  PIN la_output[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 896.000 143.890 900.000 ;
    END
  END la_output[106]
  PIN la_output[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 896.000 631.490 900.000 ;
    END
  END la_output[107]
  PIN la_output[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 896.000 142.050 900.000 ;
    END
  END la_output[108]
  PIN la_output[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.050 896.000 633.330 900.000 ;
    END
  END la_output[109]
  PIN la_output[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 896.000 140.210 900.000 ;
    END
  END la_output[10]
  PIN la_output[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 896.000 635.170 900.000 ;
    END
  END la_output[110]
  PIN la_output[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 896.000 138.370 900.000 ;
    END
  END la_output[111]
  PIN la_output[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.730 896.000 637.010 900.000 ;
    END
  END la_output[112]
  PIN la_output[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 896.000 136.530 900.000 ;
    END
  END la_output[113]
  PIN la_output[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 896.000 638.850 900.000 ;
    END
  END la_output[114]
  PIN la_output[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 896.000 134.690 900.000 ;
    END
  END la_output[115]
  PIN la_output[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 896.000 640.690 900.000 ;
    END
  END la_output[116]
  PIN la_output[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 896.000 132.850 900.000 ;
    END
  END la_output[117]
  PIN la_output[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.250 896.000 642.530 900.000 ;
    END
  END la_output[118]
  PIN la_output[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 896.000 131.010 900.000 ;
    END
  END la_output[119]
  PIN la_output[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 896.000 644.370 900.000 ;
    END
  END la_output[11]
  PIN la_output[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 896.000 129.170 900.000 ;
    END
  END la_output[120]
  PIN la_output[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 896.000 646.210 900.000 ;
    END
  END la_output[121]
  PIN la_output[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 896.000 127.330 900.000 ;
    END
  END la_output[122]
  PIN la_output[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.770 896.000 648.050 900.000 ;
    END
  END la_output[123]
  PIN la_output[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 896.000 125.490 900.000 ;
    END
  END la_output[124]
  PIN la_output[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 896.000 649.890 900.000 ;
    END
  END la_output[125]
  PIN la_output[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 896.000 123.650 900.000 ;
    END
  END la_output[126]
  PIN la_output[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.450 896.000 651.730 900.000 ;
    END
  END la_output[127]
  PIN la_output[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 896.000 121.810 900.000 ;
    END
  END la_output[12]
  PIN la_output[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 896.000 653.570 900.000 ;
    END
  END la_output[13]
  PIN la_output[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 896.000 119.970 900.000 ;
    END
  END la_output[14]
  PIN la_output[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.130 896.000 655.410 900.000 ;
    END
  END la_output[15]
  PIN la_output[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 896.000 118.130 900.000 ;
    END
  END la_output[16]
  PIN la_output[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 896.000 657.250 900.000 ;
    END
  END la_output[17]
  PIN la_output[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 896.000 116.290 900.000 ;
    END
  END la_output[18]
  PIN la_output[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.810 896.000 659.090 900.000 ;
    END
  END la_output[19]
  PIN la_output[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 896.000 114.450 900.000 ;
    END
  END la_output[1]
  PIN la_output[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 896.000 660.930 900.000 ;
    END
  END la_output[20]
  PIN la_output[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 896.000 112.610 900.000 ;
    END
  END la_output[21]
  PIN la_output[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 896.000 662.770 900.000 ;
    END
  END la_output[22]
  PIN la_output[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 896.000 110.770 900.000 ;
    END
  END la_output[23]
  PIN la_output[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.330 896.000 664.610 900.000 ;
    END
  END la_output[24]
  PIN la_output[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 896.000 108.930 900.000 ;
    END
  END la_output[25]
  PIN la_output[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.170 896.000 666.450 900.000 ;
    END
  END la_output[26]
  PIN la_output[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 896.000 107.090 900.000 ;
    END
  END la_output[27]
  PIN la_output[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.010 896.000 668.290 900.000 ;
    END
  END la_output[28]
  PIN la_output[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 896.000 105.250 900.000 ;
    END
  END la_output[29]
  PIN la_output[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 896.000 670.130 900.000 ;
    END
  END la_output[2]
  PIN la_output[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 896.000 103.410 900.000 ;
    END
  END la_output[30]
  PIN la_output[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.690 896.000 671.970 900.000 ;
    END
  END la_output[31]
  PIN la_output[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 896.000 101.570 900.000 ;
    END
  END la_output[32]
  PIN la_output[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 896.000 673.810 900.000 ;
    END
  END la_output[33]
  PIN la_output[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 896.000 99.730 900.000 ;
    END
  END la_output[34]
  PIN la_output[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.370 896.000 675.650 900.000 ;
    END
  END la_output[35]
  PIN la_output[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 896.000 97.890 900.000 ;
    END
  END la_output[36]
  PIN la_output[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.210 896.000 677.490 900.000 ;
    END
  END la_output[37]
  PIN la_output[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 896.000 96.050 900.000 ;
    END
  END la_output[38]
  PIN la_output[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 896.000 679.330 900.000 ;
    END
  END la_output[39]
  PIN la_output[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 896.000 94.210 900.000 ;
    END
  END la_output[3]
  PIN la_output[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.890 896.000 681.170 900.000 ;
    END
  END la_output[40]
  PIN la_output[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 896.000 92.370 900.000 ;
    END
  END la_output[41]
  PIN la_output[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 896.000 683.010 900.000 ;
    END
  END la_output[42]
  PIN la_output[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 896.000 90.530 900.000 ;
    END
  END la_output[43]
  PIN la_output[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.570 896.000 684.850 900.000 ;
    END
  END la_output[44]
  PIN la_output[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 896.000 88.690 900.000 ;
    END
  END la_output[45]
  PIN la_output[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 896.000 686.690 900.000 ;
    END
  END la_output[46]
  PIN la_output[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 896.000 86.850 900.000 ;
    END
  END la_output[47]
  PIN la_output[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 896.000 688.530 900.000 ;
    END
  END la_output[48]
  PIN la_output[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 896.000 85.010 900.000 ;
    END
  END la_output[49]
  PIN la_output[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 896.000 690.370 900.000 ;
    END
  END la_output[4]
  PIN la_output[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 896.000 83.170 900.000 ;
    END
  END la_output[50]
  PIN la_output[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.930 896.000 692.210 900.000 ;
    END
  END la_output[51]
  PIN la_output[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 896.000 81.330 900.000 ;
    END
  END la_output[52]
  PIN la_output[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 896.000 694.050 900.000 ;
    END
  END la_output[53]
  PIN la_output[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 896.000 79.490 900.000 ;
    END
  END la_output[54]
  PIN la_output[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 896.000 695.890 900.000 ;
    END
  END la_output[55]
  PIN la_output[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 896.000 77.650 900.000 ;
    END
  END la_output[56]
  PIN la_output[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 896.000 697.730 900.000 ;
    END
  END la_output[57]
  PIN la_output[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 896.000 75.810 900.000 ;
    END
  END la_output[58]
  PIN la_output[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 896.000 699.570 900.000 ;
    END
  END la_output[59]
  PIN la_output[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 896.000 73.970 900.000 ;
    END
  END la_output[5]
  PIN la_output[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.130 896.000 701.410 900.000 ;
    END
  END la_output[60]
  PIN la_output[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 896.000 72.130 900.000 ;
    END
  END la_output[61]
  PIN la_output[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.970 896.000 703.250 900.000 ;
    END
  END la_output[62]
  PIN la_output[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 896.000 70.290 900.000 ;
    END
  END la_output[63]
  PIN la_output[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.810 896.000 705.090 900.000 ;
    END
  END la_output[64]
  PIN la_output[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 896.000 68.450 900.000 ;
    END
  END la_output[65]
  PIN la_output[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.650 896.000 706.930 900.000 ;
    END
  END la_output[66]
  PIN la_output[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 896.000 66.610 900.000 ;
    END
  END la_output[67]
  PIN la_output[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 896.000 708.770 900.000 ;
    END
  END la_output[68]
  PIN la_output[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 896.000 64.770 900.000 ;
    END
  END la_output[69]
  PIN la_output[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 896.000 710.610 900.000 ;
    END
  END la_output[6]
  PIN la_output[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 896.000 62.930 900.000 ;
    END
  END la_output[70]
  PIN la_output[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 896.000 712.450 900.000 ;
    END
  END la_output[71]
  PIN la_output[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 896.000 61.090 900.000 ;
    END
  END la_output[72]
  PIN la_output[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.010 896.000 714.290 900.000 ;
    END
  END la_output[73]
  PIN la_output[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 896.000 716.130 900.000 ;
    END
  END la_output[74]
  PIN la_output[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 896.000 57.410 900.000 ;
    END
  END la_output[75]
  PIN la_output[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 896.000 717.970 900.000 ;
    END
  END la_output[76]
  PIN la_output[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 896.000 55.570 900.000 ;
    END
  END la_output[77]
  PIN la_output[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.530 896.000 719.810 900.000 ;
    END
  END la_output[78]
  PIN la_output[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 896.000 53.730 900.000 ;
    END
  END la_output[79]
  PIN la_output[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 896.000 721.650 900.000 ;
    END
  END la_output[7]
  PIN la_output[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 896.000 51.890 900.000 ;
    END
  END la_output[80]
  PIN la_output[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 896.000 723.490 900.000 ;
    END
  END la_output[81]
  PIN la_output[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 896.000 50.050 900.000 ;
    END
  END la_output[82]
  PIN la_output[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 896.000 725.330 900.000 ;
    END
  END la_output[83]
  PIN la_output[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 896.000 48.210 900.000 ;
    END
  END la_output[84]
  PIN la_output[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.890 896.000 727.170 900.000 ;
    END
  END la_output[85]
  PIN la_output[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 896.000 46.370 900.000 ;
    END
  END la_output[86]
  PIN la_output[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.730 896.000 729.010 900.000 ;
    END
  END la_output[87]
  PIN la_output[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 896.000 44.530 900.000 ;
    END
  END la_output[88]
  PIN la_output[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.570 896.000 730.850 900.000 ;
    END
  END la_output[89]
  PIN la_output[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 896.000 42.690 900.000 ;
    END
  END la_output[8]
  PIN la_output[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.410 896.000 732.690 900.000 ;
    END
  END la_output[90]
  PIN la_output[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 896.000 40.850 900.000 ;
    END
  END la_output[91]
  PIN la_output[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 896.000 734.530 900.000 ;
    END
  END la_output[92]
  PIN la_output[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 896.000 39.010 900.000 ;
    END
  END la_output[93]
  PIN la_output[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.090 896.000 736.370 900.000 ;
    END
  END la_output[94]
  PIN la_output[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 896.000 37.170 900.000 ;
    END
  END la_output[95]
  PIN la_output[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 896.000 738.210 900.000 ;
    END
  END la_output[96]
  PIN la_output[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 896.000 35.330 900.000 ;
    END
  END la_output[97]
  PIN la_output[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.770 896.000 740.050 900.000 ;
    END
  END la_output[98]
  PIN la_output[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 896.000 33.490 900.000 ;
    END
  END la_output[99]
  PIN la_output[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 896.000 741.890 900.000 ;
    END
  END la_output[9]
  PIN mask_rev[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 136.040 2150.000 136.640 ;
    END
  END mask_rev[0]
  PIN mask_rev[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 133.320 2150.000 133.920 ;
    END
  END mask_rev[10]
  PIN mask_rev[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 138.760 2150.000 139.360 ;
    END
  END mask_rev[11]
  PIN mask_rev[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 130.600 2150.000 131.200 ;
    END
  END mask_rev[12]
  PIN mask_rev[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 141.480 2150.000 142.080 ;
    END
  END mask_rev[13]
  PIN mask_rev[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 127.880 2150.000 128.480 ;
    END
  END mask_rev[14]
  PIN mask_rev[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 144.200 2150.000 144.800 ;
    END
  END mask_rev[15]
  PIN mask_rev[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 125.160 2150.000 125.760 ;
    END
  END mask_rev[16]
  PIN mask_rev[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 146.920 2150.000 147.520 ;
    END
  END mask_rev[17]
  PIN mask_rev[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 122.440 2150.000 123.040 ;
    END
  END mask_rev[18]
  PIN mask_rev[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 149.640 2150.000 150.240 ;
    END
  END mask_rev[19]
  PIN mask_rev[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 119.720 2150.000 120.320 ;
    END
  END mask_rev[1]
  PIN mask_rev[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 152.360 2150.000 152.960 ;
    END
  END mask_rev[20]
  PIN mask_rev[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 117.000 2150.000 117.600 ;
    END
  END mask_rev[21]
  PIN mask_rev[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 155.080 2150.000 155.680 ;
    END
  END mask_rev[22]
  PIN mask_rev[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 114.280 2150.000 114.880 ;
    END
  END mask_rev[23]
  PIN mask_rev[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 157.800 2150.000 158.400 ;
    END
  END mask_rev[24]
  PIN mask_rev[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 111.560 2150.000 112.160 ;
    END
  END mask_rev[25]
  PIN mask_rev[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 160.520 2150.000 161.120 ;
    END
  END mask_rev[26]
  PIN mask_rev[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 108.840 2150.000 109.440 ;
    END
  END mask_rev[27]
  PIN mask_rev[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 163.240 2150.000 163.840 ;
    END
  END mask_rev[28]
  PIN mask_rev[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 106.120 2150.000 106.720 ;
    END
  END mask_rev[29]
  PIN mask_rev[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 165.960 2150.000 166.560 ;
    END
  END mask_rev[2]
  PIN mask_rev[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 103.400 2150.000 104.000 ;
    END
  END mask_rev[30]
  PIN mask_rev[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 168.680 2150.000 169.280 ;
    END
  END mask_rev[31]
  PIN mask_rev[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 100.680 2150.000 101.280 ;
    END
  END mask_rev[3]
  PIN mask_rev[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 171.400 2150.000 172.000 ;
    END
  END mask_rev[4]
  PIN mask_rev[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 97.960 2150.000 98.560 ;
    END
  END mask_rev[5]
  PIN mask_rev[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 174.120 2150.000 174.720 ;
    END
  END mask_rev[6]
  PIN mask_rev[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 95.240 2150.000 95.840 ;
    END
  END mask_rev[7]
  PIN mask_rev[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 176.840 2150.000 177.440 ;
    END
  END mask_rev[8]
  PIN mask_rev[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 92.520 2150.000 93.120 ;
    END
  END mask_rev[9]
  PIN mgmt_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END mgmt_addr[0]
  PIN mgmt_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END mgmt_addr[1]
  PIN mgmt_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END mgmt_addr[2]
  PIN mgmt_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END mgmt_addr[3]
  PIN mgmt_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END mgmt_addr[4]
  PIN mgmt_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END mgmt_addr[5]
  PIN mgmt_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END mgmt_addr[6]
  PIN mgmt_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END mgmt_addr[7]
  PIN mgmt_addr_ro[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END mgmt_addr_ro[0]
  PIN mgmt_addr_ro[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END mgmt_addr_ro[1]
  PIN mgmt_addr_ro[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END mgmt_addr_ro[2]
  PIN mgmt_addr_ro[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END mgmt_addr_ro[3]
  PIN mgmt_addr_ro[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END mgmt_addr_ro[4]
  PIN mgmt_addr_ro[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END mgmt_addr_ro[5]
  PIN mgmt_addr_ro[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END mgmt_addr_ro[6]
  PIN mgmt_addr_ro[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END mgmt_addr_ro[7]
  PIN mgmt_ena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END mgmt_ena[0]
  PIN mgmt_ena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END mgmt_ena[1]
  PIN mgmt_ena_ro
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END mgmt_ena_ro
  PIN mgmt_in_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 340.040 2150.000 340.640 ;
    END
  END mgmt_in_data[0]
  PIN mgmt_in_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END mgmt_in_data[10]
  PIN mgmt_in_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END mgmt_in_data[11]
  PIN mgmt_in_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END mgmt_in_data[12]
  PIN mgmt_in_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END mgmt_in_data[13]
  PIN mgmt_in_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END mgmt_in_data[14]
  PIN mgmt_in_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END mgmt_in_data[15]
  PIN mgmt_in_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END mgmt_in_data[16]
  PIN mgmt_in_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END mgmt_in_data[17]
  PIN mgmt_in_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END mgmt_in_data[18]
  PIN mgmt_in_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END mgmt_in_data[19]
  PIN mgmt_in_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 563.080 2150.000 563.680 ;
    END
  END mgmt_in_data[1]
  PIN mgmt_in_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END mgmt_in_data[20]
  PIN mgmt_in_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END mgmt_in_data[21]
  PIN mgmt_in_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END mgmt_in_data[22]
  PIN mgmt_in_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END mgmt_in_data[23]
  PIN mgmt_in_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END mgmt_in_data[24]
  PIN mgmt_in_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END mgmt_in_data[25]
  PIN mgmt_in_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END mgmt_in_data[26]
  PIN mgmt_in_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END mgmt_in_data[27]
  PIN mgmt_in_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END mgmt_in_data[28]
  PIN mgmt_in_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END mgmt_in_data[29]
  PIN mgmt_in_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END mgmt_in_data[2]
  PIN mgmt_in_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END mgmt_in_data[30]
  PIN mgmt_in_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END mgmt_in_data[31]
  PIN mgmt_in_data[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END mgmt_in_data[32]
  PIN mgmt_in_data[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END mgmt_in_data[33]
  PIN mgmt_in_data[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END mgmt_in_data[34]
  PIN mgmt_in_data[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END mgmt_in_data[35]
  PIN mgmt_in_data[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END mgmt_in_data[36]
  PIN mgmt_in_data[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END mgmt_in_data[37]
  PIN mgmt_in_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END mgmt_in_data[3]
  PIN mgmt_in_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END mgmt_in_data[4]
  PIN mgmt_in_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END mgmt_in_data[5]
  PIN mgmt_in_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END mgmt_in_data[6]
  PIN mgmt_in_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END mgmt_in_data[7]
  PIN mgmt_in_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END mgmt_in_data[8]
  PIN mgmt_in_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END mgmt_in_data[9]
  PIN mgmt_out_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END mgmt_out_data[0]
  PIN mgmt_out_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2145.530 896.000 2145.810 900.000 ;
    END
  END mgmt_out_data[10]
  PIN mgmt_out_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 894.920 2150.000 895.520 ;
    END
  END mgmt_out_data[11]
  PIN mgmt_out_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2143.690 896.000 2143.970 900.000 ;
    END
  END mgmt_out_data[12]
  PIN mgmt_out_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 892.200 2150.000 892.800 ;
    END
  END mgmt_out_data[13]
  PIN mgmt_out_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2141.850 896.000 2142.130 900.000 ;
    END
  END mgmt_out_data[14]
  PIN mgmt_out_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1692.890 896.000 1693.170 900.000 ;
    END
  END mgmt_out_data[15]
  PIN mgmt_out_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.290 896.000 1435.570 900.000 ;
    END
  END mgmt_out_data[16]
  PIN mgmt_out_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.730 896.000 1051.010 900.000 ;
    END
  END mgmt_out_data[17]
  PIN mgmt_out_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.450 896.000 743.730 900.000 ;
    END
  END mgmt_out_data[18]
  PIN mgmt_out_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 896.000 745.570 900.000 ;
    END
  END mgmt_out_data[19]
  PIN mgmt_out_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END mgmt_out_data[1]
  PIN mgmt_out_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 896.000 31.650 900.000 ;
    END
  END mgmt_out_data[20]
  PIN mgmt_out_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 896.000 4.050 900.000 ;
    END
  END mgmt_out_data[21]
  PIN mgmt_out_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.920 4.000 895.520 ;
    END
  END mgmt_out_data[22]
  PIN mgmt_out_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 896.000 5.890 900.000 ;
    END
  END mgmt_out_data[23]
  PIN mgmt_out_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.200 4.000 892.800 ;
    END
  END mgmt_out_data[24]
  PIN mgmt_out_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 896.000 7.730 900.000 ;
    END
  END mgmt_out_data[25]
  PIN mgmt_out_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 896.000 9.570 900.000 ;
    END
  END mgmt_out_data[26]
  PIN mgmt_out_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 889.480 4.000 890.080 ;
    END
  END mgmt_out_data[27]
  PIN mgmt_out_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 896.000 11.410 900.000 ;
    END
  END mgmt_out_data[28]
  PIN mgmt_out_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 886.760 4.000 887.360 ;
    END
  END mgmt_out_data[29]
  PIN mgmt_out_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 786.120 2150.000 786.720 ;
    END
  END mgmt_out_data[2]
  PIN mgmt_out_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 896.000 13.250 900.000 ;
    END
  END mgmt_out_data[30]
  PIN mgmt_out_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 896.000 15.090 900.000 ;
    END
  END mgmt_out_data[31]
  PIN mgmt_out_data[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END mgmt_out_data[32]
  PIN mgmt_out_data[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 896.000 16.930 900.000 ;
    END
  END mgmt_out_data[33]
  PIN mgmt_out_data[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 881.320 4.000 881.920 ;
    END
  END mgmt_out_data[34]
  PIN mgmt_out_data[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 896.000 18.770 900.000 ;
    END
  END mgmt_out_data[35]
  PIN mgmt_out_data[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 896.000 20.610 900.000 ;
    END
  END mgmt_out_data[36]
  PIN mgmt_out_data[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 745.320 4.000 745.920 ;
    END
  END mgmt_out_data[37]
  PIN mgmt_out_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2140.010 896.000 2140.290 900.000 ;
    END
  END mgmt_out_data[3]
  PIN mgmt_out_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 889.480 2150.000 890.080 ;
    END
  END mgmt_out_data[4]
  PIN mgmt_out_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2138.170 896.000 2138.450 900.000 ;
    END
  END mgmt_out_data[5]
  PIN mgmt_out_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 886.760 2150.000 887.360 ;
    END
  END mgmt_out_data[6]
  PIN mgmt_out_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.330 896.000 2136.610 900.000 ;
    END
  END mgmt_out_data[7]
  PIN mgmt_out_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2134.490 896.000 2134.770 900.000 ;
    END
  END mgmt_out_data[8]
  PIN mgmt_out_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 884.040 2150.000 884.640 ;
    END
  END mgmt_out_data[9]
  PIN mgmt_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END mgmt_rdata[0]
  PIN mgmt_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END mgmt_rdata[10]
  PIN mgmt_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END mgmt_rdata[11]
  PIN mgmt_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END mgmt_rdata[12]
  PIN mgmt_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END mgmt_rdata[13]
  PIN mgmt_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END mgmt_rdata[14]
  PIN mgmt_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END mgmt_rdata[15]
  PIN mgmt_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END mgmt_rdata[16]
  PIN mgmt_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END mgmt_rdata[17]
  PIN mgmt_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END mgmt_rdata[18]
  PIN mgmt_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END mgmt_rdata[19]
  PIN mgmt_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END mgmt_rdata[1]
  PIN mgmt_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END mgmt_rdata[20]
  PIN mgmt_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END mgmt_rdata[21]
  PIN mgmt_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END mgmt_rdata[22]
  PIN mgmt_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END mgmt_rdata[23]
  PIN mgmt_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END mgmt_rdata[24]
  PIN mgmt_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END mgmt_rdata[25]
  PIN mgmt_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END mgmt_rdata[26]
  PIN mgmt_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END mgmt_rdata[27]
  PIN mgmt_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END mgmt_rdata[28]
  PIN mgmt_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END mgmt_rdata[29]
  PIN mgmt_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END mgmt_rdata[2]
  PIN mgmt_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END mgmt_rdata[30]
  PIN mgmt_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END mgmt_rdata[31]
  PIN mgmt_rdata[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END mgmt_rdata[32]
  PIN mgmt_rdata[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END mgmt_rdata[33]
  PIN mgmt_rdata[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END mgmt_rdata[34]
  PIN mgmt_rdata[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END mgmt_rdata[35]
  PIN mgmt_rdata[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END mgmt_rdata[36]
  PIN mgmt_rdata[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END mgmt_rdata[37]
  PIN mgmt_rdata[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END mgmt_rdata[38]
  PIN mgmt_rdata[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END mgmt_rdata[39]
  PIN mgmt_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END mgmt_rdata[3]
  PIN mgmt_rdata[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END mgmt_rdata[40]
  PIN mgmt_rdata[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END mgmt_rdata[41]
  PIN mgmt_rdata[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END mgmt_rdata[42]
  PIN mgmt_rdata[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END mgmt_rdata[43]
  PIN mgmt_rdata[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END mgmt_rdata[44]
  PIN mgmt_rdata[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END mgmt_rdata[45]
  PIN mgmt_rdata[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END mgmt_rdata[46]
  PIN mgmt_rdata[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END mgmt_rdata[47]
  PIN mgmt_rdata[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END mgmt_rdata[48]
  PIN mgmt_rdata[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END mgmt_rdata[49]
  PIN mgmt_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END mgmt_rdata[4]
  PIN mgmt_rdata[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END mgmt_rdata[50]
  PIN mgmt_rdata[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END mgmt_rdata[51]
  PIN mgmt_rdata[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END mgmt_rdata[52]
  PIN mgmt_rdata[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END mgmt_rdata[53]
  PIN mgmt_rdata[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END mgmt_rdata[54]
  PIN mgmt_rdata[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END mgmt_rdata[55]
  PIN mgmt_rdata[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END mgmt_rdata[56]
  PIN mgmt_rdata[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END mgmt_rdata[57]
  PIN mgmt_rdata[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END mgmt_rdata[58]
  PIN mgmt_rdata[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END mgmt_rdata[59]
  PIN mgmt_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END mgmt_rdata[5]
  PIN mgmt_rdata[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END mgmt_rdata[60]
  PIN mgmt_rdata[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END mgmt_rdata[61]
  PIN mgmt_rdata[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END mgmt_rdata[62]
  PIN mgmt_rdata[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END mgmt_rdata[63]
  PIN mgmt_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END mgmt_rdata[6]
  PIN mgmt_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END mgmt_rdata[7]
  PIN mgmt_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END mgmt_rdata[8]
  PIN mgmt_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END mgmt_rdata[9]
  PIN mgmt_rdata_ro[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END mgmt_rdata_ro[0]
  PIN mgmt_rdata_ro[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END mgmt_rdata_ro[10]
  PIN mgmt_rdata_ro[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END mgmt_rdata_ro[11]
  PIN mgmt_rdata_ro[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END mgmt_rdata_ro[12]
  PIN mgmt_rdata_ro[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END mgmt_rdata_ro[13]
  PIN mgmt_rdata_ro[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END mgmt_rdata_ro[14]
  PIN mgmt_rdata_ro[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END mgmt_rdata_ro[15]
  PIN mgmt_rdata_ro[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END mgmt_rdata_ro[16]
  PIN mgmt_rdata_ro[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END mgmt_rdata_ro[17]
  PIN mgmt_rdata_ro[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END mgmt_rdata_ro[18]
  PIN mgmt_rdata_ro[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END mgmt_rdata_ro[19]
  PIN mgmt_rdata_ro[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END mgmt_rdata_ro[1]
  PIN mgmt_rdata_ro[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END mgmt_rdata_ro[20]
  PIN mgmt_rdata_ro[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END mgmt_rdata_ro[21]
  PIN mgmt_rdata_ro[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END mgmt_rdata_ro[22]
  PIN mgmt_rdata_ro[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END mgmt_rdata_ro[23]
  PIN mgmt_rdata_ro[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END mgmt_rdata_ro[24]
  PIN mgmt_rdata_ro[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END mgmt_rdata_ro[25]
  PIN mgmt_rdata_ro[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END mgmt_rdata_ro[26]
  PIN mgmt_rdata_ro[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END mgmt_rdata_ro[27]
  PIN mgmt_rdata_ro[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END mgmt_rdata_ro[28]
  PIN mgmt_rdata_ro[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END mgmt_rdata_ro[29]
  PIN mgmt_rdata_ro[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END mgmt_rdata_ro[2]
  PIN mgmt_rdata_ro[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END mgmt_rdata_ro[30]
  PIN mgmt_rdata_ro[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END mgmt_rdata_ro[31]
  PIN mgmt_rdata_ro[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END mgmt_rdata_ro[3]
  PIN mgmt_rdata_ro[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END mgmt_rdata_ro[4]
  PIN mgmt_rdata_ro[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END mgmt_rdata_ro[5]
  PIN mgmt_rdata_ro[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END mgmt_rdata_ro[6]
  PIN mgmt_rdata_ro[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END mgmt_rdata_ro[7]
  PIN mgmt_rdata_ro[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END mgmt_rdata_ro[8]
  PIN mgmt_rdata_ro[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END mgmt_rdata_ro[9]
  PIN mgmt_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END mgmt_wdata[0]
  PIN mgmt_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END mgmt_wdata[10]
  PIN mgmt_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END mgmt_wdata[11]
  PIN mgmt_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END mgmt_wdata[12]
  PIN mgmt_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END mgmt_wdata[13]
  PIN mgmt_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END mgmt_wdata[14]
  PIN mgmt_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END mgmt_wdata[15]
  PIN mgmt_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END mgmt_wdata[16]
  PIN mgmt_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END mgmt_wdata[17]
  PIN mgmt_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END mgmt_wdata[18]
  PIN mgmt_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END mgmt_wdata[19]
  PIN mgmt_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END mgmt_wdata[1]
  PIN mgmt_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END mgmt_wdata[20]
  PIN mgmt_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END mgmt_wdata[21]
  PIN mgmt_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END mgmt_wdata[22]
  PIN mgmt_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END mgmt_wdata[23]
  PIN mgmt_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END mgmt_wdata[24]
  PIN mgmt_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END mgmt_wdata[25]
  PIN mgmt_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END mgmt_wdata[26]
  PIN mgmt_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END mgmt_wdata[27]
  PIN mgmt_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END mgmt_wdata[28]
  PIN mgmt_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END mgmt_wdata[29]
  PIN mgmt_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END mgmt_wdata[2]
  PIN mgmt_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END mgmt_wdata[30]
  PIN mgmt_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END mgmt_wdata[31]
  PIN mgmt_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END mgmt_wdata[3]
  PIN mgmt_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END mgmt_wdata[4]
  PIN mgmt_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END mgmt_wdata[5]
  PIN mgmt_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END mgmt_wdata[6]
  PIN mgmt_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END mgmt_wdata[7]
  PIN mgmt_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END mgmt_wdata[8]
  PIN mgmt_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END mgmt_wdata[9]
  PIN mgmt_wen[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END mgmt_wen[0]
  PIN mgmt_wen[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END mgmt_wen[1]
  PIN mgmt_wen_mask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END mgmt_wen_mask[0]
  PIN mgmt_wen_mask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END mgmt_wen_mask[1]
  PIN mgmt_wen_mask[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END mgmt_wen_mask[2]
  PIN mgmt_wen_mask[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END mgmt_wen_mask[3]
  PIN mgmt_wen_mask[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END mgmt_wen_mask[4]
  PIN mgmt_wen_mask[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END mgmt_wen_mask[5]
  PIN mgmt_wen_mask[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END mgmt_wen_mask[6]
  PIN mgmt_wen_mask[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END mgmt_wen_mask[7]
  PIN mprj2_vcc_pwrgood
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 896.000 29.810 900.000 ;
    END
  END mprj2_vcc_pwrgood
  PIN mprj2_vdd_pwrgood
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 896.000 27.970 900.000 ;
    END
  END mprj2_vdd_pwrgood
  PIN mprj_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 878.600 4.000 879.200 ;
    END
  END mprj_ack_i
  PIN mprj_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 896.000 747.410 900.000 ;
    END
  END mprj_adr_o[0]
  PIN mprj_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 896.000 26.130 900.000 ;
    END
  END mprj_adr_o[10]
  PIN mprj_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.970 896.000 749.250 900.000 ;
    END
  END mprj_adr_o[11]
  PIN mprj_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 896.000 24.290 900.000 ;
    END
  END mprj_adr_o[12]
  PIN mprj_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 896.000 751.090 900.000 ;
    END
  END mprj_adr_o[13]
  PIN mprj_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 896.000 22.450 900.000 ;
    END
  END mprj_adr_o[14]
  PIN mprj_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 896.000 752.930 900.000 ;
    END
  END mprj_adr_o[15]
  PIN mprj_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 896.000 754.770 900.000 ;
    END
  END mprj_adr_o[16]
  PIN mprj_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.330 896.000 756.610 900.000 ;
    END
  END mprj_adr_o[17]
  PIN mprj_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 896.000 758.450 900.000 ;
    END
  END mprj_adr_o[18]
  PIN mprj_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 896.000 760.290 900.000 ;
    END
  END mprj_adr_o[19]
  PIN mprj_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.850 896.000 762.130 900.000 ;
    END
  END mprj_adr_o[1]
  PIN mprj_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 896.000 763.970 900.000 ;
    END
  END mprj_adr_o[20]
  PIN mprj_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.530 896.000 765.810 900.000 ;
    END
  END mprj_adr_o[21]
  PIN mprj_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 896.000 767.650 900.000 ;
    END
  END mprj_adr_o[22]
  PIN mprj_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.210 896.000 769.490 900.000 ;
    END
  END mprj_adr_o[23]
  PIN mprj_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.050 896.000 771.330 900.000 ;
    END
  END mprj_adr_o[24]
  PIN mprj_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 896.000 773.170 900.000 ;
    END
  END mprj_adr_o[25]
  PIN mprj_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.730 896.000 775.010 900.000 ;
    END
  END mprj_adr_o[26]
  PIN mprj_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 896.000 776.850 900.000 ;
    END
  END mprj_adr_o[27]
  PIN mprj_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.410 896.000 778.690 900.000 ;
    END
  END mprj_adr_o[28]
  PIN mprj_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.250 896.000 780.530 900.000 ;
    END
  END mprj_adr_o[29]
  PIN mprj_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 896.000 782.370 900.000 ;
    END
  END mprj_adr_o[2]
  PIN mprj_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.930 896.000 784.210 900.000 ;
    END
  END mprj_adr_o[30]
  PIN mprj_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 896.000 786.050 900.000 ;
    END
  END mprj_adr_o[31]
  PIN mprj_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.610 896.000 787.890 900.000 ;
    END
  END mprj_adr_o[3]
  PIN mprj_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 896.000 789.730 900.000 ;
    END
  END mprj_adr_o[4]
  PIN mprj_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.290 896.000 791.570 900.000 ;
    END
  END mprj_adr_o[5]
  PIN mprj_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 896.000 793.410 900.000 ;
    END
  END mprj_adr_o[6]
  PIN mprj_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.970 896.000 795.250 900.000 ;
    END
  END mprj_adr_o[7]
  PIN mprj_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.810 896.000 797.090 900.000 ;
    END
  END mprj_adr_o[8]
  PIN mprj_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 896.000 798.930 900.000 ;
    END
  END mprj_adr_o[9]
  PIN mprj_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 875.880 4.000 876.480 ;
    END
  END mprj_cyc_o
  PIN mprj_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.160 4.000 873.760 ;
    END
  END mprj_dat_i[0]
  PIN mprj_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END mprj_dat_i[10]
  PIN mprj_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.720 4.000 868.320 ;
    END
  END mprj_dat_i[11]
  PIN mprj_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 865.000 4.000 865.600 ;
    END
  END mprj_dat_i[12]
  PIN mprj_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 862.280 4.000 862.880 ;
    END
  END mprj_dat_i[13]
  PIN mprj_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 859.560 4.000 860.160 ;
    END
  END mprj_dat_i[14]
  PIN mprj_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END mprj_dat_i[15]
  PIN mprj_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 854.120 4.000 854.720 ;
    END
  END mprj_dat_i[16]
  PIN mprj_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 851.400 4.000 852.000 ;
    END
  END mprj_dat_i[17]
  PIN mprj_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 848.680 4.000 849.280 ;
    END
  END mprj_dat_i[18]
  PIN mprj_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 845.960 4.000 846.560 ;
    END
  END mprj_dat_i[19]
  PIN mprj_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END mprj_dat_i[1]
  PIN mprj_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 840.520 4.000 841.120 ;
    END
  END mprj_dat_i[20]
  PIN mprj_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 837.800 4.000 838.400 ;
    END
  END mprj_dat_i[21]
  PIN mprj_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 835.080 4.000 835.680 ;
    END
  END mprj_dat_i[22]
  PIN mprj_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 832.360 4.000 832.960 ;
    END
  END mprj_dat_i[23]
  PIN mprj_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END mprj_dat_i[24]
  PIN mprj_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.920 4.000 827.520 ;
    END
  END mprj_dat_i[25]
  PIN mprj_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 824.200 4.000 824.800 ;
    END
  END mprj_dat_i[26]
  PIN mprj_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 821.480 4.000 822.080 ;
    END
  END mprj_dat_i[27]
  PIN mprj_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 818.760 4.000 819.360 ;
    END
  END mprj_dat_i[28]
  PIN mprj_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 816.040 4.000 816.640 ;
    END
  END mprj_dat_i[29]
  PIN mprj_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 813.320 4.000 813.920 ;
    END
  END mprj_dat_i[2]
  PIN mprj_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 810.600 4.000 811.200 ;
    END
  END mprj_dat_i[30]
  PIN mprj_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.880 4.000 808.480 ;
    END
  END mprj_dat_i[31]
  PIN mprj_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.160 4.000 805.760 ;
    END
  END mprj_dat_i[3]
  PIN mprj_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.440 4.000 803.040 ;
    END
  END mprj_dat_i[4]
  PIN mprj_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.720 4.000 800.320 ;
    END
  END mprj_dat_i[5]
  PIN mprj_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.000 4.000 797.600 ;
    END
  END mprj_dat_i[6]
  PIN mprj_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 794.280 4.000 794.880 ;
    END
  END mprj_dat_i[7]
  PIN mprj_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 791.560 4.000 792.160 ;
    END
  END mprj_dat_i[8]
  PIN mprj_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END mprj_dat_i[9]
  PIN mprj_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.490 896.000 800.770 900.000 ;
    END
  END mprj_dat_o[0]
  PIN mprj_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.330 896.000 802.610 900.000 ;
    END
  END mprj_dat_o[10]
  PIN mprj_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.170 896.000 804.450 900.000 ;
    END
  END mprj_dat_o[11]
  PIN mprj_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.010 896.000 806.290 900.000 ;
    END
  END mprj_dat_o[12]
  PIN mprj_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.850 896.000 808.130 900.000 ;
    END
  END mprj_dat_o[13]
  PIN mprj_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.690 896.000 809.970 900.000 ;
    END
  END mprj_dat_o[14]
  PIN mprj_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 896.000 811.810 900.000 ;
    END
  END mprj_dat_o[15]
  PIN mprj_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.370 896.000 813.650 900.000 ;
    END
  END mprj_dat_o[16]
  PIN mprj_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 896.000 815.490 900.000 ;
    END
  END mprj_dat_o[17]
  PIN mprj_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.050 896.000 817.330 900.000 ;
    END
  END mprj_dat_o[18]
  PIN mprj_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.890 896.000 819.170 900.000 ;
    END
  END mprj_dat_o[19]
  PIN mprj_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.730 896.000 821.010 900.000 ;
    END
  END mprj_dat_o[1]
  PIN mprj_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.570 896.000 822.850 900.000 ;
    END
  END mprj_dat_o[20]
  PIN mprj_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 896.000 824.690 900.000 ;
    END
  END mprj_dat_o[21]
  PIN mprj_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.250 896.000 826.530 900.000 ;
    END
  END mprj_dat_o[22]
  PIN mprj_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 896.000 828.370 900.000 ;
    END
  END mprj_dat_o[23]
  PIN mprj_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.930 896.000 830.210 900.000 ;
    END
  END mprj_dat_o[24]
  PIN mprj_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.770 896.000 832.050 900.000 ;
    END
  END mprj_dat_o[25]
  PIN mprj_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.610 896.000 833.890 900.000 ;
    END
  END mprj_dat_o[26]
  PIN mprj_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.450 896.000 835.730 900.000 ;
    END
  END mprj_dat_o[27]
  PIN mprj_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 896.000 837.570 900.000 ;
    END
  END mprj_dat_o[28]
  PIN mprj_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.130 896.000 839.410 900.000 ;
    END
  END mprj_dat_o[29]
  PIN mprj_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.970 896.000 841.250 900.000 ;
    END
  END mprj_dat_o[2]
  PIN mprj_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.810 896.000 843.090 900.000 ;
    END
  END mprj_dat_o[30]
  PIN mprj_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.650 896.000 844.930 900.000 ;
    END
  END mprj_dat_o[31]
  PIN mprj_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.490 896.000 846.770 900.000 ;
    END
  END mprj_dat_o[3]
  PIN mprj_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.330 896.000 848.610 900.000 ;
    END
  END mprj_dat_o[4]
  PIN mprj_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 896.000 850.450 900.000 ;
    END
  END mprj_dat_o[5]
  PIN mprj_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.010 896.000 852.290 900.000 ;
    END
  END mprj_dat_o[6]
  PIN mprj_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.850 896.000 854.130 900.000 ;
    END
  END mprj_dat_o[7]
  PIN mprj_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 896.000 855.970 900.000 ;
    END
  END mprj_dat_o[8]
  PIN mprj_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.530 896.000 857.810 900.000 ;
    END
  END mprj_dat_o[9]
  PIN mprj_io_loader_clock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.770 896.000 1476.050 900.000 ;
    END
  END mprj_io_loader_clock
  PIN mprj_io_loader_data
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 331.880 2150.000 332.480 ;
    END
  END mprj_io_loader_data
  PIN mprj_io_loader_resetn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1499.690 896.000 1499.970 900.000 ;
    END
  END mprj_io_loader_resetn
  PIN mprj_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.370 896.000 859.650 900.000 ;
    END
  END mprj_sel_o[0]
  PIN mprj_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.210 896.000 861.490 900.000 ;
    END
  END mprj_sel_o[1]
  PIN mprj_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 896.000 863.330 900.000 ;
    END
  END mprj_sel_o[2]
  PIN mprj_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.890 896.000 865.170 900.000 ;
    END
  END mprj_sel_o[3]
  PIN mprj_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.730 896.000 867.010 900.000 ;
    END
  END mprj_stb_o
  PIN mprj_vcc_pwrgood
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.570 896.000 868.850 900.000 ;
    END
  END mprj_vcc_pwrgood
  PIN mprj_vdd_pwrgood
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.410 896.000 870.690 900.000 ;
    END
  END mprj_vdd_pwrgood
  PIN mprj_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 896.000 872.530 900.000 ;
    END
  END mprj_we_o
  PIN porb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 253.000 2150.000 253.600 ;
    END
  END porb
  PIN pwr_ctrl_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END pwr_ctrl_out[0]
  PIN pwr_ctrl_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END pwr_ctrl_out[1]
  PIN pwr_ctrl_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END pwr_ctrl_out[2]
  PIN pwr_ctrl_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END pwr_ctrl_out[3]
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END resetb
  PIN sdo_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 560.360 2150.000 560.960 ;
    END
  END sdo_out
  PIN sdo_outenb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 565.800 2150.000 566.400 ;
    END
  END sdo_outenb
  PIN user_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.090 896.000 874.370 900.000 ;
    END
  END user_clk
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2121.040 10.640 2122.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2071.040 10.640 2072.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2021.040 10.640 2022.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1971.040 10.640 1972.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1921.040 10.640 1922.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1871.040 220.840 1872.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1821.040 220.840 1822.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1771.040 220.840 1772.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1721.040 220.840 1722.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1671.040 10.640 1672.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1621.040 10.640 1622.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1571.040 10.640 1572.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1521.040 10.640 1522.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1471.040 10.640 1472.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1421.040 10.640 1422.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1371.040 10.640 1372.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1321.040 10.640 1322.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1271.040 10.640 1272.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1221.040 10.640 1222.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1171.040 10.640 1172.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1121.040 10.640 1122.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1071.040 10.640 1072.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1021.040 686.160 1022.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 971.040 686.160 972.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 921.040 686.160 922.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 871.040 686.160 872.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 821.040 686.160 822.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 771.040 686.160 772.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 721.040 686.160 722.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 671.040 686.160 672.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 621.040 686.160 622.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 571.040 686.160 572.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 521.040 686.160 522.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 471.040 686.160 472.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 421.040 686.160 422.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 371.040 686.160 372.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 321.040 686.160 322.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 271.040 10.640 272.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 221.040 10.640 222.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 121.040 10.640 122.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 71.040 10.640 72.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 886.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1021.040 10.640 1022.640 151.640 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 971.040 10.640 972.640 151.640 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 921.040 10.640 922.640 151.640 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 871.040 10.640 872.640 151.640 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 821.040 10.640 822.640 151.640 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 771.040 10.640 772.640 151.640 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 721.040 10.640 722.640 151.640 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 671.040 10.640 672.640 151.640 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 621.040 10.640 622.640 151.640 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 571.040 10.640 572.640 151.640 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 521.040 10.640 522.640 151.640 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 151.640 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 421.040 10.640 422.640 151.640 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 371.040 10.640 372.640 151.640 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 151.640 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 792.390 2144.060 793.990 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 639.210 2144.060 640.810 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 486.030 2144.060 487.630 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 332.850 2144.060 334.450 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 179.670 2144.060 181.270 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 2144.060 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2096.040 10.640 2097.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2046.040 10.640 2047.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1996.040 10.640 1997.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1946.040 10.640 1947.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1896.040 220.840 1897.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1846.040 220.840 1847.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1796.040 220.840 1797.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1746.040 220.840 1747.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1696.040 220.840 1697.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1646.040 10.640 1647.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1596.040 10.640 1597.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1546.040 10.640 1547.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1496.040 10.640 1497.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1446.040 10.640 1447.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1396.040 10.640 1397.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1346.040 10.640 1347.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1296.040 10.640 1297.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1246.040 10.640 1247.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1196.040 10.640 1197.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1146.040 10.640 1147.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1096.040 10.640 1097.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1046.040 686.160 1047.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 996.040 686.160 997.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 946.040 686.160 947.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 896.040 686.160 897.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 846.040 686.160 847.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 796.040 686.160 797.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 746.040 686.160 747.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 696.040 686.160 697.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 646.040 686.160 647.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 596.040 686.160 597.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 546.040 686.160 547.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 496.040 686.160 497.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 446.040 686.160 447.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 396.040 686.160 397.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 346.040 686.160 347.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 296.040 10.640 297.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 246.040 10.640 247.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 196.040 10.640 197.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 146.040 10.640 147.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.040 10.640 97.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 46.040 10.640 47.640 886.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1046.040 10.640 1047.640 151.640 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 996.040 10.640 997.640 151.640 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 946.040 10.640 947.640 151.640 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 896.040 10.640 897.640 151.640 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 846.040 10.640 847.640 151.640 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 796.040 10.640 797.640 151.640 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 746.040 10.640 747.640 151.640 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 696.040 10.640 697.640 151.640 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 646.040 10.640 647.640 151.640 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 596.040 10.640 597.640 151.640 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 546.040 10.640 547.640 151.640 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 496.040 10.640 497.640 151.640 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 446.040 10.640 447.640 151.640 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 396.040 10.640 397.640 151.640 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 346.040 10.640 347.640 151.640 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 868.980 2144.060 870.580 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 715.800 2144.060 717.400 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 562.620 2144.060 564.220 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 409.440 2144.060 411.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 256.260 2144.060 257.860 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 2144.060 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2144.060 896.155 ;
      LAYER met1 ;
        RECT 2.830 4.460 2145.830 898.580 ;
      LAYER met2 ;
        RECT 2.860 895.720 3.490 898.610 ;
        RECT 4.330 895.720 5.330 898.610 ;
        RECT 6.170 895.720 7.170 898.610 ;
        RECT 8.010 895.720 9.010 898.610 ;
        RECT 9.850 895.720 10.850 898.610 ;
        RECT 11.690 895.720 12.690 898.610 ;
        RECT 13.530 895.720 14.530 898.610 ;
        RECT 15.370 895.720 16.370 898.610 ;
        RECT 17.210 895.720 18.210 898.610 ;
        RECT 19.050 895.720 20.050 898.610 ;
        RECT 20.890 895.720 21.890 898.610 ;
        RECT 22.730 895.720 23.730 898.610 ;
        RECT 24.570 895.720 25.570 898.610 ;
        RECT 26.410 895.720 27.410 898.610 ;
        RECT 28.250 895.720 29.250 898.610 ;
        RECT 30.090 895.720 31.090 898.610 ;
        RECT 31.930 895.720 32.930 898.610 ;
        RECT 33.770 895.720 34.770 898.610 ;
        RECT 35.610 895.720 36.610 898.610 ;
        RECT 37.450 895.720 38.450 898.610 ;
        RECT 39.290 895.720 40.290 898.610 ;
        RECT 41.130 895.720 42.130 898.610 ;
        RECT 42.970 895.720 43.970 898.610 ;
        RECT 44.810 895.720 45.810 898.610 ;
        RECT 46.650 895.720 47.650 898.610 ;
        RECT 48.490 895.720 49.490 898.610 ;
        RECT 50.330 895.720 51.330 898.610 ;
        RECT 52.170 895.720 53.170 898.610 ;
        RECT 54.010 895.720 55.010 898.610 ;
        RECT 55.850 895.720 56.850 898.610 ;
        RECT 57.690 895.720 58.690 898.610 ;
        RECT 59.530 895.720 60.530 898.610 ;
        RECT 61.370 895.720 62.370 898.610 ;
        RECT 63.210 895.720 64.210 898.610 ;
        RECT 65.050 895.720 66.050 898.610 ;
        RECT 66.890 895.720 67.890 898.610 ;
        RECT 68.730 895.720 69.730 898.610 ;
        RECT 70.570 895.720 71.570 898.610 ;
        RECT 72.410 895.720 73.410 898.610 ;
        RECT 74.250 895.720 75.250 898.610 ;
        RECT 76.090 895.720 77.090 898.610 ;
        RECT 77.930 895.720 78.930 898.610 ;
        RECT 79.770 895.720 80.770 898.610 ;
        RECT 81.610 895.720 82.610 898.610 ;
        RECT 83.450 895.720 84.450 898.610 ;
        RECT 85.290 895.720 86.290 898.610 ;
        RECT 87.130 895.720 88.130 898.610 ;
        RECT 88.970 895.720 89.970 898.610 ;
        RECT 90.810 895.720 91.810 898.610 ;
        RECT 92.650 895.720 93.650 898.610 ;
        RECT 94.490 895.720 95.490 898.610 ;
        RECT 96.330 895.720 97.330 898.610 ;
        RECT 98.170 895.720 99.170 898.610 ;
        RECT 100.010 895.720 101.010 898.610 ;
        RECT 101.850 895.720 102.850 898.610 ;
        RECT 103.690 895.720 104.690 898.610 ;
        RECT 105.530 895.720 106.530 898.610 ;
        RECT 107.370 895.720 108.370 898.610 ;
        RECT 109.210 895.720 110.210 898.610 ;
        RECT 111.050 895.720 112.050 898.610 ;
        RECT 112.890 895.720 113.890 898.610 ;
        RECT 114.730 895.720 115.730 898.610 ;
        RECT 116.570 895.720 117.570 898.610 ;
        RECT 118.410 895.720 119.410 898.610 ;
        RECT 120.250 895.720 121.250 898.610 ;
        RECT 122.090 895.720 123.090 898.610 ;
        RECT 123.930 895.720 124.930 898.610 ;
        RECT 125.770 895.720 126.770 898.610 ;
        RECT 127.610 895.720 128.610 898.610 ;
        RECT 129.450 895.720 130.450 898.610 ;
        RECT 131.290 895.720 132.290 898.610 ;
        RECT 133.130 895.720 134.130 898.610 ;
        RECT 134.970 895.720 135.970 898.610 ;
        RECT 136.810 895.720 137.810 898.610 ;
        RECT 138.650 895.720 139.650 898.610 ;
        RECT 140.490 895.720 141.490 898.610 ;
        RECT 142.330 895.720 143.330 898.610 ;
        RECT 144.170 895.720 145.170 898.610 ;
        RECT 146.010 895.720 147.010 898.610 ;
        RECT 147.850 895.720 148.850 898.610 ;
        RECT 149.690 895.720 150.690 898.610 ;
        RECT 151.530 895.720 152.530 898.610 ;
        RECT 153.370 895.720 154.370 898.610 ;
        RECT 155.210 895.720 156.210 898.610 ;
        RECT 157.050 895.720 158.050 898.610 ;
        RECT 158.890 895.720 159.890 898.610 ;
        RECT 160.730 895.720 161.730 898.610 ;
        RECT 162.570 895.720 163.570 898.610 ;
        RECT 164.410 895.720 165.410 898.610 ;
        RECT 166.250 895.720 167.250 898.610 ;
        RECT 168.090 895.720 169.090 898.610 ;
        RECT 169.930 895.720 170.930 898.610 ;
        RECT 171.770 895.720 172.770 898.610 ;
        RECT 173.610 895.720 174.610 898.610 ;
        RECT 175.450 895.720 176.450 898.610 ;
        RECT 177.290 895.720 178.290 898.610 ;
        RECT 179.130 895.720 180.130 898.610 ;
        RECT 180.970 895.720 181.970 898.610 ;
        RECT 182.810 895.720 183.810 898.610 ;
        RECT 184.650 895.720 185.650 898.610 ;
        RECT 186.490 895.720 187.490 898.610 ;
        RECT 188.330 895.720 189.330 898.610 ;
        RECT 190.170 895.720 191.170 898.610 ;
        RECT 192.010 895.720 193.010 898.610 ;
        RECT 193.850 895.720 194.850 898.610 ;
        RECT 195.690 895.720 196.690 898.610 ;
        RECT 197.530 895.720 198.530 898.610 ;
        RECT 199.370 895.720 200.370 898.610 ;
        RECT 201.210 895.720 202.210 898.610 ;
        RECT 203.050 895.720 204.050 898.610 ;
        RECT 204.890 895.720 205.890 898.610 ;
        RECT 206.730 895.720 207.730 898.610 ;
        RECT 208.570 895.720 209.570 898.610 ;
        RECT 210.410 895.720 211.410 898.610 ;
        RECT 212.250 895.720 213.250 898.610 ;
        RECT 214.090 895.720 215.090 898.610 ;
        RECT 215.930 895.720 216.930 898.610 ;
        RECT 217.770 895.720 218.770 898.610 ;
        RECT 219.610 895.720 220.610 898.610 ;
        RECT 221.450 895.720 222.450 898.610 ;
        RECT 223.290 895.720 224.290 898.610 ;
        RECT 225.130 895.720 226.130 898.610 ;
        RECT 226.970 895.720 227.970 898.610 ;
        RECT 228.810 895.720 229.810 898.610 ;
        RECT 230.650 895.720 231.650 898.610 ;
        RECT 232.490 895.720 233.490 898.610 ;
        RECT 234.330 895.720 235.330 898.610 ;
        RECT 236.170 895.720 237.170 898.610 ;
        RECT 238.010 895.720 239.010 898.610 ;
        RECT 239.850 895.720 240.850 898.610 ;
        RECT 241.690 895.720 242.690 898.610 ;
        RECT 243.530 895.720 244.530 898.610 ;
        RECT 245.370 895.720 246.370 898.610 ;
        RECT 247.210 895.720 248.210 898.610 ;
        RECT 249.050 895.720 250.050 898.610 ;
        RECT 250.890 895.720 251.890 898.610 ;
        RECT 252.730 895.720 253.730 898.610 ;
        RECT 254.570 895.720 255.570 898.610 ;
        RECT 256.410 895.720 257.410 898.610 ;
        RECT 258.250 895.720 259.250 898.610 ;
        RECT 260.090 895.720 261.090 898.610 ;
        RECT 261.930 895.720 262.930 898.610 ;
        RECT 263.770 895.720 264.770 898.610 ;
        RECT 265.610 895.720 266.610 898.610 ;
        RECT 267.450 895.720 268.450 898.610 ;
        RECT 269.290 895.720 270.290 898.610 ;
        RECT 271.130 895.720 272.130 898.610 ;
        RECT 272.970 895.720 273.970 898.610 ;
        RECT 274.810 895.720 275.810 898.610 ;
        RECT 276.650 895.720 277.650 898.610 ;
        RECT 278.490 895.720 279.490 898.610 ;
        RECT 280.330 895.720 281.330 898.610 ;
        RECT 282.170 895.720 283.170 898.610 ;
        RECT 284.010 895.720 285.010 898.610 ;
        RECT 285.850 895.720 286.850 898.610 ;
        RECT 287.690 895.720 288.690 898.610 ;
        RECT 289.530 895.720 290.530 898.610 ;
        RECT 291.370 895.720 292.370 898.610 ;
        RECT 293.210 895.720 294.210 898.610 ;
        RECT 295.050 895.720 296.050 898.610 ;
        RECT 296.890 895.720 297.890 898.610 ;
        RECT 298.730 895.720 299.730 898.610 ;
        RECT 300.570 895.720 301.570 898.610 ;
        RECT 302.410 895.720 303.410 898.610 ;
        RECT 304.250 895.720 305.250 898.610 ;
        RECT 306.090 895.720 307.090 898.610 ;
        RECT 307.930 895.720 308.930 898.610 ;
        RECT 309.770 895.720 310.770 898.610 ;
        RECT 311.610 895.720 312.610 898.610 ;
        RECT 313.450 895.720 314.450 898.610 ;
        RECT 315.290 895.720 316.290 898.610 ;
        RECT 317.130 895.720 318.130 898.610 ;
        RECT 318.970 895.720 319.970 898.610 ;
        RECT 320.810 895.720 321.810 898.610 ;
        RECT 322.650 895.720 323.650 898.610 ;
        RECT 324.490 895.720 325.490 898.610 ;
        RECT 326.330 895.720 327.330 898.610 ;
        RECT 328.170 895.720 329.170 898.610 ;
        RECT 330.010 895.720 331.010 898.610 ;
        RECT 331.850 895.720 332.850 898.610 ;
        RECT 333.690 895.720 334.690 898.610 ;
        RECT 335.530 895.720 336.530 898.610 ;
        RECT 337.370 895.720 338.370 898.610 ;
        RECT 339.210 895.720 340.210 898.610 ;
        RECT 341.050 895.720 342.050 898.610 ;
        RECT 342.890 895.720 343.890 898.610 ;
        RECT 344.730 895.720 345.730 898.610 ;
        RECT 346.570 895.720 347.570 898.610 ;
        RECT 348.410 895.720 349.410 898.610 ;
        RECT 350.250 895.720 351.250 898.610 ;
        RECT 352.090 895.720 353.090 898.610 ;
        RECT 353.930 895.720 354.930 898.610 ;
        RECT 355.770 895.720 356.770 898.610 ;
        RECT 357.610 895.720 358.610 898.610 ;
        RECT 359.450 895.720 360.450 898.610 ;
        RECT 361.290 895.720 362.290 898.610 ;
        RECT 363.130 895.720 364.130 898.610 ;
        RECT 364.970 895.720 365.970 898.610 ;
        RECT 366.810 895.720 367.810 898.610 ;
        RECT 368.650 895.720 369.650 898.610 ;
        RECT 370.490 895.720 371.490 898.610 ;
        RECT 372.330 895.720 373.330 898.610 ;
        RECT 374.170 895.720 375.170 898.610 ;
        RECT 376.010 895.720 377.010 898.610 ;
        RECT 377.850 895.720 378.850 898.610 ;
        RECT 379.690 895.720 380.690 898.610 ;
        RECT 381.530 895.720 382.530 898.610 ;
        RECT 383.370 895.720 384.370 898.610 ;
        RECT 385.210 895.720 386.210 898.610 ;
        RECT 387.050 895.720 388.050 898.610 ;
        RECT 388.890 895.720 389.890 898.610 ;
        RECT 390.730 895.720 391.730 898.610 ;
        RECT 392.570 895.720 393.570 898.610 ;
        RECT 394.410 895.720 395.410 898.610 ;
        RECT 396.250 895.720 397.250 898.610 ;
        RECT 398.090 895.720 399.090 898.610 ;
        RECT 399.930 895.720 400.930 898.610 ;
        RECT 401.770 895.720 402.770 898.610 ;
        RECT 403.610 895.720 404.610 898.610 ;
        RECT 405.450 895.720 406.450 898.610 ;
        RECT 407.290 895.720 408.290 898.610 ;
        RECT 409.130 895.720 410.130 898.610 ;
        RECT 410.970 895.720 411.970 898.610 ;
        RECT 412.810 895.720 413.810 898.610 ;
        RECT 414.650 895.720 415.650 898.610 ;
        RECT 416.490 895.720 417.490 898.610 ;
        RECT 418.330 895.720 419.330 898.610 ;
        RECT 420.170 895.720 421.170 898.610 ;
        RECT 422.010 895.720 423.010 898.610 ;
        RECT 423.850 895.720 424.850 898.610 ;
        RECT 425.690 895.720 426.690 898.610 ;
        RECT 427.530 895.720 428.530 898.610 ;
        RECT 429.370 895.720 430.370 898.610 ;
        RECT 431.210 895.720 432.210 898.610 ;
        RECT 433.050 895.720 434.050 898.610 ;
        RECT 434.890 895.720 435.890 898.610 ;
        RECT 436.730 895.720 437.730 898.610 ;
        RECT 438.570 895.720 439.570 898.610 ;
        RECT 440.410 895.720 441.410 898.610 ;
        RECT 442.250 895.720 443.250 898.610 ;
        RECT 444.090 895.720 445.090 898.610 ;
        RECT 445.930 895.720 446.930 898.610 ;
        RECT 447.770 895.720 448.770 898.610 ;
        RECT 449.610 895.720 450.610 898.610 ;
        RECT 451.450 895.720 452.450 898.610 ;
        RECT 453.290 895.720 454.290 898.610 ;
        RECT 455.130 895.720 456.130 898.610 ;
        RECT 456.970 895.720 457.970 898.610 ;
        RECT 458.810 895.720 459.810 898.610 ;
        RECT 460.650 895.720 461.650 898.610 ;
        RECT 462.490 895.720 463.490 898.610 ;
        RECT 464.330 895.720 465.330 898.610 ;
        RECT 466.170 895.720 467.170 898.610 ;
        RECT 468.010 895.720 469.010 898.610 ;
        RECT 469.850 895.720 470.850 898.610 ;
        RECT 471.690 895.720 472.690 898.610 ;
        RECT 473.530 895.720 474.530 898.610 ;
        RECT 475.370 895.720 476.370 898.610 ;
        RECT 477.210 895.720 478.210 898.610 ;
        RECT 479.050 895.720 480.050 898.610 ;
        RECT 480.890 895.720 481.890 898.610 ;
        RECT 482.730 895.720 483.730 898.610 ;
        RECT 484.570 895.720 485.570 898.610 ;
        RECT 486.410 895.720 487.410 898.610 ;
        RECT 488.250 895.720 489.250 898.610 ;
        RECT 490.090 895.720 491.090 898.610 ;
        RECT 491.930 895.720 492.930 898.610 ;
        RECT 493.770 895.720 494.770 898.610 ;
        RECT 495.610 895.720 496.610 898.610 ;
        RECT 497.450 895.720 498.450 898.610 ;
        RECT 499.290 895.720 500.290 898.610 ;
        RECT 501.130 895.720 502.130 898.610 ;
        RECT 502.970 895.720 503.970 898.610 ;
        RECT 504.810 895.720 505.810 898.610 ;
        RECT 506.650 895.720 507.650 898.610 ;
        RECT 508.490 895.720 509.490 898.610 ;
        RECT 510.330 895.720 511.330 898.610 ;
        RECT 512.170 895.720 513.170 898.610 ;
        RECT 514.010 895.720 515.010 898.610 ;
        RECT 515.850 895.720 516.850 898.610 ;
        RECT 517.690 895.720 518.690 898.610 ;
        RECT 519.530 895.720 520.530 898.610 ;
        RECT 521.370 895.720 522.370 898.610 ;
        RECT 523.210 895.720 524.210 898.610 ;
        RECT 525.050 895.720 526.050 898.610 ;
        RECT 526.890 895.720 527.890 898.610 ;
        RECT 528.730 895.720 529.730 898.610 ;
        RECT 530.570 895.720 531.570 898.610 ;
        RECT 532.410 895.720 533.410 898.610 ;
        RECT 534.250 895.720 535.250 898.610 ;
        RECT 536.090 895.720 537.090 898.610 ;
        RECT 537.930 895.720 538.930 898.610 ;
        RECT 539.770 895.720 540.770 898.610 ;
        RECT 541.610 895.720 542.610 898.610 ;
        RECT 543.450 895.720 544.450 898.610 ;
        RECT 545.290 895.720 546.290 898.610 ;
        RECT 547.130 895.720 548.130 898.610 ;
        RECT 548.970 895.720 549.970 898.610 ;
        RECT 550.810 895.720 551.810 898.610 ;
        RECT 552.650 895.720 553.650 898.610 ;
        RECT 554.490 895.720 555.490 898.610 ;
        RECT 556.330 895.720 557.330 898.610 ;
        RECT 558.170 895.720 559.170 898.610 ;
        RECT 560.010 895.720 561.010 898.610 ;
        RECT 561.850 895.720 562.850 898.610 ;
        RECT 563.690 895.720 564.690 898.610 ;
        RECT 565.530 895.720 566.530 898.610 ;
        RECT 567.370 895.720 568.370 898.610 ;
        RECT 569.210 895.720 570.210 898.610 ;
        RECT 571.050 895.720 572.050 898.610 ;
        RECT 572.890 895.720 573.890 898.610 ;
        RECT 574.730 895.720 575.730 898.610 ;
        RECT 576.570 895.720 577.570 898.610 ;
        RECT 578.410 895.720 579.410 898.610 ;
        RECT 580.250 895.720 581.250 898.610 ;
        RECT 582.090 895.720 583.090 898.610 ;
        RECT 583.930 895.720 584.930 898.610 ;
        RECT 585.770 895.720 586.770 898.610 ;
        RECT 587.610 895.720 588.610 898.610 ;
        RECT 589.450 895.720 590.450 898.610 ;
        RECT 591.290 895.720 592.290 898.610 ;
        RECT 593.130 895.720 594.130 898.610 ;
        RECT 594.970 895.720 595.970 898.610 ;
        RECT 596.810 895.720 597.810 898.610 ;
        RECT 598.650 895.720 599.650 898.610 ;
        RECT 600.490 895.720 601.490 898.610 ;
        RECT 602.330 895.720 603.330 898.610 ;
        RECT 604.170 895.720 605.170 898.610 ;
        RECT 606.010 895.720 607.010 898.610 ;
        RECT 607.850 895.720 608.850 898.610 ;
        RECT 609.690 895.720 610.690 898.610 ;
        RECT 611.530 895.720 612.530 898.610 ;
        RECT 613.370 895.720 614.370 898.610 ;
        RECT 615.210 895.720 616.210 898.610 ;
        RECT 617.050 895.720 618.050 898.610 ;
        RECT 618.890 895.720 619.890 898.610 ;
        RECT 620.730 895.720 621.730 898.610 ;
        RECT 622.570 895.720 623.570 898.610 ;
        RECT 624.410 895.720 625.410 898.610 ;
        RECT 626.250 895.720 627.250 898.610 ;
        RECT 628.090 895.720 629.090 898.610 ;
        RECT 629.930 895.720 630.930 898.610 ;
        RECT 631.770 895.720 632.770 898.610 ;
        RECT 633.610 895.720 634.610 898.610 ;
        RECT 635.450 895.720 636.450 898.610 ;
        RECT 637.290 895.720 638.290 898.610 ;
        RECT 639.130 895.720 640.130 898.610 ;
        RECT 640.970 895.720 641.970 898.610 ;
        RECT 642.810 895.720 643.810 898.610 ;
        RECT 644.650 895.720 645.650 898.610 ;
        RECT 646.490 895.720 647.490 898.610 ;
        RECT 648.330 895.720 649.330 898.610 ;
        RECT 650.170 895.720 651.170 898.610 ;
        RECT 652.010 895.720 653.010 898.610 ;
        RECT 653.850 895.720 654.850 898.610 ;
        RECT 655.690 895.720 656.690 898.610 ;
        RECT 657.530 895.720 658.530 898.610 ;
        RECT 659.370 895.720 660.370 898.610 ;
        RECT 661.210 895.720 662.210 898.610 ;
        RECT 663.050 895.720 664.050 898.610 ;
        RECT 664.890 895.720 665.890 898.610 ;
        RECT 666.730 895.720 667.730 898.610 ;
        RECT 668.570 895.720 669.570 898.610 ;
        RECT 670.410 895.720 671.410 898.610 ;
        RECT 672.250 895.720 673.250 898.610 ;
        RECT 674.090 895.720 675.090 898.610 ;
        RECT 675.930 895.720 676.930 898.610 ;
        RECT 677.770 895.720 678.770 898.610 ;
        RECT 679.610 895.720 680.610 898.610 ;
        RECT 681.450 895.720 682.450 898.610 ;
        RECT 683.290 895.720 684.290 898.610 ;
        RECT 685.130 895.720 686.130 898.610 ;
        RECT 686.970 895.720 687.970 898.610 ;
        RECT 688.810 895.720 689.810 898.610 ;
        RECT 690.650 895.720 691.650 898.610 ;
        RECT 692.490 895.720 693.490 898.610 ;
        RECT 694.330 895.720 695.330 898.610 ;
        RECT 696.170 895.720 697.170 898.610 ;
        RECT 698.010 895.720 699.010 898.610 ;
        RECT 699.850 895.720 700.850 898.610 ;
        RECT 701.690 895.720 702.690 898.610 ;
        RECT 703.530 895.720 704.530 898.610 ;
        RECT 705.370 895.720 706.370 898.610 ;
        RECT 707.210 895.720 708.210 898.610 ;
        RECT 709.050 895.720 710.050 898.610 ;
        RECT 710.890 895.720 711.890 898.610 ;
        RECT 712.730 895.720 713.730 898.610 ;
        RECT 714.570 895.720 715.570 898.610 ;
        RECT 716.410 895.720 717.410 898.610 ;
        RECT 718.250 895.720 719.250 898.610 ;
        RECT 720.090 895.720 721.090 898.610 ;
        RECT 721.930 895.720 722.930 898.610 ;
        RECT 723.770 895.720 724.770 898.610 ;
        RECT 725.610 895.720 726.610 898.610 ;
        RECT 727.450 895.720 728.450 898.610 ;
        RECT 729.290 895.720 730.290 898.610 ;
        RECT 731.130 895.720 732.130 898.610 ;
        RECT 732.970 895.720 733.970 898.610 ;
        RECT 734.810 895.720 735.810 898.610 ;
        RECT 736.650 895.720 737.650 898.610 ;
        RECT 738.490 895.720 739.490 898.610 ;
        RECT 740.330 895.720 741.330 898.610 ;
        RECT 742.170 895.720 743.170 898.610 ;
        RECT 744.010 895.720 745.010 898.610 ;
        RECT 745.850 895.720 746.850 898.610 ;
        RECT 747.690 895.720 748.690 898.610 ;
        RECT 749.530 895.720 750.530 898.610 ;
        RECT 751.370 895.720 752.370 898.610 ;
        RECT 753.210 895.720 754.210 898.610 ;
        RECT 755.050 895.720 756.050 898.610 ;
        RECT 756.890 895.720 757.890 898.610 ;
        RECT 758.730 895.720 759.730 898.610 ;
        RECT 760.570 895.720 761.570 898.610 ;
        RECT 762.410 895.720 763.410 898.610 ;
        RECT 764.250 895.720 765.250 898.610 ;
        RECT 766.090 895.720 767.090 898.610 ;
        RECT 767.930 895.720 768.930 898.610 ;
        RECT 769.770 895.720 770.770 898.610 ;
        RECT 771.610 895.720 772.610 898.610 ;
        RECT 773.450 895.720 774.450 898.610 ;
        RECT 775.290 895.720 776.290 898.610 ;
        RECT 777.130 895.720 778.130 898.610 ;
        RECT 778.970 895.720 779.970 898.610 ;
        RECT 780.810 895.720 781.810 898.610 ;
        RECT 782.650 895.720 783.650 898.610 ;
        RECT 784.490 895.720 785.490 898.610 ;
        RECT 786.330 895.720 787.330 898.610 ;
        RECT 788.170 895.720 789.170 898.610 ;
        RECT 790.010 895.720 791.010 898.610 ;
        RECT 791.850 895.720 792.850 898.610 ;
        RECT 793.690 895.720 794.690 898.610 ;
        RECT 795.530 895.720 796.530 898.610 ;
        RECT 797.370 895.720 798.370 898.610 ;
        RECT 799.210 895.720 800.210 898.610 ;
        RECT 801.050 895.720 802.050 898.610 ;
        RECT 802.890 895.720 803.890 898.610 ;
        RECT 804.730 895.720 805.730 898.610 ;
        RECT 806.570 895.720 807.570 898.610 ;
        RECT 808.410 895.720 809.410 898.610 ;
        RECT 810.250 895.720 811.250 898.610 ;
        RECT 812.090 895.720 813.090 898.610 ;
        RECT 813.930 895.720 814.930 898.610 ;
        RECT 815.770 895.720 816.770 898.610 ;
        RECT 817.610 895.720 818.610 898.610 ;
        RECT 819.450 895.720 820.450 898.610 ;
        RECT 821.290 895.720 822.290 898.610 ;
        RECT 823.130 895.720 824.130 898.610 ;
        RECT 824.970 895.720 825.970 898.610 ;
        RECT 826.810 895.720 827.810 898.610 ;
        RECT 828.650 895.720 829.650 898.610 ;
        RECT 830.490 895.720 831.490 898.610 ;
        RECT 832.330 895.720 833.330 898.610 ;
        RECT 834.170 895.720 835.170 898.610 ;
        RECT 836.010 895.720 837.010 898.610 ;
        RECT 837.850 895.720 838.850 898.610 ;
        RECT 839.690 895.720 840.690 898.610 ;
        RECT 841.530 895.720 842.530 898.610 ;
        RECT 843.370 895.720 844.370 898.610 ;
        RECT 845.210 895.720 846.210 898.610 ;
        RECT 847.050 895.720 848.050 898.610 ;
        RECT 848.890 895.720 849.890 898.610 ;
        RECT 850.730 895.720 851.730 898.610 ;
        RECT 852.570 895.720 853.570 898.610 ;
        RECT 854.410 895.720 855.410 898.610 ;
        RECT 856.250 895.720 857.250 898.610 ;
        RECT 858.090 895.720 859.090 898.610 ;
        RECT 859.930 895.720 860.930 898.610 ;
        RECT 861.770 895.720 862.770 898.610 ;
        RECT 863.610 895.720 864.610 898.610 ;
        RECT 865.450 895.720 866.450 898.610 ;
        RECT 867.290 895.720 868.290 898.610 ;
        RECT 869.130 895.720 870.130 898.610 ;
        RECT 870.970 895.720 871.970 898.610 ;
        RECT 872.810 895.720 873.810 898.610 ;
        RECT 874.650 895.720 1050.450 898.610 ;
        RECT 1051.290 895.720 1435.010 898.610 ;
        RECT 1435.850 895.720 1475.490 898.610 ;
        RECT 1476.330 895.720 1499.410 898.610 ;
        RECT 1500.250 895.720 1692.610 898.610 ;
        RECT 1693.450 895.720 2134.210 898.610 ;
        RECT 2135.050 895.720 2136.050 898.610 ;
        RECT 2136.890 895.720 2137.890 898.610 ;
        RECT 2138.730 895.720 2139.730 898.610 ;
        RECT 2140.570 895.720 2141.570 898.610 ;
        RECT 2142.410 895.720 2143.410 898.610 ;
        RECT 2144.250 895.720 2145.250 898.610 ;
        RECT 2.860 4.280 2145.800 895.720 ;
        RECT 3.410 4.000 3.490 4.280 ;
        RECT 4.330 4.000 4.410 4.280 ;
        RECT 5.250 4.000 5.330 4.280 ;
        RECT 6.170 4.000 6.250 4.280 ;
        RECT 7.090 4.000 7.170 4.280 ;
        RECT 8.010 4.000 8.090 4.280 ;
        RECT 8.930 4.000 9.010 4.280 ;
        RECT 9.850 4.000 9.930 4.280 ;
        RECT 10.770 4.000 10.850 4.280 ;
        RECT 11.690 4.000 11.770 4.280 ;
        RECT 12.610 4.000 12.690 4.280 ;
        RECT 13.530 4.000 13.610 4.280 ;
        RECT 14.450 4.000 14.530 4.280 ;
        RECT 15.370 4.000 15.450 4.280 ;
        RECT 16.290 4.000 16.370 4.280 ;
        RECT 17.210 4.000 17.290 4.280 ;
        RECT 18.130 4.000 18.210 4.280 ;
        RECT 19.050 4.000 19.130 4.280 ;
        RECT 19.970 4.000 20.050 4.280 ;
        RECT 20.890 4.000 20.970 4.280 ;
        RECT 21.810 4.000 21.890 4.280 ;
        RECT 22.730 4.000 22.810 4.280 ;
        RECT 23.650 4.000 23.730 4.280 ;
        RECT 24.570 4.000 24.650 4.280 ;
        RECT 25.490 4.000 25.570 4.280 ;
        RECT 26.410 4.000 26.490 4.280 ;
        RECT 27.330 4.000 27.410 4.280 ;
        RECT 28.250 4.000 28.330 4.280 ;
        RECT 29.170 4.000 29.250 4.280 ;
        RECT 30.090 4.000 30.170 4.280 ;
        RECT 31.010 4.000 31.090 4.280 ;
        RECT 31.930 4.000 32.010 4.280 ;
        RECT 32.850 4.000 32.930 4.280 ;
        RECT 33.770 4.000 33.850 4.280 ;
        RECT 34.690 4.000 34.770 4.280 ;
        RECT 35.610 4.000 35.690 4.280 ;
        RECT 36.530 4.000 36.610 4.280 ;
        RECT 37.450 4.000 37.530 4.280 ;
        RECT 38.370 4.000 38.450 4.280 ;
        RECT 39.290 4.000 39.370 4.280 ;
        RECT 40.210 4.000 40.290 4.280 ;
        RECT 41.130 4.000 41.210 4.280 ;
        RECT 42.050 4.000 42.130 4.280 ;
        RECT 42.970 4.000 43.050 4.280 ;
        RECT 43.890 4.000 43.970 4.280 ;
        RECT 44.810 4.000 44.890 4.280 ;
        RECT 45.730 4.000 45.810 4.280 ;
        RECT 46.650 4.000 46.730 4.280 ;
        RECT 47.570 4.000 47.650 4.280 ;
        RECT 48.490 4.000 48.570 4.280 ;
        RECT 49.410 4.000 49.490 4.280 ;
        RECT 50.330 4.000 50.410 4.280 ;
        RECT 51.250 4.000 51.330 4.280 ;
        RECT 52.170 4.000 52.250 4.280 ;
        RECT 53.090 4.000 53.170 4.280 ;
        RECT 54.010 4.000 54.090 4.280 ;
        RECT 54.930 4.000 55.010 4.280 ;
        RECT 55.850 4.000 55.930 4.280 ;
        RECT 56.770 4.000 56.850 4.280 ;
        RECT 57.690 4.000 57.770 4.280 ;
        RECT 58.610 4.000 58.690 4.280 ;
        RECT 59.530 4.000 59.610 4.280 ;
        RECT 60.450 4.000 60.530 4.280 ;
        RECT 61.370 4.000 61.450 4.280 ;
        RECT 62.290 4.000 62.370 4.280 ;
        RECT 63.210 4.000 63.290 4.280 ;
        RECT 64.130 4.000 64.210 4.280 ;
        RECT 65.050 4.000 65.130 4.280 ;
        RECT 65.970 4.000 66.050 4.280 ;
        RECT 66.890 4.000 66.970 4.280 ;
        RECT 67.810 4.000 67.890 4.280 ;
        RECT 68.730 4.000 68.810 4.280 ;
        RECT 69.650 4.000 69.730 4.280 ;
        RECT 70.570 4.000 70.650 4.280 ;
        RECT 71.490 4.000 71.570 4.280 ;
        RECT 72.410 4.000 72.490 4.280 ;
        RECT 73.330 4.000 73.410 4.280 ;
        RECT 74.250 4.000 74.330 4.280 ;
        RECT 75.170 4.000 75.250 4.280 ;
        RECT 76.090 4.000 76.170 4.280 ;
        RECT 77.010 4.000 77.090 4.280 ;
        RECT 77.930 4.000 78.010 4.280 ;
        RECT 78.850 4.000 78.930 4.280 ;
        RECT 79.770 4.000 79.850 4.280 ;
        RECT 80.690 4.000 81.690 4.280 ;
        RECT 82.530 4.000 83.530 4.280 ;
        RECT 84.370 4.000 85.370 4.280 ;
        RECT 86.210 4.000 87.210 4.280 ;
        RECT 88.050 4.000 89.050 4.280 ;
        RECT 89.890 4.000 90.890 4.280 ;
        RECT 91.730 4.000 92.730 4.280 ;
        RECT 93.570 4.000 94.570 4.280 ;
        RECT 95.410 4.000 96.410 4.280 ;
        RECT 97.250 4.000 98.250 4.280 ;
        RECT 99.090 4.000 100.090 4.280 ;
        RECT 100.930 4.000 101.930 4.280 ;
        RECT 102.770 4.000 103.770 4.280 ;
        RECT 104.610 4.000 105.610 4.280 ;
        RECT 106.450 4.000 107.450 4.280 ;
        RECT 108.290 4.000 109.290 4.280 ;
        RECT 110.130 4.000 111.130 4.280 ;
        RECT 111.970 4.000 112.970 4.280 ;
        RECT 113.810 4.000 114.810 4.280 ;
        RECT 115.650 4.000 116.650 4.280 ;
        RECT 117.490 4.000 118.490 4.280 ;
        RECT 119.330 4.000 120.330 4.280 ;
        RECT 121.170 4.000 122.170 4.280 ;
        RECT 123.010 4.000 124.010 4.280 ;
        RECT 124.850 4.000 125.850 4.280 ;
        RECT 126.690 4.000 127.690 4.280 ;
        RECT 128.530 4.000 129.530 4.280 ;
        RECT 130.370 4.000 131.370 4.280 ;
        RECT 132.210 4.000 133.210 4.280 ;
        RECT 134.050 4.000 135.050 4.280 ;
        RECT 135.890 4.000 136.890 4.280 ;
        RECT 137.730 4.000 138.730 4.280 ;
        RECT 139.570 4.000 140.570 4.280 ;
        RECT 141.410 4.000 142.410 4.280 ;
        RECT 143.250 4.000 144.250 4.280 ;
        RECT 145.090 4.000 146.090 4.280 ;
        RECT 146.930 4.000 147.930 4.280 ;
        RECT 148.770 4.000 149.770 4.280 ;
        RECT 150.610 4.000 151.610 4.280 ;
        RECT 152.450 4.000 153.450 4.280 ;
        RECT 154.290 4.000 155.290 4.280 ;
        RECT 156.130 4.000 157.130 4.280 ;
        RECT 157.970 4.000 158.970 4.280 ;
        RECT 159.810 4.000 160.810 4.280 ;
        RECT 161.650 4.000 162.650 4.280 ;
        RECT 163.490 4.000 164.490 4.280 ;
        RECT 165.330 4.000 166.330 4.280 ;
        RECT 167.170 4.000 168.170 4.280 ;
        RECT 169.010 4.000 2145.800 4.280 ;
      LAYER met3 ;
        RECT 4.400 894.520 2145.600 895.385 ;
        RECT 3.990 893.200 2146.050 894.520 ;
        RECT 4.400 891.800 2145.600 893.200 ;
        RECT 3.990 890.480 2146.050 891.800 ;
        RECT 4.400 889.080 2145.600 890.480 ;
        RECT 3.990 887.760 2146.050 889.080 ;
        RECT 4.400 886.360 2145.600 887.760 ;
        RECT 3.990 885.040 2146.050 886.360 ;
        RECT 4.400 883.640 2145.600 885.040 ;
        RECT 3.990 882.320 2146.050 883.640 ;
        RECT 4.400 880.920 2146.050 882.320 ;
        RECT 3.990 879.600 2146.050 880.920 ;
        RECT 4.400 878.200 2146.050 879.600 ;
        RECT 3.990 876.880 2146.050 878.200 ;
        RECT 4.400 875.480 2146.050 876.880 ;
        RECT 3.990 874.160 2146.050 875.480 ;
        RECT 4.400 872.760 2146.050 874.160 ;
        RECT 3.990 871.440 2146.050 872.760 ;
        RECT 4.400 870.040 2146.050 871.440 ;
        RECT 3.990 868.720 2146.050 870.040 ;
        RECT 4.400 867.320 2146.050 868.720 ;
        RECT 3.990 866.000 2146.050 867.320 ;
        RECT 4.400 864.600 2146.050 866.000 ;
        RECT 3.990 863.280 2146.050 864.600 ;
        RECT 4.400 861.880 2146.050 863.280 ;
        RECT 3.990 860.560 2146.050 861.880 ;
        RECT 4.400 859.160 2146.050 860.560 ;
        RECT 3.990 857.840 2146.050 859.160 ;
        RECT 4.400 856.440 2146.050 857.840 ;
        RECT 3.990 855.120 2146.050 856.440 ;
        RECT 4.400 853.720 2146.050 855.120 ;
        RECT 3.990 852.400 2146.050 853.720 ;
        RECT 4.400 851.000 2146.050 852.400 ;
        RECT 3.990 849.680 2146.050 851.000 ;
        RECT 4.400 848.280 2146.050 849.680 ;
        RECT 3.990 846.960 2146.050 848.280 ;
        RECT 4.400 845.560 2146.050 846.960 ;
        RECT 3.990 844.240 2146.050 845.560 ;
        RECT 4.400 842.840 2146.050 844.240 ;
        RECT 3.990 841.520 2146.050 842.840 ;
        RECT 4.400 840.120 2146.050 841.520 ;
        RECT 3.990 838.800 2146.050 840.120 ;
        RECT 4.400 837.400 2146.050 838.800 ;
        RECT 3.990 836.080 2146.050 837.400 ;
        RECT 4.400 834.680 2146.050 836.080 ;
        RECT 3.990 833.360 2146.050 834.680 ;
        RECT 4.400 831.960 2146.050 833.360 ;
        RECT 3.990 830.640 2146.050 831.960 ;
        RECT 4.400 829.240 2146.050 830.640 ;
        RECT 3.990 827.920 2146.050 829.240 ;
        RECT 4.400 826.520 2146.050 827.920 ;
        RECT 3.990 825.200 2146.050 826.520 ;
        RECT 4.400 823.800 2146.050 825.200 ;
        RECT 3.990 822.480 2146.050 823.800 ;
        RECT 4.400 821.080 2146.050 822.480 ;
        RECT 3.990 819.760 2146.050 821.080 ;
        RECT 4.400 818.360 2146.050 819.760 ;
        RECT 3.990 817.040 2146.050 818.360 ;
        RECT 4.400 815.640 2146.050 817.040 ;
        RECT 3.990 814.320 2146.050 815.640 ;
        RECT 4.400 812.920 2146.050 814.320 ;
        RECT 3.990 811.600 2146.050 812.920 ;
        RECT 4.400 810.200 2146.050 811.600 ;
        RECT 3.990 808.880 2146.050 810.200 ;
        RECT 4.400 807.480 2146.050 808.880 ;
        RECT 3.990 806.160 2146.050 807.480 ;
        RECT 4.400 804.760 2146.050 806.160 ;
        RECT 3.990 803.440 2146.050 804.760 ;
        RECT 4.400 802.040 2146.050 803.440 ;
        RECT 3.990 800.720 2146.050 802.040 ;
        RECT 4.400 799.320 2146.050 800.720 ;
        RECT 3.990 798.000 2146.050 799.320 ;
        RECT 4.400 796.600 2146.050 798.000 ;
        RECT 3.990 795.280 2146.050 796.600 ;
        RECT 4.400 793.880 2146.050 795.280 ;
        RECT 3.990 792.560 2146.050 793.880 ;
        RECT 4.400 791.160 2146.050 792.560 ;
        RECT 3.990 789.840 2146.050 791.160 ;
        RECT 4.400 788.440 2146.050 789.840 ;
        RECT 3.990 787.120 2146.050 788.440 ;
        RECT 3.990 785.720 2145.600 787.120 ;
        RECT 3.990 746.320 2146.050 785.720 ;
        RECT 4.400 744.920 2146.050 746.320 ;
        RECT 3.990 566.800 2146.050 744.920 ;
        RECT 3.990 565.400 2145.600 566.800 ;
        RECT 3.990 564.080 2146.050 565.400 ;
        RECT 3.990 562.680 2145.600 564.080 ;
        RECT 3.990 561.360 2146.050 562.680 ;
        RECT 3.990 559.960 2145.600 561.360 ;
        RECT 3.990 341.040 2146.050 559.960 ;
        RECT 3.990 339.640 2145.600 341.040 ;
        RECT 3.990 338.320 2146.050 339.640 ;
        RECT 3.990 336.920 2145.600 338.320 ;
        RECT 3.990 335.600 2146.050 336.920 ;
        RECT 3.990 334.200 2145.600 335.600 ;
        RECT 3.990 332.880 2146.050 334.200 ;
        RECT 3.990 331.480 2145.600 332.880 ;
        RECT 3.990 254.000 2146.050 331.480 ;
        RECT 3.990 252.600 2145.600 254.000 ;
        RECT 3.990 243.120 2146.050 252.600 ;
        RECT 4.400 241.720 2146.050 243.120 ;
        RECT 3.990 240.400 2146.050 241.720 ;
        RECT 4.400 239.000 2146.050 240.400 ;
        RECT 3.990 237.680 2146.050 239.000 ;
        RECT 4.400 236.280 2146.050 237.680 ;
        RECT 3.990 234.960 2146.050 236.280 ;
        RECT 4.400 233.560 2146.050 234.960 ;
        RECT 3.990 232.240 2146.050 233.560 ;
        RECT 4.400 230.840 2146.050 232.240 ;
        RECT 3.990 229.520 2146.050 230.840 ;
        RECT 4.400 228.120 2146.050 229.520 ;
        RECT 3.990 226.800 2146.050 228.120 ;
        RECT 4.400 225.400 2146.050 226.800 ;
        RECT 3.990 224.080 2146.050 225.400 ;
        RECT 4.400 222.680 2146.050 224.080 ;
        RECT 3.990 221.360 2146.050 222.680 ;
        RECT 4.400 219.960 2146.050 221.360 ;
        RECT 3.990 218.640 2146.050 219.960 ;
        RECT 4.400 217.240 2146.050 218.640 ;
        RECT 3.990 215.920 2146.050 217.240 ;
        RECT 4.400 214.520 2146.050 215.920 ;
        RECT 3.990 213.200 2146.050 214.520 ;
        RECT 4.400 211.800 2146.050 213.200 ;
        RECT 3.990 210.480 2146.050 211.800 ;
        RECT 4.400 209.080 2146.050 210.480 ;
        RECT 3.990 207.760 2146.050 209.080 ;
        RECT 4.400 206.360 2146.050 207.760 ;
        RECT 3.990 205.040 2146.050 206.360 ;
        RECT 4.400 203.640 2146.050 205.040 ;
        RECT 3.990 202.320 2146.050 203.640 ;
        RECT 4.400 200.920 2146.050 202.320 ;
        RECT 3.990 199.600 2146.050 200.920 ;
        RECT 4.400 198.200 2146.050 199.600 ;
        RECT 3.990 196.880 2146.050 198.200 ;
        RECT 4.400 195.480 2146.050 196.880 ;
        RECT 3.990 194.160 2146.050 195.480 ;
        RECT 4.400 192.760 2146.050 194.160 ;
        RECT 3.990 191.440 2146.050 192.760 ;
        RECT 4.400 190.040 2146.050 191.440 ;
        RECT 3.990 188.720 2146.050 190.040 ;
        RECT 4.400 187.320 2146.050 188.720 ;
        RECT 3.990 186.000 2146.050 187.320 ;
        RECT 4.400 184.600 2146.050 186.000 ;
        RECT 3.990 183.280 2146.050 184.600 ;
        RECT 4.400 181.880 2146.050 183.280 ;
        RECT 3.990 180.560 2146.050 181.880 ;
        RECT 4.400 179.160 2146.050 180.560 ;
        RECT 3.990 177.840 2146.050 179.160 ;
        RECT 4.400 176.440 2145.600 177.840 ;
        RECT 3.990 175.120 2146.050 176.440 ;
        RECT 4.400 173.720 2145.600 175.120 ;
        RECT 3.990 172.400 2146.050 173.720 ;
        RECT 4.400 171.000 2145.600 172.400 ;
        RECT 3.990 169.680 2146.050 171.000 ;
        RECT 4.400 168.280 2145.600 169.680 ;
        RECT 3.990 166.960 2146.050 168.280 ;
        RECT 4.400 165.560 2145.600 166.960 ;
        RECT 3.990 164.240 2146.050 165.560 ;
        RECT 4.400 162.840 2145.600 164.240 ;
        RECT 3.990 161.520 2146.050 162.840 ;
        RECT 4.400 160.120 2145.600 161.520 ;
        RECT 3.990 158.800 2146.050 160.120 ;
        RECT 4.400 157.400 2145.600 158.800 ;
        RECT 3.990 156.080 2146.050 157.400 ;
        RECT 4.400 154.680 2145.600 156.080 ;
        RECT 3.990 153.360 2146.050 154.680 ;
        RECT 4.400 151.960 2145.600 153.360 ;
        RECT 3.990 150.640 2146.050 151.960 ;
        RECT 4.400 149.240 2145.600 150.640 ;
        RECT 3.990 147.920 2146.050 149.240 ;
        RECT 4.400 146.520 2145.600 147.920 ;
        RECT 3.990 145.200 2146.050 146.520 ;
        RECT 4.400 143.800 2145.600 145.200 ;
        RECT 3.990 142.480 2146.050 143.800 ;
        RECT 4.400 141.080 2145.600 142.480 ;
        RECT 3.990 139.760 2146.050 141.080 ;
        RECT 4.400 138.360 2145.600 139.760 ;
        RECT 3.990 137.040 2146.050 138.360 ;
        RECT 4.400 135.640 2145.600 137.040 ;
        RECT 3.990 134.320 2146.050 135.640 ;
        RECT 4.400 132.920 2145.600 134.320 ;
        RECT 3.990 131.600 2146.050 132.920 ;
        RECT 4.400 130.200 2145.600 131.600 ;
        RECT 3.990 128.880 2146.050 130.200 ;
        RECT 4.400 127.480 2145.600 128.880 ;
        RECT 3.990 126.160 2146.050 127.480 ;
        RECT 4.400 124.760 2145.600 126.160 ;
        RECT 3.990 123.440 2146.050 124.760 ;
        RECT 4.400 122.040 2145.600 123.440 ;
        RECT 3.990 120.720 2146.050 122.040 ;
        RECT 4.400 119.320 2145.600 120.720 ;
        RECT 3.990 118.000 2146.050 119.320 ;
        RECT 4.400 116.600 2145.600 118.000 ;
        RECT 3.990 115.280 2146.050 116.600 ;
        RECT 4.400 113.880 2145.600 115.280 ;
        RECT 3.990 112.560 2146.050 113.880 ;
        RECT 4.400 111.160 2145.600 112.560 ;
        RECT 3.990 109.840 2146.050 111.160 ;
        RECT 4.400 108.440 2145.600 109.840 ;
        RECT 3.990 107.120 2146.050 108.440 ;
        RECT 4.400 105.720 2145.600 107.120 ;
        RECT 3.990 104.400 2146.050 105.720 ;
        RECT 4.400 103.000 2145.600 104.400 ;
        RECT 3.990 101.680 2146.050 103.000 ;
        RECT 4.400 100.280 2145.600 101.680 ;
        RECT 3.990 98.960 2146.050 100.280 ;
        RECT 4.400 97.560 2145.600 98.960 ;
        RECT 3.990 96.240 2146.050 97.560 ;
        RECT 4.400 94.840 2145.600 96.240 ;
        RECT 3.990 93.520 2146.050 94.840 ;
        RECT 4.400 92.120 2145.600 93.520 ;
        RECT 3.990 90.800 2146.050 92.120 ;
        RECT 4.400 89.400 2146.050 90.800 ;
        RECT 3.990 88.080 2146.050 89.400 ;
        RECT 4.400 86.680 2146.050 88.080 ;
        RECT 3.990 85.360 2146.050 86.680 ;
        RECT 4.400 83.960 2146.050 85.360 ;
        RECT 3.990 82.640 2146.050 83.960 ;
        RECT 4.400 81.240 2146.050 82.640 ;
        RECT 3.990 79.920 2146.050 81.240 ;
        RECT 4.400 78.520 2146.050 79.920 ;
        RECT 3.990 77.200 2146.050 78.520 ;
        RECT 4.400 75.800 2146.050 77.200 ;
        RECT 3.990 74.480 2146.050 75.800 ;
        RECT 4.400 73.080 2146.050 74.480 ;
        RECT 3.990 71.760 2146.050 73.080 ;
        RECT 4.400 70.360 2146.050 71.760 ;
        RECT 3.990 69.040 2146.050 70.360 ;
        RECT 4.400 67.640 2146.050 69.040 ;
        RECT 3.990 66.320 2146.050 67.640 ;
        RECT 4.400 64.920 2146.050 66.320 ;
        RECT 3.990 63.600 2146.050 64.920 ;
        RECT 4.400 62.200 2146.050 63.600 ;
        RECT 3.990 60.880 2146.050 62.200 ;
        RECT 4.400 59.480 2146.050 60.880 ;
        RECT 3.990 58.160 2146.050 59.480 ;
        RECT 4.400 56.760 2146.050 58.160 ;
        RECT 3.990 55.440 2146.050 56.760 ;
        RECT 4.400 54.040 2146.050 55.440 ;
        RECT 3.990 52.720 2146.050 54.040 ;
        RECT 4.400 51.320 2146.050 52.720 ;
        RECT 3.990 50.000 2146.050 51.320 ;
        RECT 4.400 48.600 2146.050 50.000 ;
        RECT 3.990 47.280 2146.050 48.600 ;
        RECT 4.400 45.880 2146.050 47.280 ;
        RECT 3.990 44.560 2146.050 45.880 ;
        RECT 4.400 43.160 2146.050 44.560 ;
        RECT 3.990 41.840 2146.050 43.160 ;
        RECT 4.400 40.440 2146.050 41.840 ;
        RECT 3.990 39.120 2146.050 40.440 ;
        RECT 4.400 37.720 2146.050 39.120 ;
        RECT 3.990 36.400 2146.050 37.720 ;
        RECT 4.400 35.000 2146.050 36.400 ;
        RECT 3.990 33.680 2146.050 35.000 ;
        RECT 4.400 32.280 2146.050 33.680 ;
        RECT 3.990 30.960 2146.050 32.280 ;
        RECT 4.400 29.560 2146.050 30.960 ;
        RECT 3.990 28.240 2146.050 29.560 ;
        RECT 4.400 26.840 2146.050 28.240 ;
        RECT 3.990 25.520 2146.050 26.840 ;
        RECT 4.400 24.120 2146.050 25.520 ;
        RECT 3.990 22.800 2146.050 24.120 ;
        RECT 4.400 21.400 2146.050 22.800 ;
        RECT 3.990 20.080 2146.050 21.400 ;
        RECT 4.400 18.680 2146.050 20.080 ;
        RECT 3.990 17.360 2146.050 18.680 ;
        RECT 4.400 15.960 2146.050 17.360 ;
        RECT 3.990 14.640 2146.050 15.960 ;
        RECT 4.400 13.240 2146.050 14.640 ;
        RECT 3.990 11.920 2146.050 13.240 ;
        RECT 4.400 10.520 2146.050 11.920 ;
        RECT 3.990 9.200 2146.050 10.520 ;
        RECT 4.400 7.800 2146.050 9.200 ;
        RECT 3.990 6.480 2146.050 7.800 ;
        RECT 4.400 5.080 2146.050 6.480 ;
        RECT 3.990 4.255 2146.050 5.080 ;
      LAYER met4 ;
        RECT 15.935 887.360 2128.585 893.345 ;
        RECT 15.935 10.240 20.640 887.360 ;
        RECT 23.040 10.240 45.640 887.360 ;
        RECT 48.040 10.240 70.640 887.360 ;
        RECT 73.040 10.240 95.640 887.360 ;
        RECT 98.040 10.240 120.640 887.360 ;
        RECT 123.040 10.240 145.640 887.360 ;
        RECT 148.040 10.240 170.640 887.360 ;
        RECT 173.040 10.240 195.640 887.360 ;
        RECT 198.040 10.240 220.640 887.360 ;
        RECT 223.040 10.240 245.640 887.360 ;
        RECT 248.040 10.240 270.640 887.360 ;
        RECT 273.040 10.240 295.640 887.360 ;
        RECT 298.040 685.760 320.640 887.360 ;
        RECT 323.040 685.760 345.640 887.360 ;
        RECT 348.040 685.760 370.640 887.360 ;
        RECT 373.040 685.760 395.640 887.360 ;
        RECT 398.040 685.760 420.640 887.360 ;
        RECT 423.040 685.760 445.640 887.360 ;
        RECT 448.040 685.760 470.640 887.360 ;
        RECT 473.040 685.760 495.640 887.360 ;
        RECT 498.040 685.760 520.640 887.360 ;
        RECT 523.040 685.760 545.640 887.360 ;
        RECT 548.040 685.760 570.640 887.360 ;
        RECT 573.040 685.760 595.640 887.360 ;
        RECT 598.040 685.760 620.640 887.360 ;
        RECT 623.040 685.760 645.640 887.360 ;
        RECT 648.040 685.760 670.640 887.360 ;
        RECT 673.040 685.760 695.640 887.360 ;
        RECT 698.040 685.760 720.640 887.360 ;
        RECT 723.040 685.760 745.640 887.360 ;
        RECT 748.040 685.760 770.640 887.360 ;
        RECT 773.040 685.760 795.640 887.360 ;
        RECT 798.040 685.760 820.640 887.360 ;
        RECT 823.040 685.760 845.640 887.360 ;
        RECT 848.040 685.760 870.640 887.360 ;
        RECT 873.040 685.760 895.640 887.360 ;
        RECT 898.040 685.760 920.640 887.360 ;
        RECT 923.040 685.760 945.640 887.360 ;
        RECT 948.040 685.760 970.640 887.360 ;
        RECT 973.040 685.760 995.640 887.360 ;
        RECT 998.040 685.760 1020.640 887.360 ;
        RECT 1023.040 685.760 1045.640 887.360 ;
        RECT 1048.040 685.760 1070.640 887.360 ;
        RECT 298.040 152.040 1070.640 685.760 ;
        RECT 298.040 10.240 320.640 152.040 ;
        RECT 323.040 10.240 345.640 152.040 ;
        RECT 348.040 10.240 370.640 152.040 ;
        RECT 373.040 10.240 395.640 152.040 ;
        RECT 398.040 10.240 420.640 152.040 ;
        RECT 423.040 10.240 445.640 152.040 ;
        RECT 448.040 10.240 470.640 152.040 ;
        RECT 473.040 10.240 495.640 152.040 ;
        RECT 498.040 10.240 520.640 152.040 ;
        RECT 523.040 10.240 545.640 152.040 ;
        RECT 548.040 10.240 570.640 152.040 ;
        RECT 573.040 10.240 595.640 152.040 ;
        RECT 598.040 10.240 620.640 152.040 ;
        RECT 623.040 10.240 645.640 152.040 ;
        RECT 648.040 10.240 670.640 152.040 ;
        RECT 673.040 10.240 695.640 152.040 ;
        RECT 698.040 10.240 720.640 152.040 ;
        RECT 723.040 10.240 745.640 152.040 ;
        RECT 748.040 10.240 770.640 152.040 ;
        RECT 773.040 10.240 795.640 152.040 ;
        RECT 798.040 10.240 820.640 152.040 ;
        RECT 823.040 10.240 845.640 152.040 ;
        RECT 848.040 10.240 870.640 152.040 ;
        RECT 873.040 10.240 895.640 152.040 ;
        RECT 898.040 10.240 920.640 152.040 ;
        RECT 923.040 10.240 945.640 152.040 ;
        RECT 948.040 10.240 970.640 152.040 ;
        RECT 973.040 10.240 995.640 152.040 ;
        RECT 998.040 10.240 1020.640 152.040 ;
        RECT 1023.040 10.240 1045.640 152.040 ;
        RECT 1048.040 10.240 1070.640 152.040 ;
        RECT 1073.040 10.240 1095.640 887.360 ;
        RECT 1098.040 10.240 1120.640 887.360 ;
        RECT 1123.040 10.240 1145.640 887.360 ;
        RECT 1148.040 10.240 1170.640 887.360 ;
        RECT 1173.040 10.240 1195.640 887.360 ;
        RECT 1198.040 10.240 1220.640 887.360 ;
        RECT 1223.040 10.240 1245.640 887.360 ;
        RECT 1248.040 10.240 1270.640 887.360 ;
        RECT 1273.040 10.240 1295.640 887.360 ;
        RECT 1298.040 10.240 1320.640 887.360 ;
        RECT 1323.040 10.240 1345.640 887.360 ;
        RECT 1348.040 10.240 1370.640 887.360 ;
        RECT 1373.040 10.240 1395.640 887.360 ;
        RECT 1398.040 10.240 1420.640 887.360 ;
        RECT 1423.040 10.240 1445.640 887.360 ;
        RECT 1448.040 10.240 1470.640 887.360 ;
        RECT 1473.040 10.240 1495.640 887.360 ;
        RECT 1498.040 10.240 1520.640 887.360 ;
        RECT 1523.040 10.240 1545.640 887.360 ;
        RECT 1548.040 10.240 1570.640 887.360 ;
        RECT 1573.040 10.240 1595.640 887.360 ;
        RECT 1598.040 10.240 1620.640 887.360 ;
        RECT 1623.040 10.240 1645.640 887.360 ;
        RECT 1648.040 10.240 1670.640 887.360 ;
        RECT 1673.040 220.440 1695.640 887.360 ;
        RECT 1698.040 220.440 1720.640 887.360 ;
        RECT 1723.040 220.440 1745.640 887.360 ;
        RECT 1748.040 220.440 1770.640 887.360 ;
        RECT 1773.040 220.440 1795.640 887.360 ;
        RECT 1798.040 220.440 1820.640 887.360 ;
        RECT 1823.040 220.440 1845.640 887.360 ;
        RECT 1848.040 220.440 1870.640 887.360 ;
        RECT 1873.040 220.440 1895.640 887.360 ;
        RECT 1898.040 220.440 1920.640 887.360 ;
        RECT 1673.040 10.240 1920.640 220.440 ;
        RECT 1923.040 10.240 1945.640 887.360 ;
        RECT 1948.040 10.240 1970.640 887.360 ;
        RECT 1973.040 10.240 1995.640 887.360 ;
        RECT 1998.040 10.240 2020.640 887.360 ;
        RECT 2023.040 10.240 2045.640 887.360 ;
        RECT 2048.040 10.240 2070.640 887.360 ;
        RECT 2073.040 10.240 2095.640 887.360 ;
        RECT 2098.040 10.240 2120.640 887.360 ;
        RECT 2123.040 10.240 2128.585 887.360 ;
        RECT 15.935 4.255 2128.585 10.240 ;
      LAYER met5 ;
        RECT 303.260 872.180 1750.180 876.300 ;
        RECT 303.260 795.590 1750.180 867.380 ;
        RECT 303.260 719.000 1750.180 790.790 ;
        RECT 303.260 642.410 1750.180 714.200 ;
        RECT 303.260 565.820 1750.180 637.610 ;
        RECT 303.260 489.230 1750.180 561.020 ;
        RECT 303.260 412.640 1750.180 484.430 ;
        RECT 303.260 336.050 1750.180 407.840 ;
        RECT 303.260 259.460 1750.180 331.250 ;
        RECT 303.260 235.500 1750.180 254.660 ;
  END
END mgmt_core
END LIBRARY

