magic
tech sky130A
magscale 1 2
timestamp 1607567184
<< obsli1 >>
rect 1104 221 198812 10591
<< obsm1 >>
rect 198 8 199810 10600
<< metal2 >>
rect 202 10200 258 11400
rect 570 10200 626 11400
rect 1030 10200 1086 11400
rect 1490 10200 1546 11400
rect 1858 10200 1914 11400
rect 2318 10200 2374 11400
rect 2778 10200 2834 11400
rect 3238 10200 3294 11400
rect 3606 10200 3662 11400
rect 4066 10200 4122 11400
rect 4526 10200 4582 11400
rect 4986 10200 5042 11400
rect 5354 10200 5410 11400
rect 5814 10200 5870 11400
rect 6274 10200 6330 11400
rect 6734 10200 6790 11400
rect 7102 10200 7158 11400
rect 7562 10200 7618 11400
rect 8022 10200 8078 11400
rect 8390 10200 8446 11400
rect 8850 10200 8906 11400
rect 9310 10200 9366 11400
rect 9770 10200 9826 11400
rect 10138 10200 10194 11400
rect 10598 10200 10654 11400
rect 11058 10200 11114 11400
rect 11518 10200 11574 11400
rect 11886 10200 11942 11400
rect 12346 10200 12402 11400
rect 12806 10200 12862 11400
rect 13266 10200 13322 11400
rect 13634 10200 13690 11400
rect 14094 10200 14150 11400
rect 14554 10200 14610 11400
rect 15014 10200 15070 11400
rect 15382 10200 15438 11400
rect 15842 10200 15898 11400
rect 16302 10200 16358 11400
rect 16670 10200 16726 11400
rect 17130 10200 17186 11400
rect 17590 10200 17646 11400
rect 18050 10200 18106 11400
rect 18418 10200 18474 11400
rect 18878 10200 18934 11400
rect 19338 10200 19394 11400
rect 19798 10200 19854 11400
rect 20166 10200 20222 11400
rect 20626 10200 20682 11400
rect 21086 10200 21142 11400
rect 21546 10200 21602 11400
rect 21914 10200 21970 11400
rect 22374 10200 22430 11400
rect 22834 10200 22890 11400
rect 23294 10200 23350 11400
rect 23662 10200 23718 11400
rect 24122 10200 24178 11400
rect 24582 10200 24638 11400
rect 24950 10200 25006 11400
rect 25410 10200 25466 11400
rect 25870 10200 25926 11400
rect 26330 10200 26386 11400
rect 26698 10200 26754 11400
rect 27158 10200 27214 11400
rect 27618 10200 27674 11400
rect 28078 10200 28134 11400
rect 28446 10200 28502 11400
rect 28906 10200 28962 11400
rect 29366 10200 29422 11400
rect 29826 10200 29882 11400
rect 30194 10200 30250 11400
rect 30654 10200 30710 11400
rect 31114 10200 31170 11400
rect 31574 10200 31630 11400
rect 31942 10200 31998 11400
rect 32402 10200 32458 11400
rect 32862 10200 32918 11400
rect 33230 10200 33286 11400
rect 33690 10200 33746 11400
rect 34150 10200 34206 11400
rect 34610 10200 34666 11400
rect 34978 10200 35034 11400
rect 35438 10200 35494 11400
rect 35898 10200 35954 11400
rect 36358 10200 36414 11400
rect 36726 10200 36782 11400
rect 37186 10200 37242 11400
rect 37646 10200 37702 11400
rect 38106 10200 38162 11400
rect 38474 10200 38530 11400
rect 38934 10200 38990 11400
rect 39394 10200 39450 11400
rect 39854 10200 39910 11400
rect 40222 10200 40278 11400
rect 40682 10200 40738 11400
rect 41142 10200 41198 11400
rect 41510 10200 41566 11400
rect 41970 10200 42026 11400
rect 42430 10200 42486 11400
rect 42890 10200 42946 11400
rect 43258 10200 43314 11400
rect 43718 10200 43774 11400
rect 44178 10200 44234 11400
rect 44638 10200 44694 11400
rect 45006 10200 45062 11400
rect 45466 10200 45522 11400
rect 45926 10200 45982 11400
rect 46386 10200 46442 11400
rect 46754 10200 46810 11400
rect 47214 10200 47270 11400
rect 47674 10200 47730 11400
rect 48134 10200 48190 11400
rect 48502 10200 48558 11400
rect 48962 10200 49018 11400
rect 49422 10200 49478 11400
rect 49790 10200 49846 11400
rect 50250 10200 50306 11400
rect 50710 10200 50766 11400
rect 51170 10200 51226 11400
rect 51538 10200 51594 11400
rect 51998 10200 52054 11400
rect 52458 10200 52514 11400
rect 52918 10200 52974 11400
rect 53286 10200 53342 11400
rect 53746 10200 53802 11400
rect 54206 10200 54262 11400
rect 54666 10200 54722 11400
rect 55034 10200 55090 11400
rect 55494 10200 55550 11400
rect 55954 10200 56010 11400
rect 56322 10200 56378 11400
rect 56782 10200 56838 11400
rect 57242 10200 57298 11400
rect 57702 10200 57758 11400
rect 58070 10200 58126 11400
rect 58530 10200 58586 11400
rect 58990 10200 59046 11400
rect 59450 10200 59506 11400
rect 59818 10200 59874 11400
rect 60278 10200 60334 11400
rect 60738 10200 60794 11400
rect 61198 10200 61254 11400
rect 61566 10200 61622 11400
rect 62026 10200 62082 11400
rect 62486 10200 62542 11400
rect 62946 10200 63002 11400
rect 63314 10200 63370 11400
rect 63774 10200 63830 11400
rect 64234 10200 64290 11400
rect 64602 10200 64658 11400
rect 65062 10200 65118 11400
rect 65522 10200 65578 11400
rect 65982 10200 66038 11400
rect 66350 10200 66406 11400
rect 66810 10200 66866 11400
rect 67270 10200 67326 11400
rect 67730 10200 67786 11400
rect 68098 10200 68154 11400
rect 68558 10200 68614 11400
rect 69018 10200 69074 11400
rect 69478 10200 69534 11400
rect 69846 10200 69902 11400
rect 70306 10200 70362 11400
rect 70766 10200 70822 11400
rect 71226 10200 71282 11400
rect 71594 10200 71650 11400
rect 72054 10200 72110 11400
rect 72514 10200 72570 11400
rect 72882 10200 72938 11400
rect 73342 10200 73398 11400
rect 73802 10200 73858 11400
rect 74262 10200 74318 11400
rect 74630 10200 74686 11400
rect 75090 10200 75146 11400
rect 75550 10200 75606 11400
rect 76010 10200 76066 11400
rect 76378 10200 76434 11400
rect 76838 10200 76894 11400
rect 77298 10200 77354 11400
rect 77758 10200 77814 11400
rect 78126 10200 78182 11400
rect 78586 10200 78642 11400
rect 79046 10200 79102 11400
rect 79506 10200 79562 11400
rect 79874 10200 79930 11400
rect 80334 10200 80390 11400
rect 80794 10200 80850 11400
rect 81162 10200 81218 11400
rect 81622 10200 81678 11400
rect 82082 10200 82138 11400
rect 82542 10200 82598 11400
rect 82910 10200 82966 11400
rect 83370 10200 83426 11400
rect 83830 10200 83886 11400
rect 84290 10200 84346 11400
rect 84658 10200 84714 11400
rect 85118 10200 85174 11400
rect 85578 10200 85634 11400
rect 86038 10200 86094 11400
rect 86406 10200 86462 11400
rect 86866 10200 86922 11400
rect 87326 10200 87382 11400
rect 87786 10200 87842 11400
rect 88154 10200 88210 11400
rect 88614 10200 88670 11400
rect 89074 10200 89130 11400
rect 89442 10200 89498 11400
rect 89902 10200 89958 11400
rect 90362 10200 90418 11400
rect 90822 10200 90878 11400
rect 91190 10200 91246 11400
rect 91650 10200 91706 11400
rect 92110 10200 92166 11400
rect 92570 10200 92626 11400
rect 92938 10200 92994 11400
rect 93398 10200 93454 11400
rect 93858 10200 93914 11400
rect 94318 10200 94374 11400
rect 94686 10200 94742 11400
rect 95146 10200 95202 11400
rect 95606 10200 95662 11400
rect 96066 10200 96122 11400
rect 96434 10200 96490 11400
rect 96894 10200 96950 11400
rect 97354 10200 97410 11400
rect 97722 10200 97778 11400
rect 98182 10200 98238 11400
rect 98642 10200 98698 11400
rect 99102 10200 99158 11400
rect 99470 10200 99526 11400
rect 99930 10200 99986 11400
rect 100390 10200 100446 11400
rect 100850 10200 100906 11400
rect 101218 10200 101274 11400
rect 101678 10200 101734 11400
rect 102138 10200 102194 11400
rect 102598 10200 102654 11400
rect 102966 10200 103022 11400
rect 103426 10200 103482 11400
rect 103886 10200 103942 11400
rect 104254 10200 104310 11400
rect 104714 10200 104770 11400
rect 105174 10200 105230 11400
rect 105634 10200 105690 11400
rect 106002 10200 106058 11400
rect 106462 10200 106518 11400
rect 106922 10200 106978 11400
rect 107382 10200 107438 11400
rect 107750 10200 107806 11400
rect 108210 10200 108266 11400
rect 108670 10200 108726 11400
rect 109130 10200 109186 11400
rect 109498 10200 109554 11400
rect 109958 10200 110014 11400
rect 110418 10200 110474 11400
rect 110878 10200 110934 11400
rect 111246 10200 111302 11400
rect 111706 10200 111762 11400
rect 112166 10200 112222 11400
rect 112534 10200 112590 11400
rect 112994 10200 113050 11400
rect 113454 10200 113510 11400
rect 113914 10200 113970 11400
rect 114282 10200 114338 11400
rect 114742 10200 114798 11400
rect 115202 10200 115258 11400
rect 115662 10200 115718 11400
rect 116030 10200 116086 11400
rect 116490 10200 116546 11400
rect 116950 10200 117006 11400
rect 117410 10200 117466 11400
rect 117778 10200 117834 11400
rect 118238 10200 118294 11400
rect 118698 10200 118754 11400
rect 119158 10200 119214 11400
rect 119526 10200 119582 11400
rect 119986 10200 120042 11400
rect 120446 10200 120502 11400
rect 120814 10200 120870 11400
rect 121274 10200 121330 11400
rect 121734 10200 121790 11400
rect 122194 10200 122250 11400
rect 122562 10200 122618 11400
rect 123022 10200 123078 11400
rect 123482 10200 123538 11400
rect 123942 10200 123998 11400
rect 124310 10200 124366 11400
rect 124770 10200 124826 11400
rect 125230 10200 125286 11400
rect 125690 10200 125746 11400
rect 126058 10200 126114 11400
rect 126518 10200 126574 11400
rect 126978 10200 127034 11400
rect 127438 10200 127494 11400
rect 127806 10200 127862 11400
rect 128266 10200 128322 11400
rect 128726 10200 128782 11400
rect 129094 10200 129150 11400
rect 129554 10200 129610 11400
rect 130014 10200 130070 11400
rect 130474 10200 130530 11400
rect 130842 10200 130898 11400
rect 131302 10200 131358 11400
rect 131762 10200 131818 11400
rect 132222 10200 132278 11400
rect 132590 10200 132646 11400
rect 133050 10200 133106 11400
rect 133510 10200 133566 11400
rect 133970 10200 134026 11400
rect 134338 10200 134394 11400
rect 134798 10200 134854 11400
rect 135258 10200 135314 11400
rect 135718 10200 135774 11400
rect 136086 10200 136142 11400
rect 136546 10200 136602 11400
rect 137006 10200 137062 11400
rect 137374 10200 137430 11400
rect 137834 10200 137890 11400
rect 138294 10200 138350 11400
rect 138754 10200 138810 11400
rect 139122 10200 139178 11400
rect 139582 10200 139638 11400
rect 140042 10200 140098 11400
rect 140502 10200 140558 11400
rect 140870 10200 140926 11400
rect 141330 10200 141386 11400
rect 141790 10200 141846 11400
rect 142250 10200 142306 11400
rect 142618 10200 142674 11400
rect 143078 10200 143134 11400
rect 143538 10200 143594 11400
rect 143998 10200 144054 11400
rect 144366 10200 144422 11400
rect 144826 10200 144882 11400
rect 145286 10200 145342 11400
rect 145654 10200 145710 11400
rect 146114 10200 146170 11400
rect 146574 10200 146630 11400
rect 147034 10200 147090 11400
rect 147402 10200 147458 11400
rect 147862 10200 147918 11400
rect 148322 10200 148378 11400
rect 148782 10200 148838 11400
rect 149150 10200 149206 11400
rect 149610 10200 149666 11400
rect 150070 10200 150126 11400
rect 150530 10200 150586 11400
rect 150898 10200 150954 11400
rect 151358 10200 151414 11400
rect 151818 10200 151874 11400
rect 152186 10200 152242 11400
rect 152646 10200 152702 11400
rect 153106 10200 153162 11400
rect 153566 10200 153622 11400
rect 153934 10200 153990 11400
rect 154394 10200 154450 11400
rect 154854 10200 154910 11400
rect 155314 10200 155370 11400
rect 155682 10200 155738 11400
rect 156142 10200 156198 11400
rect 156602 10200 156658 11400
rect 157062 10200 157118 11400
rect 157430 10200 157486 11400
rect 157890 10200 157946 11400
rect 158350 10200 158406 11400
rect 158810 10200 158866 11400
rect 159178 10200 159234 11400
rect 159638 10200 159694 11400
rect 160098 10200 160154 11400
rect 160466 10200 160522 11400
rect 160926 10200 160982 11400
rect 161386 10200 161442 11400
rect 161846 10200 161902 11400
rect 162214 10200 162270 11400
rect 162674 10200 162730 11400
rect 163134 10200 163190 11400
rect 163594 10200 163650 11400
rect 163962 10200 164018 11400
rect 164422 10200 164478 11400
rect 164882 10200 164938 11400
rect 165342 10200 165398 11400
rect 165710 10200 165766 11400
rect 166170 10200 166226 11400
rect 166630 10200 166686 11400
rect 167090 10200 167146 11400
rect 167458 10200 167514 11400
rect 167918 10200 167974 11400
rect 168378 10200 168434 11400
rect 168746 10200 168802 11400
rect 169206 10200 169262 11400
rect 169666 10200 169722 11400
rect 170126 10200 170182 11400
rect 170494 10200 170550 11400
rect 170954 10200 171010 11400
rect 171414 10200 171470 11400
rect 171874 10200 171930 11400
rect 172242 10200 172298 11400
rect 172702 10200 172758 11400
rect 173162 10200 173218 11400
rect 173622 10200 173678 11400
rect 173990 10200 174046 11400
rect 174450 10200 174506 11400
rect 174910 10200 174966 11400
rect 175370 10200 175426 11400
rect 175738 10200 175794 11400
rect 176198 10200 176254 11400
rect 176658 10200 176714 11400
rect 177026 10200 177082 11400
rect 177486 10200 177542 11400
rect 177946 10200 178002 11400
rect 178406 10200 178462 11400
rect 178774 10200 178830 11400
rect 179234 10200 179290 11400
rect 179694 10200 179750 11400
rect 180154 10200 180210 11400
rect 180522 10200 180578 11400
rect 180982 10200 181038 11400
rect 181442 10200 181498 11400
rect 181902 10200 181958 11400
rect 182270 10200 182326 11400
rect 182730 10200 182786 11400
rect 183190 10200 183246 11400
rect 183650 10200 183706 11400
rect 184018 10200 184074 11400
rect 184478 10200 184534 11400
rect 184938 10200 184994 11400
rect 185306 10200 185362 11400
rect 185766 10200 185822 11400
rect 186226 10200 186282 11400
rect 186686 10200 186742 11400
rect 187054 10200 187110 11400
rect 187514 10200 187570 11400
rect 187974 10200 188030 11400
rect 188434 10200 188490 11400
rect 188802 10200 188858 11400
rect 189262 10200 189318 11400
rect 189722 10200 189778 11400
rect 190182 10200 190238 11400
rect 190550 10200 190606 11400
rect 191010 10200 191066 11400
rect 191470 10200 191526 11400
rect 191930 10200 191986 11400
rect 192298 10200 192354 11400
rect 192758 10200 192814 11400
rect 193218 10200 193274 11400
rect 193586 10200 193642 11400
rect 194046 10200 194102 11400
rect 194506 10200 194562 11400
rect 194966 10200 195022 11400
rect 195334 10200 195390 11400
rect 195794 10200 195850 11400
rect 196254 10200 196310 11400
rect 196714 10200 196770 11400
rect 197082 10200 197138 11400
rect 197542 10200 197598 11400
rect 198002 10200 198058 11400
rect 198462 10200 198518 11400
rect 198830 10200 198886 11400
rect 199290 10200 199346 11400
rect 199750 10200 199806 11400
rect 202 -400 258 800
rect 570 -400 626 800
rect 1030 -400 1086 800
rect 1490 -400 1546 800
rect 1858 -400 1914 800
rect 2318 -400 2374 800
rect 2778 -400 2834 800
rect 3238 -400 3294 800
rect 3606 -400 3662 800
rect 4066 -400 4122 800
rect 4526 -400 4582 800
rect 4986 -400 5042 800
rect 5354 -400 5410 800
rect 5814 -400 5870 800
rect 6274 -400 6330 800
rect 6734 -400 6790 800
rect 7102 -400 7158 800
rect 7562 -400 7618 800
rect 8022 -400 8078 800
rect 8390 -400 8446 800
rect 8850 -400 8906 800
rect 9310 -400 9366 800
rect 9770 -400 9826 800
rect 10138 -400 10194 800
rect 10598 -400 10654 800
rect 11058 -400 11114 800
rect 11518 -400 11574 800
rect 11886 -400 11942 800
rect 12346 -400 12402 800
rect 12806 -400 12862 800
rect 13266 -400 13322 800
rect 13634 -400 13690 800
rect 14094 -400 14150 800
rect 14554 -400 14610 800
rect 15014 -400 15070 800
rect 15382 -400 15438 800
rect 15842 -400 15898 800
rect 16302 -400 16358 800
rect 16670 -400 16726 800
rect 17130 -400 17186 800
rect 17590 -400 17646 800
rect 18050 -400 18106 800
rect 18418 -400 18474 800
rect 18878 -400 18934 800
rect 19338 -400 19394 800
rect 19798 -400 19854 800
rect 20166 -400 20222 800
rect 20626 -400 20682 800
rect 21086 -400 21142 800
rect 21546 -400 21602 800
rect 21914 -400 21970 800
rect 22374 -400 22430 800
rect 22834 -400 22890 800
rect 23294 -400 23350 800
rect 23662 -400 23718 800
rect 24122 -400 24178 800
rect 24582 -400 24638 800
rect 24950 -400 25006 800
rect 25410 -400 25466 800
rect 25870 -400 25926 800
rect 26330 -400 26386 800
rect 26698 -400 26754 800
rect 27158 -400 27214 800
rect 27618 -400 27674 800
rect 28078 -400 28134 800
rect 28446 -400 28502 800
rect 28906 -400 28962 800
rect 29366 -400 29422 800
rect 29826 -400 29882 800
rect 30194 -400 30250 800
rect 30654 -400 30710 800
rect 31114 -400 31170 800
rect 31574 -400 31630 800
rect 31942 -400 31998 800
rect 32402 -400 32458 800
rect 32862 -400 32918 800
rect 33230 -400 33286 800
rect 33690 -400 33746 800
rect 34150 -400 34206 800
rect 34610 -400 34666 800
rect 34978 -400 35034 800
rect 35438 -400 35494 800
rect 35898 -400 35954 800
rect 36358 -400 36414 800
rect 36726 -400 36782 800
rect 37186 -400 37242 800
rect 37646 -400 37702 800
rect 38106 -400 38162 800
rect 38474 -400 38530 800
rect 38934 -400 38990 800
rect 39394 -400 39450 800
rect 39854 -400 39910 800
rect 40222 -400 40278 800
rect 40682 -400 40738 800
rect 41142 -400 41198 800
rect 41510 -400 41566 800
rect 41970 -400 42026 800
rect 42430 -400 42486 800
rect 42890 -400 42946 800
rect 43258 -400 43314 800
rect 43718 -400 43774 800
rect 44178 -400 44234 800
rect 44638 -400 44694 800
rect 45006 -400 45062 800
rect 45466 -400 45522 800
rect 45926 -400 45982 800
rect 46386 -400 46442 800
rect 46754 -400 46810 800
rect 47214 -400 47270 800
rect 47674 -400 47730 800
rect 48134 -400 48190 800
rect 48502 -400 48558 800
rect 48962 -400 49018 800
rect 49422 -400 49478 800
rect 49790 -400 49846 800
rect 50250 -400 50306 800
rect 50710 -400 50766 800
rect 51170 -400 51226 800
rect 51538 -400 51594 800
rect 51998 -400 52054 800
rect 52458 -400 52514 800
rect 52918 -400 52974 800
rect 53286 -400 53342 800
rect 53746 -400 53802 800
rect 54206 -400 54262 800
rect 54666 -400 54722 800
rect 55034 -400 55090 800
rect 55494 -400 55550 800
rect 55954 -400 56010 800
rect 56322 -400 56378 800
rect 56782 -400 56838 800
rect 57242 -400 57298 800
rect 57702 -400 57758 800
rect 58070 -400 58126 800
rect 58530 -400 58586 800
rect 58990 -400 59046 800
rect 59450 -400 59506 800
rect 59818 -400 59874 800
rect 60278 -400 60334 800
rect 60738 -400 60794 800
rect 61198 -400 61254 800
rect 61566 -400 61622 800
rect 62026 -400 62082 800
rect 62486 -400 62542 800
rect 62946 -400 63002 800
rect 63314 -400 63370 800
rect 63774 -400 63830 800
rect 64234 -400 64290 800
rect 64602 -400 64658 800
rect 65062 -400 65118 800
rect 65522 -400 65578 800
rect 65982 -400 66038 800
rect 66350 -400 66406 800
rect 66810 -400 66866 800
rect 67270 -400 67326 800
rect 67730 -400 67786 800
rect 68098 -400 68154 800
rect 68558 -400 68614 800
rect 69018 -400 69074 800
rect 69478 -400 69534 800
rect 69846 -400 69902 800
rect 70306 -400 70362 800
rect 70766 -400 70822 800
rect 71226 -400 71282 800
rect 71594 -400 71650 800
rect 72054 -400 72110 800
rect 72514 -400 72570 800
rect 72882 -400 72938 800
rect 73342 -400 73398 800
rect 73802 -400 73858 800
rect 74262 -400 74318 800
rect 74630 -400 74686 800
rect 75090 -400 75146 800
rect 75550 -400 75606 800
rect 76010 -400 76066 800
rect 76378 -400 76434 800
rect 76838 -400 76894 800
rect 77298 -400 77354 800
rect 77758 -400 77814 800
rect 78126 -400 78182 800
rect 78586 -400 78642 800
rect 79046 -400 79102 800
rect 79506 -400 79562 800
rect 79874 -400 79930 800
rect 80334 -400 80390 800
rect 80794 -400 80850 800
rect 81162 -400 81218 800
rect 81622 -400 81678 800
rect 82082 -400 82138 800
rect 82542 -400 82598 800
rect 82910 -400 82966 800
rect 83370 -400 83426 800
rect 83830 -400 83886 800
rect 84290 -400 84346 800
rect 84658 -400 84714 800
rect 85118 -400 85174 800
rect 85578 -400 85634 800
rect 86038 -400 86094 800
rect 86406 -400 86462 800
rect 86866 -400 86922 800
rect 87326 -400 87382 800
rect 87786 -400 87842 800
rect 88154 -400 88210 800
rect 88614 -400 88670 800
rect 89074 -400 89130 800
rect 89442 -400 89498 800
rect 89902 -400 89958 800
rect 90362 -400 90418 800
rect 90822 -400 90878 800
rect 91190 -400 91246 800
rect 91650 -400 91706 800
rect 92110 -400 92166 800
rect 92570 -400 92626 800
rect 92938 -400 92994 800
rect 93398 -400 93454 800
rect 93858 -400 93914 800
rect 94318 -400 94374 800
rect 94686 -400 94742 800
rect 95146 -400 95202 800
rect 95606 -400 95662 800
rect 96066 -400 96122 800
rect 96434 -400 96490 800
rect 96894 -400 96950 800
rect 97354 -400 97410 800
rect 97722 -400 97778 800
rect 98182 -400 98238 800
rect 98642 -400 98698 800
rect 99102 -400 99158 800
rect 99470 -400 99526 800
rect 99930 -400 99986 800
rect 100390 -400 100446 800
rect 100850 -400 100906 800
rect 101218 -400 101274 800
rect 101678 -400 101734 800
rect 102138 -400 102194 800
rect 102598 -400 102654 800
rect 102966 -400 103022 800
rect 103426 -400 103482 800
rect 103886 -400 103942 800
rect 104254 -400 104310 800
rect 104714 -400 104770 800
rect 105174 -400 105230 800
rect 105634 -400 105690 800
rect 106002 -400 106058 800
rect 106462 -400 106518 800
rect 106922 -400 106978 800
rect 107382 -400 107438 800
rect 107750 -400 107806 800
rect 108210 -400 108266 800
rect 108670 -400 108726 800
rect 109130 -400 109186 800
rect 109498 -400 109554 800
rect 109958 -400 110014 800
rect 110418 -400 110474 800
rect 110878 -400 110934 800
rect 111246 -400 111302 800
rect 111706 -400 111762 800
rect 112166 -400 112222 800
rect 112534 -400 112590 800
rect 112994 -400 113050 800
rect 113454 -400 113510 800
rect 113914 -400 113970 800
rect 114282 -400 114338 800
rect 114742 -400 114798 800
rect 115202 -400 115258 800
rect 115662 -400 115718 800
rect 116030 -400 116086 800
rect 116490 -400 116546 800
rect 116950 -400 117006 800
rect 117410 -400 117466 800
rect 117778 -400 117834 800
rect 118238 -400 118294 800
rect 118698 -400 118754 800
rect 119158 -400 119214 800
rect 119526 -400 119582 800
rect 119986 -400 120042 800
rect 120446 -400 120502 800
rect 120814 -400 120870 800
rect 121274 -400 121330 800
rect 121734 -400 121790 800
rect 122194 -400 122250 800
rect 122562 -400 122618 800
rect 123022 -400 123078 800
rect 123482 -400 123538 800
rect 123942 -400 123998 800
rect 124310 -400 124366 800
rect 124770 -400 124826 800
rect 125230 -400 125286 800
rect 125690 -400 125746 800
rect 126058 -400 126114 800
rect 126518 -400 126574 800
rect 126978 -400 127034 800
rect 127438 -400 127494 800
rect 127806 -400 127862 800
rect 128266 -400 128322 800
rect 128726 -400 128782 800
rect 129094 -400 129150 800
rect 129554 -400 129610 800
rect 130014 -400 130070 800
rect 130474 -400 130530 800
rect 130842 -400 130898 800
rect 131302 -400 131358 800
rect 131762 -400 131818 800
rect 132222 -400 132278 800
rect 132590 -400 132646 800
rect 133050 -400 133106 800
rect 133510 -400 133566 800
rect 133970 -400 134026 800
rect 134338 -400 134394 800
rect 134798 -400 134854 800
rect 135258 -400 135314 800
rect 135718 -400 135774 800
rect 136086 -400 136142 800
rect 136546 -400 136602 800
rect 137006 -400 137062 800
rect 137374 -400 137430 800
rect 137834 -400 137890 800
rect 138294 -400 138350 800
rect 138754 -400 138810 800
rect 139122 -400 139178 800
rect 139582 -400 139638 800
rect 140042 -400 140098 800
rect 140502 -400 140558 800
rect 140870 -400 140926 800
rect 141330 -400 141386 800
rect 141790 -400 141846 800
rect 142250 -400 142306 800
rect 142618 -400 142674 800
rect 143078 -400 143134 800
rect 143538 -400 143594 800
rect 143998 -400 144054 800
rect 144366 -400 144422 800
rect 144826 -400 144882 800
rect 145286 -400 145342 800
rect 145654 -400 145710 800
rect 146114 -400 146170 800
rect 146574 -400 146630 800
rect 147034 -400 147090 800
rect 147402 -400 147458 800
rect 147862 -400 147918 800
rect 148322 -400 148378 800
rect 148782 -400 148838 800
rect 149150 -400 149206 800
rect 149610 -400 149666 800
rect 150070 -400 150126 800
rect 150530 -400 150586 800
rect 150898 -400 150954 800
rect 151358 -400 151414 800
rect 151818 -400 151874 800
rect 152186 -400 152242 800
rect 152646 -400 152702 800
rect 153106 -400 153162 800
rect 153566 -400 153622 800
rect 153934 -400 153990 800
rect 154394 -400 154450 800
rect 154854 -400 154910 800
rect 155314 -400 155370 800
rect 155682 -400 155738 800
rect 156142 -400 156198 800
rect 156602 -400 156658 800
rect 157062 -400 157118 800
rect 157430 -400 157486 800
rect 157890 -400 157946 800
rect 158350 -400 158406 800
rect 158810 -400 158866 800
rect 159178 -400 159234 800
rect 159638 -400 159694 800
rect 160098 -400 160154 800
rect 160466 -400 160522 800
rect 160926 -400 160982 800
rect 161386 -400 161442 800
rect 161846 -400 161902 800
rect 162214 -400 162270 800
rect 162674 -400 162730 800
rect 163134 -400 163190 800
rect 163594 -400 163650 800
rect 163962 -400 164018 800
rect 164422 -400 164478 800
rect 164882 -400 164938 800
rect 165342 -400 165398 800
rect 165710 -400 165766 800
rect 166170 -400 166226 800
rect 166630 -400 166686 800
rect 167090 -400 167146 800
rect 167458 -400 167514 800
rect 167918 -400 167974 800
rect 168378 -400 168434 800
rect 168746 -400 168802 800
rect 169206 -400 169262 800
rect 169666 -400 169722 800
rect 170126 -400 170182 800
rect 170494 -400 170550 800
rect 170954 -400 171010 800
rect 171414 -400 171470 800
rect 171874 -400 171930 800
rect 172242 -400 172298 800
rect 172702 -400 172758 800
rect 173162 -400 173218 800
rect 173622 -400 173678 800
rect 173990 -400 174046 800
rect 174450 -400 174506 800
rect 174910 -400 174966 800
rect 175370 -400 175426 800
rect 175738 -400 175794 800
rect 176198 -400 176254 800
rect 176658 -400 176714 800
rect 177026 -400 177082 800
rect 177486 -400 177542 800
rect 177946 -400 178002 800
rect 178406 -400 178462 800
rect 178774 -400 178830 800
rect 179234 -400 179290 800
rect 179694 -400 179750 800
rect 180154 -400 180210 800
rect 180522 -400 180578 800
rect 180982 -400 181038 800
rect 181442 -400 181498 800
rect 181902 -400 181958 800
rect 182270 -400 182326 800
rect 182730 -400 182786 800
rect 183190 -400 183246 800
rect 183650 -400 183706 800
rect 184018 -400 184074 800
rect 184478 -400 184534 800
rect 184938 -400 184994 800
rect 185306 -400 185362 800
rect 185766 -400 185822 800
rect 186226 -400 186282 800
rect 186686 -400 186742 800
rect 187054 -400 187110 800
rect 187514 -400 187570 800
rect 187974 -400 188030 800
rect 188434 -400 188490 800
rect 188802 -400 188858 800
rect 189262 -400 189318 800
rect 189722 -400 189778 800
rect 190182 -400 190238 800
rect 190550 -400 190606 800
rect 191010 -400 191066 800
rect 191470 -400 191526 800
rect 191930 -400 191986 800
rect 192298 -400 192354 800
rect 192758 -400 192814 800
rect 193218 -400 193274 800
rect 193586 -400 193642 800
rect 194046 -400 194102 800
rect 194506 -400 194562 800
rect 194966 -400 195022 800
rect 195334 -400 195390 800
rect 195794 -400 195850 800
rect 196254 -400 196310 800
rect 196714 -400 196770 800
rect 197082 -400 197138 800
rect 197542 -400 197598 800
rect 198002 -400 198058 800
rect 198462 -400 198518 800
rect 198830 -400 198886 800
rect 199290 -400 199346 800
rect 199750 -400 199806 800
<< obsm2 >>
rect 314 10144 514 10606
rect 682 10144 974 10606
rect 1142 10144 1434 10606
rect 1602 10144 1802 10606
rect 1970 10144 2262 10606
rect 2430 10144 2722 10606
rect 2890 10144 3182 10606
rect 3350 10144 3550 10606
rect 3718 10144 4010 10606
rect 4178 10144 4470 10606
rect 4638 10144 4930 10606
rect 5098 10144 5298 10606
rect 5466 10144 5758 10606
rect 5926 10144 6218 10606
rect 6386 10144 6678 10606
rect 6846 10144 7046 10606
rect 7214 10144 7506 10606
rect 7674 10144 7966 10606
rect 8134 10144 8334 10606
rect 8502 10144 8794 10606
rect 8962 10144 9254 10606
rect 9422 10144 9714 10606
rect 9882 10144 10082 10606
rect 10250 10144 10542 10606
rect 10710 10144 11002 10606
rect 11170 10144 11462 10606
rect 11630 10144 11830 10606
rect 11998 10144 12290 10606
rect 12458 10144 12750 10606
rect 12918 10144 13210 10606
rect 13378 10144 13578 10606
rect 13746 10144 14038 10606
rect 14206 10144 14498 10606
rect 14666 10144 14958 10606
rect 15126 10144 15326 10606
rect 15494 10144 15786 10606
rect 15954 10144 16246 10606
rect 16414 10144 16614 10606
rect 16782 10144 17074 10606
rect 17242 10144 17534 10606
rect 17702 10144 17994 10606
rect 18162 10144 18362 10606
rect 18530 10144 18822 10606
rect 18990 10144 19282 10606
rect 19450 10144 19742 10606
rect 19910 10144 20110 10606
rect 20278 10144 20570 10606
rect 20738 10144 21030 10606
rect 21198 10144 21490 10606
rect 21658 10144 21858 10606
rect 22026 10144 22318 10606
rect 22486 10144 22778 10606
rect 22946 10144 23238 10606
rect 23406 10144 23606 10606
rect 23774 10144 24066 10606
rect 24234 10144 24526 10606
rect 24694 10144 24894 10606
rect 25062 10144 25354 10606
rect 25522 10144 25814 10606
rect 25982 10144 26274 10606
rect 26442 10144 26642 10606
rect 26810 10144 27102 10606
rect 27270 10144 27562 10606
rect 27730 10144 28022 10606
rect 28190 10144 28390 10606
rect 28558 10144 28850 10606
rect 29018 10144 29310 10606
rect 29478 10144 29770 10606
rect 29938 10144 30138 10606
rect 30306 10144 30598 10606
rect 30766 10144 31058 10606
rect 31226 10144 31518 10606
rect 31686 10144 31886 10606
rect 32054 10144 32346 10606
rect 32514 10144 32806 10606
rect 32974 10144 33174 10606
rect 33342 10144 33634 10606
rect 33802 10144 34094 10606
rect 34262 10144 34554 10606
rect 34722 10144 34922 10606
rect 35090 10144 35382 10606
rect 35550 10144 35842 10606
rect 36010 10144 36302 10606
rect 36470 10144 36670 10606
rect 36838 10144 37130 10606
rect 37298 10144 37590 10606
rect 37758 10144 38050 10606
rect 38218 10144 38418 10606
rect 38586 10144 38878 10606
rect 39046 10144 39338 10606
rect 39506 10144 39798 10606
rect 39966 10144 40166 10606
rect 40334 10144 40626 10606
rect 40794 10144 41086 10606
rect 41254 10144 41454 10606
rect 41622 10144 41914 10606
rect 42082 10144 42374 10606
rect 42542 10144 42834 10606
rect 43002 10144 43202 10606
rect 43370 10144 43662 10606
rect 43830 10144 44122 10606
rect 44290 10144 44582 10606
rect 44750 10144 44950 10606
rect 45118 10144 45410 10606
rect 45578 10144 45870 10606
rect 46038 10144 46330 10606
rect 46498 10144 46698 10606
rect 46866 10144 47158 10606
rect 47326 10144 47618 10606
rect 47786 10144 48078 10606
rect 48246 10144 48446 10606
rect 48614 10144 48906 10606
rect 49074 10144 49366 10606
rect 49534 10144 49734 10606
rect 49902 10144 50194 10606
rect 50362 10144 50654 10606
rect 50822 10144 51114 10606
rect 51282 10144 51482 10606
rect 51650 10144 51942 10606
rect 52110 10144 52402 10606
rect 52570 10144 52862 10606
rect 53030 10144 53230 10606
rect 53398 10144 53690 10606
rect 53858 10144 54150 10606
rect 54318 10144 54610 10606
rect 54778 10144 54978 10606
rect 55146 10144 55438 10606
rect 55606 10144 55898 10606
rect 56066 10144 56266 10606
rect 56434 10144 56726 10606
rect 56894 10144 57186 10606
rect 57354 10144 57646 10606
rect 57814 10144 58014 10606
rect 58182 10144 58474 10606
rect 58642 10144 58934 10606
rect 59102 10144 59394 10606
rect 59562 10144 59762 10606
rect 59930 10144 60222 10606
rect 60390 10144 60682 10606
rect 60850 10144 61142 10606
rect 61310 10144 61510 10606
rect 61678 10144 61970 10606
rect 62138 10144 62430 10606
rect 62598 10144 62890 10606
rect 63058 10144 63258 10606
rect 63426 10144 63718 10606
rect 63886 10144 64178 10606
rect 64346 10144 64546 10606
rect 64714 10144 65006 10606
rect 65174 10144 65466 10606
rect 65634 10144 65926 10606
rect 66094 10144 66294 10606
rect 66462 10144 66754 10606
rect 66922 10144 67214 10606
rect 67382 10144 67674 10606
rect 67842 10144 68042 10606
rect 68210 10144 68502 10606
rect 68670 10144 68962 10606
rect 69130 10144 69422 10606
rect 69590 10144 69790 10606
rect 69958 10144 70250 10606
rect 70418 10144 70710 10606
rect 70878 10144 71170 10606
rect 71338 10144 71538 10606
rect 71706 10144 71998 10606
rect 72166 10144 72458 10606
rect 72626 10144 72826 10606
rect 72994 10144 73286 10606
rect 73454 10144 73746 10606
rect 73914 10144 74206 10606
rect 74374 10144 74574 10606
rect 74742 10144 75034 10606
rect 75202 10144 75494 10606
rect 75662 10144 75954 10606
rect 76122 10144 76322 10606
rect 76490 10144 76782 10606
rect 76950 10144 77242 10606
rect 77410 10144 77702 10606
rect 77870 10144 78070 10606
rect 78238 10144 78530 10606
rect 78698 10144 78990 10606
rect 79158 10144 79450 10606
rect 79618 10144 79818 10606
rect 79986 10144 80278 10606
rect 80446 10144 80738 10606
rect 80906 10144 81106 10606
rect 81274 10144 81566 10606
rect 81734 10144 82026 10606
rect 82194 10144 82486 10606
rect 82654 10144 82854 10606
rect 83022 10144 83314 10606
rect 83482 10144 83774 10606
rect 83942 10144 84234 10606
rect 84402 10144 84602 10606
rect 84770 10144 85062 10606
rect 85230 10144 85522 10606
rect 85690 10144 85982 10606
rect 86150 10144 86350 10606
rect 86518 10144 86810 10606
rect 86978 10144 87270 10606
rect 87438 10144 87730 10606
rect 87898 10144 88098 10606
rect 88266 10144 88558 10606
rect 88726 10144 89018 10606
rect 89186 10144 89386 10606
rect 89554 10144 89846 10606
rect 90014 10144 90306 10606
rect 90474 10144 90766 10606
rect 90934 10144 91134 10606
rect 91302 10144 91594 10606
rect 91762 10144 92054 10606
rect 92222 10144 92514 10606
rect 92682 10144 92882 10606
rect 93050 10144 93342 10606
rect 93510 10144 93802 10606
rect 93970 10144 94262 10606
rect 94430 10144 94630 10606
rect 94798 10144 95090 10606
rect 95258 10144 95550 10606
rect 95718 10144 96010 10606
rect 96178 10144 96378 10606
rect 96546 10144 96838 10606
rect 97006 10144 97298 10606
rect 97466 10144 97666 10606
rect 97834 10144 98126 10606
rect 98294 10144 98586 10606
rect 98754 10144 99046 10606
rect 99214 10144 99414 10606
rect 99582 10144 99874 10606
rect 100042 10144 100334 10606
rect 100502 10144 100794 10606
rect 100962 10144 101162 10606
rect 101330 10144 101622 10606
rect 101790 10144 102082 10606
rect 102250 10144 102542 10606
rect 102710 10144 102910 10606
rect 103078 10144 103370 10606
rect 103538 10144 103830 10606
rect 103998 10144 104198 10606
rect 104366 10144 104658 10606
rect 104826 10144 105118 10606
rect 105286 10144 105578 10606
rect 105746 10144 105946 10606
rect 106114 10144 106406 10606
rect 106574 10144 106866 10606
rect 107034 10144 107326 10606
rect 107494 10144 107694 10606
rect 107862 10144 108154 10606
rect 108322 10144 108614 10606
rect 108782 10144 109074 10606
rect 109242 10144 109442 10606
rect 109610 10144 109902 10606
rect 110070 10144 110362 10606
rect 110530 10144 110822 10606
rect 110990 10144 111190 10606
rect 111358 10144 111650 10606
rect 111818 10144 112110 10606
rect 112278 10144 112478 10606
rect 112646 10144 112938 10606
rect 113106 10144 113398 10606
rect 113566 10144 113858 10606
rect 114026 10144 114226 10606
rect 114394 10144 114686 10606
rect 114854 10144 115146 10606
rect 115314 10144 115606 10606
rect 115774 10144 115974 10606
rect 116142 10144 116434 10606
rect 116602 10144 116894 10606
rect 117062 10144 117354 10606
rect 117522 10144 117722 10606
rect 117890 10144 118182 10606
rect 118350 10144 118642 10606
rect 118810 10144 119102 10606
rect 119270 10144 119470 10606
rect 119638 10144 119930 10606
rect 120098 10144 120390 10606
rect 120558 10144 120758 10606
rect 120926 10144 121218 10606
rect 121386 10144 121678 10606
rect 121846 10144 122138 10606
rect 122306 10144 122506 10606
rect 122674 10144 122966 10606
rect 123134 10144 123426 10606
rect 123594 10144 123886 10606
rect 124054 10144 124254 10606
rect 124422 10144 124714 10606
rect 124882 10144 125174 10606
rect 125342 10144 125634 10606
rect 125802 10144 126002 10606
rect 126170 10144 126462 10606
rect 126630 10144 126922 10606
rect 127090 10144 127382 10606
rect 127550 10144 127750 10606
rect 127918 10144 128210 10606
rect 128378 10144 128670 10606
rect 128838 10144 129038 10606
rect 129206 10144 129498 10606
rect 129666 10144 129958 10606
rect 130126 10144 130418 10606
rect 130586 10144 130786 10606
rect 130954 10144 131246 10606
rect 131414 10144 131706 10606
rect 131874 10144 132166 10606
rect 132334 10144 132534 10606
rect 132702 10144 132994 10606
rect 133162 10144 133454 10606
rect 133622 10144 133914 10606
rect 134082 10144 134282 10606
rect 134450 10144 134742 10606
rect 134910 10144 135202 10606
rect 135370 10144 135662 10606
rect 135830 10144 136030 10606
rect 136198 10144 136490 10606
rect 136658 10144 136950 10606
rect 137118 10144 137318 10606
rect 137486 10144 137778 10606
rect 137946 10144 138238 10606
rect 138406 10144 138698 10606
rect 138866 10144 139066 10606
rect 139234 10144 139526 10606
rect 139694 10144 139986 10606
rect 140154 10144 140446 10606
rect 140614 10144 140814 10606
rect 140982 10144 141274 10606
rect 141442 10144 141734 10606
rect 141902 10144 142194 10606
rect 142362 10144 142562 10606
rect 142730 10144 143022 10606
rect 143190 10144 143482 10606
rect 143650 10144 143942 10606
rect 144110 10144 144310 10606
rect 144478 10144 144770 10606
rect 144938 10144 145230 10606
rect 145398 10144 145598 10606
rect 145766 10144 146058 10606
rect 146226 10144 146518 10606
rect 146686 10144 146978 10606
rect 147146 10144 147346 10606
rect 147514 10144 147806 10606
rect 147974 10144 148266 10606
rect 148434 10144 148726 10606
rect 148894 10144 149094 10606
rect 149262 10144 149554 10606
rect 149722 10144 150014 10606
rect 150182 10144 150474 10606
rect 150642 10144 150842 10606
rect 151010 10144 151302 10606
rect 151470 10144 151762 10606
rect 151930 10144 152130 10606
rect 152298 10144 152590 10606
rect 152758 10144 153050 10606
rect 153218 10144 153510 10606
rect 153678 10144 153878 10606
rect 154046 10144 154338 10606
rect 154506 10144 154798 10606
rect 154966 10144 155258 10606
rect 155426 10144 155626 10606
rect 155794 10144 156086 10606
rect 156254 10144 156546 10606
rect 156714 10144 157006 10606
rect 157174 10144 157374 10606
rect 157542 10144 157834 10606
rect 158002 10144 158294 10606
rect 158462 10144 158754 10606
rect 158922 10144 159122 10606
rect 159290 10144 159582 10606
rect 159750 10144 160042 10606
rect 160210 10144 160410 10606
rect 160578 10144 160870 10606
rect 161038 10144 161330 10606
rect 161498 10144 161790 10606
rect 161958 10144 162158 10606
rect 162326 10144 162618 10606
rect 162786 10144 163078 10606
rect 163246 10144 163538 10606
rect 163706 10144 163906 10606
rect 164074 10144 164366 10606
rect 164534 10144 164826 10606
rect 164994 10144 165286 10606
rect 165454 10144 165654 10606
rect 165822 10144 166114 10606
rect 166282 10144 166574 10606
rect 166742 10144 167034 10606
rect 167202 10144 167402 10606
rect 167570 10144 167862 10606
rect 168030 10144 168322 10606
rect 168490 10144 168690 10606
rect 168858 10144 169150 10606
rect 169318 10144 169610 10606
rect 169778 10144 170070 10606
rect 170238 10144 170438 10606
rect 170606 10144 170898 10606
rect 171066 10144 171358 10606
rect 171526 10144 171818 10606
rect 171986 10144 172186 10606
rect 172354 10144 172646 10606
rect 172814 10144 173106 10606
rect 173274 10144 173566 10606
rect 173734 10144 173934 10606
rect 174102 10144 174394 10606
rect 174562 10144 174854 10606
rect 175022 10144 175314 10606
rect 175482 10144 175682 10606
rect 175850 10144 176142 10606
rect 176310 10144 176602 10606
rect 176770 10144 176970 10606
rect 177138 10144 177430 10606
rect 177598 10144 177890 10606
rect 178058 10144 178350 10606
rect 178518 10144 178718 10606
rect 178886 10144 179178 10606
rect 179346 10144 179638 10606
rect 179806 10144 180098 10606
rect 180266 10144 180466 10606
rect 180634 10144 180926 10606
rect 181094 10144 181386 10606
rect 181554 10144 181846 10606
rect 182014 10144 182214 10606
rect 182382 10144 182674 10606
rect 182842 10144 183134 10606
rect 183302 10144 183594 10606
rect 183762 10144 183962 10606
rect 184130 10144 184422 10606
rect 184590 10144 184882 10606
rect 185050 10144 185250 10606
rect 185418 10144 185710 10606
rect 185878 10144 186170 10606
rect 186338 10144 186630 10606
rect 186798 10144 186998 10606
rect 187166 10144 187458 10606
rect 187626 10144 187918 10606
rect 188086 10144 188378 10606
rect 188546 10144 188746 10606
rect 188914 10144 189206 10606
rect 189374 10144 189666 10606
rect 189834 10144 190126 10606
rect 190294 10144 190494 10606
rect 190662 10144 190954 10606
rect 191122 10144 191414 10606
rect 191582 10144 191874 10606
rect 192042 10144 192242 10606
rect 192410 10144 192702 10606
rect 192870 10144 193162 10606
rect 193330 10144 193530 10606
rect 193698 10144 193990 10606
rect 194158 10144 194450 10606
rect 194618 10144 194910 10606
rect 195078 10144 195278 10606
rect 195446 10144 195738 10606
rect 195906 10144 196198 10606
rect 196366 10144 196658 10606
rect 196826 10144 197026 10606
rect 197194 10144 197486 10606
rect 197654 10144 197946 10606
rect 198114 10144 198406 10606
rect 198574 10144 198774 10606
rect 198942 10144 199234 10606
rect 199402 10144 199694 10606
rect 204 856 199804 10144
rect 314 2 514 856
rect 682 2 974 856
rect 1142 2 1434 856
rect 1602 2 1802 856
rect 1970 2 2262 856
rect 2430 2 2722 856
rect 2890 2 3182 856
rect 3350 2 3550 856
rect 3718 2 4010 856
rect 4178 2 4470 856
rect 4638 2 4930 856
rect 5098 2 5298 856
rect 5466 2 5758 856
rect 5926 2 6218 856
rect 6386 2 6678 856
rect 6846 2 7046 856
rect 7214 2 7506 856
rect 7674 2 7966 856
rect 8134 2 8334 856
rect 8502 2 8794 856
rect 8962 2 9254 856
rect 9422 2 9714 856
rect 9882 2 10082 856
rect 10250 2 10542 856
rect 10710 2 11002 856
rect 11170 2 11462 856
rect 11630 2 11830 856
rect 11998 2 12290 856
rect 12458 2 12750 856
rect 12918 2 13210 856
rect 13378 2 13578 856
rect 13746 2 14038 856
rect 14206 2 14498 856
rect 14666 2 14958 856
rect 15126 2 15326 856
rect 15494 2 15786 856
rect 15954 2 16246 856
rect 16414 2 16614 856
rect 16782 2 17074 856
rect 17242 2 17534 856
rect 17702 2 17994 856
rect 18162 2 18362 856
rect 18530 2 18822 856
rect 18990 2 19282 856
rect 19450 2 19742 856
rect 19910 2 20110 856
rect 20278 2 20570 856
rect 20738 2 21030 856
rect 21198 2 21490 856
rect 21658 2 21858 856
rect 22026 2 22318 856
rect 22486 2 22778 856
rect 22946 2 23238 856
rect 23406 2 23606 856
rect 23774 2 24066 856
rect 24234 2 24526 856
rect 24694 2 24894 856
rect 25062 2 25354 856
rect 25522 2 25814 856
rect 25982 2 26274 856
rect 26442 2 26642 856
rect 26810 2 27102 856
rect 27270 2 27562 856
rect 27730 2 28022 856
rect 28190 2 28390 856
rect 28558 2 28850 856
rect 29018 2 29310 856
rect 29478 2 29770 856
rect 29938 2 30138 856
rect 30306 2 30598 856
rect 30766 2 31058 856
rect 31226 2 31518 856
rect 31686 2 31886 856
rect 32054 2 32346 856
rect 32514 2 32806 856
rect 32974 2 33174 856
rect 33342 2 33634 856
rect 33802 2 34094 856
rect 34262 2 34554 856
rect 34722 2 34922 856
rect 35090 2 35382 856
rect 35550 2 35842 856
rect 36010 2 36302 856
rect 36470 2 36670 856
rect 36838 2 37130 856
rect 37298 2 37590 856
rect 37758 2 38050 856
rect 38218 2 38418 856
rect 38586 2 38878 856
rect 39046 2 39338 856
rect 39506 2 39798 856
rect 39966 2 40166 856
rect 40334 2 40626 856
rect 40794 2 41086 856
rect 41254 2 41454 856
rect 41622 2 41914 856
rect 42082 2 42374 856
rect 42542 2 42834 856
rect 43002 2 43202 856
rect 43370 2 43662 856
rect 43830 2 44122 856
rect 44290 2 44582 856
rect 44750 2 44950 856
rect 45118 2 45410 856
rect 45578 2 45870 856
rect 46038 2 46330 856
rect 46498 2 46698 856
rect 46866 2 47158 856
rect 47326 2 47618 856
rect 47786 2 48078 856
rect 48246 2 48446 856
rect 48614 2 48906 856
rect 49074 2 49366 856
rect 49534 2 49734 856
rect 49902 2 50194 856
rect 50362 2 50654 856
rect 50822 2 51114 856
rect 51282 2 51482 856
rect 51650 2 51942 856
rect 52110 2 52402 856
rect 52570 2 52862 856
rect 53030 2 53230 856
rect 53398 2 53690 856
rect 53858 2 54150 856
rect 54318 2 54610 856
rect 54778 2 54978 856
rect 55146 2 55438 856
rect 55606 2 55898 856
rect 56066 2 56266 856
rect 56434 2 56726 856
rect 56894 2 57186 856
rect 57354 2 57646 856
rect 57814 2 58014 856
rect 58182 2 58474 856
rect 58642 2 58934 856
rect 59102 2 59394 856
rect 59562 2 59762 856
rect 59930 2 60222 856
rect 60390 2 60682 856
rect 60850 2 61142 856
rect 61310 2 61510 856
rect 61678 2 61970 856
rect 62138 2 62430 856
rect 62598 2 62890 856
rect 63058 2 63258 856
rect 63426 2 63718 856
rect 63886 2 64178 856
rect 64346 2 64546 856
rect 64714 2 65006 856
rect 65174 2 65466 856
rect 65634 2 65926 856
rect 66094 2 66294 856
rect 66462 2 66754 856
rect 66922 2 67214 856
rect 67382 2 67674 856
rect 67842 2 68042 856
rect 68210 2 68502 856
rect 68670 2 68962 856
rect 69130 2 69422 856
rect 69590 2 69790 856
rect 69958 2 70250 856
rect 70418 2 70710 856
rect 70878 2 71170 856
rect 71338 2 71538 856
rect 71706 2 71998 856
rect 72166 2 72458 856
rect 72626 2 72826 856
rect 72994 2 73286 856
rect 73454 2 73746 856
rect 73914 2 74206 856
rect 74374 2 74574 856
rect 74742 2 75034 856
rect 75202 2 75494 856
rect 75662 2 75954 856
rect 76122 2 76322 856
rect 76490 2 76782 856
rect 76950 2 77242 856
rect 77410 2 77702 856
rect 77870 2 78070 856
rect 78238 2 78530 856
rect 78698 2 78990 856
rect 79158 2 79450 856
rect 79618 2 79818 856
rect 79986 2 80278 856
rect 80446 2 80738 856
rect 80906 2 81106 856
rect 81274 2 81566 856
rect 81734 2 82026 856
rect 82194 2 82486 856
rect 82654 2 82854 856
rect 83022 2 83314 856
rect 83482 2 83774 856
rect 83942 2 84234 856
rect 84402 2 84602 856
rect 84770 2 85062 856
rect 85230 2 85522 856
rect 85690 2 85982 856
rect 86150 2 86350 856
rect 86518 2 86810 856
rect 86978 2 87270 856
rect 87438 2 87730 856
rect 87898 2 88098 856
rect 88266 2 88558 856
rect 88726 2 89018 856
rect 89186 2 89386 856
rect 89554 2 89846 856
rect 90014 2 90306 856
rect 90474 2 90766 856
rect 90934 2 91134 856
rect 91302 2 91594 856
rect 91762 2 92054 856
rect 92222 2 92514 856
rect 92682 2 92882 856
rect 93050 2 93342 856
rect 93510 2 93802 856
rect 93970 2 94262 856
rect 94430 2 94630 856
rect 94798 2 95090 856
rect 95258 2 95550 856
rect 95718 2 96010 856
rect 96178 2 96378 856
rect 96546 2 96838 856
rect 97006 2 97298 856
rect 97466 2 97666 856
rect 97834 2 98126 856
rect 98294 2 98586 856
rect 98754 2 99046 856
rect 99214 2 99414 856
rect 99582 2 99874 856
rect 100042 2 100334 856
rect 100502 2 100794 856
rect 100962 2 101162 856
rect 101330 2 101622 856
rect 101790 2 102082 856
rect 102250 2 102542 856
rect 102710 2 102910 856
rect 103078 2 103370 856
rect 103538 2 103830 856
rect 103998 2 104198 856
rect 104366 2 104658 856
rect 104826 2 105118 856
rect 105286 2 105578 856
rect 105746 2 105946 856
rect 106114 2 106406 856
rect 106574 2 106866 856
rect 107034 2 107326 856
rect 107494 2 107694 856
rect 107862 2 108154 856
rect 108322 2 108614 856
rect 108782 2 109074 856
rect 109242 2 109442 856
rect 109610 2 109902 856
rect 110070 2 110362 856
rect 110530 2 110822 856
rect 110990 2 111190 856
rect 111358 2 111650 856
rect 111818 2 112110 856
rect 112278 2 112478 856
rect 112646 2 112938 856
rect 113106 2 113398 856
rect 113566 2 113858 856
rect 114026 2 114226 856
rect 114394 2 114686 856
rect 114854 2 115146 856
rect 115314 2 115606 856
rect 115774 2 115974 856
rect 116142 2 116434 856
rect 116602 2 116894 856
rect 117062 2 117354 856
rect 117522 2 117722 856
rect 117890 2 118182 856
rect 118350 2 118642 856
rect 118810 2 119102 856
rect 119270 2 119470 856
rect 119638 2 119930 856
rect 120098 2 120390 856
rect 120558 2 120758 856
rect 120926 2 121218 856
rect 121386 2 121678 856
rect 121846 2 122138 856
rect 122306 2 122506 856
rect 122674 2 122966 856
rect 123134 2 123426 856
rect 123594 2 123886 856
rect 124054 2 124254 856
rect 124422 2 124714 856
rect 124882 2 125174 856
rect 125342 2 125634 856
rect 125802 2 126002 856
rect 126170 2 126462 856
rect 126630 2 126922 856
rect 127090 2 127382 856
rect 127550 2 127750 856
rect 127918 2 128210 856
rect 128378 2 128670 856
rect 128838 2 129038 856
rect 129206 2 129498 856
rect 129666 2 129958 856
rect 130126 2 130418 856
rect 130586 2 130786 856
rect 130954 2 131246 856
rect 131414 2 131706 856
rect 131874 2 132166 856
rect 132334 2 132534 856
rect 132702 2 132994 856
rect 133162 2 133454 856
rect 133622 2 133914 856
rect 134082 2 134282 856
rect 134450 2 134742 856
rect 134910 2 135202 856
rect 135370 2 135662 856
rect 135830 2 136030 856
rect 136198 2 136490 856
rect 136658 2 136950 856
rect 137118 2 137318 856
rect 137486 2 137778 856
rect 137946 2 138238 856
rect 138406 2 138698 856
rect 138866 2 139066 856
rect 139234 2 139526 856
rect 139694 2 139986 856
rect 140154 2 140446 856
rect 140614 2 140814 856
rect 140982 2 141274 856
rect 141442 2 141734 856
rect 141902 2 142194 856
rect 142362 2 142562 856
rect 142730 2 143022 856
rect 143190 2 143482 856
rect 143650 2 143942 856
rect 144110 2 144310 856
rect 144478 2 144770 856
rect 144938 2 145230 856
rect 145398 2 145598 856
rect 145766 2 146058 856
rect 146226 2 146518 856
rect 146686 2 146978 856
rect 147146 2 147346 856
rect 147514 2 147806 856
rect 147974 2 148266 856
rect 148434 2 148726 856
rect 148894 2 149094 856
rect 149262 2 149554 856
rect 149722 2 150014 856
rect 150182 2 150474 856
rect 150642 2 150842 856
rect 151010 2 151302 856
rect 151470 2 151762 856
rect 151930 2 152130 856
rect 152298 2 152590 856
rect 152758 2 153050 856
rect 153218 2 153510 856
rect 153678 2 153878 856
rect 154046 2 154338 856
rect 154506 2 154798 856
rect 154966 2 155258 856
rect 155426 2 155626 856
rect 155794 2 156086 856
rect 156254 2 156546 856
rect 156714 2 157006 856
rect 157174 2 157374 856
rect 157542 2 157834 856
rect 158002 2 158294 856
rect 158462 2 158754 856
rect 158922 2 159122 856
rect 159290 2 159582 856
rect 159750 2 160042 856
rect 160210 2 160410 856
rect 160578 2 160870 856
rect 161038 2 161330 856
rect 161498 2 161790 856
rect 161958 2 162158 856
rect 162326 2 162618 856
rect 162786 2 163078 856
rect 163246 2 163538 856
rect 163706 2 163906 856
rect 164074 2 164366 856
rect 164534 2 164826 856
rect 164994 2 165286 856
rect 165454 2 165654 856
rect 165822 2 166114 856
rect 166282 2 166574 856
rect 166742 2 167034 856
rect 167202 2 167402 856
rect 167570 2 167862 856
rect 168030 2 168322 856
rect 168490 2 168690 856
rect 168858 2 169150 856
rect 169318 2 169610 856
rect 169778 2 170070 856
rect 170238 2 170438 856
rect 170606 2 170898 856
rect 171066 2 171358 856
rect 171526 2 171818 856
rect 171986 2 172186 856
rect 172354 2 172646 856
rect 172814 2 173106 856
rect 173274 2 173566 856
rect 173734 2 173934 856
rect 174102 2 174394 856
rect 174562 2 174854 856
rect 175022 2 175314 856
rect 175482 2 175682 856
rect 175850 2 176142 856
rect 176310 2 176602 856
rect 176770 2 176970 856
rect 177138 2 177430 856
rect 177598 2 177890 856
rect 178058 2 178350 856
rect 178518 2 178718 856
rect 178886 2 179178 856
rect 179346 2 179638 856
rect 179806 2 180098 856
rect 180266 2 180466 856
rect 180634 2 180926 856
rect 181094 2 181386 856
rect 181554 2 181846 856
rect 182014 2 182214 856
rect 182382 2 182674 856
rect 182842 2 183134 856
rect 183302 2 183594 856
rect 183762 2 183962 856
rect 184130 2 184422 856
rect 184590 2 184882 856
rect 185050 2 185250 856
rect 185418 2 185710 856
rect 185878 2 186170 856
rect 186338 2 186630 856
rect 186798 2 186998 856
rect 187166 2 187458 856
rect 187626 2 187918 856
rect 188086 2 188378 856
rect 188546 2 188746 856
rect 188914 2 189206 856
rect 189374 2 189666 856
rect 189834 2 190126 856
rect 190294 2 190494 856
rect 190662 2 190954 856
rect 191122 2 191414 856
rect 191582 2 191874 856
rect 192042 2 192242 856
rect 192410 2 192702 856
rect 192870 2 193162 856
rect 193330 2 193530 856
rect 193698 2 193990 856
rect 194158 2 194450 856
rect 194618 2 194910 856
rect 195078 2 195278 856
rect 195446 2 195738 856
rect 195906 2 196198 856
rect 196366 2 196658 856
rect 196826 2 197026 856
rect 197194 2 197486 856
rect 197654 2 197946 856
rect 198114 2 198406 856
rect 198574 2 198774 856
rect 198942 2 199234 856
rect 199402 2 199694 856
<< metal3 >>
rect -1586 12422 201502 12482
rect -1446 12282 201362 12342
rect -1306 12142 201222 12202
rect -1166 12002 201082 12062
rect -1026 11862 200942 11922
rect -886 11722 200802 11782
rect -746 11582 200662 11642
rect -606 11442 200522 11502
rect -466 11302 200382 11362
rect -326 11162 200242 11222
rect -400 9120 800 9240
rect -400 5448 800 5568
rect -400 1776 800 1896
rect -326 -342 200242 -282
rect -466 -482 200382 -422
rect -606 -622 200522 -562
rect -746 -762 200662 -702
rect -886 -902 200802 -842
rect -1026 -1042 200942 -982
rect -1166 -1182 201082 -1122
rect -1306 -1322 201222 -1262
rect -1446 -1462 201362 -1402
rect -1586 -1602 201502 -1542
<< obsm3 >>
rect 0 9320 200000 11000
rect 880 9040 200000 9320
rect 0 5648 200000 9040
rect 880 5368 200000 5648
rect 0 1976 200000 5368
rect 880 1696 200000 1976
rect 0 0 200000 1696
<< metal4 >>
rect -1586 -1602 -1526 12482
rect -1446 -1462 -1386 12342
rect -1306 -1322 -1246 12202
rect -1166 -1182 -1106 12062
rect -1026 -1042 -966 11922
rect -886 -902 -826 11782
rect -746 -762 -686 11642
rect -606 -622 -546 11502
rect -466 -482 -406 11362
rect -326 -342 -266 11222
rect 4074 -482 4134 11362
rect 4474 -762 4534 11642
rect 4874 -1042 4934 11922
rect 5274 -1322 5334 12202
rect 5674 -1602 5734 12482
rect 24074 -482 24134 11362
rect 24474 -762 24534 11642
rect 24874 -1042 24934 11922
rect 25274 -1322 25334 12202
rect 25674 -1602 25734 12482
rect 44074 -482 44134 11362
rect 44474 -762 44534 11642
rect 44874 -1042 44934 11922
rect 45274 -1322 45334 12202
rect 45674 -1602 45734 12482
rect 64074 -482 64134 11362
rect 64474 -762 64534 11642
rect 64874 -1042 64934 11922
rect 65274 -1322 65334 12202
rect 65674 -1602 65734 12482
rect 84074 -482 84134 11362
rect 84474 -762 84534 11642
rect 84874 -1042 84934 11922
rect 85274 -1322 85334 12202
rect 85674 -1602 85734 12482
rect 104074 -482 104134 11362
rect 104474 -762 104534 11642
rect 104874 -1042 104934 11922
rect 105274 -1322 105334 12202
rect 105674 -1602 105734 12482
rect 124074 -482 124134 11362
rect 124474 -762 124534 11642
rect 124874 -1042 124934 11922
rect 125274 -1322 125334 12202
rect 125674 -1602 125734 12482
rect 144074 -482 144134 11362
rect 144474 -762 144534 11642
rect 144874 -1042 144934 11922
rect 145274 -1322 145334 12202
rect 145674 -1602 145734 12482
rect 164074 -482 164134 11362
rect 164474 -762 164534 11642
rect 164874 -1042 164934 11922
rect 165274 -1322 165334 12202
rect 165674 -1602 165734 12482
rect 184074 -482 184134 11362
rect 184474 -762 184534 11642
rect 184874 -1042 184934 11922
rect 185274 -1322 185334 12202
rect 185674 -1602 185734 12482
rect 200182 -342 200242 11222
rect 200322 -482 200382 11362
rect 200462 -622 200522 11502
rect 200602 -762 200662 11642
rect 200742 -902 200802 11782
rect 200882 -1042 200942 11922
rect 201022 -1182 201082 12062
rect 201162 -1322 201222 12202
rect 201302 -1462 201362 12342
rect 201442 -1602 201502 12482
<< obsm4 >>
rect 0 0 3994 11000
rect 4214 0 4394 11000
rect 4614 0 4794 11000
rect 5014 0 5194 11000
rect 5414 0 5594 11000
rect 5814 0 23994 11000
rect 24214 0 24394 11000
rect 24614 0 24794 11000
rect 25014 0 25194 11000
rect 25414 0 25594 11000
rect 25814 0 43994 11000
rect 44214 0 44394 11000
rect 44614 0 44794 11000
rect 45014 0 45194 11000
rect 45414 0 45594 11000
rect 45814 0 63994 11000
rect 64214 0 64394 11000
rect 64614 0 64794 11000
rect 65014 0 65194 11000
rect 65414 0 65594 11000
rect 65814 0 83994 11000
rect 84214 0 84394 11000
rect 84614 0 84794 11000
rect 85014 0 85194 11000
rect 85414 0 85594 11000
rect 85814 0 103994 11000
rect 104214 0 104394 11000
rect 104614 0 104794 11000
rect 105014 0 105194 11000
rect 105414 0 105594 11000
rect 105814 0 123994 11000
rect 124214 0 124394 11000
rect 124614 0 124794 11000
rect 125014 0 125194 11000
rect 125414 0 125594 11000
rect 125814 0 143994 11000
rect 144214 0 144394 11000
rect 144614 0 144794 11000
rect 145014 0 145194 11000
rect 145414 0 145594 11000
rect 145814 0 163994 11000
rect 164214 0 164394 11000
rect 164614 0 164794 11000
rect 165014 0 165194 11000
rect 165414 0 165594 11000
rect 165814 0 183994 11000
rect 184214 0 184394 11000
rect 184614 0 184794 11000
rect 185014 0 185194 11000
rect 185414 0 185594 11000
rect 185814 0 200000 11000
<< labels >>
rlabel metal3 s -400 1776 800 1896 6 caravel_clk
port 1 nsew signal input
rlabel metal3 s -400 5448 800 5568 6 caravel_clk2
port 2 nsew signal input
rlabel metal3 s -400 9120 800 9240 6 caravel_rstn
port 3 nsew signal input
rlabel metal2 s 1858 10200 1914 11400 6 la_data_in_core[0]
port 4 nsew signal output
rlabel metal2 s 45466 10200 45522 11400 6 la_data_in_core[100]
port 5 nsew signal output
rlabel metal2 s 45926 10200 45982 11400 6 la_data_in_core[101]
port 6 nsew signal output
rlabel metal2 s 46386 10200 46442 11400 6 la_data_in_core[102]
port 7 nsew signal output
rlabel metal2 s 46754 10200 46810 11400 6 la_data_in_core[103]
port 8 nsew signal output
rlabel metal2 s 47214 10200 47270 11400 6 la_data_in_core[104]
port 9 nsew signal output
rlabel metal2 s 47674 10200 47730 11400 6 la_data_in_core[105]
port 10 nsew signal output
rlabel metal2 s 48134 10200 48190 11400 6 la_data_in_core[106]
port 11 nsew signal output
rlabel metal2 s 48502 10200 48558 11400 6 la_data_in_core[107]
port 12 nsew signal output
rlabel metal2 s 48962 10200 49018 11400 6 la_data_in_core[108]
port 13 nsew signal output
rlabel metal2 s 49422 10200 49478 11400 6 la_data_in_core[109]
port 14 nsew signal output
rlabel metal2 s 6274 10200 6330 11400 6 la_data_in_core[10]
port 15 nsew signal output
rlabel metal2 s 49790 10200 49846 11400 6 la_data_in_core[110]
port 16 nsew signal output
rlabel metal2 s 50250 10200 50306 11400 6 la_data_in_core[111]
port 17 nsew signal output
rlabel metal2 s 50710 10200 50766 11400 6 la_data_in_core[112]
port 18 nsew signal output
rlabel metal2 s 51170 10200 51226 11400 6 la_data_in_core[113]
port 19 nsew signal output
rlabel metal2 s 51538 10200 51594 11400 6 la_data_in_core[114]
port 20 nsew signal output
rlabel metal2 s 51998 10200 52054 11400 6 la_data_in_core[115]
port 21 nsew signal output
rlabel metal2 s 52458 10200 52514 11400 6 la_data_in_core[116]
port 22 nsew signal output
rlabel metal2 s 52918 10200 52974 11400 6 la_data_in_core[117]
port 23 nsew signal output
rlabel metal2 s 53286 10200 53342 11400 6 la_data_in_core[118]
port 24 nsew signal output
rlabel metal2 s 53746 10200 53802 11400 6 la_data_in_core[119]
port 25 nsew signal output
rlabel metal2 s 6734 10200 6790 11400 6 la_data_in_core[11]
port 26 nsew signal output
rlabel metal2 s 54206 10200 54262 11400 6 la_data_in_core[120]
port 27 nsew signal output
rlabel metal2 s 54666 10200 54722 11400 6 la_data_in_core[121]
port 28 nsew signal output
rlabel metal2 s 55034 10200 55090 11400 6 la_data_in_core[122]
port 29 nsew signal output
rlabel metal2 s 55494 10200 55550 11400 6 la_data_in_core[123]
port 30 nsew signal output
rlabel metal2 s 55954 10200 56010 11400 6 la_data_in_core[124]
port 31 nsew signal output
rlabel metal2 s 56322 10200 56378 11400 6 la_data_in_core[125]
port 32 nsew signal output
rlabel metal2 s 56782 10200 56838 11400 6 la_data_in_core[126]
port 33 nsew signal output
rlabel metal2 s 57242 10200 57298 11400 6 la_data_in_core[127]
port 34 nsew signal output
rlabel metal2 s 7102 10200 7158 11400 6 la_data_in_core[12]
port 35 nsew signal output
rlabel metal2 s 7562 10200 7618 11400 6 la_data_in_core[13]
port 36 nsew signal output
rlabel metal2 s 8022 10200 8078 11400 6 la_data_in_core[14]
port 37 nsew signal output
rlabel metal2 s 8390 10200 8446 11400 6 la_data_in_core[15]
port 38 nsew signal output
rlabel metal2 s 8850 10200 8906 11400 6 la_data_in_core[16]
port 39 nsew signal output
rlabel metal2 s 9310 10200 9366 11400 6 la_data_in_core[17]
port 40 nsew signal output
rlabel metal2 s 9770 10200 9826 11400 6 la_data_in_core[18]
port 41 nsew signal output
rlabel metal2 s 10138 10200 10194 11400 6 la_data_in_core[19]
port 42 nsew signal output
rlabel metal2 s 2318 10200 2374 11400 6 la_data_in_core[1]
port 43 nsew signal output
rlabel metal2 s 10598 10200 10654 11400 6 la_data_in_core[20]
port 44 nsew signal output
rlabel metal2 s 11058 10200 11114 11400 6 la_data_in_core[21]
port 45 nsew signal output
rlabel metal2 s 11518 10200 11574 11400 6 la_data_in_core[22]
port 46 nsew signal output
rlabel metal2 s 11886 10200 11942 11400 6 la_data_in_core[23]
port 47 nsew signal output
rlabel metal2 s 12346 10200 12402 11400 6 la_data_in_core[24]
port 48 nsew signal output
rlabel metal2 s 12806 10200 12862 11400 6 la_data_in_core[25]
port 49 nsew signal output
rlabel metal2 s 13266 10200 13322 11400 6 la_data_in_core[26]
port 50 nsew signal output
rlabel metal2 s 13634 10200 13690 11400 6 la_data_in_core[27]
port 51 nsew signal output
rlabel metal2 s 14094 10200 14150 11400 6 la_data_in_core[28]
port 52 nsew signal output
rlabel metal2 s 14554 10200 14610 11400 6 la_data_in_core[29]
port 53 nsew signal output
rlabel metal2 s 2778 10200 2834 11400 6 la_data_in_core[2]
port 54 nsew signal output
rlabel metal2 s 15014 10200 15070 11400 6 la_data_in_core[30]
port 55 nsew signal output
rlabel metal2 s 15382 10200 15438 11400 6 la_data_in_core[31]
port 56 nsew signal output
rlabel metal2 s 15842 10200 15898 11400 6 la_data_in_core[32]
port 57 nsew signal output
rlabel metal2 s 16302 10200 16358 11400 6 la_data_in_core[33]
port 58 nsew signal output
rlabel metal2 s 16670 10200 16726 11400 6 la_data_in_core[34]
port 59 nsew signal output
rlabel metal2 s 17130 10200 17186 11400 6 la_data_in_core[35]
port 60 nsew signal output
rlabel metal2 s 17590 10200 17646 11400 6 la_data_in_core[36]
port 61 nsew signal output
rlabel metal2 s 18050 10200 18106 11400 6 la_data_in_core[37]
port 62 nsew signal output
rlabel metal2 s 18418 10200 18474 11400 6 la_data_in_core[38]
port 63 nsew signal output
rlabel metal2 s 18878 10200 18934 11400 6 la_data_in_core[39]
port 64 nsew signal output
rlabel metal2 s 3238 10200 3294 11400 6 la_data_in_core[3]
port 65 nsew signal output
rlabel metal2 s 19338 10200 19394 11400 6 la_data_in_core[40]
port 66 nsew signal output
rlabel metal2 s 19798 10200 19854 11400 6 la_data_in_core[41]
port 67 nsew signal output
rlabel metal2 s 20166 10200 20222 11400 6 la_data_in_core[42]
port 68 nsew signal output
rlabel metal2 s 20626 10200 20682 11400 6 la_data_in_core[43]
port 69 nsew signal output
rlabel metal2 s 21086 10200 21142 11400 6 la_data_in_core[44]
port 70 nsew signal output
rlabel metal2 s 21546 10200 21602 11400 6 la_data_in_core[45]
port 71 nsew signal output
rlabel metal2 s 21914 10200 21970 11400 6 la_data_in_core[46]
port 72 nsew signal output
rlabel metal2 s 22374 10200 22430 11400 6 la_data_in_core[47]
port 73 nsew signal output
rlabel metal2 s 22834 10200 22890 11400 6 la_data_in_core[48]
port 74 nsew signal output
rlabel metal2 s 23294 10200 23350 11400 6 la_data_in_core[49]
port 75 nsew signal output
rlabel metal2 s 3606 10200 3662 11400 6 la_data_in_core[4]
port 76 nsew signal output
rlabel metal2 s 23662 10200 23718 11400 6 la_data_in_core[50]
port 77 nsew signal output
rlabel metal2 s 24122 10200 24178 11400 6 la_data_in_core[51]
port 78 nsew signal output
rlabel metal2 s 24582 10200 24638 11400 6 la_data_in_core[52]
port 79 nsew signal output
rlabel metal2 s 24950 10200 25006 11400 6 la_data_in_core[53]
port 80 nsew signal output
rlabel metal2 s 25410 10200 25466 11400 6 la_data_in_core[54]
port 81 nsew signal output
rlabel metal2 s 25870 10200 25926 11400 6 la_data_in_core[55]
port 82 nsew signal output
rlabel metal2 s 26330 10200 26386 11400 6 la_data_in_core[56]
port 83 nsew signal output
rlabel metal2 s 26698 10200 26754 11400 6 la_data_in_core[57]
port 84 nsew signal output
rlabel metal2 s 27158 10200 27214 11400 6 la_data_in_core[58]
port 85 nsew signal output
rlabel metal2 s 27618 10200 27674 11400 6 la_data_in_core[59]
port 86 nsew signal output
rlabel metal2 s 4066 10200 4122 11400 6 la_data_in_core[5]
port 87 nsew signal output
rlabel metal2 s 28078 10200 28134 11400 6 la_data_in_core[60]
port 88 nsew signal output
rlabel metal2 s 28446 10200 28502 11400 6 la_data_in_core[61]
port 89 nsew signal output
rlabel metal2 s 28906 10200 28962 11400 6 la_data_in_core[62]
port 90 nsew signal output
rlabel metal2 s 29366 10200 29422 11400 6 la_data_in_core[63]
port 91 nsew signal output
rlabel metal2 s 29826 10200 29882 11400 6 la_data_in_core[64]
port 92 nsew signal output
rlabel metal2 s 30194 10200 30250 11400 6 la_data_in_core[65]
port 93 nsew signal output
rlabel metal2 s 30654 10200 30710 11400 6 la_data_in_core[66]
port 94 nsew signal output
rlabel metal2 s 31114 10200 31170 11400 6 la_data_in_core[67]
port 95 nsew signal output
rlabel metal2 s 31574 10200 31630 11400 6 la_data_in_core[68]
port 96 nsew signal output
rlabel metal2 s 31942 10200 31998 11400 6 la_data_in_core[69]
port 97 nsew signal output
rlabel metal2 s 4526 10200 4582 11400 6 la_data_in_core[6]
port 98 nsew signal output
rlabel metal2 s 32402 10200 32458 11400 6 la_data_in_core[70]
port 99 nsew signal output
rlabel metal2 s 32862 10200 32918 11400 6 la_data_in_core[71]
port 100 nsew signal output
rlabel metal2 s 33230 10200 33286 11400 6 la_data_in_core[72]
port 101 nsew signal output
rlabel metal2 s 33690 10200 33746 11400 6 la_data_in_core[73]
port 102 nsew signal output
rlabel metal2 s 34150 10200 34206 11400 6 la_data_in_core[74]
port 103 nsew signal output
rlabel metal2 s 34610 10200 34666 11400 6 la_data_in_core[75]
port 104 nsew signal output
rlabel metal2 s 34978 10200 35034 11400 6 la_data_in_core[76]
port 105 nsew signal output
rlabel metal2 s 35438 10200 35494 11400 6 la_data_in_core[77]
port 106 nsew signal output
rlabel metal2 s 35898 10200 35954 11400 6 la_data_in_core[78]
port 107 nsew signal output
rlabel metal2 s 36358 10200 36414 11400 6 la_data_in_core[79]
port 108 nsew signal output
rlabel metal2 s 4986 10200 5042 11400 6 la_data_in_core[7]
port 109 nsew signal output
rlabel metal2 s 36726 10200 36782 11400 6 la_data_in_core[80]
port 110 nsew signal output
rlabel metal2 s 37186 10200 37242 11400 6 la_data_in_core[81]
port 111 nsew signal output
rlabel metal2 s 37646 10200 37702 11400 6 la_data_in_core[82]
port 112 nsew signal output
rlabel metal2 s 38106 10200 38162 11400 6 la_data_in_core[83]
port 113 nsew signal output
rlabel metal2 s 38474 10200 38530 11400 6 la_data_in_core[84]
port 114 nsew signal output
rlabel metal2 s 38934 10200 38990 11400 6 la_data_in_core[85]
port 115 nsew signal output
rlabel metal2 s 39394 10200 39450 11400 6 la_data_in_core[86]
port 116 nsew signal output
rlabel metal2 s 39854 10200 39910 11400 6 la_data_in_core[87]
port 117 nsew signal output
rlabel metal2 s 40222 10200 40278 11400 6 la_data_in_core[88]
port 118 nsew signal output
rlabel metal2 s 40682 10200 40738 11400 6 la_data_in_core[89]
port 119 nsew signal output
rlabel metal2 s 5354 10200 5410 11400 6 la_data_in_core[8]
port 120 nsew signal output
rlabel metal2 s 41142 10200 41198 11400 6 la_data_in_core[90]
port 121 nsew signal output
rlabel metal2 s 41510 10200 41566 11400 6 la_data_in_core[91]
port 122 nsew signal output
rlabel metal2 s 41970 10200 42026 11400 6 la_data_in_core[92]
port 123 nsew signal output
rlabel metal2 s 42430 10200 42486 11400 6 la_data_in_core[93]
port 124 nsew signal output
rlabel metal2 s 42890 10200 42946 11400 6 la_data_in_core[94]
port 125 nsew signal output
rlabel metal2 s 43258 10200 43314 11400 6 la_data_in_core[95]
port 126 nsew signal output
rlabel metal2 s 43718 10200 43774 11400 6 la_data_in_core[96]
port 127 nsew signal output
rlabel metal2 s 44178 10200 44234 11400 6 la_data_in_core[97]
port 128 nsew signal output
rlabel metal2 s 44638 10200 44694 11400 6 la_data_in_core[98]
port 129 nsew signal output
rlabel metal2 s 45006 10200 45062 11400 6 la_data_in_core[99]
port 130 nsew signal output
rlabel metal2 s 5814 10200 5870 11400 6 la_data_in_core[9]
port 131 nsew signal output
rlabel metal2 s 55954 -400 56010 800 6 la_data_in_mprj[0]
port 132 nsew signal output
rlabel metal2 s 99470 -400 99526 800 6 la_data_in_mprj[100]
port 133 nsew signal output
rlabel metal2 s 99930 -400 99986 800 6 la_data_in_mprj[101]
port 134 nsew signal output
rlabel metal2 s 100390 -400 100446 800 6 la_data_in_mprj[102]
port 135 nsew signal output
rlabel metal2 s 100850 -400 100906 800 6 la_data_in_mprj[103]
port 136 nsew signal output
rlabel metal2 s 101218 -400 101274 800 6 la_data_in_mprj[104]
port 137 nsew signal output
rlabel metal2 s 101678 -400 101734 800 6 la_data_in_mprj[105]
port 138 nsew signal output
rlabel metal2 s 102138 -400 102194 800 6 la_data_in_mprj[106]
port 139 nsew signal output
rlabel metal2 s 102598 -400 102654 800 6 la_data_in_mprj[107]
port 140 nsew signal output
rlabel metal2 s 102966 -400 103022 800 6 la_data_in_mprj[108]
port 141 nsew signal output
rlabel metal2 s 103426 -400 103482 800 6 la_data_in_mprj[109]
port 142 nsew signal output
rlabel metal2 s 60278 -400 60334 800 6 la_data_in_mprj[10]
port 143 nsew signal output
rlabel metal2 s 103886 -400 103942 800 6 la_data_in_mprj[110]
port 144 nsew signal output
rlabel metal2 s 104254 -400 104310 800 6 la_data_in_mprj[111]
port 145 nsew signal output
rlabel metal2 s 104714 -400 104770 800 6 la_data_in_mprj[112]
port 146 nsew signal output
rlabel metal2 s 105174 -400 105230 800 6 la_data_in_mprj[113]
port 147 nsew signal output
rlabel metal2 s 105634 -400 105690 800 6 la_data_in_mprj[114]
port 148 nsew signal output
rlabel metal2 s 106002 -400 106058 800 6 la_data_in_mprj[115]
port 149 nsew signal output
rlabel metal2 s 106462 -400 106518 800 6 la_data_in_mprj[116]
port 150 nsew signal output
rlabel metal2 s 106922 -400 106978 800 6 la_data_in_mprj[117]
port 151 nsew signal output
rlabel metal2 s 107382 -400 107438 800 6 la_data_in_mprj[118]
port 152 nsew signal output
rlabel metal2 s 107750 -400 107806 800 6 la_data_in_mprj[119]
port 153 nsew signal output
rlabel metal2 s 60738 -400 60794 800 6 la_data_in_mprj[11]
port 154 nsew signal output
rlabel metal2 s 108210 -400 108266 800 6 la_data_in_mprj[120]
port 155 nsew signal output
rlabel metal2 s 108670 -400 108726 800 6 la_data_in_mprj[121]
port 156 nsew signal output
rlabel metal2 s 109130 -400 109186 800 6 la_data_in_mprj[122]
port 157 nsew signal output
rlabel metal2 s 109498 -400 109554 800 6 la_data_in_mprj[123]
port 158 nsew signal output
rlabel metal2 s 109958 -400 110014 800 6 la_data_in_mprj[124]
port 159 nsew signal output
rlabel metal2 s 110418 -400 110474 800 6 la_data_in_mprj[125]
port 160 nsew signal output
rlabel metal2 s 110878 -400 110934 800 6 la_data_in_mprj[126]
port 161 nsew signal output
rlabel metal2 s 111246 -400 111302 800 6 la_data_in_mprj[127]
port 162 nsew signal output
rlabel metal2 s 61198 -400 61254 800 6 la_data_in_mprj[12]
port 163 nsew signal output
rlabel metal2 s 61566 -400 61622 800 6 la_data_in_mprj[13]
port 164 nsew signal output
rlabel metal2 s 62026 -400 62082 800 6 la_data_in_mprj[14]
port 165 nsew signal output
rlabel metal2 s 62486 -400 62542 800 6 la_data_in_mprj[15]
port 166 nsew signal output
rlabel metal2 s 62946 -400 63002 800 6 la_data_in_mprj[16]
port 167 nsew signal output
rlabel metal2 s 63314 -400 63370 800 6 la_data_in_mprj[17]
port 168 nsew signal output
rlabel metal2 s 63774 -400 63830 800 6 la_data_in_mprj[18]
port 169 nsew signal output
rlabel metal2 s 64234 -400 64290 800 6 la_data_in_mprj[19]
port 170 nsew signal output
rlabel metal2 s 56322 -400 56378 800 6 la_data_in_mprj[1]
port 171 nsew signal output
rlabel metal2 s 64602 -400 64658 800 6 la_data_in_mprj[20]
port 172 nsew signal output
rlabel metal2 s 65062 -400 65118 800 6 la_data_in_mprj[21]
port 173 nsew signal output
rlabel metal2 s 65522 -400 65578 800 6 la_data_in_mprj[22]
port 174 nsew signal output
rlabel metal2 s 65982 -400 66038 800 6 la_data_in_mprj[23]
port 175 nsew signal output
rlabel metal2 s 66350 -400 66406 800 6 la_data_in_mprj[24]
port 176 nsew signal output
rlabel metal2 s 66810 -400 66866 800 6 la_data_in_mprj[25]
port 177 nsew signal output
rlabel metal2 s 67270 -400 67326 800 6 la_data_in_mprj[26]
port 178 nsew signal output
rlabel metal2 s 67730 -400 67786 800 6 la_data_in_mprj[27]
port 179 nsew signal output
rlabel metal2 s 68098 -400 68154 800 6 la_data_in_mprj[28]
port 180 nsew signal output
rlabel metal2 s 68558 -400 68614 800 6 la_data_in_mprj[29]
port 181 nsew signal output
rlabel metal2 s 56782 -400 56838 800 6 la_data_in_mprj[2]
port 182 nsew signal output
rlabel metal2 s 69018 -400 69074 800 6 la_data_in_mprj[30]
port 183 nsew signal output
rlabel metal2 s 69478 -400 69534 800 6 la_data_in_mprj[31]
port 184 nsew signal output
rlabel metal2 s 69846 -400 69902 800 6 la_data_in_mprj[32]
port 185 nsew signal output
rlabel metal2 s 70306 -400 70362 800 6 la_data_in_mprj[33]
port 186 nsew signal output
rlabel metal2 s 70766 -400 70822 800 6 la_data_in_mprj[34]
port 187 nsew signal output
rlabel metal2 s 71226 -400 71282 800 6 la_data_in_mprj[35]
port 188 nsew signal output
rlabel metal2 s 71594 -400 71650 800 6 la_data_in_mprj[36]
port 189 nsew signal output
rlabel metal2 s 72054 -400 72110 800 6 la_data_in_mprj[37]
port 190 nsew signal output
rlabel metal2 s 72514 -400 72570 800 6 la_data_in_mprj[38]
port 191 nsew signal output
rlabel metal2 s 72882 -400 72938 800 6 la_data_in_mprj[39]
port 192 nsew signal output
rlabel metal2 s 57242 -400 57298 800 6 la_data_in_mprj[3]
port 193 nsew signal output
rlabel metal2 s 73342 -400 73398 800 6 la_data_in_mprj[40]
port 194 nsew signal output
rlabel metal2 s 73802 -400 73858 800 6 la_data_in_mprj[41]
port 195 nsew signal output
rlabel metal2 s 74262 -400 74318 800 6 la_data_in_mprj[42]
port 196 nsew signal output
rlabel metal2 s 74630 -400 74686 800 6 la_data_in_mprj[43]
port 197 nsew signal output
rlabel metal2 s 75090 -400 75146 800 6 la_data_in_mprj[44]
port 198 nsew signal output
rlabel metal2 s 75550 -400 75606 800 6 la_data_in_mprj[45]
port 199 nsew signal output
rlabel metal2 s 76010 -400 76066 800 6 la_data_in_mprj[46]
port 200 nsew signal output
rlabel metal2 s 76378 -400 76434 800 6 la_data_in_mprj[47]
port 201 nsew signal output
rlabel metal2 s 76838 -400 76894 800 6 la_data_in_mprj[48]
port 202 nsew signal output
rlabel metal2 s 77298 -400 77354 800 6 la_data_in_mprj[49]
port 203 nsew signal output
rlabel metal2 s 57702 -400 57758 800 6 la_data_in_mprj[4]
port 204 nsew signal output
rlabel metal2 s 77758 -400 77814 800 6 la_data_in_mprj[50]
port 205 nsew signal output
rlabel metal2 s 78126 -400 78182 800 6 la_data_in_mprj[51]
port 206 nsew signal output
rlabel metal2 s 78586 -400 78642 800 6 la_data_in_mprj[52]
port 207 nsew signal output
rlabel metal2 s 79046 -400 79102 800 6 la_data_in_mprj[53]
port 208 nsew signal output
rlabel metal2 s 79506 -400 79562 800 6 la_data_in_mprj[54]
port 209 nsew signal output
rlabel metal2 s 79874 -400 79930 800 6 la_data_in_mprj[55]
port 210 nsew signal output
rlabel metal2 s 80334 -400 80390 800 6 la_data_in_mprj[56]
port 211 nsew signal output
rlabel metal2 s 80794 -400 80850 800 6 la_data_in_mprj[57]
port 212 nsew signal output
rlabel metal2 s 81162 -400 81218 800 6 la_data_in_mprj[58]
port 213 nsew signal output
rlabel metal2 s 81622 -400 81678 800 6 la_data_in_mprj[59]
port 214 nsew signal output
rlabel metal2 s 58070 -400 58126 800 6 la_data_in_mprj[5]
port 215 nsew signal output
rlabel metal2 s 82082 -400 82138 800 6 la_data_in_mprj[60]
port 216 nsew signal output
rlabel metal2 s 82542 -400 82598 800 6 la_data_in_mprj[61]
port 217 nsew signal output
rlabel metal2 s 82910 -400 82966 800 6 la_data_in_mprj[62]
port 218 nsew signal output
rlabel metal2 s 83370 -400 83426 800 6 la_data_in_mprj[63]
port 219 nsew signal output
rlabel metal2 s 83830 -400 83886 800 6 la_data_in_mprj[64]
port 220 nsew signal output
rlabel metal2 s 84290 -400 84346 800 6 la_data_in_mprj[65]
port 221 nsew signal output
rlabel metal2 s 84658 -400 84714 800 6 la_data_in_mprj[66]
port 222 nsew signal output
rlabel metal2 s 85118 -400 85174 800 6 la_data_in_mprj[67]
port 223 nsew signal output
rlabel metal2 s 85578 -400 85634 800 6 la_data_in_mprj[68]
port 224 nsew signal output
rlabel metal2 s 86038 -400 86094 800 6 la_data_in_mprj[69]
port 225 nsew signal output
rlabel metal2 s 58530 -400 58586 800 6 la_data_in_mprj[6]
port 226 nsew signal output
rlabel metal2 s 86406 -400 86462 800 6 la_data_in_mprj[70]
port 227 nsew signal output
rlabel metal2 s 86866 -400 86922 800 6 la_data_in_mprj[71]
port 228 nsew signal output
rlabel metal2 s 87326 -400 87382 800 6 la_data_in_mprj[72]
port 229 nsew signal output
rlabel metal2 s 87786 -400 87842 800 6 la_data_in_mprj[73]
port 230 nsew signal output
rlabel metal2 s 88154 -400 88210 800 6 la_data_in_mprj[74]
port 231 nsew signal output
rlabel metal2 s 88614 -400 88670 800 6 la_data_in_mprj[75]
port 232 nsew signal output
rlabel metal2 s 89074 -400 89130 800 6 la_data_in_mprj[76]
port 233 nsew signal output
rlabel metal2 s 89442 -400 89498 800 6 la_data_in_mprj[77]
port 234 nsew signal output
rlabel metal2 s 89902 -400 89958 800 6 la_data_in_mprj[78]
port 235 nsew signal output
rlabel metal2 s 90362 -400 90418 800 6 la_data_in_mprj[79]
port 236 nsew signal output
rlabel metal2 s 58990 -400 59046 800 6 la_data_in_mprj[7]
port 237 nsew signal output
rlabel metal2 s 90822 -400 90878 800 6 la_data_in_mprj[80]
port 238 nsew signal output
rlabel metal2 s 91190 -400 91246 800 6 la_data_in_mprj[81]
port 239 nsew signal output
rlabel metal2 s 91650 -400 91706 800 6 la_data_in_mprj[82]
port 240 nsew signal output
rlabel metal2 s 92110 -400 92166 800 6 la_data_in_mprj[83]
port 241 nsew signal output
rlabel metal2 s 92570 -400 92626 800 6 la_data_in_mprj[84]
port 242 nsew signal output
rlabel metal2 s 92938 -400 92994 800 6 la_data_in_mprj[85]
port 243 nsew signal output
rlabel metal2 s 93398 -400 93454 800 6 la_data_in_mprj[86]
port 244 nsew signal output
rlabel metal2 s 93858 -400 93914 800 6 la_data_in_mprj[87]
port 245 nsew signal output
rlabel metal2 s 94318 -400 94374 800 6 la_data_in_mprj[88]
port 246 nsew signal output
rlabel metal2 s 94686 -400 94742 800 6 la_data_in_mprj[89]
port 247 nsew signal output
rlabel metal2 s 59450 -400 59506 800 6 la_data_in_mprj[8]
port 248 nsew signal output
rlabel metal2 s 95146 -400 95202 800 6 la_data_in_mprj[90]
port 249 nsew signal output
rlabel metal2 s 95606 -400 95662 800 6 la_data_in_mprj[91]
port 250 nsew signal output
rlabel metal2 s 96066 -400 96122 800 6 la_data_in_mprj[92]
port 251 nsew signal output
rlabel metal2 s 96434 -400 96490 800 6 la_data_in_mprj[93]
port 252 nsew signal output
rlabel metal2 s 96894 -400 96950 800 6 la_data_in_mprj[94]
port 253 nsew signal output
rlabel metal2 s 97354 -400 97410 800 6 la_data_in_mprj[95]
port 254 nsew signal output
rlabel metal2 s 97722 -400 97778 800 6 la_data_in_mprj[96]
port 255 nsew signal output
rlabel metal2 s 98182 -400 98238 800 6 la_data_in_mprj[97]
port 256 nsew signal output
rlabel metal2 s 98642 -400 98698 800 6 la_data_in_mprj[98]
port 257 nsew signal output
rlabel metal2 s 99102 -400 99158 800 6 la_data_in_mprj[99]
port 258 nsew signal output
rlabel metal2 s 59818 -400 59874 800 6 la_data_in_mprj[9]
port 259 nsew signal output
rlabel metal2 s 57702 10200 57758 11400 6 la_data_out_core[0]
port 260 nsew signal input
rlabel metal2 s 101218 10200 101274 11400 6 la_data_out_core[100]
port 261 nsew signal input
rlabel metal2 s 101678 10200 101734 11400 6 la_data_out_core[101]
port 262 nsew signal input
rlabel metal2 s 102138 10200 102194 11400 6 la_data_out_core[102]
port 263 nsew signal input
rlabel metal2 s 102598 10200 102654 11400 6 la_data_out_core[103]
port 264 nsew signal input
rlabel metal2 s 102966 10200 103022 11400 6 la_data_out_core[104]
port 265 nsew signal input
rlabel metal2 s 103426 10200 103482 11400 6 la_data_out_core[105]
port 266 nsew signal input
rlabel metal2 s 103886 10200 103942 11400 6 la_data_out_core[106]
port 267 nsew signal input
rlabel metal2 s 104254 10200 104310 11400 6 la_data_out_core[107]
port 268 nsew signal input
rlabel metal2 s 104714 10200 104770 11400 6 la_data_out_core[108]
port 269 nsew signal input
rlabel metal2 s 105174 10200 105230 11400 6 la_data_out_core[109]
port 270 nsew signal input
rlabel metal2 s 62026 10200 62082 11400 6 la_data_out_core[10]
port 271 nsew signal input
rlabel metal2 s 105634 10200 105690 11400 6 la_data_out_core[110]
port 272 nsew signal input
rlabel metal2 s 106002 10200 106058 11400 6 la_data_out_core[111]
port 273 nsew signal input
rlabel metal2 s 106462 10200 106518 11400 6 la_data_out_core[112]
port 274 nsew signal input
rlabel metal2 s 106922 10200 106978 11400 6 la_data_out_core[113]
port 275 nsew signal input
rlabel metal2 s 107382 10200 107438 11400 6 la_data_out_core[114]
port 276 nsew signal input
rlabel metal2 s 107750 10200 107806 11400 6 la_data_out_core[115]
port 277 nsew signal input
rlabel metal2 s 108210 10200 108266 11400 6 la_data_out_core[116]
port 278 nsew signal input
rlabel metal2 s 108670 10200 108726 11400 6 la_data_out_core[117]
port 279 nsew signal input
rlabel metal2 s 109130 10200 109186 11400 6 la_data_out_core[118]
port 280 nsew signal input
rlabel metal2 s 109498 10200 109554 11400 6 la_data_out_core[119]
port 281 nsew signal input
rlabel metal2 s 62486 10200 62542 11400 6 la_data_out_core[11]
port 282 nsew signal input
rlabel metal2 s 109958 10200 110014 11400 6 la_data_out_core[120]
port 283 nsew signal input
rlabel metal2 s 110418 10200 110474 11400 6 la_data_out_core[121]
port 284 nsew signal input
rlabel metal2 s 110878 10200 110934 11400 6 la_data_out_core[122]
port 285 nsew signal input
rlabel metal2 s 111246 10200 111302 11400 6 la_data_out_core[123]
port 286 nsew signal input
rlabel metal2 s 111706 10200 111762 11400 6 la_data_out_core[124]
port 287 nsew signal input
rlabel metal2 s 112166 10200 112222 11400 6 la_data_out_core[125]
port 288 nsew signal input
rlabel metal2 s 112534 10200 112590 11400 6 la_data_out_core[126]
port 289 nsew signal input
rlabel metal2 s 112994 10200 113050 11400 6 la_data_out_core[127]
port 290 nsew signal input
rlabel metal2 s 62946 10200 63002 11400 6 la_data_out_core[12]
port 291 nsew signal input
rlabel metal2 s 63314 10200 63370 11400 6 la_data_out_core[13]
port 292 nsew signal input
rlabel metal2 s 63774 10200 63830 11400 6 la_data_out_core[14]
port 293 nsew signal input
rlabel metal2 s 64234 10200 64290 11400 6 la_data_out_core[15]
port 294 nsew signal input
rlabel metal2 s 64602 10200 64658 11400 6 la_data_out_core[16]
port 295 nsew signal input
rlabel metal2 s 65062 10200 65118 11400 6 la_data_out_core[17]
port 296 nsew signal input
rlabel metal2 s 65522 10200 65578 11400 6 la_data_out_core[18]
port 297 nsew signal input
rlabel metal2 s 65982 10200 66038 11400 6 la_data_out_core[19]
port 298 nsew signal input
rlabel metal2 s 58070 10200 58126 11400 6 la_data_out_core[1]
port 299 nsew signal input
rlabel metal2 s 66350 10200 66406 11400 6 la_data_out_core[20]
port 300 nsew signal input
rlabel metal2 s 66810 10200 66866 11400 6 la_data_out_core[21]
port 301 nsew signal input
rlabel metal2 s 67270 10200 67326 11400 6 la_data_out_core[22]
port 302 nsew signal input
rlabel metal2 s 67730 10200 67786 11400 6 la_data_out_core[23]
port 303 nsew signal input
rlabel metal2 s 68098 10200 68154 11400 6 la_data_out_core[24]
port 304 nsew signal input
rlabel metal2 s 68558 10200 68614 11400 6 la_data_out_core[25]
port 305 nsew signal input
rlabel metal2 s 69018 10200 69074 11400 6 la_data_out_core[26]
port 306 nsew signal input
rlabel metal2 s 69478 10200 69534 11400 6 la_data_out_core[27]
port 307 nsew signal input
rlabel metal2 s 69846 10200 69902 11400 6 la_data_out_core[28]
port 308 nsew signal input
rlabel metal2 s 70306 10200 70362 11400 6 la_data_out_core[29]
port 309 nsew signal input
rlabel metal2 s 58530 10200 58586 11400 6 la_data_out_core[2]
port 310 nsew signal input
rlabel metal2 s 70766 10200 70822 11400 6 la_data_out_core[30]
port 311 nsew signal input
rlabel metal2 s 71226 10200 71282 11400 6 la_data_out_core[31]
port 312 nsew signal input
rlabel metal2 s 71594 10200 71650 11400 6 la_data_out_core[32]
port 313 nsew signal input
rlabel metal2 s 72054 10200 72110 11400 6 la_data_out_core[33]
port 314 nsew signal input
rlabel metal2 s 72514 10200 72570 11400 6 la_data_out_core[34]
port 315 nsew signal input
rlabel metal2 s 72882 10200 72938 11400 6 la_data_out_core[35]
port 316 nsew signal input
rlabel metal2 s 73342 10200 73398 11400 6 la_data_out_core[36]
port 317 nsew signal input
rlabel metal2 s 73802 10200 73858 11400 6 la_data_out_core[37]
port 318 nsew signal input
rlabel metal2 s 74262 10200 74318 11400 6 la_data_out_core[38]
port 319 nsew signal input
rlabel metal2 s 74630 10200 74686 11400 6 la_data_out_core[39]
port 320 nsew signal input
rlabel metal2 s 58990 10200 59046 11400 6 la_data_out_core[3]
port 321 nsew signal input
rlabel metal2 s 75090 10200 75146 11400 6 la_data_out_core[40]
port 322 nsew signal input
rlabel metal2 s 75550 10200 75606 11400 6 la_data_out_core[41]
port 323 nsew signal input
rlabel metal2 s 76010 10200 76066 11400 6 la_data_out_core[42]
port 324 nsew signal input
rlabel metal2 s 76378 10200 76434 11400 6 la_data_out_core[43]
port 325 nsew signal input
rlabel metal2 s 76838 10200 76894 11400 6 la_data_out_core[44]
port 326 nsew signal input
rlabel metal2 s 77298 10200 77354 11400 6 la_data_out_core[45]
port 327 nsew signal input
rlabel metal2 s 77758 10200 77814 11400 6 la_data_out_core[46]
port 328 nsew signal input
rlabel metal2 s 78126 10200 78182 11400 6 la_data_out_core[47]
port 329 nsew signal input
rlabel metal2 s 78586 10200 78642 11400 6 la_data_out_core[48]
port 330 nsew signal input
rlabel metal2 s 79046 10200 79102 11400 6 la_data_out_core[49]
port 331 nsew signal input
rlabel metal2 s 59450 10200 59506 11400 6 la_data_out_core[4]
port 332 nsew signal input
rlabel metal2 s 79506 10200 79562 11400 6 la_data_out_core[50]
port 333 nsew signal input
rlabel metal2 s 79874 10200 79930 11400 6 la_data_out_core[51]
port 334 nsew signal input
rlabel metal2 s 80334 10200 80390 11400 6 la_data_out_core[52]
port 335 nsew signal input
rlabel metal2 s 80794 10200 80850 11400 6 la_data_out_core[53]
port 336 nsew signal input
rlabel metal2 s 81162 10200 81218 11400 6 la_data_out_core[54]
port 337 nsew signal input
rlabel metal2 s 81622 10200 81678 11400 6 la_data_out_core[55]
port 338 nsew signal input
rlabel metal2 s 82082 10200 82138 11400 6 la_data_out_core[56]
port 339 nsew signal input
rlabel metal2 s 82542 10200 82598 11400 6 la_data_out_core[57]
port 340 nsew signal input
rlabel metal2 s 82910 10200 82966 11400 6 la_data_out_core[58]
port 341 nsew signal input
rlabel metal2 s 83370 10200 83426 11400 6 la_data_out_core[59]
port 342 nsew signal input
rlabel metal2 s 59818 10200 59874 11400 6 la_data_out_core[5]
port 343 nsew signal input
rlabel metal2 s 83830 10200 83886 11400 6 la_data_out_core[60]
port 344 nsew signal input
rlabel metal2 s 84290 10200 84346 11400 6 la_data_out_core[61]
port 345 nsew signal input
rlabel metal2 s 84658 10200 84714 11400 6 la_data_out_core[62]
port 346 nsew signal input
rlabel metal2 s 85118 10200 85174 11400 6 la_data_out_core[63]
port 347 nsew signal input
rlabel metal2 s 85578 10200 85634 11400 6 la_data_out_core[64]
port 348 nsew signal input
rlabel metal2 s 86038 10200 86094 11400 6 la_data_out_core[65]
port 349 nsew signal input
rlabel metal2 s 86406 10200 86462 11400 6 la_data_out_core[66]
port 350 nsew signal input
rlabel metal2 s 86866 10200 86922 11400 6 la_data_out_core[67]
port 351 nsew signal input
rlabel metal2 s 87326 10200 87382 11400 6 la_data_out_core[68]
port 352 nsew signal input
rlabel metal2 s 87786 10200 87842 11400 6 la_data_out_core[69]
port 353 nsew signal input
rlabel metal2 s 60278 10200 60334 11400 6 la_data_out_core[6]
port 354 nsew signal input
rlabel metal2 s 88154 10200 88210 11400 6 la_data_out_core[70]
port 355 nsew signal input
rlabel metal2 s 88614 10200 88670 11400 6 la_data_out_core[71]
port 356 nsew signal input
rlabel metal2 s 89074 10200 89130 11400 6 la_data_out_core[72]
port 357 nsew signal input
rlabel metal2 s 89442 10200 89498 11400 6 la_data_out_core[73]
port 358 nsew signal input
rlabel metal2 s 89902 10200 89958 11400 6 la_data_out_core[74]
port 359 nsew signal input
rlabel metal2 s 90362 10200 90418 11400 6 la_data_out_core[75]
port 360 nsew signal input
rlabel metal2 s 90822 10200 90878 11400 6 la_data_out_core[76]
port 361 nsew signal input
rlabel metal2 s 91190 10200 91246 11400 6 la_data_out_core[77]
port 362 nsew signal input
rlabel metal2 s 91650 10200 91706 11400 6 la_data_out_core[78]
port 363 nsew signal input
rlabel metal2 s 92110 10200 92166 11400 6 la_data_out_core[79]
port 364 nsew signal input
rlabel metal2 s 60738 10200 60794 11400 6 la_data_out_core[7]
port 365 nsew signal input
rlabel metal2 s 92570 10200 92626 11400 6 la_data_out_core[80]
port 366 nsew signal input
rlabel metal2 s 92938 10200 92994 11400 6 la_data_out_core[81]
port 367 nsew signal input
rlabel metal2 s 93398 10200 93454 11400 6 la_data_out_core[82]
port 368 nsew signal input
rlabel metal2 s 93858 10200 93914 11400 6 la_data_out_core[83]
port 369 nsew signal input
rlabel metal2 s 94318 10200 94374 11400 6 la_data_out_core[84]
port 370 nsew signal input
rlabel metal2 s 94686 10200 94742 11400 6 la_data_out_core[85]
port 371 nsew signal input
rlabel metal2 s 95146 10200 95202 11400 6 la_data_out_core[86]
port 372 nsew signal input
rlabel metal2 s 95606 10200 95662 11400 6 la_data_out_core[87]
port 373 nsew signal input
rlabel metal2 s 96066 10200 96122 11400 6 la_data_out_core[88]
port 374 nsew signal input
rlabel metal2 s 96434 10200 96490 11400 6 la_data_out_core[89]
port 375 nsew signal input
rlabel metal2 s 61198 10200 61254 11400 6 la_data_out_core[8]
port 376 nsew signal input
rlabel metal2 s 96894 10200 96950 11400 6 la_data_out_core[90]
port 377 nsew signal input
rlabel metal2 s 97354 10200 97410 11400 6 la_data_out_core[91]
port 378 nsew signal input
rlabel metal2 s 97722 10200 97778 11400 6 la_data_out_core[92]
port 379 nsew signal input
rlabel metal2 s 98182 10200 98238 11400 6 la_data_out_core[93]
port 380 nsew signal input
rlabel metal2 s 98642 10200 98698 11400 6 la_data_out_core[94]
port 381 nsew signal input
rlabel metal2 s 99102 10200 99158 11400 6 la_data_out_core[95]
port 382 nsew signal input
rlabel metal2 s 99470 10200 99526 11400 6 la_data_out_core[96]
port 383 nsew signal input
rlabel metal2 s 99930 10200 99986 11400 6 la_data_out_core[97]
port 384 nsew signal input
rlabel metal2 s 100390 10200 100446 11400 6 la_data_out_core[98]
port 385 nsew signal input
rlabel metal2 s 100850 10200 100906 11400 6 la_data_out_core[99]
port 386 nsew signal input
rlabel metal2 s 61566 10200 61622 11400 6 la_data_out_core[9]
port 387 nsew signal input
rlabel metal2 s 202 -400 258 800 6 la_data_out_mprj[0]
port 388 nsew signal input
rlabel metal2 s 43718 -400 43774 800 6 la_data_out_mprj[100]
port 389 nsew signal input
rlabel metal2 s 44178 -400 44234 800 6 la_data_out_mprj[101]
port 390 nsew signal input
rlabel metal2 s 44638 -400 44694 800 6 la_data_out_mprj[102]
port 391 nsew signal input
rlabel metal2 s 45006 -400 45062 800 6 la_data_out_mprj[103]
port 392 nsew signal input
rlabel metal2 s 45466 -400 45522 800 6 la_data_out_mprj[104]
port 393 nsew signal input
rlabel metal2 s 45926 -400 45982 800 6 la_data_out_mprj[105]
port 394 nsew signal input
rlabel metal2 s 46386 -400 46442 800 6 la_data_out_mprj[106]
port 395 nsew signal input
rlabel metal2 s 46754 -400 46810 800 6 la_data_out_mprj[107]
port 396 nsew signal input
rlabel metal2 s 47214 -400 47270 800 6 la_data_out_mprj[108]
port 397 nsew signal input
rlabel metal2 s 47674 -400 47730 800 6 la_data_out_mprj[109]
port 398 nsew signal input
rlabel metal2 s 4526 -400 4582 800 6 la_data_out_mprj[10]
port 399 nsew signal input
rlabel metal2 s 48134 -400 48190 800 6 la_data_out_mprj[110]
port 400 nsew signal input
rlabel metal2 s 48502 -400 48558 800 6 la_data_out_mprj[111]
port 401 nsew signal input
rlabel metal2 s 48962 -400 49018 800 6 la_data_out_mprj[112]
port 402 nsew signal input
rlabel metal2 s 49422 -400 49478 800 6 la_data_out_mprj[113]
port 403 nsew signal input
rlabel metal2 s 49790 -400 49846 800 6 la_data_out_mprj[114]
port 404 nsew signal input
rlabel metal2 s 50250 -400 50306 800 6 la_data_out_mprj[115]
port 405 nsew signal input
rlabel metal2 s 50710 -400 50766 800 6 la_data_out_mprj[116]
port 406 nsew signal input
rlabel metal2 s 51170 -400 51226 800 6 la_data_out_mprj[117]
port 407 nsew signal input
rlabel metal2 s 51538 -400 51594 800 6 la_data_out_mprj[118]
port 408 nsew signal input
rlabel metal2 s 51998 -400 52054 800 6 la_data_out_mprj[119]
port 409 nsew signal input
rlabel metal2 s 4986 -400 5042 800 6 la_data_out_mprj[11]
port 410 nsew signal input
rlabel metal2 s 52458 -400 52514 800 6 la_data_out_mprj[120]
port 411 nsew signal input
rlabel metal2 s 52918 -400 52974 800 6 la_data_out_mprj[121]
port 412 nsew signal input
rlabel metal2 s 53286 -400 53342 800 6 la_data_out_mprj[122]
port 413 nsew signal input
rlabel metal2 s 53746 -400 53802 800 6 la_data_out_mprj[123]
port 414 nsew signal input
rlabel metal2 s 54206 -400 54262 800 6 la_data_out_mprj[124]
port 415 nsew signal input
rlabel metal2 s 54666 -400 54722 800 6 la_data_out_mprj[125]
port 416 nsew signal input
rlabel metal2 s 55034 -400 55090 800 6 la_data_out_mprj[126]
port 417 nsew signal input
rlabel metal2 s 55494 -400 55550 800 6 la_data_out_mprj[127]
port 418 nsew signal input
rlabel metal2 s 5354 -400 5410 800 6 la_data_out_mprj[12]
port 419 nsew signal input
rlabel metal2 s 5814 -400 5870 800 6 la_data_out_mprj[13]
port 420 nsew signal input
rlabel metal2 s 6274 -400 6330 800 6 la_data_out_mprj[14]
port 421 nsew signal input
rlabel metal2 s 6734 -400 6790 800 6 la_data_out_mprj[15]
port 422 nsew signal input
rlabel metal2 s 7102 -400 7158 800 6 la_data_out_mprj[16]
port 423 nsew signal input
rlabel metal2 s 7562 -400 7618 800 6 la_data_out_mprj[17]
port 424 nsew signal input
rlabel metal2 s 8022 -400 8078 800 6 la_data_out_mprj[18]
port 425 nsew signal input
rlabel metal2 s 8390 -400 8446 800 6 la_data_out_mprj[19]
port 426 nsew signal input
rlabel metal2 s 570 -400 626 800 6 la_data_out_mprj[1]
port 427 nsew signal input
rlabel metal2 s 8850 -400 8906 800 6 la_data_out_mprj[20]
port 428 nsew signal input
rlabel metal2 s 9310 -400 9366 800 6 la_data_out_mprj[21]
port 429 nsew signal input
rlabel metal2 s 9770 -400 9826 800 6 la_data_out_mprj[22]
port 430 nsew signal input
rlabel metal2 s 10138 -400 10194 800 6 la_data_out_mprj[23]
port 431 nsew signal input
rlabel metal2 s 10598 -400 10654 800 6 la_data_out_mprj[24]
port 432 nsew signal input
rlabel metal2 s 11058 -400 11114 800 6 la_data_out_mprj[25]
port 433 nsew signal input
rlabel metal2 s 11518 -400 11574 800 6 la_data_out_mprj[26]
port 434 nsew signal input
rlabel metal2 s 11886 -400 11942 800 6 la_data_out_mprj[27]
port 435 nsew signal input
rlabel metal2 s 12346 -400 12402 800 6 la_data_out_mprj[28]
port 436 nsew signal input
rlabel metal2 s 12806 -400 12862 800 6 la_data_out_mprj[29]
port 437 nsew signal input
rlabel metal2 s 1030 -400 1086 800 6 la_data_out_mprj[2]
port 438 nsew signal input
rlabel metal2 s 13266 -400 13322 800 6 la_data_out_mprj[30]
port 439 nsew signal input
rlabel metal2 s 13634 -400 13690 800 6 la_data_out_mprj[31]
port 440 nsew signal input
rlabel metal2 s 14094 -400 14150 800 6 la_data_out_mprj[32]
port 441 nsew signal input
rlabel metal2 s 14554 -400 14610 800 6 la_data_out_mprj[33]
port 442 nsew signal input
rlabel metal2 s 15014 -400 15070 800 6 la_data_out_mprj[34]
port 443 nsew signal input
rlabel metal2 s 15382 -400 15438 800 6 la_data_out_mprj[35]
port 444 nsew signal input
rlabel metal2 s 15842 -400 15898 800 6 la_data_out_mprj[36]
port 445 nsew signal input
rlabel metal2 s 16302 -400 16358 800 6 la_data_out_mprj[37]
port 446 nsew signal input
rlabel metal2 s 16670 -400 16726 800 6 la_data_out_mprj[38]
port 447 nsew signal input
rlabel metal2 s 17130 -400 17186 800 6 la_data_out_mprj[39]
port 448 nsew signal input
rlabel metal2 s 1490 -400 1546 800 6 la_data_out_mprj[3]
port 449 nsew signal input
rlabel metal2 s 17590 -400 17646 800 6 la_data_out_mprj[40]
port 450 nsew signal input
rlabel metal2 s 18050 -400 18106 800 6 la_data_out_mprj[41]
port 451 nsew signal input
rlabel metal2 s 18418 -400 18474 800 6 la_data_out_mprj[42]
port 452 nsew signal input
rlabel metal2 s 18878 -400 18934 800 6 la_data_out_mprj[43]
port 453 nsew signal input
rlabel metal2 s 19338 -400 19394 800 6 la_data_out_mprj[44]
port 454 nsew signal input
rlabel metal2 s 19798 -400 19854 800 6 la_data_out_mprj[45]
port 455 nsew signal input
rlabel metal2 s 20166 -400 20222 800 6 la_data_out_mprj[46]
port 456 nsew signal input
rlabel metal2 s 20626 -400 20682 800 6 la_data_out_mprj[47]
port 457 nsew signal input
rlabel metal2 s 21086 -400 21142 800 6 la_data_out_mprj[48]
port 458 nsew signal input
rlabel metal2 s 21546 -400 21602 800 6 la_data_out_mprj[49]
port 459 nsew signal input
rlabel metal2 s 1858 -400 1914 800 6 la_data_out_mprj[4]
port 460 nsew signal input
rlabel metal2 s 21914 -400 21970 800 6 la_data_out_mprj[50]
port 461 nsew signal input
rlabel metal2 s 22374 -400 22430 800 6 la_data_out_mprj[51]
port 462 nsew signal input
rlabel metal2 s 22834 -400 22890 800 6 la_data_out_mprj[52]
port 463 nsew signal input
rlabel metal2 s 23294 -400 23350 800 6 la_data_out_mprj[53]
port 464 nsew signal input
rlabel metal2 s 23662 -400 23718 800 6 la_data_out_mprj[54]
port 465 nsew signal input
rlabel metal2 s 24122 -400 24178 800 6 la_data_out_mprj[55]
port 466 nsew signal input
rlabel metal2 s 24582 -400 24638 800 6 la_data_out_mprj[56]
port 467 nsew signal input
rlabel metal2 s 24950 -400 25006 800 6 la_data_out_mprj[57]
port 468 nsew signal input
rlabel metal2 s 25410 -400 25466 800 6 la_data_out_mprj[58]
port 469 nsew signal input
rlabel metal2 s 25870 -400 25926 800 6 la_data_out_mprj[59]
port 470 nsew signal input
rlabel metal2 s 2318 -400 2374 800 6 la_data_out_mprj[5]
port 471 nsew signal input
rlabel metal2 s 26330 -400 26386 800 6 la_data_out_mprj[60]
port 472 nsew signal input
rlabel metal2 s 26698 -400 26754 800 6 la_data_out_mprj[61]
port 473 nsew signal input
rlabel metal2 s 27158 -400 27214 800 6 la_data_out_mprj[62]
port 474 nsew signal input
rlabel metal2 s 27618 -400 27674 800 6 la_data_out_mprj[63]
port 475 nsew signal input
rlabel metal2 s 28078 -400 28134 800 6 la_data_out_mprj[64]
port 476 nsew signal input
rlabel metal2 s 28446 -400 28502 800 6 la_data_out_mprj[65]
port 477 nsew signal input
rlabel metal2 s 28906 -400 28962 800 6 la_data_out_mprj[66]
port 478 nsew signal input
rlabel metal2 s 29366 -400 29422 800 6 la_data_out_mprj[67]
port 479 nsew signal input
rlabel metal2 s 29826 -400 29882 800 6 la_data_out_mprj[68]
port 480 nsew signal input
rlabel metal2 s 30194 -400 30250 800 6 la_data_out_mprj[69]
port 481 nsew signal input
rlabel metal2 s 2778 -400 2834 800 6 la_data_out_mprj[6]
port 482 nsew signal input
rlabel metal2 s 30654 -400 30710 800 6 la_data_out_mprj[70]
port 483 nsew signal input
rlabel metal2 s 31114 -400 31170 800 6 la_data_out_mprj[71]
port 484 nsew signal input
rlabel metal2 s 31574 -400 31630 800 6 la_data_out_mprj[72]
port 485 nsew signal input
rlabel metal2 s 31942 -400 31998 800 6 la_data_out_mprj[73]
port 486 nsew signal input
rlabel metal2 s 32402 -400 32458 800 6 la_data_out_mprj[74]
port 487 nsew signal input
rlabel metal2 s 32862 -400 32918 800 6 la_data_out_mprj[75]
port 488 nsew signal input
rlabel metal2 s 33230 -400 33286 800 6 la_data_out_mprj[76]
port 489 nsew signal input
rlabel metal2 s 33690 -400 33746 800 6 la_data_out_mprj[77]
port 490 nsew signal input
rlabel metal2 s 34150 -400 34206 800 6 la_data_out_mprj[78]
port 491 nsew signal input
rlabel metal2 s 34610 -400 34666 800 6 la_data_out_mprj[79]
port 492 nsew signal input
rlabel metal2 s 3238 -400 3294 800 6 la_data_out_mprj[7]
port 493 nsew signal input
rlabel metal2 s 34978 -400 35034 800 6 la_data_out_mprj[80]
port 494 nsew signal input
rlabel metal2 s 35438 -400 35494 800 6 la_data_out_mprj[81]
port 495 nsew signal input
rlabel metal2 s 35898 -400 35954 800 6 la_data_out_mprj[82]
port 496 nsew signal input
rlabel metal2 s 36358 -400 36414 800 6 la_data_out_mprj[83]
port 497 nsew signal input
rlabel metal2 s 36726 -400 36782 800 6 la_data_out_mprj[84]
port 498 nsew signal input
rlabel metal2 s 37186 -400 37242 800 6 la_data_out_mprj[85]
port 499 nsew signal input
rlabel metal2 s 37646 -400 37702 800 6 la_data_out_mprj[86]
port 500 nsew signal input
rlabel metal2 s 38106 -400 38162 800 6 la_data_out_mprj[87]
port 501 nsew signal input
rlabel metal2 s 38474 -400 38530 800 6 la_data_out_mprj[88]
port 502 nsew signal input
rlabel metal2 s 38934 -400 38990 800 6 la_data_out_mprj[89]
port 503 nsew signal input
rlabel metal2 s 3606 -400 3662 800 6 la_data_out_mprj[8]
port 504 nsew signal input
rlabel metal2 s 39394 -400 39450 800 6 la_data_out_mprj[90]
port 505 nsew signal input
rlabel metal2 s 39854 -400 39910 800 6 la_data_out_mprj[91]
port 506 nsew signal input
rlabel metal2 s 40222 -400 40278 800 6 la_data_out_mprj[92]
port 507 nsew signal input
rlabel metal2 s 40682 -400 40738 800 6 la_data_out_mprj[93]
port 508 nsew signal input
rlabel metal2 s 41142 -400 41198 800 6 la_data_out_mprj[94]
port 509 nsew signal input
rlabel metal2 s 41510 -400 41566 800 6 la_data_out_mprj[95]
port 510 nsew signal input
rlabel metal2 s 41970 -400 42026 800 6 la_data_out_mprj[96]
port 511 nsew signal input
rlabel metal2 s 42430 -400 42486 800 6 la_data_out_mprj[97]
port 512 nsew signal input
rlabel metal2 s 42890 -400 42946 800 6 la_data_out_mprj[98]
port 513 nsew signal input
rlabel metal2 s 43258 -400 43314 800 6 la_data_out_mprj[99]
port 514 nsew signal input
rlabel metal2 s 4066 -400 4122 800 6 la_data_out_mprj[9]
port 515 nsew signal input
rlabel metal2 s 113454 10200 113510 11400 6 la_oen_core[0]
port 516 nsew signal output
rlabel metal2 s 157062 10200 157118 11400 6 la_oen_core[100]
port 517 nsew signal output
rlabel metal2 s 157430 10200 157486 11400 6 la_oen_core[101]
port 518 nsew signal output
rlabel metal2 s 157890 10200 157946 11400 6 la_oen_core[102]
port 519 nsew signal output
rlabel metal2 s 158350 10200 158406 11400 6 la_oen_core[103]
port 520 nsew signal output
rlabel metal2 s 158810 10200 158866 11400 6 la_oen_core[104]
port 521 nsew signal output
rlabel metal2 s 159178 10200 159234 11400 6 la_oen_core[105]
port 522 nsew signal output
rlabel metal2 s 159638 10200 159694 11400 6 la_oen_core[106]
port 523 nsew signal output
rlabel metal2 s 160098 10200 160154 11400 6 la_oen_core[107]
port 524 nsew signal output
rlabel metal2 s 160466 10200 160522 11400 6 la_oen_core[108]
port 525 nsew signal output
rlabel metal2 s 160926 10200 160982 11400 6 la_oen_core[109]
port 526 nsew signal output
rlabel metal2 s 117778 10200 117834 11400 6 la_oen_core[10]
port 527 nsew signal output
rlabel metal2 s 161386 10200 161442 11400 6 la_oen_core[110]
port 528 nsew signal output
rlabel metal2 s 161846 10200 161902 11400 6 la_oen_core[111]
port 529 nsew signal output
rlabel metal2 s 162214 10200 162270 11400 6 la_oen_core[112]
port 530 nsew signal output
rlabel metal2 s 162674 10200 162730 11400 6 la_oen_core[113]
port 531 nsew signal output
rlabel metal2 s 163134 10200 163190 11400 6 la_oen_core[114]
port 532 nsew signal output
rlabel metal2 s 163594 10200 163650 11400 6 la_oen_core[115]
port 533 nsew signal output
rlabel metal2 s 163962 10200 164018 11400 6 la_oen_core[116]
port 534 nsew signal output
rlabel metal2 s 164422 10200 164478 11400 6 la_oen_core[117]
port 535 nsew signal output
rlabel metal2 s 164882 10200 164938 11400 6 la_oen_core[118]
port 536 nsew signal output
rlabel metal2 s 165342 10200 165398 11400 6 la_oen_core[119]
port 537 nsew signal output
rlabel metal2 s 118238 10200 118294 11400 6 la_oen_core[11]
port 538 nsew signal output
rlabel metal2 s 165710 10200 165766 11400 6 la_oen_core[120]
port 539 nsew signal output
rlabel metal2 s 166170 10200 166226 11400 6 la_oen_core[121]
port 540 nsew signal output
rlabel metal2 s 166630 10200 166686 11400 6 la_oen_core[122]
port 541 nsew signal output
rlabel metal2 s 167090 10200 167146 11400 6 la_oen_core[123]
port 542 nsew signal output
rlabel metal2 s 167458 10200 167514 11400 6 la_oen_core[124]
port 543 nsew signal output
rlabel metal2 s 167918 10200 167974 11400 6 la_oen_core[125]
port 544 nsew signal output
rlabel metal2 s 168378 10200 168434 11400 6 la_oen_core[126]
port 545 nsew signal output
rlabel metal2 s 168746 10200 168802 11400 6 la_oen_core[127]
port 546 nsew signal output
rlabel metal2 s 118698 10200 118754 11400 6 la_oen_core[12]
port 547 nsew signal output
rlabel metal2 s 119158 10200 119214 11400 6 la_oen_core[13]
port 548 nsew signal output
rlabel metal2 s 119526 10200 119582 11400 6 la_oen_core[14]
port 549 nsew signal output
rlabel metal2 s 119986 10200 120042 11400 6 la_oen_core[15]
port 550 nsew signal output
rlabel metal2 s 120446 10200 120502 11400 6 la_oen_core[16]
port 551 nsew signal output
rlabel metal2 s 120814 10200 120870 11400 6 la_oen_core[17]
port 552 nsew signal output
rlabel metal2 s 121274 10200 121330 11400 6 la_oen_core[18]
port 553 nsew signal output
rlabel metal2 s 121734 10200 121790 11400 6 la_oen_core[19]
port 554 nsew signal output
rlabel metal2 s 113914 10200 113970 11400 6 la_oen_core[1]
port 555 nsew signal output
rlabel metal2 s 122194 10200 122250 11400 6 la_oen_core[20]
port 556 nsew signal output
rlabel metal2 s 122562 10200 122618 11400 6 la_oen_core[21]
port 557 nsew signal output
rlabel metal2 s 123022 10200 123078 11400 6 la_oen_core[22]
port 558 nsew signal output
rlabel metal2 s 123482 10200 123538 11400 6 la_oen_core[23]
port 559 nsew signal output
rlabel metal2 s 123942 10200 123998 11400 6 la_oen_core[24]
port 560 nsew signal output
rlabel metal2 s 124310 10200 124366 11400 6 la_oen_core[25]
port 561 nsew signal output
rlabel metal2 s 124770 10200 124826 11400 6 la_oen_core[26]
port 562 nsew signal output
rlabel metal2 s 125230 10200 125286 11400 6 la_oen_core[27]
port 563 nsew signal output
rlabel metal2 s 125690 10200 125746 11400 6 la_oen_core[28]
port 564 nsew signal output
rlabel metal2 s 126058 10200 126114 11400 6 la_oen_core[29]
port 565 nsew signal output
rlabel metal2 s 114282 10200 114338 11400 6 la_oen_core[2]
port 566 nsew signal output
rlabel metal2 s 126518 10200 126574 11400 6 la_oen_core[30]
port 567 nsew signal output
rlabel metal2 s 126978 10200 127034 11400 6 la_oen_core[31]
port 568 nsew signal output
rlabel metal2 s 127438 10200 127494 11400 6 la_oen_core[32]
port 569 nsew signal output
rlabel metal2 s 127806 10200 127862 11400 6 la_oen_core[33]
port 570 nsew signal output
rlabel metal2 s 128266 10200 128322 11400 6 la_oen_core[34]
port 571 nsew signal output
rlabel metal2 s 128726 10200 128782 11400 6 la_oen_core[35]
port 572 nsew signal output
rlabel metal2 s 129094 10200 129150 11400 6 la_oen_core[36]
port 573 nsew signal output
rlabel metal2 s 129554 10200 129610 11400 6 la_oen_core[37]
port 574 nsew signal output
rlabel metal2 s 130014 10200 130070 11400 6 la_oen_core[38]
port 575 nsew signal output
rlabel metal2 s 130474 10200 130530 11400 6 la_oen_core[39]
port 576 nsew signal output
rlabel metal2 s 114742 10200 114798 11400 6 la_oen_core[3]
port 577 nsew signal output
rlabel metal2 s 130842 10200 130898 11400 6 la_oen_core[40]
port 578 nsew signal output
rlabel metal2 s 131302 10200 131358 11400 6 la_oen_core[41]
port 579 nsew signal output
rlabel metal2 s 131762 10200 131818 11400 6 la_oen_core[42]
port 580 nsew signal output
rlabel metal2 s 132222 10200 132278 11400 6 la_oen_core[43]
port 581 nsew signal output
rlabel metal2 s 132590 10200 132646 11400 6 la_oen_core[44]
port 582 nsew signal output
rlabel metal2 s 133050 10200 133106 11400 6 la_oen_core[45]
port 583 nsew signal output
rlabel metal2 s 133510 10200 133566 11400 6 la_oen_core[46]
port 584 nsew signal output
rlabel metal2 s 133970 10200 134026 11400 6 la_oen_core[47]
port 585 nsew signal output
rlabel metal2 s 134338 10200 134394 11400 6 la_oen_core[48]
port 586 nsew signal output
rlabel metal2 s 134798 10200 134854 11400 6 la_oen_core[49]
port 587 nsew signal output
rlabel metal2 s 115202 10200 115258 11400 6 la_oen_core[4]
port 588 nsew signal output
rlabel metal2 s 135258 10200 135314 11400 6 la_oen_core[50]
port 589 nsew signal output
rlabel metal2 s 135718 10200 135774 11400 6 la_oen_core[51]
port 590 nsew signal output
rlabel metal2 s 136086 10200 136142 11400 6 la_oen_core[52]
port 591 nsew signal output
rlabel metal2 s 136546 10200 136602 11400 6 la_oen_core[53]
port 592 nsew signal output
rlabel metal2 s 137006 10200 137062 11400 6 la_oen_core[54]
port 593 nsew signal output
rlabel metal2 s 137374 10200 137430 11400 6 la_oen_core[55]
port 594 nsew signal output
rlabel metal2 s 137834 10200 137890 11400 6 la_oen_core[56]
port 595 nsew signal output
rlabel metal2 s 138294 10200 138350 11400 6 la_oen_core[57]
port 596 nsew signal output
rlabel metal2 s 138754 10200 138810 11400 6 la_oen_core[58]
port 597 nsew signal output
rlabel metal2 s 139122 10200 139178 11400 6 la_oen_core[59]
port 598 nsew signal output
rlabel metal2 s 115662 10200 115718 11400 6 la_oen_core[5]
port 599 nsew signal output
rlabel metal2 s 139582 10200 139638 11400 6 la_oen_core[60]
port 600 nsew signal output
rlabel metal2 s 140042 10200 140098 11400 6 la_oen_core[61]
port 601 nsew signal output
rlabel metal2 s 140502 10200 140558 11400 6 la_oen_core[62]
port 602 nsew signal output
rlabel metal2 s 140870 10200 140926 11400 6 la_oen_core[63]
port 603 nsew signal output
rlabel metal2 s 141330 10200 141386 11400 6 la_oen_core[64]
port 604 nsew signal output
rlabel metal2 s 141790 10200 141846 11400 6 la_oen_core[65]
port 605 nsew signal output
rlabel metal2 s 142250 10200 142306 11400 6 la_oen_core[66]
port 606 nsew signal output
rlabel metal2 s 142618 10200 142674 11400 6 la_oen_core[67]
port 607 nsew signal output
rlabel metal2 s 143078 10200 143134 11400 6 la_oen_core[68]
port 608 nsew signal output
rlabel metal2 s 143538 10200 143594 11400 6 la_oen_core[69]
port 609 nsew signal output
rlabel metal2 s 116030 10200 116086 11400 6 la_oen_core[6]
port 610 nsew signal output
rlabel metal2 s 143998 10200 144054 11400 6 la_oen_core[70]
port 611 nsew signal output
rlabel metal2 s 144366 10200 144422 11400 6 la_oen_core[71]
port 612 nsew signal output
rlabel metal2 s 144826 10200 144882 11400 6 la_oen_core[72]
port 613 nsew signal output
rlabel metal2 s 145286 10200 145342 11400 6 la_oen_core[73]
port 614 nsew signal output
rlabel metal2 s 145654 10200 145710 11400 6 la_oen_core[74]
port 615 nsew signal output
rlabel metal2 s 146114 10200 146170 11400 6 la_oen_core[75]
port 616 nsew signal output
rlabel metal2 s 146574 10200 146630 11400 6 la_oen_core[76]
port 617 nsew signal output
rlabel metal2 s 147034 10200 147090 11400 6 la_oen_core[77]
port 618 nsew signal output
rlabel metal2 s 147402 10200 147458 11400 6 la_oen_core[78]
port 619 nsew signal output
rlabel metal2 s 147862 10200 147918 11400 6 la_oen_core[79]
port 620 nsew signal output
rlabel metal2 s 116490 10200 116546 11400 6 la_oen_core[7]
port 621 nsew signal output
rlabel metal2 s 148322 10200 148378 11400 6 la_oen_core[80]
port 622 nsew signal output
rlabel metal2 s 148782 10200 148838 11400 6 la_oen_core[81]
port 623 nsew signal output
rlabel metal2 s 149150 10200 149206 11400 6 la_oen_core[82]
port 624 nsew signal output
rlabel metal2 s 149610 10200 149666 11400 6 la_oen_core[83]
port 625 nsew signal output
rlabel metal2 s 150070 10200 150126 11400 6 la_oen_core[84]
port 626 nsew signal output
rlabel metal2 s 150530 10200 150586 11400 6 la_oen_core[85]
port 627 nsew signal output
rlabel metal2 s 150898 10200 150954 11400 6 la_oen_core[86]
port 628 nsew signal output
rlabel metal2 s 151358 10200 151414 11400 6 la_oen_core[87]
port 629 nsew signal output
rlabel metal2 s 151818 10200 151874 11400 6 la_oen_core[88]
port 630 nsew signal output
rlabel metal2 s 152186 10200 152242 11400 6 la_oen_core[89]
port 631 nsew signal output
rlabel metal2 s 116950 10200 117006 11400 6 la_oen_core[8]
port 632 nsew signal output
rlabel metal2 s 152646 10200 152702 11400 6 la_oen_core[90]
port 633 nsew signal output
rlabel metal2 s 153106 10200 153162 11400 6 la_oen_core[91]
port 634 nsew signal output
rlabel metal2 s 153566 10200 153622 11400 6 la_oen_core[92]
port 635 nsew signal output
rlabel metal2 s 153934 10200 153990 11400 6 la_oen_core[93]
port 636 nsew signal output
rlabel metal2 s 154394 10200 154450 11400 6 la_oen_core[94]
port 637 nsew signal output
rlabel metal2 s 154854 10200 154910 11400 6 la_oen_core[95]
port 638 nsew signal output
rlabel metal2 s 155314 10200 155370 11400 6 la_oen_core[96]
port 639 nsew signal output
rlabel metal2 s 155682 10200 155738 11400 6 la_oen_core[97]
port 640 nsew signal output
rlabel metal2 s 156142 10200 156198 11400 6 la_oen_core[98]
port 641 nsew signal output
rlabel metal2 s 156602 10200 156658 11400 6 la_oen_core[99]
port 642 nsew signal output
rlabel metal2 s 117410 10200 117466 11400 6 la_oen_core[9]
port 643 nsew signal output
rlabel metal2 s 111706 -400 111762 800 6 la_oen_mprj[0]
port 644 nsew signal input
rlabel metal2 s 155314 -400 155370 800 6 la_oen_mprj[100]
port 645 nsew signal input
rlabel metal2 s 155682 -400 155738 800 6 la_oen_mprj[101]
port 646 nsew signal input
rlabel metal2 s 156142 -400 156198 800 6 la_oen_mprj[102]
port 647 nsew signal input
rlabel metal2 s 156602 -400 156658 800 6 la_oen_mprj[103]
port 648 nsew signal input
rlabel metal2 s 157062 -400 157118 800 6 la_oen_mprj[104]
port 649 nsew signal input
rlabel metal2 s 157430 -400 157486 800 6 la_oen_mprj[105]
port 650 nsew signal input
rlabel metal2 s 157890 -400 157946 800 6 la_oen_mprj[106]
port 651 nsew signal input
rlabel metal2 s 158350 -400 158406 800 6 la_oen_mprj[107]
port 652 nsew signal input
rlabel metal2 s 158810 -400 158866 800 6 la_oen_mprj[108]
port 653 nsew signal input
rlabel metal2 s 159178 -400 159234 800 6 la_oen_mprj[109]
port 654 nsew signal input
rlabel metal2 s 116030 -400 116086 800 6 la_oen_mprj[10]
port 655 nsew signal input
rlabel metal2 s 159638 -400 159694 800 6 la_oen_mprj[110]
port 656 nsew signal input
rlabel metal2 s 160098 -400 160154 800 6 la_oen_mprj[111]
port 657 nsew signal input
rlabel metal2 s 160466 -400 160522 800 6 la_oen_mprj[112]
port 658 nsew signal input
rlabel metal2 s 160926 -400 160982 800 6 la_oen_mprj[113]
port 659 nsew signal input
rlabel metal2 s 161386 -400 161442 800 6 la_oen_mprj[114]
port 660 nsew signal input
rlabel metal2 s 161846 -400 161902 800 6 la_oen_mprj[115]
port 661 nsew signal input
rlabel metal2 s 162214 -400 162270 800 6 la_oen_mprj[116]
port 662 nsew signal input
rlabel metal2 s 162674 -400 162730 800 6 la_oen_mprj[117]
port 663 nsew signal input
rlabel metal2 s 163134 -400 163190 800 6 la_oen_mprj[118]
port 664 nsew signal input
rlabel metal2 s 163594 -400 163650 800 6 la_oen_mprj[119]
port 665 nsew signal input
rlabel metal2 s 116490 -400 116546 800 6 la_oen_mprj[11]
port 666 nsew signal input
rlabel metal2 s 163962 -400 164018 800 6 la_oen_mprj[120]
port 667 nsew signal input
rlabel metal2 s 164422 -400 164478 800 6 la_oen_mprj[121]
port 668 nsew signal input
rlabel metal2 s 164882 -400 164938 800 6 la_oen_mprj[122]
port 669 nsew signal input
rlabel metal2 s 165342 -400 165398 800 6 la_oen_mprj[123]
port 670 nsew signal input
rlabel metal2 s 165710 -400 165766 800 6 la_oen_mprj[124]
port 671 nsew signal input
rlabel metal2 s 166170 -400 166226 800 6 la_oen_mprj[125]
port 672 nsew signal input
rlabel metal2 s 166630 -400 166686 800 6 la_oen_mprj[126]
port 673 nsew signal input
rlabel metal2 s 167090 -400 167146 800 6 la_oen_mprj[127]
port 674 nsew signal input
rlabel metal2 s 116950 -400 117006 800 6 la_oen_mprj[12]
port 675 nsew signal input
rlabel metal2 s 117410 -400 117466 800 6 la_oen_mprj[13]
port 676 nsew signal input
rlabel metal2 s 117778 -400 117834 800 6 la_oen_mprj[14]
port 677 nsew signal input
rlabel metal2 s 118238 -400 118294 800 6 la_oen_mprj[15]
port 678 nsew signal input
rlabel metal2 s 118698 -400 118754 800 6 la_oen_mprj[16]
port 679 nsew signal input
rlabel metal2 s 119158 -400 119214 800 6 la_oen_mprj[17]
port 680 nsew signal input
rlabel metal2 s 119526 -400 119582 800 6 la_oen_mprj[18]
port 681 nsew signal input
rlabel metal2 s 119986 -400 120042 800 6 la_oen_mprj[19]
port 682 nsew signal input
rlabel metal2 s 112166 -400 112222 800 6 la_oen_mprj[1]
port 683 nsew signal input
rlabel metal2 s 120446 -400 120502 800 6 la_oen_mprj[20]
port 684 nsew signal input
rlabel metal2 s 120814 -400 120870 800 6 la_oen_mprj[21]
port 685 nsew signal input
rlabel metal2 s 121274 -400 121330 800 6 la_oen_mprj[22]
port 686 nsew signal input
rlabel metal2 s 121734 -400 121790 800 6 la_oen_mprj[23]
port 687 nsew signal input
rlabel metal2 s 122194 -400 122250 800 6 la_oen_mprj[24]
port 688 nsew signal input
rlabel metal2 s 122562 -400 122618 800 6 la_oen_mprj[25]
port 689 nsew signal input
rlabel metal2 s 123022 -400 123078 800 6 la_oen_mprj[26]
port 690 nsew signal input
rlabel metal2 s 123482 -400 123538 800 6 la_oen_mprj[27]
port 691 nsew signal input
rlabel metal2 s 123942 -400 123998 800 6 la_oen_mprj[28]
port 692 nsew signal input
rlabel metal2 s 124310 -400 124366 800 6 la_oen_mprj[29]
port 693 nsew signal input
rlabel metal2 s 112534 -400 112590 800 6 la_oen_mprj[2]
port 694 nsew signal input
rlabel metal2 s 124770 -400 124826 800 6 la_oen_mprj[30]
port 695 nsew signal input
rlabel metal2 s 125230 -400 125286 800 6 la_oen_mprj[31]
port 696 nsew signal input
rlabel metal2 s 125690 -400 125746 800 6 la_oen_mprj[32]
port 697 nsew signal input
rlabel metal2 s 126058 -400 126114 800 6 la_oen_mprj[33]
port 698 nsew signal input
rlabel metal2 s 126518 -400 126574 800 6 la_oen_mprj[34]
port 699 nsew signal input
rlabel metal2 s 126978 -400 127034 800 6 la_oen_mprj[35]
port 700 nsew signal input
rlabel metal2 s 127438 -400 127494 800 6 la_oen_mprj[36]
port 701 nsew signal input
rlabel metal2 s 127806 -400 127862 800 6 la_oen_mprj[37]
port 702 nsew signal input
rlabel metal2 s 128266 -400 128322 800 6 la_oen_mprj[38]
port 703 nsew signal input
rlabel metal2 s 128726 -400 128782 800 6 la_oen_mprj[39]
port 704 nsew signal input
rlabel metal2 s 112994 -400 113050 800 6 la_oen_mprj[3]
port 705 nsew signal input
rlabel metal2 s 129094 -400 129150 800 6 la_oen_mprj[40]
port 706 nsew signal input
rlabel metal2 s 129554 -400 129610 800 6 la_oen_mprj[41]
port 707 nsew signal input
rlabel metal2 s 130014 -400 130070 800 6 la_oen_mprj[42]
port 708 nsew signal input
rlabel metal2 s 130474 -400 130530 800 6 la_oen_mprj[43]
port 709 nsew signal input
rlabel metal2 s 130842 -400 130898 800 6 la_oen_mprj[44]
port 710 nsew signal input
rlabel metal2 s 131302 -400 131358 800 6 la_oen_mprj[45]
port 711 nsew signal input
rlabel metal2 s 131762 -400 131818 800 6 la_oen_mprj[46]
port 712 nsew signal input
rlabel metal2 s 132222 -400 132278 800 6 la_oen_mprj[47]
port 713 nsew signal input
rlabel metal2 s 132590 -400 132646 800 6 la_oen_mprj[48]
port 714 nsew signal input
rlabel metal2 s 133050 -400 133106 800 6 la_oen_mprj[49]
port 715 nsew signal input
rlabel metal2 s 113454 -400 113510 800 6 la_oen_mprj[4]
port 716 nsew signal input
rlabel metal2 s 133510 -400 133566 800 6 la_oen_mprj[50]
port 717 nsew signal input
rlabel metal2 s 133970 -400 134026 800 6 la_oen_mprj[51]
port 718 nsew signal input
rlabel metal2 s 134338 -400 134394 800 6 la_oen_mprj[52]
port 719 nsew signal input
rlabel metal2 s 134798 -400 134854 800 6 la_oen_mprj[53]
port 720 nsew signal input
rlabel metal2 s 135258 -400 135314 800 6 la_oen_mprj[54]
port 721 nsew signal input
rlabel metal2 s 135718 -400 135774 800 6 la_oen_mprj[55]
port 722 nsew signal input
rlabel metal2 s 136086 -400 136142 800 6 la_oen_mprj[56]
port 723 nsew signal input
rlabel metal2 s 136546 -400 136602 800 6 la_oen_mprj[57]
port 724 nsew signal input
rlabel metal2 s 137006 -400 137062 800 6 la_oen_mprj[58]
port 725 nsew signal input
rlabel metal2 s 137374 -400 137430 800 6 la_oen_mprj[59]
port 726 nsew signal input
rlabel metal2 s 113914 -400 113970 800 6 la_oen_mprj[5]
port 727 nsew signal input
rlabel metal2 s 137834 -400 137890 800 6 la_oen_mprj[60]
port 728 nsew signal input
rlabel metal2 s 138294 -400 138350 800 6 la_oen_mprj[61]
port 729 nsew signal input
rlabel metal2 s 138754 -400 138810 800 6 la_oen_mprj[62]
port 730 nsew signal input
rlabel metal2 s 139122 -400 139178 800 6 la_oen_mprj[63]
port 731 nsew signal input
rlabel metal2 s 139582 -400 139638 800 6 la_oen_mprj[64]
port 732 nsew signal input
rlabel metal2 s 140042 -400 140098 800 6 la_oen_mprj[65]
port 733 nsew signal input
rlabel metal2 s 140502 -400 140558 800 6 la_oen_mprj[66]
port 734 nsew signal input
rlabel metal2 s 140870 -400 140926 800 6 la_oen_mprj[67]
port 735 nsew signal input
rlabel metal2 s 141330 -400 141386 800 6 la_oen_mprj[68]
port 736 nsew signal input
rlabel metal2 s 141790 -400 141846 800 6 la_oen_mprj[69]
port 737 nsew signal input
rlabel metal2 s 114282 -400 114338 800 6 la_oen_mprj[6]
port 738 nsew signal input
rlabel metal2 s 142250 -400 142306 800 6 la_oen_mprj[70]
port 739 nsew signal input
rlabel metal2 s 142618 -400 142674 800 6 la_oen_mprj[71]
port 740 nsew signal input
rlabel metal2 s 143078 -400 143134 800 6 la_oen_mprj[72]
port 741 nsew signal input
rlabel metal2 s 143538 -400 143594 800 6 la_oen_mprj[73]
port 742 nsew signal input
rlabel metal2 s 143998 -400 144054 800 6 la_oen_mprj[74]
port 743 nsew signal input
rlabel metal2 s 144366 -400 144422 800 6 la_oen_mprj[75]
port 744 nsew signal input
rlabel metal2 s 144826 -400 144882 800 6 la_oen_mprj[76]
port 745 nsew signal input
rlabel metal2 s 145286 -400 145342 800 6 la_oen_mprj[77]
port 746 nsew signal input
rlabel metal2 s 145654 -400 145710 800 6 la_oen_mprj[78]
port 747 nsew signal input
rlabel metal2 s 146114 -400 146170 800 6 la_oen_mprj[79]
port 748 nsew signal input
rlabel metal2 s 114742 -400 114798 800 6 la_oen_mprj[7]
port 749 nsew signal input
rlabel metal2 s 146574 -400 146630 800 6 la_oen_mprj[80]
port 750 nsew signal input
rlabel metal2 s 147034 -400 147090 800 6 la_oen_mprj[81]
port 751 nsew signal input
rlabel metal2 s 147402 -400 147458 800 6 la_oen_mprj[82]
port 752 nsew signal input
rlabel metal2 s 147862 -400 147918 800 6 la_oen_mprj[83]
port 753 nsew signal input
rlabel metal2 s 148322 -400 148378 800 6 la_oen_mprj[84]
port 754 nsew signal input
rlabel metal2 s 148782 -400 148838 800 6 la_oen_mprj[85]
port 755 nsew signal input
rlabel metal2 s 149150 -400 149206 800 6 la_oen_mprj[86]
port 756 nsew signal input
rlabel metal2 s 149610 -400 149666 800 6 la_oen_mprj[87]
port 757 nsew signal input
rlabel metal2 s 150070 -400 150126 800 6 la_oen_mprj[88]
port 758 nsew signal input
rlabel metal2 s 150530 -400 150586 800 6 la_oen_mprj[89]
port 759 nsew signal input
rlabel metal2 s 115202 -400 115258 800 6 la_oen_mprj[8]
port 760 nsew signal input
rlabel metal2 s 150898 -400 150954 800 6 la_oen_mprj[90]
port 761 nsew signal input
rlabel metal2 s 151358 -400 151414 800 6 la_oen_mprj[91]
port 762 nsew signal input
rlabel metal2 s 151818 -400 151874 800 6 la_oen_mprj[92]
port 763 nsew signal input
rlabel metal2 s 152186 -400 152242 800 6 la_oen_mprj[93]
port 764 nsew signal input
rlabel metal2 s 152646 -400 152702 800 6 la_oen_mprj[94]
port 765 nsew signal input
rlabel metal2 s 153106 -400 153162 800 6 la_oen_mprj[95]
port 766 nsew signal input
rlabel metal2 s 153566 -400 153622 800 6 la_oen_mprj[96]
port 767 nsew signal input
rlabel metal2 s 153934 -400 153990 800 6 la_oen_mprj[97]
port 768 nsew signal input
rlabel metal2 s 154394 -400 154450 800 6 la_oen_mprj[98]
port 769 nsew signal input
rlabel metal2 s 154854 -400 154910 800 6 la_oen_mprj[99]
port 770 nsew signal input
rlabel metal2 s 115662 -400 115718 800 6 la_oen_mprj[9]
port 771 nsew signal input
rlabel metal2 s 168746 -400 168802 800 6 mprj_adr_o_core[0]
port 772 nsew signal input
rlabel metal2 s 179234 -400 179290 800 6 mprj_adr_o_core[10]
port 773 nsew signal input
rlabel metal2 s 180154 -400 180210 800 6 mprj_adr_o_core[11]
port 774 nsew signal input
rlabel metal2 s 180982 -400 181038 800 6 mprj_adr_o_core[12]
port 775 nsew signal input
rlabel metal2 s 181902 -400 181958 800 6 mprj_adr_o_core[13]
port 776 nsew signal input
rlabel metal2 s 182730 -400 182786 800 6 mprj_adr_o_core[14]
port 777 nsew signal input
rlabel metal2 s 183650 -400 183706 800 6 mprj_adr_o_core[15]
port 778 nsew signal input
rlabel metal2 s 184478 -400 184534 800 6 mprj_adr_o_core[16]
port 779 nsew signal input
rlabel metal2 s 185306 -400 185362 800 6 mprj_adr_o_core[17]
port 780 nsew signal input
rlabel metal2 s 186226 -400 186282 800 6 mprj_adr_o_core[18]
port 781 nsew signal input
rlabel metal2 s 187054 -400 187110 800 6 mprj_adr_o_core[19]
port 782 nsew signal input
rlabel metal2 s 170126 -400 170182 800 6 mprj_adr_o_core[1]
port 783 nsew signal input
rlabel metal2 s 187974 -400 188030 800 6 mprj_adr_o_core[20]
port 784 nsew signal input
rlabel metal2 s 188802 -400 188858 800 6 mprj_adr_o_core[21]
port 785 nsew signal input
rlabel metal2 s 189722 -400 189778 800 6 mprj_adr_o_core[22]
port 786 nsew signal input
rlabel metal2 s 190550 -400 190606 800 6 mprj_adr_o_core[23]
port 787 nsew signal input
rlabel metal2 s 191470 -400 191526 800 6 mprj_adr_o_core[24]
port 788 nsew signal input
rlabel metal2 s 192298 -400 192354 800 6 mprj_adr_o_core[25]
port 789 nsew signal input
rlabel metal2 s 193218 -400 193274 800 6 mprj_adr_o_core[26]
port 790 nsew signal input
rlabel metal2 s 194046 -400 194102 800 6 mprj_adr_o_core[27]
port 791 nsew signal input
rlabel metal2 s 194966 -400 195022 800 6 mprj_adr_o_core[28]
port 792 nsew signal input
rlabel metal2 s 195794 -400 195850 800 6 mprj_adr_o_core[29]
port 793 nsew signal input
rlabel metal2 s 171414 -400 171470 800 6 mprj_adr_o_core[2]
port 794 nsew signal input
rlabel metal2 s 196714 -400 196770 800 6 mprj_adr_o_core[30]
port 795 nsew signal input
rlabel metal2 s 197542 -400 197598 800 6 mprj_adr_o_core[31]
port 796 nsew signal input
rlabel metal2 s 172702 -400 172758 800 6 mprj_adr_o_core[3]
port 797 nsew signal input
rlabel metal2 s 173990 -400 174046 800 6 mprj_adr_o_core[4]
port 798 nsew signal input
rlabel metal2 s 174910 -400 174966 800 6 mprj_adr_o_core[5]
port 799 nsew signal input
rlabel metal2 s 175738 -400 175794 800 6 mprj_adr_o_core[6]
port 800 nsew signal input
rlabel metal2 s 176658 -400 176714 800 6 mprj_adr_o_core[7]
port 801 nsew signal input
rlabel metal2 s 177486 -400 177542 800 6 mprj_adr_o_core[8]
port 802 nsew signal input
rlabel metal2 s 178406 -400 178462 800 6 mprj_adr_o_core[9]
port 803 nsew signal input
rlabel metal2 s 170494 10200 170550 11400 6 mprj_adr_o_user[0]
port 804 nsew signal output
rlabel metal2 s 180982 10200 181038 11400 6 mprj_adr_o_user[10]
port 805 nsew signal output
rlabel metal2 s 181902 10200 181958 11400 6 mprj_adr_o_user[11]
port 806 nsew signal output
rlabel metal2 s 182730 10200 182786 11400 6 mprj_adr_o_user[12]
port 807 nsew signal output
rlabel metal2 s 183650 10200 183706 11400 6 mprj_adr_o_user[13]
port 808 nsew signal output
rlabel metal2 s 184478 10200 184534 11400 6 mprj_adr_o_user[14]
port 809 nsew signal output
rlabel metal2 s 185306 10200 185362 11400 6 mprj_adr_o_user[15]
port 810 nsew signal output
rlabel metal2 s 186226 10200 186282 11400 6 mprj_adr_o_user[16]
port 811 nsew signal output
rlabel metal2 s 187054 10200 187110 11400 6 mprj_adr_o_user[17]
port 812 nsew signal output
rlabel metal2 s 187974 10200 188030 11400 6 mprj_adr_o_user[18]
port 813 nsew signal output
rlabel metal2 s 188802 10200 188858 11400 6 mprj_adr_o_user[19]
port 814 nsew signal output
rlabel metal2 s 171874 10200 171930 11400 6 mprj_adr_o_user[1]
port 815 nsew signal output
rlabel metal2 s 189722 10200 189778 11400 6 mprj_adr_o_user[20]
port 816 nsew signal output
rlabel metal2 s 190550 10200 190606 11400 6 mprj_adr_o_user[21]
port 817 nsew signal output
rlabel metal2 s 191470 10200 191526 11400 6 mprj_adr_o_user[22]
port 818 nsew signal output
rlabel metal2 s 192298 10200 192354 11400 6 mprj_adr_o_user[23]
port 819 nsew signal output
rlabel metal2 s 193218 10200 193274 11400 6 mprj_adr_o_user[24]
port 820 nsew signal output
rlabel metal2 s 194046 10200 194102 11400 6 mprj_adr_o_user[25]
port 821 nsew signal output
rlabel metal2 s 194966 10200 195022 11400 6 mprj_adr_o_user[26]
port 822 nsew signal output
rlabel metal2 s 195794 10200 195850 11400 6 mprj_adr_o_user[27]
port 823 nsew signal output
rlabel metal2 s 196714 10200 196770 11400 6 mprj_adr_o_user[28]
port 824 nsew signal output
rlabel metal2 s 197542 10200 197598 11400 6 mprj_adr_o_user[29]
port 825 nsew signal output
rlabel metal2 s 173162 10200 173218 11400 6 mprj_adr_o_user[2]
port 826 nsew signal output
rlabel metal2 s 198462 10200 198518 11400 6 mprj_adr_o_user[30]
port 827 nsew signal output
rlabel metal2 s 199290 10200 199346 11400 6 mprj_adr_o_user[31]
port 828 nsew signal output
rlabel metal2 s 174450 10200 174506 11400 6 mprj_adr_o_user[3]
port 829 nsew signal output
rlabel metal2 s 175738 10200 175794 11400 6 mprj_adr_o_user[4]
port 830 nsew signal output
rlabel metal2 s 176658 10200 176714 11400 6 mprj_adr_o_user[5]
port 831 nsew signal output
rlabel metal2 s 177486 10200 177542 11400 6 mprj_adr_o_user[6]
port 832 nsew signal output
rlabel metal2 s 178406 10200 178462 11400 6 mprj_adr_o_user[7]
port 833 nsew signal output
rlabel metal2 s 179234 10200 179290 11400 6 mprj_adr_o_user[8]
port 834 nsew signal output
rlabel metal2 s 180154 10200 180210 11400 6 mprj_adr_o_user[9]
port 835 nsew signal output
rlabel metal2 s 167458 -400 167514 800 6 mprj_cyc_o_core
port 836 nsew signal input
rlabel metal2 s 169206 10200 169262 11400 6 mprj_cyc_o_user
port 837 nsew signal output
rlabel metal2 s 169206 -400 169262 800 6 mprj_dat_o_core[0]
port 838 nsew signal input
rlabel metal2 s 179694 -400 179750 800 6 mprj_dat_o_core[10]
port 839 nsew signal input
rlabel metal2 s 180522 -400 180578 800 6 mprj_dat_o_core[11]
port 840 nsew signal input
rlabel metal2 s 181442 -400 181498 800 6 mprj_dat_o_core[12]
port 841 nsew signal input
rlabel metal2 s 182270 -400 182326 800 6 mprj_dat_o_core[13]
port 842 nsew signal input
rlabel metal2 s 183190 -400 183246 800 6 mprj_dat_o_core[14]
port 843 nsew signal input
rlabel metal2 s 184018 -400 184074 800 6 mprj_dat_o_core[15]
port 844 nsew signal input
rlabel metal2 s 184938 -400 184994 800 6 mprj_dat_o_core[16]
port 845 nsew signal input
rlabel metal2 s 185766 -400 185822 800 6 mprj_dat_o_core[17]
port 846 nsew signal input
rlabel metal2 s 186686 -400 186742 800 6 mprj_dat_o_core[18]
port 847 nsew signal input
rlabel metal2 s 187514 -400 187570 800 6 mprj_dat_o_core[19]
port 848 nsew signal input
rlabel metal2 s 170494 -400 170550 800 6 mprj_dat_o_core[1]
port 849 nsew signal input
rlabel metal2 s 188434 -400 188490 800 6 mprj_dat_o_core[20]
port 850 nsew signal input
rlabel metal2 s 189262 -400 189318 800 6 mprj_dat_o_core[21]
port 851 nsew signal input
rlabel metal2 s 190182 -400 190238 800 6 mprj_dat_o_core[22]
port 852 nsew signal input
rlabel metal2 s 191010 -400 191066 800 6 mprj_dat_o_core[23]
port 853 nsew signal input
rlabel metal2 s 191930 -400 191986 800 6 mprj_dat_o_core[24]
port 854 nsew signal input
rlabel metal2 s 192758 -400 192814 800 6 mprj_dat_o_core[25]
port 855 nsew signal input
rlabel metal2 s 193586 -400 193642 800 6 mprj_dat_o_core[26]
port 856 nsew signal input
rlabel metal2 s 194506 -400 194562 800 6 mprj_dat_o_core[27]
port 857 nsew signal input
rlabel metal2 s 195334 -400 195390 800 6 mprj_dat_o_core[28]
port 858 nsew signal input
rlabel metal2 s 196254 -400 196310 800 6 mprj_dat_o_core[29]
port 859 nsew signal input
rlabel metal2 s 171874 -400 171930 800 6 mprj_dat_o_core[2]
port 860 nsew signal input
rlabel metal2 s 197082 -400 197138 800 6 mprj_dat_o_core[30]
port 861 nsew signal input
rlabel metal2 s 198002 -400 198058 800 6 mprj_dat_o_core[31]
port 862 nsew signal input
rlabel metal2 s 173162 -400 173218 800 6 mprj_dat_o_core[3]
port 863 nsew signal input
rlabel metal2 s 174450 -400 174506 800 6 mprj_dat_o_core[4]
port 864 nsew signal input
rlabel metal2 s 175370 -400 175426 800 6 mprj_dat_o_core[5]
port 865 nsew signal input
rlabel metal2 s 176198 -400 176254 800 6 mprj_dat_o_core[6]
port 866 nsew signal input
rlabel metal2 s 177026 -400 177082 800 6 mprj_dat_o_core[7]
port 867 nsew signal input
rlabel metal2 s 177946 -400 178002 800 6 mprj_dat_o_core[8]
port 868 nsew signal input
rlabel metal2 s 178774 -400 178830 800 6 mprj_dat_o_core[9]
port 869 nsew signal input
rlabel metal2 s 170954 10200 171010 11400 6 mprj_dat_o_user[0]
port 870 nsew signal output
rlabel metal2 s 181442 10200 181498 11400 6 mprj_dat_o_user[10]
port 871 nsew signal output
rlabel metal2 s 182270 10200 182326 11400 6 mprj_dat_o_user[11]
port 872 nsew signal output
rlabel metal2 s 183190 10200 183246 11400 6 mprj_dat_o_user[12]
port 873 nsew signal output
rlabel metal2 s 184018 10200 184074 11400 6 mprj_dat_o_user[13]
port 874 nsew signal output
rlabel metal2 s 184938 10200 184994 11400 6 mprj_dat_o_user[14]
port 875 nsew signal output
rlabel metal2 s 185766 10200 185822 11400 6 mprj_dat_o_user[15]
port 876 nsew signal output
rlabel metal2 s 186686 10200 186742 11400 6 mprj_dat_o_user[16]
port 877 nsew signal output
rlabel metal2 s 187514 10200 187570 11400 6 mprj_dat_o_user[17]
port 878 nsew signal output
rlabel metal2 s 188434 10200 188490 11400 6 mprj_dat_o_user[18]
port 879 nsew signal output
rlabel metal2 s 189262 10200 189318 11400 6 mprj_dat_o_user[19]
port 880 nsew signal output
rlabel metal2 s 172242 10200 172298 11400 6 mprj_dat_o_user[1]
port 881 nsew signal output
rlabel metal2 s 190182 10200 190238 11400 6 mprj_dat_o_user[20]
port 882 nsew signal output
rlabel metal2 s 191010 10200 191066 11400 6 mprj_dat_o_user[21]
port 883 nsew signal output
rlabel metal2 s 191930 10200 191986 11400 6 mprj_dat_o_user[22]
port 884 nsew signal output
rlabel metal2 s 192758 10200 192814 11400 6 mprj_dat_o_user[23]
port 885 nsew signal output
rlabel metal2 s 193586 10200 193642 11400 6 mprj_dat_o_user[24]
port 886 nsew signal output
rlabel metal2 s 194506 10200 194562 11400 6 mprj_dat_o_user[25]
port 887 nsew signal output
rlabel metal2 s 195334 10200 195390 11400 6 mprj_dat_o_user[26]
port 888 nsew signal output
rlabel metal2 s 196254 10200 196310 11400 6 mprj_dat_o_user[27]
port 889 nsew signal output
rlabel metal2 s 197082 10200 197138 11400 6 mprj_dat_o_user[28]
port 890 nsew signal output
rlabel metal2 s 198002 10200 198058 11400 6 mprj_dat_o_user[29]
port 891 nsew signal output
rlabel metal2 s 173622 10200 173678 11400 6 mprj_dat_o_user[2]
port 892 nsew signal output
rlabel metal2 s 198830 10200 198886 11400 6 mprj_dat_o_user[30]
port 893 nsew signal output
rlabel metal2 s 199750 10200 199806 11400 6 mprj_dat_o_user[31]
port 894 nsew signal output
rlabel metal2 s 174910 10200 174966 11400 6 mprj_dat_o_user[3]
port 895 nsew signal output
rlabel metal2 s 176198 10200 176254 11400 6 mprj_dat_o_user[4]
port 896 nsew signal output
rlabel metal2 s 177026 10200 177082 11400 6 mprj_dat_o_user[5]
port 897 nsew signal output
rlabel metal2 s 177946 10200 178002 11400 6 mprj_dat_o_user[6]
port 898 nsew signal output
rlabel metal2 s 178774 10200 178830 11400 6 mprj_dat_o_user[7]
port 899 nsew signal output
rlabel metal2 s 179694 10200 179750 11400 6 mprj_dat_o_user[8]
port 900 nsew signal output
rlabel metal2 s 180522 10200 180578 11400 6 mprj_dat_o_user[9]
port 901 nsew signal output
rlabel metal2 s 169666 -400 169722 800 6 mprj_sel_o_core[0]
port 902 nsew signal input
rlabel metal2 s 170954 -400 171010 800 6 mprj_sel_o_core[1]
port 903 nsew signal input
rlabel metal2 s 172242 -400 172298 800 6 mprj_sel_o_core[2]
port 904 nsew signal input
rlabel metal2 s 173622 -400 173678 800 6 mprj_sel_o_core[3]
port 905 nsew signal input
rlabel metal2 s 171414 10200 171470 11400 6 mprj_sel_o_user[0]
port 906 nsew signal output
rlabel metal2 s 172702 10200 172758 11400 6 mprj_sel_o_user[1]
port 907 nsew signal output
rlabel metal2 s 173990 10200 174046 11400 6 mprj_sel_o_user[2]
port 908 nsew signal output
rlabel metal2 s 175370 10200 175426 11400 6 mprj_sel_o_user[3]
port 909 nsew signal output
rlabel metal2 s 167918 -400 167974 800 6 mprj_stb_o_core
port 910 nsew signal input
rlabel metal2 s 169666 10200 169722 11400 6 mprj_stb_o_user
port 911 nsew signal output
rlabel metal2 s 168378 -400 168434 800 6 mprj_we_o_core
port 912 nsew signal input
rlabel metal2 s 170126 10200 170182 11400 6 mprj_we_o_user
port 913 nsew signal output
rlabel metal2 s 198462 -400 198518 800 6 user1_vcc_powergood
port 914 nsew signal output
rlabel metal2 s 198830 -400 198886 800 6 user1_vdd_powergood
port 915 nsew signal output
rlabel metal2 s 199290 -400 199346 800 6 user2_vcc_powergood
port 916 nsew signal output
rlabel metal2 s 199750 -400 199806 800 6 user2_vdd_powergood
port 917 nsew signal output
rlabel metal2 s 202 10200 258 11400 6 user_clock
port 918 nsew signal output
rlabel metal2 s 570 10200 626 11400 6 user_clock2
port 919 nsew signal output
rlabel metal2 s 1030 10200 1086 11400 6 user_reset
port 920 nsew signal output
rlabel metal2 s 1490 10200 1546 11400 6 user_resetn
port 921 nsew signal output
rlabel metal3 s -326 11162 200242 11222 6 vccd1
port 922 nsew power bidirectional
rlabel metal3 s -326 -342 200242 -282 8 vccd1
port 923 nsew power bidirectional
rlabel metal4 s 164074 -482 164134 11362 6 vccd1
port 924 nsew power bidirectional
rlabel metal4 s 124074 -482 124134 11362 6 vccd1
port 925 nsew power bidirectional
rlabel metal4 s 84074 -482 84134 11362 6 vccd1
port 926 nsew power bidirectional
rlabel metal4 s 44074 -482 44134 11362 6 vccd1
port 927 nsew power bidirectional
rlabel metal4 s 4074 -482 4134 11362 6 vccd1
port 928 nsew power bidirectional
rlabel metal4 s 200182 -342 200242 11222 6 vccd1
port 929 nsew power bidirectional
rlabel metal4 s -326 -342 -266 11222 4 vccd1
port 930 nsew power bidirectional
rlabel metal3 s -466 11302 200382 11362 6 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s -466 -482 200382 -422 8 vssd1
port 932 nsew ground bidirectional
rlabel metal4 s 200322 -482 200382 11362 6 vssd1
port 933 nsew ground bidirectional
rlabel metal4 s 184074 -482 184134 11362 6 vssd1
port 934 nsew ground bidirectional
rlabel metal4 s 144074 -482 144134 11362 6 vssd1
port 935 nsew ground bidirectional
rlabel metal4 s 104074 -482 104134 11362 6 vssd1
port 936 nsew ground bidirectional
rlabel metal4 s 64074 -482 64134 11362 6 vssd1
port 937 nsew ground bidirectional
rlabel metal4 s 24074 -482 24134 11362 6 vssd1
port 938 nsew ground bidirectional
rlabel metal4 s -466 -482 -406 11362 4 vssd1
port 939 nsew ground bidirectional
rlabel metal3 s -606 11442 200522 11502 6 vccd
port 940 nsew power bidirectional
rlabel metal3 s -606 -622 200522 -562 8 vccd
port 941 nsew power bidirectional
rlabel metal4 s 164474 -762 164534 11642 6 vccd
port 942 nsew power bidirectional
rlabel metal4 s 124474 -762 124534 11642 6 vccd
port 943 nsew power bidirectional
rlabel metal4 s 84474 -762 84534 11642 6 vccd
port 944 nsew power bidirectional
rlabel metal4 s 44474 -762 44534 11642 6 vccd
port 945 nsew power bidirectional
rlabel metal4 s 4474 -762 4534 11642 6 vccd
port 946 nsew power bidirectional
rlabel metal4 s 200462 -622 200522 11502 6 vccd
port 947 nsew power bidirectional
rlabel metal4 s -606 -622 -546 11502 4 vccd
port 948 nsew power bidirectional
rlabel metal3 s -746 11582 200662 11642 6 vssd
port 949 nsew ground bidirectional
rlabel metal3 s -746 -762 200662 -702 8 vssd
port 950 nsew ground bidirectional
rlabel metal4 s 200602 -762 200662 11642 6 vssd
port 951 nsew ground bidirectional
rlabel metal4 s 184474 -762 184534 11642 6 vssd
port 952 nsew ground bidirectional
rlabel metal4 s 144474 -762 144534 11642 6 vssd
port 953 nsew ground bidirectional
rlabel metal4 s 104474 -762 104534 11642 6 vssd
port 954 nsew ground bidirectional
rlabel metal4 s 64474 -762 64534 11642 6 vssd
port 955 nsew ground bidirectional
rlabel metal4 s 24474 -762 24534 11642 6 vssd
port 956 nsew ground bidirectional
rlabel metal4 s -746 -762 -686 11642 4 vssd
port 957 nsew ground bidirectional
rlabel metal3 s -886 11722 200802 11782 6 vccd2
port 958 nsew power bidirectional
rlabel metal3 s -886 -902 200802 -842 8 vccd2
port 959 nsew power bidirectional
rlabel metal4 s 164874 -1042 164934 11922 6 vccd2
port 960 nsew power bidirectional
rlabel metal4 s 124874 -1042 124934 11922 6 vccd2
port 961 nsew power bidirectional
rlabel metal4 s 84874 -1042 84934 11922 6 vccd2
port 962 nsew power bidirectional
rlabel metal4 s 44874 -1042 44934 11922 6 vccd2
port 963 nsew power bidirectional
rlabel metal4 s 4874 -1042 4934 11922 6 vccd2
port 964 nsew power bidirectional
rlabel metal4 s 200742 -902 200802 11782 6 vccd2
port 965 nsew power bidirectional
rlabel metal4 s -886 -902 -826 11782 4 vccd2
port 966 nsew power bidirectional
rlabel metal3 s -1026 11862 200942 11922 6 vssd2
port 967 nsew ground bidirectional
rlabel metal3 s -1026 -1042 200942 -982 8 vssd2
port 968 nsew ground bidirectional
rlabel metal4 s 200882 -1042 200942 11922 6 vssd2
port 969 nsew ground bidirectional
rlabel metal4 s 184874 -1042 184934 11922 6 vssd2
port 970 nsew ground bidirectional
rlabel metal4 s 144874 -1042 144934 11922 6 vssd2
port 971 nsew ground bidirectional
rlabel metal4 s 104874 -1042 104934 11922 6 vssd2
port 972 nsew ground bidirectional
rlabel metal4 s 64874 -1042 64934 11922 6 vssd2
port 973 nsew ground bidirectional
rlabel metal4 s 24874 -1042 24934 11922 6 vssd2
port 974 nsew ground bidirectional
rlabel metal4 s -1026 -1042 -966 11922 4 vssd2
port 975 nsew ground bidirectional
rlabel metal3 s -1166 12002 201082 12062 6 vdda1
port 976 nsew power bidirectional
rlabel metal3 s -1166 -1182 201082 -1122 8 vdda1
port 977 nsew power bidirectional
rlabel metal4 s 165274 -1322 165334 12202 6 vdda1
port 978 nsew power bidirectional
rlabel metal4 s 125274 -1322 125334 12202 6 vdda1
port 979 nsew power bidirectional
rlabel metal4 s 85274 -1322 85334 12202 6 vdda1
port 980 nsew power bidirectional
rlabel metal4 s 45274 -1322 45334 12202 6 vdda1
port 981 nsew power bidirectional
rlabel metal4 s 5274 -1322 5334 12202 6 vdda1
port 982 nsew power bidirectional
rlabel metal4 s 201022 -1182 201082 12062 6 vdda1
port 983 nsew power bidirectional
rlabel metal4 s -1166 -1182 -1106 12062 4 vdda1
port 984 nsew power bidirectional
rlabel metal3 s -1306 12142 201222 12202 6 vssa1
port 985 nsew ground bidirectional
rlabel metal3 s -1306 -1322 201222 -1262 8 vssa1
port 986 nsew ground bidirectional
rlabel metal4 s 201162 -1322 201222 12202 6 vssa1
port 987 nsew ground bidirectional
rlabel metal4 s 185274 -1322 185334 12202 6 vssa1
port 988 nsew ground bidirectional
rlabel metal4 s 145274 -1322 145334 12202 6 vssa1
port 989 nsew ground bidirectional
rlabel metal4 s 105274 -1322 105334 12202 6 vssa1
port 990 nsew ground bidirectional
rlabel metal4 s 65274 -1322 65334 12202 6 vssa1
port 991 nsew ground bidirectional
rlabel metal4 s 25274 -1322 25334 12202 6 vssa1
port 992 nsew ground bidirectional
rlabel metal4 s -1306 -1322 -1246 12202 4 vssa1
port 993 nsew ground bidirectional
rlabel metal3 s -1446 12282 201362 12342 6 vdda2
port 994 nsew power bidirectional
rlabel metal3 s -1446 -1462 201362 -1402 8 vdda2
port 995 nsew power bidirectional
rlabel metal4 s 165674 -1602 165734 12482 6 vdda2
port 996 nsew power bidirectional
rlabel metal4 s 125674 -1602 125734 12482 6 vdda2
port 997 nsew power bidirectional
rlabel metal4 s 85674 -1602 85734 12482 6 vdda2
port 998 nsew power bidirectional
rlabel metal4 s 45674 -1602 45734 12482 6 vdda2
port 999 nsew power bidirectional
rlabel metal4 s 5674 -1602 5734 12482 6 vdda2
port 1000 nsew power bidirectional
rlabel metal4 s 201302 -1462 201362 12342 6 vdda2
port 1001 nsew power bidirectional
rlabel metal4 s -1446 -1462 -1386 12342 4 vdda2
port 1002 nsew power bidirectional
rlabel metal3 s -1586 12422 201502 12482 6 vssa2
port 1003 nsew ground bidirectional
rlabel metal3 s -1586 -1602 201502 -1542 8 vssa2
port 1004 nsew ground bidirectional
rlabel metal4 s 201442 -1602 201502 12482 6 vssa2
port 1005 nsew ground bidirectional
rlabel metal4 s 185674 -1602 185734 12482 6 vssa2
port 1006 nsew ground bidirectional
rlabel metal4 s 145674 -1602 145734 12482 6 vssa2
port 1007 nsew ground bidirectional
rlabel metal4 s 105674 -1602 105734 12482 6 vssa2
port 1008 nsew ground bidirectional
rlabel metal4 s 65674 -1602 65734 12482 6 vssa2
port 1009 nsew ground bidirectional
rlabel metal4 s 25674 -1602 25734 12482 6 vssa2
port 1010 nsew ground bidirectional
rlabel metal4 s -1586 -1602 -1526 12482 4 vssa2
port 1011 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 200000 11000
string LEFview TRUE
string GDS_FILE /project/openlane/mgmt_protect/runs/mgmt_protect/results/magic/mgmt_protect.gds
string GDS_END 3254710
string GDS_START 147958
<< end >>

