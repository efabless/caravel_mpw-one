magic
tech sky130A
magscale 1 2
timestamp 1625173925
<< checkpaint >>
rect 426855 1038860 447918 1043510
rect -2260 1035309 719860 1038860
rect -2260 1033509 724107 1035309
rect -2260 38357 724807 1033509
rect -2260 38047 724797 38357
rect -2260 24157 724107 38047
rect -2260 -1260 719860 24157
<< metal1 >>
rect 483664 1005153 483670 1005205
rect 483722 1005193 483728 1005205
rect 529840 1005193 529846 1005205
rect 483722 1005165 529846 1005193
rect 483722 1005153 483728 1005165
rect 529840 1005153 529846 1005165
rect 529898 1005153 529904 1005205
rect 535024 1005153 535030 1005205
rect 535082 1005193 535088 1005205
rect 561616 1005193 561622 1005205
rect 535082 1005165 561622 1005193
rect 535082 1005153 535088 1005165
rect 561616 1005153 561622 1005165
rect 561674 1005153 561680 1005205
rect 636880 1005153 636886 1005205
rect 636938 1005193 636944 1005205
rect 649360 1005193 649366 1005205
rect 636938 1005165 649366 1005193
rect 636938 1005153 636944 1005165
rect 649360 1005153 649366 1005165
rect 649418 1005153 649424 1005205
rect 529840 999381 529846 999433
rect 529898 999421 529904 999433
rect 529898 999393 529982 999421
rect 529898 999381 529904 999393
rect 529954 999347 529982 999393
rect 561616 999381 561622 999433
rect 561674 999421 561680 999433
rect 571888 999421 571894 999433
rect 561674 999393 571894 999421
rect 561674 999381 561680 999393
rect 571888 999381 571894 999393
rect 571946 999381 571952 999433
rect 532816 999347 532822 999359
rect 529954 999319 532822 999347
rect 532816 999307 532822 999319
rect 532874 999307 532880 999359
rect 484600 982817 529831 982845
rect 536290 982817 623523 982845
rect 633564 982817 647057 982845
rect 655408 892969 655414 893021
rect 655466 893009 655472 893021
rect 676240 893009 676246 893021
rect 655466 892981 676246 893009
rect 655466 892969 655472 892981
rect 676240 892969 676246 892981
rect 676298 892969 676304 893021
rect 655216 892895 655222 892947
rect 655274 892935 655280 892947
rect 676144 892935 676150 892947
rect 655274 892907 676150 892935
rect 655274 892895 655280 892907
rect 676144 892895 676150 892907
rect 676202 892895 676208 892947
rect 655120 892821 655126 892873
rect 655178 892861 655184 892873
rect 676048 892861 676054 892873
rect 655178 892833 676054 892861
rect 655178 892821 655184 892833
rect 676048 892821 676054 892833
rect 676106 892821 676112 892873
rect 673840 892377 673846 892429
rect 673898 892417 673904 892429
rect 676048 892417 676054 892429
rect 673898 892389 676054 892417
rect 673898 892377 673904 892389
rect 676048 892377 676054 892389
rect 676106 892377 676112 892429
rect 670960 891415 670966 891467
rect 671018 891455 671024 891467
rect 676048 891455 676054 891467
rect 671018 891427 676054 891455
rect 671018 891415 671024 891427
rect 676048 891415 676054 891427
rect 676106 891415 676112 891467
rect 670864 890379 670870 890431
rect 670922 890419 670928 890431
rect 676048 890419 676054 890431
rect 670922 890391 676054 890419
rect 670922 890379 670928 890391
rect 676048 890379 676054 890391
rect 676106 890379 676112 890431
rect 674032 887863 674038 887915
rect 674090 887903 674096 887915
rect 676240 887903 676246 887915
rect 674090 887875 676246 887903
rect 674090 887863 674096 887875
rect 676240 887863 676246 887875
rect 676298 887863 676304 887915
rect 674224 887123 674230 887175
rect 674282 887163 674288 887175
rect 676048 887163 676054 887175
rect 674282 887135 676054 887163
rect 674282 887123 674288 887135
rect 676048 887123 676054 887135
rect 676106 887123 676112 887175
rect 674416 887049 674422 887101
rect 674474 887089 674480 887101
rect 676240 887089 676246 887101
rect 674474 887061 676246 887089
rect 674474 887049 674480 887061
rect 676240 887049 676246 887061
rect 676298 887049 676304 887101
rect 674128 885051 674134 885103
rect 674186 885091 674192 885103
rect 676048 885091 676054 885103
rect 674186 885063 676054 885091
rect 674186 885051 674192 885063
rect 676048 885051 676054 885063
rect 676106 885051 676112 885103
rect 674320 884237 674326 884289
rect 674378 884277 674384 884289
rect 676048 884277 676054 884289
rect 674378 884249 676054 884277
rect 674378 884237 674384 884249
rect 676048 884237 676054 884249
rect 676106 884237 676112 884289
rect 674896 884163 674902 884215
rect 674954 884203 674960 884215
rect 676240 884203 676246 884215
rect 674954 884175 676246 884203
rect 674954 884163 674960 884175
rect 676240 884163 676246 884175
rect 676298 884163 676304 884215
rect 675280 883201 675286 883253
rect 675338 883241 675344 883253
rect 679984 883241 679990 883253
rect 675338 883213 679990 883241
rect 675338 883201 675344 883213
rect 679984 883201 679990 883213
rect 680042 883201 680048 883253
rect 674512 883053 674518 883105
rect 674570 883093 674576 883105
rect 680176 883093 680182 883105
rect 674570 883065 680182 883093
rect 674570 883053 674576 883065
rect 680176 883053 680182 883065
rect 680234 883053 680240 883105
rect 674992 882831 674998 882883
rect 675050 882871 675056 882883
rect 679696 882871 679702 882883
rect 675050 882843 679702 882871
rect 675050 882831 675056 882843
rect 679696 882831 679702 882843
rect 679754 882831 679760 882883
rect 674704 881499 674710 881551
rect 674762 881539 674768 881551
rect 675952 881539 675958 881551
rect 674762 881511 675958 881539
rect 674762 881499 674768 881511
rect 675952 881499 675958 881511
rect 676010 881499 676016 881551
rect 649456 881425 649462 881477
rect 649514 881465 649520 881477
rect 679696 881465 679702 881477
rect 649514 881437 679702 881465
rect 649514 881425 649520 881437
rect 679696 881425 679702 881437
rect 679754 881425 679760 881477
rect 655312 881351 655318 881403
rect 655370 881391 655376 881403
rect 675472 881391 675478 881403
rect 655370 881363 675478 881391
rect 655370 881351 655376 881363
rect 675472 881351 675478 881363
rect 675530 881351 675536 881403
rect 674800 881277 674806 881329
rect 674858 881317 674864 881329
rect 676048 881317 676054 881329
rect 674858 881289 676054 881317
rect 674858 881277 674864 881289
rect 676048 881277 676054 881289
rect 676106 881277 676112 881329
rect 674608 881203 674614 881255
rect 674666 881243 674672 881255
rect 680080 881243 680086 881255
rect 674666 881215 680086 881243
rect 674666 881203 674672 881215
rect 680080 881203 680086 881215
rect 680138 881203 680144 881255
rect 675184 880093 675190 880145
rect 675242 880133 675248 880145
rect 679792 880133 679798 880145
rect 675242 880105 679798 880133
rect 675242 880093 675248 880105
rect 679792 880093 679798 880105
rect 679850 880093 679856 880145
rect 679888 878505 679894 878517
rect 675106 878477 679894 878505
rect 675106 877999 675134 878477
rect 679888 878465 679894 878477
rect 679946 878465 679952 878517
rect 675088 877947 675094 877999
rect 675146 877947 675152 877999
rect 674992 877207 674998 877259
rect 675050 877247 675056 877259
rect 675472 877247 675478 877259
rect 675050 877219 675478 877247
rect 675050 877207 675056 877219
rect 675472 877207 675478 877219
rect 675530 877207 675536 877259
rect 674608 876689 674614 876741
rect 674666 876729 674672 876741
rect 675280 876729 675286 876741
rect 674666 876701 675286 876729
rect 674666 876689 674672 876701
rect 675280 876689 675286 876701
rect 675338 876689 675344 876741
rect 674512 876615 674518 876667
rect 674570 876655 674576 876667
rect 675376 876655 675382 876667
rect 674570 876627 675382 876655
rect 674570 876615 674576 876627
rect 675376 876615 675382 876627
rect 675434 876615 675440 876667
rect 674224 876393 674230 876445
rect 674282 876433 674288 876445
rect 674512 876433 674518 876445
rect 674282 876405 674518 876433
rect 674282 876393 674288 876405
rect 674512 876393 674518 876405
rect 674570 876393 674576 876445
rect 674032 876245 674038 876297
rect 674090 876285 674096 876297
rect 674224 876285 674230 876297
rect 674090 876257 674230 876285
rect 674090 876245 674096 876257
rect 674224 876245 674230 876257
rect 674282 876245 674288 876297
rect 674800 872989 674806 873041
rect 674858 873029 674864 873041
rect 675280 873029 675286 873041
rect 674858 873001 675286 873029
rect 674858 872989 674864 873001
rect 675280 872989 675286 873001
rect 675338 872989 675344 873041
rect 674704 872915 674710 872967
rect 674762 872955 674768 872967
rect 675184 872955 675190 872967
rect 674762 872927 675190 872955
rect 674762 872915 674768 872927
rect 675184 872915 675190 872927
rect 675242 872915 675248 872967
rect 654160 872619 654166 872671
rect 654218 872659 654224 872671
rect 675088 872659 675094 872671
rect 654218 872631 675094 872659
rect 654218 872619 654224 872631
rect 675088 872619 675094 872631
rect 675146 872619 675152 872671
rect 674608 870547 674614 870599
rect 674666 870587 674672 870599
rect 675472 870587 675478 870599
rect 674666 870559 675478 870587
rect 674666 870547 674672 870559
rect 675472 870547 675478 870559
rect 675530 870547 675536 870599
rect 674320 869733 674326 869785
rect 674378 869773 674384 869785
rect 675280 869773 675286 869785
rect 674378 869745 675286 869773
rect 674378 869733 674384 869745
rect 675280 869733 675286 869745
rect 675338 869733 675344 869785
rect 674512 869659 674518 869711
rect 674570 869699 674576 869711
rect 674992 869699 674998 869711
rect 674570 869671 674998 869699
rect 674570 869659 674576 869671
rect 674992 869659 674998 869671
rect 675050 869659 675056 869711
rect 674128 867365 674134 867417
rect 674186 867405 674192 867417
rect 675472 867405 675478 867417
rect 674186 867377 675478 867405
rect 674186 867365 674192 867377
rect 675472 867365 675478 867377
rect 675530 867365 675536 867417
rect 674224 865737 674230 865789
rect 674282 865777 674288 865789
rect 675184 865777 675190 865789
rect 674282 865749 675190 865777
rect 674282 865737 674288 865749
rect 675184 865737 675190 865749
rect 675242 865737 675248 865789
rect 653776 863961 653782 864013
rect 653834 864001 653840 864013
rect 675088 864001 675094 864013
rect 653834 863973 675094 864001
rect 653834 863961 653840 863973
rect 675088 863961 675094 863973
rect 675146 863961 675152 864013
rect 41776 817933 41782 817985
rect 41834 817973 41840 817985
rect 47440 817973 47446 817985
rect 41834 817945 47446 817973
rect 41834 817933 41840 817945
rect 47440 817933 47446 817945
rect 47498 817933 47504 817985
rect 41776 817267 41782 817319
rect 41834 817307 41840 817319
rect 44848 817307 44854 817319
rect 41834 817279 44854 817307
rect 41834 817267 41840 817279
rect 44848 817267 44854 817279
rect 44906 817267 44912 817319
rect 41584 816527 41590 816579
rect 41642 816567 41648 816579
rect 44944 816567 44950 816579
rect 41642 816539 44950 816567
rect 41642 816527 41648 816539
rect 44944 816527 44950 816539
rect 45002 816527 45008 816579
rect 41776 815787 41782 815839
rect 41834 815827 41840 815839
rect 43216 815827 43222 815839
rect 41834 815799 43222 815827
rect 41834 815787 41840 815799
rect 43216 815787 43222 815799
rect 43274 815787 43280 815839
rect 41776 814825 41782 814877
rect 41834 814865 41840 814877
rect 44656 814865 44662 814877
rect 41834 814837 44662 814865
rect 41834 814825 41840 814837
rect 44656 814825 44662 814837
rect 44714 814825 44720 814877
rect 41584 813567 41590 813619
rect 41642 813607 41648 813619
rect 44752 813607 44758 813619
rect 41642 813579 44758 813607
rect 41642 813567 41648 813579
rect 44752 813567 44758 813579
rect 44810 813567 44816 813619
rect 41584 812383 41590 812435
rect 41642 812423 41648 812435
rect 42640 812423 42646 812435
rect 41642 812395 42646 812423
rect 41642 812383 41648 812395
rect 42640 812383 42646 812395
rect 42698 812383 42704 812435
rect 41776 809423 41782 809475
rect 41834 809463 41840 809475
rect 43024 809463 43030 809475
rect 41834 809435 43030 809463
rect 41834 809423 41840 809435
rect 43024 809423 43030 809435
rect 43082 809423 43088 809475
rect 41584 807055 41590 807107
rect 41642 807095 41648 807107
rect 42928 807095 42934 807107
rect 41642 807067 42934 807095
rect 41642 807055 41648 807067
rect 42928 807055 42934 807067
rect 42986 807055 42992 807107
rect 41968 806981 41974 807033
rect 42026 807021 42032 807033
rect 43120 807021 43126 807033
rect 42026 806993 43126 807021
rect 42026 806981 42032 806993
rect 43120 806981 43126 806993
rect 43178 806981 43184 807033
rect 41584 806611 41590 806663
rect 41642 806651 41648 806663
rect 42640 806651 42646 806663
rect 41642 806623 42646 806651
rect 41642 806611 41648 806623
rect 42640 806611 42646 806623
rect 42698 806611 42704 806663
rect 41776 806389 41782 806441
rect 41834 806429 41840 806441
rect 42736 806429 42742 806441
rect 41834 806401 42742 806429
rect 41834 806389 41840 806401
rect 42736 806389 42742 806401
rect 42794 806389 42800 806441
rect 41584 805131 41590 805183
rect 41642 805171 41648 805183
rect 44560 805171 44566 805183
rect 41642 805143 44566 805171
rect 41642 805131 41648 805143
rect 44560 805131 44566 805143
rect 44618 805131 44624 805183
rect 42352 800691 42358 800743
rect 42410 800731 42416 800743
rect 57712 800731 57718 800743
rect 42410 800703 57718 800731
rect 42410 800691 42416 800703
rect 57712 800691 57718 800703
rect 57770 800691 57776 800743
rect 42448 800617 42454 800669
rect 42506 800657 42512 800669
rect 57616 800657 57622 800669
rect 42506 800629 57622 800657
rect 42506 800617 42512 800629
rect 57616 800617 57622 800629
rect 57674 800617 57680 800669
rect 41968 800173 41974 800225
rect 42026 800173 42032 800225
rect 41986 800003 42014 800173
rect 41968 799951 41974 800003
rect 42026 799951 42032 800003
rect 42352 796843 42358 796895
rect 42410 796883 42416 796895
rect 42736 796883 42742 796895
rect 42410 796855 42742 796883
rect 42410 796843 42416 796855
rect 42736 796843 42742 796855
rect 42794 796843 42800 796895
rect 42544 795067 42550 795119
rect 42602 795067 42608 795119
rect 42562 794897 42590 795067
rect 42544 794845 42550 794897
rect 42602 794845 42608 794897
rect 42448 794401 42454 794453
rect 42506 794441 42512 794453
rect 42832 794441 42838 794453
rect 42506 794413 42838 794441
rect 42506 794401 42512 794413
rect 42832 794401 42838 794413
rect 42890 794401 42896 794453
rect 42064 794253 42070 794305
rect 42122 794293 42128 794305
rect 42928 794293 42934 794305
rect 42122 794265 42934 794293
rect 42122 794253 42128 794265
rect 42928 794253 42934 794265
rect 42986 794253 42992 794305
rect 42448 793143 42454 793195
rect 42506 793183 42512 793195
rect 43024 793183 43030 793195
rect 42506 793155 43030 793183
rect 42506 793143 42512 793155
rect 43024 793143 43030 793155
rect 43082 793143 43088 793195
rect 655120 792033 655126 792085
rect 655178 792073 655184 792085
rect 675376 792073 675382 792085
rect 655178 792045 675382 792073
rect 655178 792033 655184 792045
rect 675376 792033 675382 792045
rect 675434 792033 675440 792085
rect 42160 790627 42166 790679
rect 42218 790667 42224 790679
rect 43120 790667 43126 790679
rect 42218 790639 43126 790667
rect 42218 790627 42224 790639
rect 43120 790627 43126 790639
rect 43178 790627 43184 790679
rect 42160 790109 42166 790161
rect 42218 790149 42224 790161
rect 42832 790149 42838 790161
rect 42218 790121 42838 790149
rect 42218 790109 42224 790121
rect 42832 790109 42838 790121
rect 42890 790109 42896 790161
rect 42160 789443 42166 789495
rect 42218 789483 42224 789495
rect 42736 789483 42742 789495
rect 42218 789455 42742 789483
rect 42218 789443 42224 789455
rect 42736 789443 42742 789455
rect 42794 789443 42800 789495
rect 42448 789147 42454 789199
rect 42506 789187 42512 789199
rect 58192 789187 58198 789199
rect 42506 789159 58198 789187
rect 42506 789147 42512 789159
rect 58192 789147 58198 789159
rect 58250 789147 58256 789199
rect 44944 789073 44950 789125
rect 45002 789113 45008 789125
rect 58384 789113 58390 789125
rect 45002 789085 58390 789113
rect 45002 789073 45008 789085
rect 58384 789073 58390 789085
rect 58442 789073 58448 789125
rect 42160 788703 42166 788755
rect 42218 788743 42224 788755
rect 42640 788743 42646 788755
rect 42218 788715 42646 788743
rect 42218 788703 42224 788715
rect 42640 788703 42646 788715
rect 42698 788703 42704 788755
rect 42160 787001 42166 787053
rect 42218 787041 42224 787053
rect 42544 787041 42550 787053
rect 42218 787013 42550 787041
rect 42218 787001 42224 787013
rect 42544 787001 42550 787013
rect 42602 787001 42608 787053
rect 42160 786409 42166 786461
rect 42218 786449 42224 786461
rect 42352 786449 42358 786461
rect 42218 786421 42358 786449
rect 42218 786409 42224 786421
rect 42352 786409 42358 786421
rect 42410 786409 42416 786461
rect 44848 785521 44854 785573
rect 44906 785561 44912 785573
rect 59152 785561 59158 785573
rect 44906 785533 59158 785561
rect 44906 785521 44912 785533
rect 59152 785521 59158 785533
rect 59210 785521 59216 785573
rect 47440 785373 47446 785425
rect 47498 785413 47504 785425
rect 59632 785413 59638 785425
rect 47498 785385 59638 785413
rect 47498 785373 47504 785385
rect 59632 785373 59638 785385
rect 59690 785373 59696 785425
rect 656560 783375 656566 783427
rect 656618 783415 656624 783427
rect 675184 783415 675190 783427
rect 656618 783387 675190 783415
rect 656618 783375 656624 783387
rect 675184 783375 675190 783387
rect 675242 783375 675248 783427
rect 654352 780489 654358 780541
rect 654410 780529 654416 780541
rect 675088 780529 675094 780541
rect 654410 780501 675094 780529
rect 654410 780489 654416 780501
rect 675088 780489 675094 780501
rect 675146 780489 675152 780541
rect 674896 778565 674902 778617
rect 674954 778605 674960 778617
rect 675280 778605 675286 778617
rect 674954 778577 675286 778605
rect 674954 778565 674960 778577
rect 675280 778565 675286 778577
rect 675338 778565 675344 778617
rect 674800 777307 674806 777359
rect 674858 777347 674864 777359
rect 675472 777347 675478 777359
rect 674858 777319 675478 777347
rect 674858 777307 674864 777319
rect 675472 777307 675478 777319
rect 675530 777307 675536 777359
rect 41776 774643 41782 774695
rect 41834 774683 41840 774695
rect 47440 774683 47446 774695
rect 41834 774655 47446 774683
rect 41834 774643 41840 774655
rect 47440 774643 47446 774655
rect 47498 774643 47504 774695
rect 674320 774273 674326 774325
rect 674378 774313 674384 774325
rect 675088 774313 675094 774325
rect 674378 774285 675094 774313
rect 674378 774273 674384 774285
rect 675088 774273 675094 774285
rect 675146 774273 675152 774325
rect 41584 773903 41590 773955
rect 41642 773943 41648 773955
rect 44944 773943 44950 773955
rect 41642 773915 44950 773943
rect 41642 773903 41648 773915
rect 44944 773903 44950 773915
rect 45002 773903 45008 773955
rect 41776 773459 41782 773511
rect 41834 773499 41840 773511
rect 45040 773499 45046 773511
rect 41834 773471 45046 773499
rect 41834 773459 41840 773471
rect 45040 773459 45046 773471
rect 45098 773459 45104 773511
rect 41584 773385 41590 773437
rect 41642 773425 41648 773437
rect 43216 773425 43222 773437
rect 41642 773397 43222 773425
rect 41642 773385 41648 773397
rect 43216 773385 43222 773397
rect 43274 773385 43280 773437
rect 41776 772571 41782 772623
rect 41834 772611 41840 772623
rect 43216 772611 43222 772623
rect 41834 772583 43222 772611
rect 41834 772571 41840 772583
rect 43216 772571 43222 772583
rect 43274 772571 43280 772623
rect 43120 772127 43126 772179
rect 43178 772167 43184 772179
rect 62032 772167 62038 772179
rect 43178 772139 62038 772167
rect 43178 772127 43184 772139
rect 62032 772127 62038 772139
rect 62090 772127 62096 772179
rect 41584 771905 41590 771957
rect 41642 771945 41648 771957
rect 61840 771945 61846 771957
rect 41642 771917 61846 771945
rect 41642 771905 41648 771917
rect 61840 771905 61846 771917
rect 61898 771905 61904 771957
rect 41776 767539 41782 767591
rect 41834 767579 41840 767591
rect 42736 767579 42742 767591
rect 41834 767551 42742 767579
rect 41834 767539 41840 767551
rect 42736 767539 42742 767551
rect 42794 767539 42800 767591
rect 41584 767095 41590 767147
rect 41642 767135 41648 767147
rect 42640 767135 42646 767147
rect 41642 767107 42646 767135
rect 41642 767095 41648 767107
rect 42640 767095 42646 767107
rect 42698 767095 42704 767147
rect 674416 767095 674422 767147
rect 674474 767135 674480 767147
rect 675088 767135 675094 767147
rect 674474 767107 675094 767135
rect 674474 767095 674480 767107
rect 675088 767095 675094 767107
rect 675146 767095 675152 767147
rect 41776 766577 41782 766629
rect 41834 766617 41840 766629
rect 42544 766617 42550 766629
rect 41834 766589 42550 766617
rect 41834 766577 41840 766589
rect 42544 766577 42550 766589
rect 42602 766577 42608 766629
rect 41584 765393 41590 765445
rect 41642 765433 41648 765445
rect 42832 765433 42838 765445
rect 41642 765405 42838 765433
rect 41642 765393 41648 765405
rect 42832 765393 42838 765405
rect 42890 765393 42896 765445
rect 41776 764727 41782 764779
rect 41834 764767 41840 764779
rect 42928 764767 42934 764779
rect 41834 764739 42934 764767
rect 41834 764727 41840 764739
rect 42928 764727 42934 764739
rect 42986 764727 42992 764779
rect 41584 763395 41590 763447
rect 41642 763435 41648 763447
rect 43024 763435 43030 763447
rect 41642 763407 43030 763435
rect 41642 763395 41648 763407
rect 43024 763395 43030 763407
rect 43082 763395 43088 763447
rect 42064 763247 42070 763299
rect 42122 763287 42128 763299
rect 43120 763287 43126 763299
rect 42122 763259 43126 763287
rect 42122 763247 42128 763259
rect 43120 763247 43126 763259
rect 43178 763247 43184 763299
rect 41584 761915 41590 761967
rect 41642 761955 41648 761967
rect 44848 761955 44854 761967
rect 41642 761927 44854 761955
rect 41642 761915 41648 761927
rect 44848 761915 44854 761927
rect 44906 761915 44912 761967
rect 42448 757623 42454 757675
rect 42506 757663 42512 757675
rect 43312 757663 43318 757675
rect 42506 757635 43318 757663
rect 42506 757623 42512 757635
rect 43312 757623 43318 757635
rect 43370 757623 43376 757675
rect 42448 757475 42454 757527
rect 42506 757515 42512 757527
rect 58672 757515 58678 757527
rect 42506 757487 58678 757515
rect 42506 757475 42512 757487
rect 58672 757475 58678 757487
rect 58730 757475 58736 757527
rect 43120 757253 43126 757305
rect 43178 757293 43184 757305
rect 43504 757293 43510 757305
rect 43178 757265 43510 757293
rect 43178 757253 43184 757265
rect 43504 757253 43510 757265
rect 43562 757253 43568 757305
rect 42640 757179 42646 757231
rect 42698 757219 42704 757231
rect 43408 757219 43414 757231
rect 42698 757191 43414 757219
rect 42698 757179 42704 757191
rect 43408 757179 43414 757191
rect 43466 757179 43472 757231
rect 42544 757105 42550 757157
rect 42602 757145 42608 757157
rect 43120 757145 43126 757157
rect 42602 757117 43126 757145
rect 42602 757105 42608 757117
rect 43120 757105 43126 757117
rect 43178 757105 43184 757157
rect 41872 757031 41878 757083
rect 41930 757071 41936 757083
rect 42640 757071 42646 757083
rect 41930 757043 42646 757071
rect 41930 757031 41936 757043
rect 42640 757031 42646 757043
rect 42698 757031 42704 757083
rect 41776 756957 41782 757009
rect 41834 756997 41840 757009
rect 42544 756997 42550 757009
rect 41834 756969 42550 756997
rect 41834 756957 41840 756969
rect 42544 756957 42550 756969
rect 42602 756957 42608 757009
rect 42256 756883 42262 756935
rect 42314 756923 42320 756935
rect 42314 756895 42398 756923
rect 42314 756883 42320 756895
rect 42370 756713 42398 756895
rect 42352 756661 42358 756713
rect 42410 756661 42416 756713
rect 42352 753627 42358 753679
rect 42410 753667 42416 753679
rect 42832 753667 42838 753679
rect 42410 753639 42838 753667
rect 42410 753627 42416 753639
rect 42832 753627 42838 753639
rect 42890 753627 42896 753679
rect 42832 753479 42838 753531
rect 42890 753519 42896 753531
rect 43312 753519 43318 753531
rect 42890 753491 43318 753519
rect 42890 753479 42896 753491
rect 43312 753479 43318 753491
rect 43370 753479 43376 753531
rect 42352 751777 42358 751829
rect 42410 751817 42416 751829
rect 43024 751817 43030 751829
rect 42410 751789 43030 751817
rect 42410 751777 42416 751789
rect 43024 751777 43030 751789
rect 43082 751777 43088 751829
rect 42448 751703 42454 751755
rect 42506 751743 42512 751755
rect 43312 751743 43318 751755
rect 42506 751715 43318 751743
rect 42506 751703 42512 751715
rect 43312 751703 43318 751715
rect 43370 751703 43376 751755
rect 43024 751629 43030 751681
rect 43082 751669 43088 751681
rect 43408 751669 43414 751681
rect 43082 751641 43414 751669
rect 43082 751629 43088 751641
rect 43408 751629 43414 751641
rect 43466 751629 43472 751681
rect 42448 751555 42454 751607
rect 42506 751595 42512 751607
rect 42928 751595 42934 751607
rect 42506 751567 42934 751595
rect 42506 751555 42512 751567
rect 42928 751555 42934 751567
rect 42986 751555 42992 751607
rect 42256 750593 42262 750645
rect 42314 750633 42320 750645
rect 43504 750633 43510 750645
rect 42314 750605 43510 750633
rect 42314 750593 42320 750605
rect 43504 750593 43510 750605
rect 43562 750593 43568 750645
rect 42064 749927 42070 749979
rect 42122 749967 42128 749979
rect 42736 749967 42742 749979
rect 42122 749939 42742 749967
rect 42122 749927 42128 749939
rect 42736 749927 42742 749939
rect 42794 749927 42800 749979
rect 655696 748817 655702 748869
rect 655754 748857 655760 748869
rect 675376 748857 675382 748869
rect 655754 748829 675382 748857
rect 655754 748817 655760 748829
rect 675376 748817 675382 748829
rect 675434 748817 675440 748869
rect 42064 746079 42070 746131
rect 42122 746119 42128 746131
rect 43120 746119 43126 746131
rect 42122 746091 43126 746119
rect 42122 746079 42128 746091
rect 43120 746079 43126 746091
rect 43178 746079 43184 746131
rect 42640 745931 42646 745983
rect 42698 745971 42704 745983
rect 54640 745971 54646 745983
rect 42698 745943 54646 745971
rect 42698 745931 42704 745943
rect 54640 745931 54646 745943
rect 54698 745931 54704 745983
rect 54736 745931 54742 745983
rect 54794 745971 54800 745983
rect 57616 745971 57622 745983
rect 54794 745943 57622 745971
rect 54794 745931 54800 745943
rect 57616 745931 57622 745943
rect 57674 745931 57680 745983
rect 42160 745487 42166 745539
rect 42218 745527 42224 745539
rect 43024 745527 43030 745539
rect 42218 745499 43030 745527
rect 42218 745487 42224 745499
rect 43024 745487 43030 745499
rect 43082 745487 43088 745539
rect 45040 745413 45046 745465
rect 45098 745453 45104 745465
rect 58096 745453 58102 745465
rect 45098 745425 58102 745453
rect 45098 745413 45104 745425
rect 58096 745413 58102 745425
rect 58154 745413 58160 745465
rect 43312 744969 43318 745021
rect 43370 745009 43376 745021
rect 58576 745009 58582 745021
rect 43370 744981 58582 745009
rect 43370 744969 43376 744981
rect 58576 744969 58582 744981
rect 58634 744969 58640 745021
rect 42160 743785 42166 743837
rect 42218 743825 42224 743837
rect 42832 743825 42838 743837
rect 42218 743797 42838 743825
rect 42218 743785 42224 743797
rect 42832 743785 42838 743797
rect 42890 743785 42896 743837
rect 47440 742971 47446 743023
rect 47498 743011 47504 743023
rect 59632 743011 59638 743023
rect 47498 742983 59638 743011
rect 47498 742971 47504 742983
rect 59632 742971 59638 742983
rect 59690 742971 59696 743023
rect 44944 742897 44950 742949
rect 45002 742937 45008 742949
rect 59728 742937 59734 742949
rect 45002 742909 59734 742937
rect 45002 742897 45008 742909
rect 59728 742897 59734 742909
rect 59786 742897 59792 742949
rect 674704 742749 674710 742801
rect 674762 742789 674768 742801
rect 675376 742789 675382 742801
rect 674762 742761 675382 742789
rect 674762 742749 674768 742761
rect 675376 742749 675382 742761
rect 675434 742749 675440 742801
rect 673648 737865 673654 737917
rect 673706 737905 673712 737917
rect 675376 737905 675382 737917
rect 673706 737877 675382 737905
rect 673706 737865 673712 737877
rect 675376 737865 675382 737877
rect 675434 737865 675440 737917
rect 654064 737421 654070 737473
rect 654122 737461 654128 737473
rect 674992 737461 674998 737473
rect 654122 737433 674998 737461
rect 654122 737421 654128 737433
rect 674992 737421 674998 737433
rect 675050 737421 675056 737473
rect 654160 737347 654166 737399
rect 654218 737387 654224 737399
rect 675088 737387 675094 737399
rect 654218 737359 675094 737387
rect 654218 737347 654224 737359
rect 675088 737347 675094 737359
rect 675146 737347 675152 737399
rect 675184 735719 675190 735771
rect 675242 735719 675248 735771
rect 675202 735537 675230 735719
rect 675280 735537 675286 735549
rect 675202 735509 675286 735537
rect 675280 735497 675286 735509
rect 675338 735497 675344 735549
rect 675088 733869 675094 733921
rect 675146 733909 675152 733921
rect 675376 733909 675382 733921
rect 675146 733881 675382 733909
rect 675146 733869 675152 733881
rect 675376 733869 675382 733881
rect 675434 733869 675440 733921
rect 673456 733721 673462 733773
rect 673514 733761 673520 733773
rect 675472 733761 675478 733773
rect 673514 733733 675478 733761
rect 673514 733721 673520 733733
rect 675472 733721 675478 733733
rect 675530 733721 675536 733773
rect 674224 732315 674230 732367
rect 674282 732355 674288 732367
rect 675472 732355 675478 732367
rect 674282 732327 675478 732355
rect 674282 732315 674288 732327
rect 675472 732315 675478 732327
rect 675530 732315 675536 732367
rect 674992 732019 674998 732071
rect 675050 732059 675056 732071
rect 675376 732059 675382 732071
rect 675050 732031 675382 732059
rect 675050 732019 675056 732031
rect 675376 732019 675382 732031
rect 675434 732019 675440 732071
rect 41776 731427 41782 731479
rect 41834 731467 41840 731479
rect 47536 731467 47542 731479
rect 41834 731439 47542 731467
rect 41834 731427 41840 731439
rect 47536 731427 47542 731439
rect 47594 731427 47600 731479
rect 41584 730687 41590 730739
rect 41642 730727 41648 730739
rect 44944 730727 44950 730739
rect 41642 730699 44950 730727
rect 41642 730687 41648 730699
rect 44944 730687 44950 730699
rect 45002 730687 45008 730739
rect 674704 730465 674710 730517
rect 674762 730505 674768 730517
rect 675472 730505 675478 730517
rect 674762 730477 675478 730505
rect 674762 730465 674768 730477
rect 675472 730465 675478 730477
rect 675530 730465 675536 730517
rect 41776 730317 41782 730369
rect 41834 730357 41840 730369
rect 45040 730357 45046 730369
rect 41834 730329 45046 730357
rect 41834 730317 41840 730329
rect 45040 730317 45046 730329
rect 45098 730317 45104 730369
rect 41584 730169 41590 730221
rect 41642 730209 41648 730221
rect 43216 730209 43222 730221
rect 41642 730181 43222 730209
rect 41642 730169 41648 730181
rect 43216 730169 43222 730181
rect 43274 730169 43280 730221
rect 41776 729355 41782 729407
rect 41834 729395 41840 729407
rect 43504 729395 43510 729407
rect 41834 729367 43510 729395
rect 41834 729355 41840 729367
rect 43504 729355 43510 729367
rect 43562 729355 43568 729407
rect 41776 728763 41782 728815
rect 41834 728803 41840 728815
rect 43312 728803 43318 728815
rect 41834 728775 43318 728803
rect 41834 728763 41840 728775
rect 43312 728763 43318 728775
rect 43370 728763 43376 728815
rect 40432 728689 40438 728741
rect 40490 728729 40496 728741
rect 62224 728729 62230 728741
rect 40490 728701 62230 728729
rect 40490 728689 40496 728701
rect 62224 728689 62230 728701
rect 62282 728689 62288 728741
rect 42256 728615 42262 728667
rect 42314 728655 42320 728667
rect 62416 728655 62422 728667
rect 42314 728627 62422 728655
rect 42314 728615 42320 728627
rect 62416 728615 62422 728627
rect 62474 728615 62480 728667
rect 674608 728615 674614 728667
rect 674666 728655 674672 728667
rect 675376 728655 675382 728667
rect 674666 728627 675382 728655
rect 674666 728615 674672 728627
rect 675376 728615 675382 728627
rect 675434 728615 675440 728667
rect 41776 727875 41782 727927
rect 41834 727915 41840 727927
rect 43408 727915 43414 727927
rect 41834 727887 43414 727915
rect 41834 727875 41840 727887
rect 43408 727875 43414 727887
rect 43466 727875 43472 727927
rect 41776 726543 41782 726595
rect 41834 726583 41840 726595
rect 42928 726583 42934 726595
rect 41834 726555 42934 726583
rect 41834 726543 41840 726555
rect 42928 726543 42934 726555
rect 42986 726543 42992 726595
rect 41776 726395 41782 726447
rect 41834 726435 41840 726447
rect 42832 726435 42838 726447
rect 41834 726407 42838 726435
rect 41834 726395 41840 726407
rect 42832 726395 42838 726407
rect 42890 726395 42896 726447
rect 41776 722991 41782 723043
rect 41834 723031 41840 723043
rect 43024 723031 43030 723043
rect 41834 723003 43030 723031
rect 41834 722991 41840 723003
rect 43024 722991 43030 723003
rect 43082 722991 43088 723043
rect 673840 722917 673846 722969
rect 673898 722957 673904 722969
rect 679696 722957 679702 722969
rect 673898 722929 679702 722957
rect 673898 722917 673904 722929
rect 679696 722917 679702 722929
rect 679754 722917 679760 722969
rect 41584 720919 41590 720971
rect 41642 720959 41648 720971
rect 42544 720959 42550 720971
rect 41642 720931 42550 720959
rect 41642 720919 41648 720931
rect 42544 720919 42550 720931
rect 42602 720919 42608 720971
rect 41776 720549 41782 720601
rect 41834 720589 41840 720601
rect 43120 720589 43126 720601
rect 41834 720561 43126 720589
rect 41834 720549 41840 720561
rect 43120 720549 43126 720561
rect 43178 720549 43184 720601
rect 41584 720327 41590 720379
rect 41642 720367 41648 720379
rect 42640 720367 42646 720379
rect 41642 720339 42646 720367
rect 41642 720327 41648 720339
rect 42640 720327 42646 720339
rect 42698 720327 42704 720379
rect 41776 720179 41782 720231
rect 41834 720219 41840 720231
rect 42736 720219 42742 720231
rect 41834 720191 42742 720219
rect 41834 720179 41840 720191
rect 42736 720179 42742 720191
rect 42794 720179 42800 720231
rect 41584 718699 41590 718751
rect 41642 718739 41648 718751
rect 47440 718739 47446 718751
rect 41642 718711 47446 718739
rect 41642 718699 41648 718711
rect 47440 718699 47446 718711
rect 47498 718699 47504 718751
rect 655600 714703 655606 714755
rect 655658 714743 655664 714755
rect 676240 714743 676246 714755
rect 655658 714715 676246 714743
rect 655658 714703 655664 714715
rect 676240 714703 676246 714715
rect 676298 714703 676304 714755
rect 655408 714555 655414 714607
rect 655466 714595 655472 714607
rect 676144 714595 676150 714607
rect 655466 714567 676150 714595
rect 655466 714555 655472 714567
rect 676144 714555 676150 714567
rect 676202 714555 676208 714607
rect 655216 714407 655222 714459
rect 655274 714447 655280 714459
rect 676336 714447 676342 714459
rect 655274 714419 676342 714447
rect 655274 714407 655280 714419
rect 676336 714407 676342 714419
rect 676394 714407 676400 714459
rect 42352 714259 42358 714311
rect 42410 714299 42416 714311
rect 59632 714299 59638 714311
rect 42410 714271 59638 714299
rect 42410 714259 42416 714271
rect 59632 714259 59638 714271
rect 59690 714259 59696 714311
rect 41968 713889 41974 713941
rect 42026 713929 42032 713941
rect 43216 713929 43222 713941
rect 42026 713901 43222 713929
rect 42026 713889 42032 713901
rect 43216 713889 43222 713901
rect 43274 713889 43280 713941
rect 41776 713815 41782 713867
rect 41834 713815 41840 713867
rect 41872 713815 41878 713867
rect 41930 713855 41936 713867
rect 43600 713855 43606 713867
rect 41930 713827 43606 713855
rect 41930 713815 41936 713827
rect 43600 713815 43606 713827
rect 43658 713815 43664 713867
rect 41794 713781 41822 713815
rect 41794 713753 42206 713781
rect 42178 712819 42206 713753
rect 669712 713075 669718 713127
rect 669770 713115 669776 713127
rect 670960 713115 670966 713127
rect 669770 713087 670966 713115
rect 669770 713075 669776 713087
rect 670960 713075 670966 713087
rect 671018 713115 671024 713127
rect 676048 713115 676054 713127
rect 671018 713087 676054 713115
rect 671018 713075 671024 713087
rect 676048 713075 676054 713087
rect 676106 713075 676112 713127
rect 42256 712853 42262 712905
rect 42314 712893 42320 712905
rect 42832 712893 42838 712905
rect 42314 712865 42838 712893
rect 42314 712853 42320 712865
rect 42832 712853 42838 712865
rect 42890 712853 42896 712905
rect 42178 712791 42878 712819
rect 42850 712757 42878 712791
rect 42832 712705 42838 712757
rect 42890 712705 42896 712757
rect 670672 712631 670678 712683
rect 670730 712671 670736 712683
rect 676048 712671 676054 712683
rect 670730 712643 676054 712671
rect 670730 712631 670736 712643
rect 676048 712631 676054 712643
rect 676106 712631 676112 712683
rect 669520 711891 669526 711943
rect 669578 711931 669584 711943
rect 670864 711931 670870 711943
rect 669578 711903 670870 711931
rect 669578 711891 669584 711903
rect 670864 711891 670870 711903
rect 670922 711931 670928 711943
rect 676240 711931 676246 711943
rect 670922 711903 676246 711931
rect 670922 711891 670928 711903
rect 676240 711891 676246 711903
rect 676298 711891 676304 711943
rect 42160 711669 42166 711721
rect 42218 711709 42224 711721
rect 42928 711709 42934 711721
rect 42218 711681 42934 711709
rect 42218 711669 42224 711681
rect 42928 711669 42934 711681
rect 42986 711669 42992 711721
rect 43216 711595 43222 711647
rect 43274 711595 43280 711647
rect 42256 711447 42262 711499
rect 42314 711487 42320 711499
rect 42314 711459 42398 711487
rect 42314 711447 42320 711459
rect 42370 711425 42398 711459
rect 42352 711373 42358 711425
rect 42410 711373 42416 711425
rect 43024 711373 43030 711425
rect 43082 711413 43088 711425
rect 43234 711413 43262 711595
rect 670576 711521 670582 711573
rect 670634 711561 670640 711573
rect 676048 711561 676054 711573
rect 670634 711533 676054 711561
rect 670634 711521 670640 711533
rect 676048 711521 676054 711533
rect 676106 711521 676112 711573
rect 43082 711385 43262 711413
rect 43082 711373 43088 711385
rect 43312 711373 43318 711425
rect 43370 711413 43376 711425
rect 43504 711413 43510 711425
rect 43370 711385 43510 711413
rect 43370 711373 43376 711385
rect 43504 711373 43510 711385
rect 43562 711373 43568 711425
rect 42160 711299 42166 711351
rect 42218 711339 42224 711351
rect 42218 711311 42878 711339
rect 42218 711299 42224 711311
rect 42850 711277 42878 711311
rect 42928 711299 42934 711351
rect 42986 711299 42992 711351
rect 674320 711299 674326 711351
rect 674378 711339 674384 711351
rect 676048 711339 676054 711351
rect 674378 711311 676054 711339
rect 674378 711299 674384 711311
rect 676048 711299 676054 711311
rect 676106 711299 676112 711351
rect 42832 711225 42838 711277
rect 42890 711225 42896 711277
rect 42256 711077 42262 711129
rect 42314 711117 42320 711129
rect 42946 711117 42974 711299
rect 42314 711089 42974 711117
rect 42314 711077 42320 711089
rect 42160 710855 42166 710907
rect 42218 710895 42224 710907
rect 42448 710895 42454 710907
rect 42218 710867 42454 710895
rect 42218 710855 42224 710867
rect 42448 710855 42454 710867
rect 42506 710855 42512 710907
rect 674416 710485 674422 710537
rect 674474 710525 674480 710537
rect 676048 710525 676054 710537
rect 674474 710497 676054 710525
rect 674474 710485 674480 710497
rect 676048 710485 676054 710497
rect 676106 710485 676112 710537
rect 42160 709893 42166 709945
rect 42218 709933 42224 709945
rect 42544 709933 42550 709945
rect 42218 709905 42550 709933
rect 42218 709893 42224 709905
rect 42544 709893 42550 709905
rect 42602 709893 42608 709945
rect 42064 708487 42070 708539
rect 42122 708527 42128 708539
rect 43504 708527 43510 708539
rect 42122 708499 43510 708527
rect 42122 708487 42128 708499
rect 43504 708487 43510 708499
rect 43562 708487 43568 708539
rect 675280 708413 675286 708465
rect 675338 708453 675344 708465
rect 676048 708453 676054 708465
rect 675338 708425 676054 708453
rect 675338 708413 675344 708425
rect 676048 708413 676054 708425
rect 676106 708413 676112 708465
rect 42064 708339 42070 708391
rect 42122 708379 42128 708391
rect 42736 708379 42742 708391
rect 42122 708351 42742 708379
rect 42122 708339 42128 708351
rect 42736 708339 42742 708351
rect 42794 708339 42800 708391
rect 674896 708339 674902 708391
rect 674954 708379 674960 708391
rect 676240 708379 676246 708391
rect 674954 708351 676246 708379
rect 674954 708339 674960 708351
rect 676240 708339 676246 708351
rect 676298 708339 676304 708391
rect 42256 708191 42262 708243
rect 42314 708231 42320 708243
rect 42736 708231 42742 708243
rect 42314 708203 42742 708231
rect 42314 708191 42320 708203
rect 42736 708191 42742 708203
rect 42794 708191 42800 708243
rect 42448 708043 42454 708095
rect 42506 708083 42512 708095
rect 43120 708083 43126 708095
rect 42506 708055 43126 708083
rect 42506 708043 42512 708055
rect 43120 708043 43126 708055
rect 43178 708043 43184 708095
rect 674800 708043 674806 708095
rect 674858 708083 674864 708095
rect 676048 708083 676054 708095
rect 674858 708055 676054 708083
rect 674858 708043 674864 708055
rect 676048 708043 676054 708055
rect 676106 708043 676112 708095
rect 43120 707895 43126 707947
rect 43178 707935 43184 707947
rect 43600 707935 43606 707947
rect 43178 707907 43606 707935
rect 43178 707895 43184 707907
rect 43600 707895 43606 707907
rect 43658 707895 43664 707947
rect 42448 707377 42454 707429
rect 42506 707417 42512 707429
rect 42640 707417 42646 707429
rect 42506 707389 42646 707417
rect 42506 707377 42512 707389
rect 42640 707377 42646 707389
rect 42698 707377 42704 707429
rect 42448 706711 42454 706763
rect 42506 706751 42512 706763
rect 43024 706751 43030 706763
rect 42506 706723 43030 706751
rect 42506 706711 42512 706723
rect 43024 706711 43030 706723
rect 43082 706711 43088 706763
rect 42160 704269 42166 704321
rect 42218 704309 42224 704321
rect 43120 704309 43126 704321
rect 42218 704281 43126 704309
rect 42218 704269 42224 704281
rect 43120 704269 43126 704281
rect 43178 704269 43184 704321
rect 42064 703677 42070 703729
rect 42122 703717 42128 703729
rect 42928 703717 42934 703729
rect 42122 703689 42934 703717
rect 42122 703677 42128 703689
rect 42928 703677 42934 703689
rect 42986 703677 42992 703729
rect 42256 702937 42262 702989
rect 42314 702977 42320 702989
rect 42640 702977 42646 702989
rect 42314 702949 42646 702977
rect 42314 702937 42320 702949
rect 42640 702937 42646 702949
rect 42698 702937 42704 702989
rect 42064 702863 42070 702915
rect 42122 702903 42128 702915
rect 42736 702903 42742 702915
rect 42122 702875 42742 702903
rect 42122 702863 42128 702875
rect 42736 702863 42742 702875
rect 42794 702863 42800 702915
rect 654736 702789 654742 702841
rect 654794 702829 654800 702841
rect 675376 702829 675382 702841
rect 654794 702801 675382 702829
rect 654794 702789 654800 702801
rect 675376 702789 675382 702801
rect 675434 702789 675440 702841
rect 42448 702715 42454 702767
rect 42506 702755 42512 702767
rect 58864 702755 58870 702767
rect 42506 702727 58870 702755
rect 42506 702715 42512 702727
rect 58864 702715 58870 702727
rect 58922 702715 58928 702767
rect 649456 702715 649462 702767
rect 649514 702755 649520 702767
rect 679984 702755 679990 702767
rect 649514 702727 679990 702755
rect 649514 702715 649520 702727
rect 679984 702715 679990 702727
rect 680042 702715 680048 702767
rect 43504 702641 43510 702693
rect 43562 702681 43568 702693
rect 58768 702681 58774 702693
rect 43562 702653 58774 702681
rect 43562 702641 43568 702653
rect 58768 702641 58774 702653
rect 58826 702641 58832 702693
rect 45040 702567 45046 702619
rect 45098 702607 45104 702619
rect 58672 702607 58678 702619
rect 45098 702579 58678 702607
rect 45098 702567 45104 702579
rect 58672 702567 58678 702579
rect 58730 702567 58736 702619
rect 42064 700569 42070 700621
rect 42122 700609 42128 700621
rect 42832 700609 42838 700621
rect 42122 700581 42838 700609
rect 42122 700569 42128 700581
rect 42832 700569 42838 700581
rect 42890 700569 42896 700621
rect 42160 699903 42166 699955
rect 42218 699943 42224 699955
rect 42544 699943 42550 699955
rect 42218 699915 42550 699943
rect 42218 699903 42224 699915
rect 42544 699903 42550 699915
rect 42602 699903 42608 699955
rect 670768 699829 670774 699881
rect 670826 699869 670832 699881
rect 679696 699869 679702 699881
rect 670826 699841 679702 699869
rect 670826 699829 670832 699841
rect 679696 699829 679702 699841
rect 679754 699829 679760 699881
rect 47536 699755 47542 699807
rect 47594 699795 47600 699807
rect 59248 699795 59254 699807
rect 47594 699767 59254 699795
rect 47594 699755 47600 699767
rect 59248 699755 59254 699767
rect 59306 699755 59312 699807
rect 44944 699681 44950 699733
rect 45002 699721 45008 699733
rect 58864 699721 58870 699733
rect 45002 699693 58870 699721
rect 45002 699681 45008 699693
rect 58864 699681 58870 699693
rect 58922 699681 58928 699733
rect 654160 694131 654166 694183
rect 654218 694171 654224 694183
rect 675280 694171 675286 694183
rect 654218 694143 675286 694171
rect 654218 694131 654224 694143
rect 675280 694131 675286 694143
rect 675338 694131 675344 694183
rect 673744 692873 673750 692925
rect 673802 692913 673808 692925
rect 675376 692913 675382 692925
rect 673802 692885 675382 692913
rect 673802 692873 673808 692885
rect 675376 692873 675382 692885
rect 675434 692873 675440 692925
rect 654064 691245 654070 691297
rect 654122 691285 654128 691297
rect 675088 691285 675094 691297
rect 654122 691257 675094 691285
rect 654122 691245 654128 691257
rect 675088 691245 675094 691257
rect 675146 691245 675152 691297
rect 674896 690431 674902 690483
rect 674954 690471 674960 690483
rect 675472 690471 675478 690483
rect 674954 690443 675478 690471
rect 674954 690431 674960 690443
rect 675472 690431 675478 690443
rect 675530 690431 675536 690483
rect 675184 689765 675190 689817
rect 675242 689805 675248 689817
rect 675376 689805 675382 689817
rect 675242 689777 675382 689805
rect 675242 689765 675248 689777
rect 675376 689765 675382 689777
rect 675434 689765 675440 689817
rect 674800 689099 674806 689151
rect 674858 689139 674864 689151
rect 675376 689139 675382 689151
rect 674858 689111 675382 689139
rect 674858 689099 674864 689111
rect 675376 689099 675382 689111
rect 675434 689099 675440 689151
rect 673552 688729 673558 688781
rect 673610 688769 673616 688781
rect 675472 688769 675478 688781
rect 673610 688741 675478 688769
rect 673610 688729 673616 688741
rect 675472 688729 675478 688741
rect 675530 688729 675536 688781
rect 41776 688211 41782 688263
rect 41834 688251 41840 688263
rect 50320 688251 50326 688263
rect 41834 688223 50326 688251
rect 41834 688211 41840 688223
rect 50320 688211 50326 688223
rect 50378 688211 50384 688263
rect 41584 687471 41590 687523
rect 41642 687511 41648 687523
rect 47632 687511 47638 687523
rect 41642 687483 47638 687511
rect 41642 687471 41648 687483
rect 47632 687471 47638 687483
rect 47690 687471 47696 687523
rect 41776 687175 41782 687227
rect 41834 687215 41840 687227
rect 47728 687215 47734 687227
rect 41834 687187 47734 687215
rect 41834 687175 41840 687187
rect 47728 687175 47734 687187
rect 47786 687175 47792 687227
rect 41584 686953 41590 687005
rect 41642 686993 41648 687005
rect 43312 686993 43318 687005
rect 41642 686965 43318 686993
rect 41642 686953 41648 686965
rect 43312 686953 43318 686965
rect 43370 686953 43376 687005
rect 674320 686731 674326 686783
rect 674378 686771 674384 686783
rect 675280 686771 675286 686783
rect 674378 686743 675286 686771
rect 674378 686731 674384 686743
rect 675280 686731 675286 686743
rect 675338 686731 675344 686783
rect 41584 685991 41590 686043
rect 41642 686031 41648 686043
rect 43504 686031 43510 686043
rect 41642 686003 43510 686031
rect 41642 685991 41648 686003
rect 43504 685991 43510 686003
rect 43562 685991 43568 686043
rect 41776 685325 41782 685377
rect 41834 685365 41840 685377
rect 43216 685365 43222 685377
rect 41834 685337 43222 685365
rect 41834 685325 41840 685337
rect 43216 685325 43222 685337
rect 43274 685365 43280 685377
rect 45040 685365 45046 685377
rect 43274 685337 45046 685365
rect 43274 685325 43280 685337
rect 45040 685325 45046 685337
rect 45098 685325 45104 685377
rect 41776 684141 41782 684193
rect 41834 684181 41840 684193
rect 43408 684181 43414 684193
rect 41834 684153 43414 684181
rect 41834 684141 41840 684153
rect 43408 684141 43414 684153
rect 43466 684181 43472 684193
rect 44944 684181 44950 684193
rect 43466 684153 44950 684181
rect 43466 684141 43472 684153
rect 44944 684141 44950 684153
rect 45002 684141 45008 684193
rect 674416 683623 674422 683675
rect 674474 683663 674480 683675
rect 675472 683663 675478 683675
rect 674474 683635 675478 683663
rect 674474 683623 674480 683635
rect 675472 683623 675478 683635
rect 675530 683623 675536 683675
rect 674512 682809 674518 682861
rect 674570 682849 674576 682861
rect 675184 682849 675190 682861
rect 674570 682821 675190 682849
rect 674570 682809 674576 682821
rect 675184 682809 675190 682821
rect 675242 682809 675248 682861
rect 41776 681625 41782 681677
rect 41834 681665 41840 681677
rect 42640 681665 42646 681677
rect 41834 681637 42646 681665
rect 41834 681625 41840 681637
rect 42640 681625 42646 681637
rect 42698 681625 42704 681677
rect 41776 679923 41782 679975
rect 41834 679963 41840 679975
rect 42736 679963 42742 679975
rect 41834 679935 42742 679963
rect 41834 679923 41840 679935
rect 42736 679923 42742 679935
rect 42794 679923 42800 679975
rect 41776 679701 41782 679753
rect 41834 679741 41840 679753
rect 42832 679741 42838 679753
rect 41834 679713 42838 679741
rect 41834 679701 41840 679713
rect 42832 679701 42838 679713
rect 42890 679701 42896 679753
rect 41776 677851 41782 677903
rect 41834 677891 41840 677903
rect 43120 677891 43126 677903
rect 41834 677863 43126 677891
rect 41834 677851 41840 677863
rect 43120 677851 43126 677863
rect 43178 677851 43184 677903
rect 42448 677555 42454 677607
rect 42506 677595 42512 677607
rect 42832 677595 42838 677607
rect 42506 677567 42838 677595
rect 42506 677555 42512 677567
rect 42832 677555 42838 677567
rect 42890 677555 42896 677607
rect 41776 677407 41782 677459
rect 41834 677447 41840 677459
rect 43024 677447 43030 677459
rect 41834 677419 43030 677447
rect 41834 677407 41840 677419
rect 43024 677407 43030 677419
rect 43082 677407 43088 677459
rect 41584 677259 41590 677311
rect 41642 677299 41648 677311
rect 42832 677299 42838 677311
rect 41642 677271 42838 677299
rect 41642 677259 41648 677271
rect 42832 677259 42838 677271
rect 42890 677259 42896 677311
rect 41776 677037 41782 677089
rect 41834 677077 41840 677089
rect 42640 677077 42646 677089
rect 41834 677049 42646 677077
rect 41834 677037 41840 677049
rect 42640 677037 42646 677049
rect 42698 677037 42704 677089
rect 41776 675705 41782 675757
rect 41834 675745 41840 675757
rect 47536 675745 47542 675757
rect 41834 675717 47542 675745
rect 41834 675705 41840 675717
rect 47536 675705 47542 675717
rect 47594 675705 47600 675757
rect 42448 671043 42454 671095
rect 42506 671083 42512 671095
rect 59632 671083 59638 671095
rect 42506 671055 59638 671083
rect 42506 671043 42512 671055
rect 59632 671043 59638 671055
rect 59690 671043 59696 671095
rect 42736 670895 42742 670947
rect 42794 670935 42800 670947
rect 42794 670907 42878 670935
rect 42794 670895 42800 670907
rect 42160 670747 42166 670799
rect 42218 670787 42224 670799
rect 42736 670787 42742 670799
rect 42218 670759 42742 670787
rect 42218 670747 42224 670759
rect 42736 670747 42742 670759
rect 42794 670747 42800 670799
rect 42256 670451 42262 670503
rect 42314 670451 42320 670503
rect 42274 670281 42302 670451
rect 42256 670229 42262 670281
rect 42314 670229 42320 670281
rect 42352 670229 42358 670281
rect 42410 670269 42416 670281
rect 42850 670269 42878 670907
rect 42410 670241 42878 670269
rect 42410 670229 42416 670241
rect 670768 669193 670774 669245
rect 670826 669233 670832 669245
rect 676048 669233 676054 669245
rect 670826 669205 676054 669233
rect 670826 669193 670832 669205
rect 676048 669193 676054 669205
rect 676106 669193 676112 669245
rect 42160 668527 42166 668579
rect 42218 668567 42224 668579
rect 42544 668567 42550 668579
rect 42218 668539 42550 668567
rect 42218 668527 42224 668539
rect 42544 668527 42550 668539
rect 42602 668527 42608 668579
rect 655504 668527 655510 668579
rect 655562 668567 655568 668579
rect 676144 668567 676150 668579
rect 655562 668539 676150 668567
rect 655562 668527 655568 668539
rect 676144 668527 676150 668539
rect 676202 668527 676208 668579
rect 655312 668379 655318 668431
rect 655370 668419 655376 668431
rect 676240 668419 676246 668431
rect 655370 668391 676246 668419
rect 655370 668379 655376 668391
rect 676240 668379 676246 668391
rect 676298 668379 676304 668431
rect 675088 668231 675094 668283
rect 675146 668271 675152 668283
rect 676048 668271 676054 668283
rect 675146 668243 676054 668271
rect 675146 668231 675152 668243
rect 676048 668231 676054 668243
rect 676106 668231 676112 668283
rect 655120 668157 655126 668209
rect 655178 668197 655184 668209
rect 676336 668197 676342 668209
rect 655178 668169 676342 668197
rect 655178 668157 655184 668169
rect 676336 668157 676342 668169
rect 676394 668157 676400 668209
rect 674704 668083 674710 668135
rect 674762 668123 674768 668135
rect 676048 668123 676054 668135
rect 674762 668095 676054 668123
rect 674762 668083 674768 668095
rect 676048 668083 676054 668095
rect 676106 668083 676112 668135
rect 670672 668009 670678 668061
rect 670730 668049 670736 668061
rect 675952 668049 675958 668061
rect 670730 668021 675958 668049
rect 670730 668009 670736 668021
rect 675952 668009 675958 668021
rect 676010 668009 676016 668061
rect 42160 667861 42166 667913
rect 42218 667901 42224 667913
rect 42448 667901 42454 667913
rect 42218 667873 42454 667901
rect 42218 667861 42224 667873
rect 42448 667861 42454 667873
rect 42506 667861 42512 667913
rect 670864 667639 670870 667691
rect 670922 667679 670928 667691
rect 675952 667679 675958 667691
rect 670922 667651 675958 667679
rect 670922 667639 670928 667651
rect 675952 667639 675958 667651
rect 676010 667639 676016 667691
rect 652240 666751 652246 666803
rect 652298 666791 652304 666803
rect 670576 666791 670582 666803
rect 652298 666763 670582 666791
rect 652298 666751 652304 666763
rect 670576 666751 670582 666763
rect 670634 666791 670640 666803
rect 676240 666791 676246 666803
rect 670634 666763 676246 666791
rect 670634 666751 670640 666763
rect 676240 666751 676246 666763
rect 676298 666751 676304 666803
rect 42160 666677 42166 666729
rect 42218 666717 42224 666729
rect 42832 666717 42838 666729
rect 42218 666689 42838 666717
rect 42218 666677 42224 666689
rect 42832 666677 42838 666689
rect 42890 666677 42896 666729
rect 649744 666677 649750 666729
rect 649802 666717 649808 666729
rect 670672 666717 670678 666729
rect 649802 666689 670678 666717
rect 649802 666677 649808 666689
rect 670672 666677 670678 666689
rect 670730 666677 670736 666729
rect 670960 666307 670966 666359
rect 671018 666347 671024 666359
rect 676240 666347 676246 666359
rect 671018 666319 676246 666347
rect 671018 666307 671024 666319
rect 676240 666307 676246 666319
rect 676298 666307 676304 666359
rect 42160 665271 42166 665323
rect 42218 665311 42224 665323
rect 45136 665311 45142 665323
rect 42218 665283 45142 665311
rect 42218 665271 42224 665283
rect 45136 665271 45142 665283
rect 45194 665271 45200 665323
rect 674992 665197 674998 665249
rect 675050 665237 675056 665249
rect 676240 665237 676246 665249
rect 675050 665209 676246 665237
rect 675050 665197 675056 665209
rect 676240 665197 676246 665209
rect 676298 665197 676304 665249
rect 42160 665123 42166 665175
rect 42218 665163 42224 665175
rect 42640 665163 42646 665175
rect 42218 665135 42646 665163
rect 42218 665123 42224 665135
rect 42640 665123 42646 665135
rect 42698 665123 42704 665175
rect 674608 665123 674614 665175
rect 674666 665163 674672 665175
rect 676048 665163 676054 665175
rect 674666 665135 676054 665163
rect 674666 665123 674672 665135
rect 676048 665123 676054 665135
rect 676106 665123 676112 665175
rect 42160 664827 42166 664879
rect 42218 664867 42224 664879
rect 43120 664867 43126 664879
rect 42218 664839 43126 664867
rect 42218 664827 42224 664839
rect 43120 664827 43126 664839
rect 43178 664827 43184 664879
rect 42064 664161 42070 664213
rect 42122 664201 42128 664213
rect 43024 664201 43030 664213
rect 42122 664173 43030 664201
rect 42122 664161 42128 664173
rect 43024 664161 43030 664173
rect 43082 664161 43088 664213
rect 42160 663347 42166 663399
rect 42218 663387 42224 663399
rect 42352 663387 42358 663399
rect 42218 663359 42358 663387
rect 42218 663347 42224 663359
rect 42352 663347 42358 663359
rect 42410 663347 42416 663399
rect 674224 662311 674230 662363
rect 674282 662351 674288 662363
rect 676048 662351 676054 662363
rect 674282 662323 676054 662351
rect 674282 662311 674288 662323
rect 676048 662311 676054 662323
rect 676106 662311 676112 662363
rect 42064 661053 42070 661105
rect 42122 661093 42128 661105
rect 42544 661093 42550 661105
rect 42122 661065 42550 661093
rect 42122 661053 42128 661065
rect 42544 661053 42550 661065
rect 42602 661053 42608 661105
rect 673648 660609 673654 660661
rect 673706 660649 673712 660661
rect 676048 660649 676054 660661
rect 673706 660621 676054 660649
rect 673706 660609 673712 660621
rect 676048 660609 676054 660621
rect 676106 660609 676112 660661
rect 42064 660387 42070 660439
rect 42122 660427 42128 660439
rect 42448 660427 42454 660439
rect 42122 660399 42454 660427
rect 42122 660387 42128 660399
rect 42448 660387 42454 660399
rect 42506 660387 42512 660439
rect 42160 659869 42166 659921
rect 42218 659909 42224 659921
rect 42928 659909 42934 659921
rect 42218 659881 42934 659909
rect 42218 659869 42224 659881
rect 42928 659869 42934 659881
rect 42986 659869 42992 659921
rect 673456 659869 673462 659921
rect 673514 659909 673520 659921
rect 676240 659909 676246 659921
rect 673514 659881 676246 659909
rect 673514 659869 673520 659881
rect 676240 659869 676246 659881
rect 676298 659869 676304 659921
rect 42448 659499 42454 659551
rect 42506 659539 42512 659551
rect 57712 659539 57718 659551
rect 42506 659511 57718 659539
rect 42506 659499 42512 659511
rect 57712 659499 57718 659511
rect 57770 659499 57776 659551
rect 47728 659425 47734 659477
rect 47786 659465 47792 659477
rect 59152 659465 59158 659477
rect 47786 659437 59158 659465
rect 47786 659425 47792 659437
rect 59152 659425 59158 659437
rect 59210 659425 59216 659477
rect 45136 659351 45142 659403
rect 45194 659391 45200 659403
rect 58768 659391 58774 659403
rect 45194 659363 58774 659391
rect 45194 659351 45200 659363
rect 58768 659351 58774 659363
rect 58826 659351 58832 659403
rect 42064 659055 42070 659107
rect 42122 659095 42128 659107
rect 42640 659095 42646 659107
rect 42122 659067 42646 659095
rect 42122 659055 42128 659067
rect 42640 659055 42646 659067
rect 42698 659055 42704 659107
rect 654160 656761 654166 656813
rect 654218 656801 654224 656813
rect 675376 656801 675382 656813
rect 654218 656773 675382 656801
rect 654218 656761 654224 656773
rect 675376 656761 675382 656773
rect 675434 656761 675440 656813
rect 42160 656687 42166 656739
rect 42218 656727 42224 656739
rect 42544 656727 42550 656739
rect 42218 656699 42550 656727
rect 42218 656687 42224 656699
rect 42544 656687 42550 656699
rect 42602 656687 42608 656739
rect 649552 656687 649558 656739
rect 649610 656727 649616 656739
rect 679792 656727 679798 656739
rect 649610 656699 679798 656727
rect 649610 656687 649616 656699
rect 679792 656687 679798 656699
rect 679850 656687 679856 656739
rect 50320 656613 50326 656665
rect 50378 656653 50384 656665
rect 58192 656653 58198 656665
rect 50378 656625 58198 656653
rect 50378 656613 50384 656625
rect 58192 656613 58198 656625
rect 58250 656613 58256 656665
rect 47632 656539 47638 656591
rect 47690 656579 47696 656591
rect 58384 656579 58390 656591
rect 47690 656551 58390 656579
rect 47690 656539 47696 656551
rect 58384 656539 58390 656551
rect 58442 656539 58448 656591
rect 655792 648177 655798 648229
rect 655850 648217 655856 648229
rect 675184 648217 675190 648229
rect 655850 648189 675190 648217
rect 655850 648177 655856 648189
rect 675184 648177 675190 648189
rect 675242 648177 675248 648229
rect 673840 648029 673846 648081
rect 673898 648069 673904 648081
rect 675280 648069 675286 648081
rect 673898 648041 675286 648069
rect 673898 648029 673904 648041
rect 675280 648029 675286 648041
rect 675338 648029 675344 648081
rect 655984 645143 655990 645195
rect 656042 645183 656048 645195
rect 675088 645183 675094 645195
rect 656042 645155 675094 645183
rect 656042 645143 656048 645155
rect 675088 645143 675094 645155
rect 675146 645143 675152 645195
rect 41584 644847 41590 644899
rect 41642 644887 41648 644899
rect 50320 644887 50326 644899
rect 41642 644859 50326 644887
rect 41642 644847 41648 644859
rect 50320 644847 50326 644859
rect 50378 644847 50384 644899
rect 673072 644551 673078 644603
rect 673130 644591 673136 644603
rect 675280 644591 675286 644603
rect 673130 644563 675286 644591
rect 673130 644551 673136 644563
rect 675280 644551 675286 644563
rect 675338 644551 675344 644603
rect 41584 644255 41590 644307
rect 41642 644295 41648 644307
rect 47728 644295 47734 644307
rect 41642 644267 47734 644295
rect 41642 644255 41648 644267
rect 47728 644255 47734 644267
rect 47786 644255 47792 644307
rect 41776 643959 41782 644011
rect 41834 643999 41840 644011
rect 47824 643999 47830 644011
rect 41834 643971 47830 643999
rect 41834 643959 41840 643971
rect 47824 643959 47830 643971
rect 47882 643959 47888 644011
rect 673264 643885 673270 643937
rect 673322 643925 673328 643937
rect 675280 643925 675286 643937
rect 673322 643897 675286 643925
rect 673322 643885 673328 643897
rect 675280 643885 675286 643897
rect 675338 643885 675344 643937
rect 41584 643737 41590 643789
rect 41642 643777 41648 643789
rect 43504 643777 43510 643789
rect 41642 643749 43510 643777
rect 41642 643737 41648 643749
rect 43504 643737 43510 643749
rect 43562 643737 43568 643789
rect 673168 643367 673174 643419
rect 673226 643407 673232 643419
rect 675280 643407 675286 643419
rect 673226 643379 675286 643407
rect 673226 643367 673232 643379
rect 675280 643367 675286 643379
rect 675338 643367 675344 643419
rect 41584 642775 41590 642827
rect 41642 642815 41648 642827
rect 43408 642815 43414 642827
rect 41642 642787 43414 642815
rect 41642 642775 41648 642787
rect 43408 642775 43414 642787
rect 43466 642775 43472 642827
rect 41488 642479 41494 642531
rect 41546 642519 41552 642531
rect 61936 642519 61942 642531
rect 41546 642491 61942 642519
rect 41546 642479 41552 642491
rect 61936 642479 61942 642491
rect 61994 642479 62000 642531
rect 673360 642257 673366 642309
rect 673418 642297 673424 642309
rect 675184 642297 675190 642309
rect 673418 642269 675190 642297
rect 673418 642257 673424 642269
rect 675184 642257 675190 642269
rect 675242 642257 675248 642309
rect 41584 641295 41590 641347
rect 41642 641335 41648 641347
rect 43312 641335 43318 641347
rect 41642 641307 43318 641335
rect 41642 641295 41648 641307
rect 43312 641295 43318 641307
rect 43370 641295 43376 641347
rect 41776 640555 41782 640607
rect 41834 640595 41840 640607
rect 42832 640595 42838 640607
rect 41834 640567 42838 640595
rect 41834 640555 41840 640567
rect 42832 640555 42838 640567
rect 42890 640555 42896 640607
rect 674224 639075 674230 639127
rect 674282 639115 674288 639127
rect 675088 639115 675094 639127
rect 674282 639087 675094 639115
rect 674282 639075 674288 639087
rect 675088 639075 675094 639087
rect 675146 639075 675152 639127
rect 41776 636707 41782 636759
rect 41834 636747 41840 636759
rect 43024 636747 43030 636759
rect 41834 636719 43030 636747
rect 41834 636707 41840 636719
rect 43024 636707 43030 636719
rect 43082 636707 43088 636759
rect 41776 636041 41782 636093
rect 41834 636081 41840 636093
rect 42544 636081 42550 636093
rect 41834 636053 42550 636081
rect 41834 636041 41840 636053
rect 42544 636041 42550 636053
rect 42602 636041 42608 636093
rect 41584 635375 41590 635427
rect 41642 635415 41648 635427
rect 43120 635415 43126 635427
rect 41642 635387 43126 635415
rect 41642 635375 41648 635387
rect 43120 635375 43126 635387
rect 43178 635375 43184 635427
rect 674992 635005 674998 635057
rect 675050 635045 675056 635057
rect 679696 635045 679702 635057
rect 675050 635017 679702 635045
rect 675050 635005 675056 635017
rect 679696 635005 679702 635017
rect 679754 635005 679760 635057
rect 41584 634487 41590 634539
rect 41642 634527 41648 634539
rect 42832 634527 42838 634539
rect 41642 634499 42838 634527
rect 41642 634487 41648 634499
rect 42832 634487 42838 634499
rect 42890 634487 42896 634539
rect 41584 634191 41590 634243
rect 41642 634231 41648 634243
rect 42736 634231 42742 634243
rect 41642 634203 42742 634231
rect 41642 634191 41648 634203
rect 42736 634191 42742 634203
rect 42794 634191 42800 634243
rect 41680 633895 41686 633947
rect 41738 633935 41744 633947
rect 42928 633935 42934 633947
rect 41738 633907 42934 633935
rect 41738 633895 41744 633907
rect 42928 633895 42934 633907
rect 42986 633895 42992 633947
rect 41776 632489 41782 632541
rect 41834 632529 41840 632541
rect 47632 632529 47638 632541
rect 41834 632501 47638 632529
rect 41834 632489 41840 632501
rect 47632 632489 47638 632501
rect 47690 632489 47696 632541
rect 43120 629307 43126 629359
rect 43178 629347 43184 629359
rect 43504 629347 43510 629359
rect 43178 629319 43510 629347
rect 43178 629307 43184 629319
rect 43504 629307 43510 629319
rect 43562 629307 43568 629359
rect 42928 629159 42934 629211
rect 42986 629199 42992 629211
rect 43312 629199 43318 629211
rect 42986 629171 43318 629199
rect 42986 629159 42992 629171
rect 43312 629159 43318 629171
rect 43370 629159 43376 629211
rect 674128 629085 674134 629137
rect 674186 629125 674192 629137
rect 675088 629125 675094 629137
rect 674186 629097 675094 629125
rect 674186 629085 674192 629097
rect 675088 629085 675094 629097
rect 675146 629085 675152 629137
rect 42160 628789 42166 628841
rect 42218 628829 42224 628841
rect 42832 628829 42838 628841
rect 42218 628801 42838 628829
rect 42218 628789 42224 628801
rect 42832 628789 42838 628801
rect 42890 628789 42896 628841
rect 42064 628715 42070 628767
rect 42122 628755 42128 628767
rect 42736 628755 42742 628767
rect 42122 628727 42742 628755
rect 42122 628715 42128 628727
rect 42736 628715 42742 628727
rect 42794 628715 42800 628767
rect 42160 628123 42166 628175
rect 42218 628163 42224 628175
rect 42640 628163 42646 628175
rect 42218 628135 42646 628163
rect 42218 628123 42224 628135
rect 42640 628123 42646 628135
rect 42698 628123 42704 628175
rect 42448 627975 42454 628027
rect 42506 628015 42512 628027
rect 42640 628015 42646 628027
rect 42506 627987 42646 628015
rect 42506 627975 42512 627987
rect 42640 627975 42646 627987
rect 42698 627975 42704 628027
rect 42448 627827 42454 627879
rect 42506 627867 42512 627879
rect 54640 627867 54646 627879
rect 42506 627839 54646 627867
rect 42506 627827 42512 627839
rect 54640 627827 54646 627839
rect 54698 627827 54704 627879
rect 42160 627383 42166 627435
rect 42218 627383 42224 627435
rect 42178 626535 42206 627383
rect 42256 626535 42262 626547
rect 42178 626507 42262 626535
rect 42256 626495 42262 626507
rect 42314 626495 42320 626547
rect 42352 625425 42358 625437
rect 42178 625397 42358 625425
rect 42178 625363 42206 625397
rect 42352 625385 42358 625397
rect 42410 625385 42416 625437
rect 42160 625311 42166 625363
rect 42218 625311 42224 625363
rect 42352 625237 42358 625289
rect 42410 625277 42416 625289
rect 43312 625277 43318 625289
rect 42410 625249 43318 625277
rect 42410 625237 42416 625249
rect 43312 625237 43318 625249
rect 43370 625237 43376 625289
rect 655600 624941 655606 624993
rect 655658 624981 655664 624993
rect 676240 624981 676246 624993
rect 655658 624953 676246 624981
rect 655658 624941 655664 624953
rect 676240 624941 676246 624953
rect 676298 624941 676304 624993
rect 54640 624793 54646 624845
rect 54698 624833 54704 624845
rect 58960 624833 58966 624845
rect 54698 624805 58966 624833
rect 54698 624793 54704 624805
rect 58960 624793 58966 624805
rect 59018 624793 59024 624845
rect 42160 624645 42166 624697
rect 42218 624685 42224 624697
rect 42448 624685 42454 624697
rect 42218 624657 42454 624685
rect 42218 624645 42224 624657
rect 42448 624645 42454 624657
rect 42506 624645 42512 624697
rect 42160 623461 42166 623513
rect 42218 623501 42224 623513
rect 42544 623501 42550 623513
rect 42218 623473 42550 623501
rect 42218 623461 42224 623473
rect 42544 623461 42550 623473
rect 42602 623461 42608 623513
rect 672784 623387 672790 623439
rect 672842 623427 672848 623439
rect 676048 623427 676054 623439
rect 672842 623399 676054 623427
rect 672842 623387 672848 623399
rect 676048 623387 676054 623399
rect 676106 623387 676112 623439
rect 669616 623091 669622 623143
rect 669674 623131 669680 623143
rect 670864 623131 670870 623143
rect 669674 623103 670870 623131
rect 669674 623091 669680 623103
rect 670864 623091 670870 623103
rect 670922 623131 670928 623143
rect 676048 623131 676054 623143
rect 670922 623103 676054 623131
rect 670922 623091 670928 623103
rect 676048 623091 676054 623103
rect 676106 623091 676112 623143
rect 655408 622499 655414 622551
rect 655466 622539 655472 622551
rect 676240 622539 676246 622551
rect 655466 622511 676246 622539
rect 655466 622499 655472 622511
rect 676240 622499 676246 622511
rect 676298 622499 676304 622551
rect 670768 622425 670774 622477
rect 670826 622465 670832 622477
rect 676048 622465 676054 622477
rect 670826 622437 676054 622465
rect 670826 622425 670832 622437
rect 676048 622425 676054 622437
rect 676106 622425 676112 622477
rect 655216 622351 655222 622403
rect 655274 622391 655280 622403
rect 676144 622391 676150 622403
rect 655274 622363 676150 622391
rect 655274 622351 655280 622363
rect 676144 622351 676150 622363
rect 676202 622351 676208 622403
rect 42160 622055 42166 622107
rect 42218 622095 42224 622107
rect 47920 622095 47926 622107
rect 42218 622067 47926 622095
rect 42218 622055 42224 622067
rect 47920 622055 47926 622067
rect 47978 622055 47984 622107
rect 42064 621981 42070 622033
rect 42122 622021 42128 622033
rect 42640 622021 42646 622033
rect 42122 621993 42646 622021
rect 42122 621981 42128 621993
rect 42640 621981 42646 621993
rect 42698 621981 42704 622033
rect 674512 621981 674518 622033
rect 674570 622021 674576 622033
rect 676240 622021 676246 622033
rect 674570 621993 676246 622021
rect 674570 621981 674576 621993
rect 676240 621981 676246 621993
rect 676298 621981 676304 622033
rect 670960 621907 670966 621959
rect 671018 621947 671024 621959
rect 676048 621947 676054 621959
rect 671018 621919 676054 621947
rect 671018 621907 671024 621919
rect 676048 621907 676054 621919
rect 676106 621907 676112 621959
rect 42256 621833 42262 621885
rect 42314 621873 42320 621885
rect 42640 621873 42646 621885
rect 42314 621845 42646 621873
rect 42314 621833 42320 621845
rect 42640 621833 42646 621845
rect 42698 621833 42704 621885
rect 42448 621611 42454 621663
rect 42506 621651 42512 621663
rect 42928 621651 42934 621663
rect 42506 621623 42934 621651
rect 42506 621611 42512 621623
rect 42928 621611 42934 621623
rect 42986 621611 42992 621663
rect 42352 621537 42358 621589
rect 42410 621577 42416 621589
rect 43024 621577 43030 621589
rect 42410 621549 43030 621577
rect 42410 621537 42416 621549
rect 43024 621537 43030 621549
rect 43082 621537 43088 621589
rect 42928 621463 42934 621515
rect 42986 621503 42992 621515
rect 43504 621503 43510 621515
rect 42986 621475 43510 621503
rect 42986 621463 42992 621475
rect 43504 621463 43510 621475
rect 43562 621463 43568 621515
rect 670864 621315 670870 621367
rect 670922 621355 670928 621367
rect 676048 621355 676054 621367
rect 670922 621327 676054 621355
rect 670922 621315 670928 621327
rect 676048 621315 676054 621327
rect 676106 621315 676112 621367
rect 42448 620353 42454 620405
rect 42506 620393 42512 620405
rect 43120 620393 43126 620405
rect 42506 620365 43126 620393
rect 42506 620353 42512 620365
rect 43120 620353 43126 620365
rect 43178 620353 43184 620405
rect 669808 619983 669814 620035
rect 669866 620023 669872 620035
rect 670960 620023 670966 620035
rect 669866 619995 670966 620023
rect 669866 619983 669872 619995
rect 670960 619983 670966 619995
rect 671018 619983 671024 620035
rect 674896 619021 674902 619073
rect 674954 619061 674960 619073
rect 676048 619061 676054 619073
rect 674954 619033 676054 619061
rect 674954 619021 674960 619033
rect 676048 619021 676054 619033
rect 676106 619021 676112 619073
rect 674416 618799 674422 618851
rect 674474 618839 674480 618851
rect 676240 618839 676246 618851
rect 674474 618811 676246 618839
rect 674474 618799 674480 618811
rect 676240 618799 676246 618811
rect 676298 618799 676304 618851
rect 674320 618577 674326 618629
rect 674378 618617 674384 618629
rect 676048 618617 676054 618629
rect 674378 618589 676054 618617
rect 674378 618577 674384 618589
rect 676048 618577 676054 618589
rect 676106 618577 676112 618629
rect 42256 617319 42262 617371
rect 42314 617359 42320 617371
rect 42928 617359 42934 617371
rect 42314 617331 42934 617359
rect 42314 617319 42320 617331
rect 42928 617319 42934 617331
rect 42986 617319 42992 617371
rect 42160 616653 42166 616705
rect 42218 616693 42224 616705
rect 42832 616693 42838 616705
rect 42218 616665 42838 616693
rect 42218 616653 42224 616665
rect 42832 616653 42838 616665
rect 42890 616653 42896 616705
rect 42256 616579 42262 616631
rect 42314 616619 42320 616631
rect 42736 616619 42742 616631
rect 42314 616591 42742 616619
rect 42314 616579 42320 616591
rect 42736 616579 42742 616591
rect 42794 616579 42800 616631
rect 42928 616357 42934 616409
rect 42986 616397 42992 616409
rect 58192 616397 58198 616409
rect 42986 616369 58198 616397
rect 42986 616357 42992 616369
rect 58192 616357 58198 616369
rect 58250 616357 58256 616409
rect 47824 616283 47830 616335
rect 47882 616323 47888 616335
rect 58960 616323 58966 616335
rect 47882 616295 58966 616323
rect 47882 616283 47888 616295
rect 58960 616283 58966 616295
rect 59018 616283 59024 616335
rect 674800 616283 674806 616335
rect 674858 616323 674864 616335
rect 676048 616323 676054 616335
rect 674858 616295 676054 616323
rect 674858 616283 674864 616295
rect 676048 616283 676054 616295
rect 676106 616283 676112 616335
rect 47920 616209 47926 616261
rect 47978 616249 47984 616261
rect 59632 616249 59638 616261
rect 47978 616221 59638 616249
rect 47978 616209 47984 616221
rect 59632 616209 59638 616221
rect 59690 616209 59696 616261
rect 673744 615617 673750 615669
rect 673802 615657 673808 615669
rect 676240 615657 676246 615669
rect 673802 615629 676246 615657
rect 673802 615617 673808 615629
rect 676240 615617 676246 615629
rect 676298 615617 676304 615669
rect 673552 614433 673558 614485
rect 673610 614473 673616 614485
rect 676048 614473 676054 614485
rect 673610 614445 676054 614473
rect 673610 614433 673616 614445
rect 676048 614433 676054 614445
rect 676106 614433 676112 614485
rect 655792 613471 655798 613523
rect 655850 613511 655856 613523
rect 675376 613511 675382 613523
rect 655850 613483 675382 613511
rect 655850 613471 655856 613483
rect 675376 613471 675382 613483
rect 675434 613471 675440 613523
rect 50320 613397 50326 613449
rect 50378 613437 50384 613449
rect 59632 613437 59638 613449
rect 50378 613409 59638 613437
rect 50378 613397 50384 613409
rect 59632 613397 59638 613409
rect 59690 613397 59696 613449
rect 47728 613323 47734 613375
rect 47786 613363 47792 613375
rect 59536 613363 59542 613375
rect 47786 613335 59542 613363
rect 47786 613323 47792 613335
rect 59536 613323 59542 613335
rect 59594 613323 59600 613375
rect 42064 612805 42070 612857
rect 42122 612845 42128 612857
rect 42832 612845 42838 612857
rect 42122 612817 42838 612845
rect 42122 612805 42128 612817
rect 42832 612805 42838 612817
rect 42890 612805 42896 612857
rect 649648 610585 649654 610637
rect 649706 610625 649712 610637
rect 679984 610625 679990 610637
rect 649706 610597 679990 610625
rect 649706 610585 649712 610597
rect 679984 610585 679990 610597
rect 680042 610585 680048 610637
rect 673744 603259 673750 603311
rect 673802 603299 673808 603311
rect 675376 603299 675382 603311
rect 673802 603271 675382 603299
rect 673802 603259 673808 603271
rect 675376 603259 675382 603271
rect 675434 603259 675440 603311
rect 673648 602667 673654 602719
rect 673706 602707 673712 602719
rect 675376 602707 675382 602719
rect 673706 602679 675382 602707
rect 673706 602667 673712 602679
rect 675376 602667 675382 602679
rect 675434 602667 675440 602719
rect 656560 602075 656566 602127
rect 656618 602115 656624 602127
rect 674896 602115 674902 602127
rect 656618 602087 674902 602115
rect 656618 602075 656624 602087
rect 674896 602075 674902 602087
rect 674954 602075 674960 602127
rect 653968 602001 653974 602053
rect 654026 602041 654032 602053
rect 674992 602041 674998 602053
rect 654026 602013 674998 602041
rect 654026 602001 654032 602013
rect 674992 602001 674998 602013
rect 675050 602001 675056 602053
rect 41584 601631 41590 601683
rect 41642 601671 41648 601683
rect 50320 601671 50326 601683
rect 41642 601643 50326 601671
rect 41642 601631 41648 601643
rect 50320 601631 50326 601643
rect 50378 601631 50384 601683
rect 41776 601335 41782 601387
rect 41834 601375 41840 601387
rect 47728 601375 47734 601387
rect 41834 601347 47734 601375
rect 41834 601335 41840 601347
rect 47728 601335 47734 601347
rect 47786 601335 47792 601387
rect 41776 600743 41782 600795
rect 41834 600783 41840 600795
rect 47824 600783 47830 600795
rect 41834 600755 47830 600783
rect 41834 600743 41840 600755
rect 47824 600743 47830 600755
rect 47882 600743 47888 600795
rect 41776 600373 41782 600425
rect 41834 600413 41840 600425
rect 43312 600413 43318 600425
rect 41834 600385 43318 600413
rect 41834 600373 41840 600385
rect 43312 600373 43318 600385
rect 43370 600373 43376 600425
rect 41776 599781 41782 599833
rect 41834 599821 41840 599833
rect 43600 599821 43606 599833
rect 41834 599793 43606 599821
rect 41834 599781 41840 599793
rect 43600 599781 43606 599793
rect 43658 599781 43664 599833
rect 673456 599781 673462 599833
rect 673514 599821 673520 599833
rect 675376 599821 675382 599833
rect 673514 599793 675382 599821
rect 673514 599781 673520 599793
rect 675376 599781 675382 599793
rect 675434 599781 675440 599833
rect 41776 599263 41782 599315
rect 41834 599303 41840 599315
rect 43408 599303 43414 599315
rect 41834 599275 43414 599303
rect 41834 599263 41840 599275
rect 43408 599263 43414 599275
rect 43466 599263 43472 599315
rect 673552 599263 673558 599315
rect 673610 599303 673616 599315
rect 675088 599303 675094 599315
rect 673610 599275 675094 599303
rect 673610 599263 673616 599275
rect 675088 599263 675094 599275
rect 675146 599263 675152 599315
rect 39856 599041 39862 599093
rect 39914 599081 39920 599093
rect 41680 599081 41686 599093
rect 39914 599053 41686 599081
rect 39914 599041 39920 599053
rect 41680 599041 41686 599053
rect 41738 599041 41744 599093
rect 672880 598375 672886 598427
rect 672938 598415 672944 598427
rect 675184 598415 675190 598427
rect 672938 598387 675190 598415
rect 672938 598375 672944 598387
rect 675184 598375 675190 598387
rect 675242 598375 675248 598427
rect 41776 598301 41782 598353
rect 41834 598341 41840 598353
rect 43504 598341 43510 598353
rect 41834 598313 43510 598341
rect 41834 598301 41840 598313
rect 43504 598301 43510 598313
rect 43562 598301 43568 598353
rect 41776 597857 41782 597909
rect 41834 597897 41840 597909
rect 43216 597897 43222 597909
rect 41834 597869 43222 597897
rect 41834 597857 41840 597869
rect 43216 597857 43222 597869
rect 43274 597857 43280 597909
rect 41584 596599 41590 596651
rect 41642 596639 41648 596651
rect 42736 596639 42742 596651
rect 41642 596611 42742 596639
rect 41642 596599 41648 596611
rect 42736 596599 42742 596611
rect 42794 596599 42800 596651
rect 672976 596525 672982 596577
rect 673034 596565 673040 596577
rect 675088 596565 675094 596577
rect 673034 596537 675094 596565
rect 673034 596525 673040 596537
rect 675088 596525 675094 596537
rect 675146 596525 675152 596577
rect 43216 596155 43222 596207
rect 43274 596195 43280 596207
rect 45136 596195 45142 596207
rect 43274 596167 45142 596195
rect 43274 596155 43280 596167
rect 45136 596155 45142 596167
rect 45194 596155 45200 596207
rect 41584 595045 41590 595097
rect 41642 595085 41648 595097
rect 43120 595085 43126 595097
rect 41642 595057 43126 595085
rect 41642 595045 41648 595057
rect 43120 595045 43126 595057
rect 43178 595045 43184 595097
rect 41776 594897 41782 594949
rect 41834 594937 41840 594949
rect 42928 594937 42934 594949
rect 41834 594909 42934 594937
rect 41834 594897 41840 594909
rect 42928 594897 42934 594909
rect 42986 594897 42992 594949
rect 41584 593639 41590 593691
rect 41642 593679 41648 593691
rect 42832 593679 42838 593691
rect 41642 593651 42838 593679
rect 41642 593639 41648 593651
rect 42832 593639 42838 593651
rect 42890 593639 42896 593691
rect 41680 592159 41686 592211
rect 41738 592199 41744 592211
rect 42640 592199 42646 592211
rect 41738 592171 42646 592199
rect 41738 592159 41744 592171
rect 42640 592159 42646 592171
rect 42698 592159 42704 592211
rect 41968 590827 41974 590879
rect 42026 590867 42032 590879
rect 43024 590867 43030 590879
rect 42026 590839 43030 590867
rect 42026 590827 42032 590839
rect 43024 590827 43030 590839
rect 43082 590827 43088 590879
rect 41584 590679 41590 590731
rect 41642 590719 41648 590731
rect 42544 590719 42550 590731
rect 41642 590691 42550 590719
rect 41642 590679 41648 590691
rect 42544 590679 42550 590691
rect 42602 590679 42608 590731
rect 672784 590309 672790 590361
rect 672842 590349 672848 590361
rect 679696 590349 679702 590361
rect 672842 590321 679702 590349
rect 672842 590309 672848 590321
rect 679696 590309 679702 590321
rect 679754 590309 679760 590361
rect 42160 587571 42166 587623
rect 42218 587611 42224 587623
rect 43120 587611 43126 587623
rect 42218 587583 43126 587611
rect 42218 587571 42224 587583
rect 43120 587571 43126 587583
rect 43178 587571 43184 587623
rect 41584 587497 41590 587549
rect 41642 587537 41648 587549
rect 56080 587537 56086 587549
rect 41642 587509 56086 587537
rect 41642 587497 41648 587509
rect 56080 587497 56086 587509
rect 56138 587497 56144 587549
rect 42448 587423 42454 587475
rect 42506 587463 42512 587475
rect 42736 587463 42742 587475
rect 42506 587435 42742 587463
rect 42506 587423 42512 587435
rect 42736 587423 42742 587435
rect 42794 587423 42800 587475
rect 42832 587423 42838 587475
rect 42890 587463 42896 587475
rect 43312 587463 43318 587475
rect 42890 587435 43318 587463
rect 42890 587423 42896 587435
rect 43312 587423 43318 587435
rect 43370 587423 43376 587475
rect 41872 587053 41878 587105
rect 41930 587093 41936 587105
rect 43120 587093 43126 587105
rect 41930 587065 43126 587093
rect 41930 587053 41936 587065
rect 43120 587053 43126 587065
rect 43178 587053 43184 587105
rect 674608 586387 674614 586439
rect 674666 586427 674672 586439
rect 675088 586427 675094 586439
rect 674666 586399 675094 586427
rect 674666 586387 674672 586399
rect 675088 586387 675094 586399
rect 675146 586387 675152 586439
rect 42736 585795 42742 585847
rect 42794 585835 42800 585847
rect 43216 585835 43222 585847
rect 42794 585807 43222 585835
rect 42794 585795 42800 585807
rect 43216 585795 43222 585807
rect 43274 585795 43280 585847
rect 42256 585055 42262 585107
rect 42314 585095 42320 585107
rect 42544 585095 42550 585107
rect 42314 585067 42550 585095
rect 42314 585055 42320 585067
rect 42544 585055 42550 585067
rect 42602 585055 42608 585107
rect 42352 584907 42358 584959
rect 42410 584947 42416 584959
rect 43024 584947 43030 584959
rect 42410 584919 43030 584947
rect 42410 584907 42416 584919
rect 43024 584907 43030 584919
rect 43082 584907 43088 584959
rect 42448 584685 42454 584737
rect 42506 584725 42512 584737
rect 58960 584725 58966 584737
rect 42506 584697 58966 584725
rect 42506 584685 42512 584697
rect 58960 584685 58966 584697
rect 59018 584685 59024 584737
rect 41776 584167 41782 584219
rect 41834 584167 41840 584219
rect 42064 584167 42070 584219
rect 42122 584207 42128 584219
rect 42640 584207 42646 584219
rect 42122 584179 42646 584207
rect 42122 584167 42128 584179
rect 42640 584167 42646 584179
rect 42698 584167 42704 584219
rect 41794 583997 41822 584167
rect 41776 583945 41782 583997
rect 41834 583945 41840 583997
rect 42256 582243 42262 582295
rect 42314 582283 42320 582295
rect 42314 582255 42398 582283
rect 42314 582243 42320 582255
rect 42370 582073 42398 582255
rect 42352 582021 42358 582073
rect 42410 582021 42416 582073
rect 42352 581059 42358 581111
rect 42410 581059 42416 581111
rect 42370 580741 42398 581059
rect 42352 580689 42358 580741
rect 42410 580689 42416 580741
rect 42352 579875 42358 579927
rect 42410 579915 42416 579927
rect 42410 579887 42590 579915
rect 42410 579875 42416 579887
rect 42562 579853 42590 579887
rect 42544 579801 42550 579853
rect 42602 579801 42608 579853
rect 42448 578987 42454 579039
rect 42506 579027 42512 579039
rect 47920 579027 47926 579039
rect 42506 578999 47926 579027
rect 42506 578987 42512 578999
rect 47920 578987 47926 578999
rect 47978 578987 47984 579039
rect 42352 578913 42358 578965
rect 42410 578953 42416 578965
rect 42928 578953 42934 578965
rect 42410 578925 42934 578953
rect 42410 578913 42416 578925
rect 42928 578913 42934 578925
rect 42986 578913 42992 578965
rect 42928 578765 42934 578817
rect 42986 578805 42992 578817
rect 43312 578805 43318 578817
rect 42986 578777 43318 578805
rect 42986 578765 42992 578777
rect 43312 578765 43318 578777
rect 43370 578765 43376 578817
rect 42256 578543 42262 578595
rect 42314 578583 42320 578595
rect 42736 578583 42742 578595
rect 42314 578555 42742 578583
rect 42314 578543 42320 578555
rect 42736 578543 42742 578555
rect 42794 578543 42800 578595
rect 42256 577729 42262 577781
rect 42314 577769 42320 577781
rect 42832 577769 42838 577781
rect 42314 577741 42838 577769
rect 42314 577729 42320 577741
rect 42832 577729 42838 577741
rect 42890 577729 42896 577781
rect 42448 576619 42454 576671
rect 42506 576659 42512 576671
rect 43024 576659 43030 576671
rect 42506 576631 43030 576659
rect 42506 576619 42512 576631
rect 43024 576619 43030 576631
rect 43082 576619 43088 576671
rect 655504 576619 655510 576671
rect 655562 576659 655568 576671
rect 676240 576659 676246 576671
rect 655562 576631 676246 576659
rect 655562 576619 655568 576631
rect 676240 576619 676246 576631
rect 676298 576619 676304 576671
rect 655312 576471 655318 576523
rect 655370 576511 655376 576523
rect 676144 576511 676150 576523
rect 655370 576483 676150 576511
rect 655370 576471 655376 576483
rect 676144 576471 676150 576483
rect 676202 576471 676208 576523
rect 655120 576323 655126 576375
rect 655178 576363 655184 576375
rect 676336 576363 676342 576375
rect 655178 576335 676342 576363
rect 655178 576323 655184 576335
rect 676336 576323 676342 576335
rect 676394 576323 676400 576375
rect 672784 576175 672790 576227
rect 672842 576215 672848 576227
rect 676240 576215 676246 576227
rect 672842 576187 676246 576215
rect 672842 576175 672848 576187
rect 676240 576175 676246 576187
rect 676298 576175 676304 576227
rect 674224 575953 674230 576005
rect 674282 575993 674288 576005
rect 676048 575993 676054 576005
rect 674282 575965 676054 575993
rect 674282 575953 674288 575965
rect 676048 575953 676054 575965
rect 676106 575953 676112 576005
rect 670768 575879 670774 575931
rect 670826 575919 670832 575931
rect 675952 575919 675958 575931
rect 670826 575891 675958 575919
rect 670826 575879 670832 575891
rect 675952 575879 675958 575891
rect 676010 575879 676016 575931
rect 672592 575435 672598 575487
rect 672650 575475 672656 575487
rect 675952 575475 675958 575487
rect 672650 575447 675958 575475
rect 672650 575435 672656 575447
rect 675952 575435 675958 575447
rect 676010 575435 676016 575487
rect 670864 574917 670870 574969
rect 670922 574957 670928 574969
rect 675952 574957 675958 574969
rect 670922 574929 675958 574957
rect 670922 574917 670928 574929
rect 675952 574917 675958 574929
rect 676010 574917 676016 574969
rect 672688 574103 672694 574155
rect 672746 574143 672752 574155
rect 676240 574143 676246 574155
rect 672746 574115 676246 574143
rect 672746 574103 672752 574115
rect 676240 574103 676246 574115
rect 676298 574103 676304 574155
rect 42064 573215 42070 573267
rect 42122 573255 42128 573267
rect 42928 573255 42934 573267
rect 42122 573227 42934 573255
rect 42122 573215 42128 573227
rect 42928 573215 42934 573227
rect 42986 573215 42992 573267
rect 669904 573215 669910 573267
rect 669962 573255 669968 573267
rect 670864 573255 670870 573267
rect 669962 573227 670870 573255
rect 669962 573215 669968 573227
rect 670864 573215 670870 573227
rect 670922 573215 670928 573267
rect 42448 573141 42454 573193
rect 42506 573181 42512 573193
rect 58192 573181 58198 573193
rect 42506 573153 58198 573181
rect 42506 573141 42512 573153
rect 58192 573141 58198 573153
rect 58250 573141 58256 573193
rect 670096 573141 670102 573193
rect 670154 573181 670160 573193
rect 670768 573181 670774 573193
rect 670154 573153 670774 573181
rect 670154 573141 670160 573153
rect 670768 573141 670774 573153
rect 670826 573141 670832 573193
rect 47824 573067 47830 573119
rect 47882 573107 47888 573119
rect 58960 573107 58966 573119
rect 47882 573079 58966 573107
rect 47882 573067 47888 573079
rect 58960 573067 58966 573079
rect 59018 573067 59024 573119
rect 674128 573067 674134 573119
rect 674186 573107 674192 573119
rect 676048 573107 676054 573119
rect 674186 573079 676054 573107
rect 674186 573067 674192 573079
rect 676048 573067 676054 573079
rect 676106 573067 676112 573119
rect 47920 572993 47926 573045
rect 47978 573033 47984 573045
rect 59632 573033 59638 573045
rect 47978 573005 59638 573033
rect 47978 572993 47984 573005
rect 59632 572993 59638 573005
rect 59690 572993 59696 573045
rect 42160 572623 42166 572675
rect 42218 572663 42224 572675
rect 42832 572663 42838 572675
rect 42218 572635 42838 572663
rect 42218 572623 42224 572635
rect 42832 572623 42838 572635
rect 42890 572623 42896 572675
rect 42064 570995 42070 571047
rect 42122 571035 42128 571047
rect 43120 571035 43126 571047
rect 42122 571007 43126 571035
rect 42122 570995 42128 571007
rect 43120 570995 43126 571007
rect 43178 570995 43184 571047
rect 42352 570403 42358 570455
rect 42410 570443 42416 570455
rect 42544 570443 42550 570455
rect 42410 570415 42550 570443
rect 42410 570403 42416 570415
rect 42544 570403 42550 570415
rect 42602 570403 42608 570455
rect 50320 570181 50326 570233
rect 50378 570221 50384 570233
rect 59344 570221 59350 570233
rect 50378 570193 59350 570221
rect 50378 570181 50384 570193
rect 59344 570181 59350 570193
rect 59402 570181 59408 570233
rect 47728 570107 47734 570159
rect 47786 570147 47792 570159
rect 59536 570147 59542 570159
rect 47786 570119 59542 570147
rect 47786 570107 47792 570119
rect 59536 570107 59542 570119
rect 59594 570107 59600 570159
rect 673360 569515 673366 569567
rect 673418 569555 673424 569567
rect 676048 569555 676054 569567
rect 673418 569527 676054 569555
rect 673418 569515 673424 569527
rect 676048 569515 676054 569527
rect 676106 569515 676112 569567
rect 673264 569145 673270 569197
rect 673322 569185 673328 569197
rect 676240 569185 676246 569197
rect 673322 569157 676246 569185
rect 673322 569145 673328 569157
rect 676240 569145 676246 569157
rect 676298 569145 676304 569197
rect 673840 568405 673846 568457
rect 673898 568445 673904 568457
rect 676048 568445 676054 568457
rect 673898 568417 676054 568445
rect 673898 568405 673904 568417
rect 676048 568405 676054 568417
rect 676106 568405 676112 568457
rect 673072 567961 673078 568013
rect 673130 568001 673136 568013
rect 676048 568001 676054 568013
rect 673130 567973 676054 568001
rect 673130 567961 673136 567973
rect 676048 567961 676054 567973
rect 676106 567961 676112 568013
rect 673168 567665 673174 567717
rect 673226 567705 673232 567717
rect 676240 567705 676246 567717
rect 673226 567677 676246 567705
rect 673226 567665 673232 567677
rect 676240 567665 676246 567677
rect 676298 567665 676304 567717
rect 655696 567443 655702 567495
rect 655754 567483 655760 567495
rect 675376 567483 675382 567495
rect 655754 567455 675382 567483
rect 655754 567443 655760 567455
rect 675376 567443 675382 567455
rect 675434 567443 675440 567495
rect 649840 564483 649846 564535
rect 649898 564523 649904 564535
rect 679792 564523 679798 564535
rect 649898 564495 679798 564523
rect 649898 564483 649904 564495
rect 679792 564483 679798 564495
rect 679850 564483 679856 564535
rect 674032 559525 674038 559577
rect 674090 559565 674096 559577
rect 675376 559565 675382 559577
rect 674090 559537 675382 559565
rect 674090 559525 674096 559537
rect 675376 559525 675382 559537
rect 675434 559525 675440 559577
rect 656560 558785 656566 558837
rect 656618 558825 656624 558837
rect 675184 558825 675190 558837
rect 656618 558797 675190 558825
rect 656618 558785 656624 558797
rect 675184 558785 675190 558797
rect 675242 558785 675248 558837
rect 674800 558045 674806 558097
rect 674858 558085 674864 558097
rect 675376 558085 675382 558097
rect 674858 558057 675382 558085
rect 674858 558045 674864 558057
rect 675376 558045 675382 558057
rect 675434 558045 675440 558097
rect 654160 555825 654166 555877
rect 654218 555865 654224 555877
rect 675088 555865 675094 555877
rect 654218 555837 675094 555865
rect 654218 555825 654224 555837
rect 675088 555825 675094 555837
rect 675146 555825 675152 555877
rect 674320 555233 674326 555285
rect 674378 555273 674384 555285
rect 675472 555273 675478 555285
rect 674378 555245 675478 555273
rect 674378 555233 674384 555245
rect 675472 555233 675478 555245
rect 675530 555233 675536 555285
rect 674992 553753 674998 553805
rect 675050 553793 675056 553805
rect 675472 553793 675478 553805
rect 675050 553765 675478 553793
rect 675050 553753 675056 553765
rect 675472 553753 675478 553765
rect 675530 553753 675536 553805
rect 673840 553309 673846 553361
rect 673898 553349 673904 553361
rect 675376 553349 675382 553361
rect 673898 553321 675382 553349
rect 673898 553309 673904 553321
rect 675376 553309 675382 553321
rect 675434 553309 675440 553361
rect 674224 551903 674230 551955
rect 674282 551943 674288 551955
rect 675472 551943 675478 551955
rect 674282 551915 675478 551943
rect 674282 551903 674288 551915
rect 675472 551903 675478 551915
rect 675530 551903 675536 551955
rect 674512 548869 674518 548921
rect 674570 548909 674576 548921
rect 675088 548909 675094 548921
rect 674570 548881 675094 548909
rect 674570 548869 674576 548881
rect 675088 548869 675094 548881
rect 675146 548869 675152 548921
rect 672784 547167 672790 547219
rect 672842 547207 672848 547219
rect 679696 547207 679702 547219
rect 672842 547179 679702 547207
rect 672842 547167 672848 547179
rect 679696 547167 679702 547179
rect 679754 547167 679760 547219
rect 674416 543615 674422 543667
rect 674474 543655 674480 543667
rect 675088 543655 675094 543667
rect 674474 543627 675094 543655
rect 674474 543615 674480 543627
rect 675088 543615 675094 543627
rect 675146 543615 675152 543667
rect 42352 541543 42358 541595
rect 42410 541583 42416 541595
rect 57712 541583 57718 541595
rect 42410 541555 57718 541583
rect 42410 541543 42416 541555
rect 57712 541543 57718 541555
rect 57770 541543 57776 541595
rect 42448 541469 42454 541521
rect 42506 541509 42512 541521
rect 57616 541509 57622 541521
rect 42506 541481 57622 541509
rect 42506 541469 42512 541481
rect 57616 541469 57622 541481
rect 57674 541469 57680 541521
rect 655600 533403 655606 533455
rect 655658 533443 655664 533455
rect 676048 533443 676054 533455
rect 655658 533415 676054 533443
rect 655658 533403 655664 533415
rect 676048 533403 676054 533415
rect 676106 533403 676112 533455
rect 655408 533255 655414 533307
rect 655466 533295 655472 533307
rect 676240 533295 676246 533307
rect 655466 533267 676246 533295
rect 655466 533255 655472 533267
rect 676240 533255 676246 533267
rect 676298 533255 676304 533307
rect 655216 533107 655222 533159
rect 655274 533147 655280 533159
rect 676144 533147 676150 533159
rect 655274 533119 676150 533147
rect 655274 533107 655280 533119
rect 676144 533107 676150 533119
rect 676202 533107 676208 533159
rect 674704 532737 674710 532789
rect 674762 532777 674768 532789
rect 676048 532777 676054 532789
rect 674762 532749 676054 532777
rect 674762 532737 674768 532749
rect 676048 532737 676054 532749
rect 676106 532737 676112 532789
rect 672592 532663 672598 532715
rect 672650 532703 672656 532715
rect 675952 532703 675958 532715
rect 672650 532675 675958 532703
rect 672650 532663 672656 532675
rect 675952 532663 675958 532675
rect 676010 532663 676016 532715
rect 672400 531479 672406 531531
rect 672458 531519 672464 531531
rect 672688 531519 672694 531531
rect 672458 531491 672694 531519
rect 672458 531479 672464 531491
rect 672688 531479 672694 531491
rect 672746 531519 672752 531531
rect 676240 531519 676246 531531
rect 672746 531491 676246 531519
rect 672746 531479 672752 531491
rect 676240 531479 676246 531491
rect 676298 531479 676304 531531
rect 42544 529925 42550 529977
rect 42602 529965 42608 529977
rect 58192 529965 58198 529977
rect 42602 529937 58198 529965
rect 42602 529925 42608 529937
rect 58192 529925 58198 529937
rect 58250 529925 58256 529977
rect 674608 529851 674614 529903
rect 674666 529891 674672 529903
rect 676048 529891 676054 529903
rect 674666 529863 676054 529891
rect 674666 529851 674672 529863
rect 676048 529851 676054 529863
rect 676106 529851 676112 529903
rect 673744 526669 673750 526721
rect 673802 526709 673808 526721
rect 676048 526709 676054 526721
rect 673802 526681 676054 526709
rect 673802 526669 673808 526681
rect 676048 526669 676054 526681
rect 676106 526669 676112 526721
rect 672976 526299 672982 526351
rect 673034 526339 673040 526351
rect 676048 526339 676054 526351
rect 673034 526311 676054 526339
rect 673034 526299 673040 526311
rect 676048 526299 676054 526311
rect 676106 526299 676112 526351
rect 673552 525929 673558 525981
rect 673610 525969 673616 525981
rect 676240 525969 676246 525981
rect 673610 525941 676246 525969
rect 673610 525929 673616 525941
rect 676240 525929 676246 525941
rect 676298 525929 676304 525981
rect 42064 525707 42070 525759
rect 42122 525747 42128 525759
rect 42544 525747 42550 525759
rect 42122 525719 42550 525747
rect 42122 525707 42128 525719
rect 42544 525707 42550 525719
rect 42602 525707 42608 525759
rect 673648 525189 673654 525241
rect 673706 525229 673712 525241
rect 676048 525229 676054 525241
rect 673706 525201 676054 525229
rect 673706 525189 673712 525201
rect 676048 525189 676054 525201
rect 676106 525189 676112 525241
rect 673456 524819 673462 524871
rect 673514 524859 673520 524871
rect 676048 524859 676054 524871
rect 673514 524831 676054 524859
rect 673514 524819 673520 524831
rect 676048 524819 676054 524831
rect 676106 524819 676112 524871
rect 672880 524449 672886 524501
rect 672938 524489 672944 524501
rect 676240 524489 676246 524501
rect 672938 524461 676246 524489
rect 672938 524449 672944 524461
rect 676240 524449 676246 524461
rect 676298 524449 676304 524501
rect 50320 524301 50326 524353
rect 50378 524341 50384 524353
rect 58576 524341 58582 524353
rect 50378 524313 58582 524341
rect 50378 524301 50384 524313
rect 58576 524301 58582 524313
rect 58634 524301 58640 524353
rect 47728 524227 47734 524279
rect 47786 524267 47792 524279
rect 59344 524267 59350 524279
rect 47786 524239 59350 524267
rect 47786 524227 47792 524239
rect 59344 524227 59350 524239
rect 59402 524227 59408 524279
rect 42256 522229 42262 522281
rect 42314 522269 42320 522281
rect 42448 522269 42454 522281
rect 42314 522241 42454 522269
rect 42314 522229 42320 522241
rect 42448 522229 42454 522241
rect 42506 522229 42512 522281
rect 649936 521267 649942 521319
rect 649994 521307 650000 521319
rect 679792 521307 679798 521319
rect 649994 521279 679798 521307
rect 649994 521267 650000 521279
rect 679792 521267 679798 521279
rect 679850 521267 679856 521319
rect 676528 498253 676534 498305
rect 676586 498293 676592 498305
rect 679696 498293 679702 498305
rect 676586 498265 679702 498293
rect 676586 498253 676592 498265
rect 679696 498253 679702 498265
rect 679754 498253 679760 498305
rect 655504 490039 655510 490091
rect 655562 490079 655568 490091
rect 676240 490079 676246 490091
rect 655562 490051 676246 490079
rect 655562 490039 655568 490051
rect 676240 490039 676246 490051
rect 676298 490039 676304 490091
rect 655312 489891 655318 489943
rect 655370 489931 655376 489943
rect 676240 489931 676246 489943
rect 655370 489903 676246 489931
rect 655370 489891 655376 489903
rect 676240 489891 676246 489903
rect 676298 489891 676304 489943
rect 655120 489743 655126 489795
rect 655178 489783 655184 489795
rect 676144 489783 676150 489795
rect 655178 489755 676150 489783
rect 655178 489743 655184 489755
rect 676144 489743 676150 489755
rect 676202 489743 676208 489795
rect 676240 488707 676246 488759
rect 676298 488747 676304 488759
rect 676720 488747 676726 488759
rect 676298 488719 676726 488747
rect 676298 488707 676304 488719
rect 676720 488707 676726 488719
rect 676778 488707 676784 488759
rect 670288 488115 670294 488167
rect 670346 488155 670352 488167
rect 676048 488155 676054 488167
rect 670346 488127 676054 488155
rect 670346 488115 670352 488127
rect 676048 488115 676054 488127
rect 676106 488155 676112 488167
rect 676624 488155 676630 488167
rect 676106 488127 676630 488155
rect 676106 488115 676112 488127
rect 676624 488115 676630 488127
rect 676682 488115 676688 488167
rect 670480 487079 670486 487131
rect 670538 487119 670544 487131
rect 676240 487119 676246 487131
rect 670538 487091 676246 487119
rect 670538 487079 670544 487091
rect 676240 487079 676246 487091
rect 676298 487079 676304 487131
rect 672496 486783 672502 486835
rect 672554 486823 672560 486835
rect 676048 486823 676054 486835
rect 672554 486795 676054 486823
rect 672554 486783 672560 486795
rect 676048 486783 676054 486795
rect 676106 486783 676112 486835
rect 674512 486635 674518 486687
rect 674570 486675 674576 486687
rect 676048 486675 676054 486687
rect 674570 486647 676054 486675
rect 674570 486635 674576 486647
rect 676048 486635 676054 486647
rect 676106 486635 676112 486687
rect 674032 486561 674038 486613
rect 674090 486601 674096 486613
rect 676240 486601 676246 486613
rect 674090 486573 676246 486601
rect 674090 486561 674096 486573
rect 676240 486561 676246 486573
rect 676298 486561 676304 486613
rect 674320 485673 674326 485725
rect 674378 485713 674384 485725
rect 676048 485713 676054 485725
rect 674378 485685 676054 485713
rect 674378 485673 674384 485685
rect 676048 485673 676054 485685
rect 676106 485673 676112 485725
rect 674800 483749 674806 483801
rect 674858 483789 674864 483801
rect 676048 483789 676054 483801
rect 674858 483761 676054 483789
rect 674858 483749 674864 483761
rect 676048 483749 676054 483761
rect 676106 483749 676112 483801
rect 674416 483675 674422 483727
rect 674474 483715 674480 483727
rect 675952 483715 675958 483727
rect 674474 483687 675958 483715
rect 674474 483675 674480 483687
rect 675952 483675 675958 483687
rect 676010 483675 676016 483727
rect 674992 483601 674998 483653
rect 675050 483641 675056 483653
rect 676240 483641 676246 483653
rect 675050 483613 676246 483641
rect 675050 483601 675056 483613
rect 676240 483601 676246 483613
rect 676298 483601 676304 483653
rect 674224 482121 674230 482173
rect 674282 482161 674288 482173
rect 676048 482161 676054 482173
rect 674282 482133 676054 482161
rect 674282 482121 674288 482133
rect 676048 482121 676054 482133
rect 676106 482121 676112 482173
rect 673840 480049 673846 480101
rect 673898 480089 673904 480101
rect 676240 480089 676246 480101
rect 673898 480061 676246 480089
rect 673898 480049 673904 480061
rect 676240 480049 676246 480061
rect 676298 480049 676304 480101
rect 650032 478125 650038 478177
rect 650090 478165 650096 478177
rect 679888 478165 679894 478177
rect 650090 478137 679894 478165
rect 650090 478125 650096 478137
rect 679888 478125 679894 478137
rect 679946 478125 679952 478177
rect 41863 476105 41915 476111
rect 50320 476093 50326 476105
rect 41915 476065 50326 476093
rect 50320 476053 50326 476065
rect 50378 476053 50384 476105
rect 41863 476047 41915 476053
rect 41844 475535 41850 475587
rect 41902 475575 41908 475587
rect 47728 475575 47734 475587
rect 41902 475547 47734 475575
rect 41902 475535 41908 475547
rect 47728 475535 47734 475547
rect 47786 475535 47792 475587
rect 42035 474573 42041 474625
rect 42093 474613 42099 474625
rect 43600 474613 43606 474625
rect 42093 474585 43606 474613
rect 42093 474573 42099 474585
rect 43600 474573 43606 474585
rect 43658 474573 43664 474625
rect 41776 472353 41782 472405
rect 41834 472393 41840 472405
rect 58960 472393 58966 472405
rect 41834 472365 58966 472393
rect 41834 472353 41840 472365
rect 58960 472353 58966 472365
rect 59018 472353 59024 472405
rect 41776 463547 41782 463599
rect 41834 463587 41840 463599
rect 47728 463587 47734 463599
rect 41834 463559 47734 463587
rect 41834 463547 41840 463559
rect 47728 463547 47734 463559
rect 47786 463547 47792 463599
rect 34480 463103 34486 463155
rect 34538 463143 34544 463155
rect 41776 463143 41782 463155
rect 34538 463115 41782 463143
rect 34538 463103 34544 463115
rect 41776 463103 41782 463115
rect 41834 463103 41840 463155
rect 673840 440607 673846 440659
rect 673898 440647 673904 440659
rect 675280 440647 675286 440659
rect 673898 440619 675286 440647
rect 673898 440607 673904 440619
rect 675280 440607 675286 440619
rect 675338 440607 675344 440659
rect 39664 437835 39670 437847
rect 38722 437807 39670 437835
rect 25840 437721 25846 437773
rect 25898 437761 25904 437773
rect 38722 437761 38750 437807
rect 39664 437795 39670 437807
rect 39722 437835 39728 437847
rect 62512 437835 62518 437847
rect 39722 437807 62518 437835
rect 39722 437795 39728 437807
rect 62512 437795 62518 437807
rect 62570 437795 62576 437847
rect 25898 437733 38750 437761
rect 25898 437721 25904 437733
rect 670960 434909 670966 434961
rect 671018 434949 671024 434961
rect 672496 434949 672502 434961
rect 671018 434921 672502 434949
rect 671018 434909 671024 434921
rect 672496 434909 672502 434921
rect 672554 434909 672560 434961
rect 41584 428443 41590 428495
rect 41642 428483 41648 428495
rect 48016 428483 48022 428495
rect 41642 428455 48022 428483
rect 41642 428443 41648 428455
rect 48016 428443 48022 428455
rect 48074 428443 48080 428495
rect 41776 428073 41782 428125
rect 41834 428113 41840 428125
rect 47920 428113 47926 428125
rect 41834 428085 47926 428113
rect 41834 428073 41840 428085
rect 47920 428073 47926 428085
rect 47978 428073 47984 428125
rect 39760 427629 39766 427681
rect 39818 427669 39824 427681
rect 41584 427669 41590 427681
rect 39818 427641 41590 427669
rect 39818 427629 39824 427641
rect 41584 427629 41590 427641
rect 41642 427629 41648 427681
rect 41776 427555 41782 427607
rect 41834 427595 41840 427607
rect 48112 427595 48118 427607
rect 41834 427567 48118 427595
rect 41834 427555 41840 427567
rect 48112 427555 48118 427567
rect 48170 427555 48176 427607
rect 41776 426519 41782 426571
rect 41834 426559 41840 426571
rect 43216 426559 43222 426571
rect 41834 426531 43222 426559
rect 41834 426519 41840 426531
rect 43216 426519 43222 426531
rect 43274 426519 43280 426571
rect 41584 424965 41590 425017
rect 41642 425005 41648 425017
rect 41642 424977 49113 425005
rect 41642 424965 41648 424977
rect 49085 423405 49113 424977
rect 62608 423405 62614 423417
rect 49085 423377 62614 423405
rect 62608 423365 62614 423377
rect 62666 423365 62672 423417
rect 40144 419119 40150 419171
rect 40202 419159 40208 419171
rect 42448 419159 42454 419171
rect 40202 419131 42454 419159
rect 40202 419119 40208 419131
rect 42448 419119 42454 419131
rect 42506 419119 42512 419171
rect 39952 419045 39958 419097
rect 40010 419085 40016 419097
rect 42928 419085 42934 419097
rect 40010 419057 42934 419085
rect 40010 419045 40016 419057
rect 42928 419045 42934 419057
rect 42986 419045 42992 419097
rect 39856 418971 39862 419023
rect 39914 419011 39920 419023
rect 43024 419011 43030 419023
rect 39914 418983 43030 419011
rect 39914 418971 39920 418983
rect 43024 418971 43030 418983
rect 43082 418971 43088 419023
rect 41584 418083 41590 418135
rect 41642 418123 41648 418135
rect 42736 418123 42742 418135
rect 41642 418095 42742 418123
rect 41642 418083 41648 418095
rect 42736 418083 42742 418095
rect 42794 418083 42800 418135
rect 34480 417713 34486 417765
rect 34538 417753 34544 417765
rect 42352 417753 42358 417765
rect 34538 417725 42358 417753
rect 34538 417713 34544 417725
rect 42352 417713 42358 417725
rect 42410 417713 42416 417765
rect 41776 417195 41782 417247
rect 41834 417235 41840 417247
rect 42832 417235 42838 417247
rect 41834 417207 42838 417235
rect 41834 417195 41840 417207
rect 42832 417195 42838 417207
rect 42890 417195 42896 417247
rect 41584 416455 41590 416507
rect 41642 416495 41648 416507
rect 42640 416495 42646 416507
rect 41642 416467 42646 416495
rect 41642 416455 41648 416467
rect 42640 416455 42646 416467
rect 42698 416455 42704 416507
rect 41776 416085 41782 416137
rect 41834 416125 41840 416137
rect 47824 416125 47830 416137
rect 41834 416097 47830 416125
rect 41834 416085 41840 416097
rect 47824 416085 47830 416097
rect 47882 416085 47888 416137
rect 42160 409453 42166 409505
rect 42218 409493 42224 409505
rect 42448 409493 42454 409505
rect 42218 409465 42454 409493
rect 42218 409453 42224 409465
rect 42448 409453 42454 409465
rect 42506 409453 42512 409505
rect 42352 408121 42358 408173
rect 42410 408161 42416 408173
rect 42832 408161 42838 408173
rect 42410 408133 42838 408161
rect 42410 408121 42416 408133
rect 42832 408121 42838 408133
rect 42890 408121 42896 408173
rect 42160 408047 42166 408099
rect 42218 408087 42224 408099
rect 42544 408087 42550 408099
rect 42218 408059 42550 408087
rect 42218 408047 42224 408059
rect 42544 408047 42550 408059
rect 42602 408047 42608 408099
rect 42064 407973 42070 408025
rect 42122 408013 42128 408025
rect 42448 408013 42454 408025
rect 42122 407985 42454 408013
rect 42122 407973 42128 407985
rect 42448 407973 42454 407985
rect 42506 407973 42512 408025
rect 42064 407455 42070 407507
rect 42122 407495 42128 407507
rect 42736 407495 42742 407507
rect 42122 407467 42742 407495
rect 42122 407455 42128 407467
rect 42736 407455 42742 407467
rect 42794 407455 42800 407507
rect 42160 407011 42166 407063
rect 42218 407051 42224 407063
rect 42640 407051 42646 407063
rect 42218 407023 42646 407051
rect 42218 407011 42224 407023
rect 42640 407011 42646 407023
rect 42698 407011 42704 407063
rect 42256 406049 42262 406101
rect 42314 406089 42320 406101
rect 58480 406089 58486 406101
rect 42314 406061 58486 406089
rect 42314 406049 42320 406061
rect 58480 406049 58486 406061
rect 58538 406049 58544 406101
rect 42160 403163 42166 403215
rect 42218 403203 42224 403215
rect 43024 403203 43030 403215
rect 42218 403175 43030 403203
rect 42218 403163 42224 403175
rect 43024 403163 43030 403175
rect 43082 403163 43088 403215
rect 42448 403015 42454 403067
rect 42506 403055 42512 403067
rect 58768 403055 58774 403067
rect 42506 403027 58774 403055
rect 42506 403015 42512 403027
rect 58768 403015 58774 403027
rect 58826 403015 58832 403067
rect 673744 400573 673750 400625
rect 673802 400613 673808 400625
rect 675952 400613 675958 400625
rect 673802 400585 675958 400613
rect 673802 400573 673808 400585
rect 675952 400573 675958 400585
rect 676010 400573 676016 400625
rect 655504 400499 655510 400551
rect 655562 400539 655568 400551
rect 676048 400539 676054 400551
rect 655562 400511 676054 400539
rect 655562 400499 655568 400511
rect 676048 400499 676054 400511
rect 676106 400499 676112 400551
rect 655312 400425 655318 400477
rect 655370 400465 655376 400477
rect 676240 400465 676246 400477
rect 655370 400437 676246 400465
rect 655370 400425 655376 400437
rect 676240 400425 676246 400437
rect 676298 400425 676304 400477
rect 655120 400351 655126 400403
rect 655178 400391 655184 400403
rect 676144 400391 676150 400403
rect 655178 400363 676150 400391
rect 655178 400351 655184 400363
rect 676144 400351 676150 400363
rect 676202 400351 676208 400403
rect 48016 400277 48022 400329
rect 48074 400317 48080 400329
rect 58192 400317 58198 400329
rect 48074 400289 58198 400317
rect 48074 400277 48080 400289
rect 58192 400277 58198 400289
rect 58250 400277 58256 400329
rect 672496 400277 672502 400329
rect 672554 400317 672560 400329
rect 673840 400317 673846 400329
rect 672554 400289 673846 400317
rect 672554 400277 672560 400289
rect 673840 400277 673846 400289
rect 673898 400317 673904 400329
rect 676240 400317 676246 400329
rect 673898 400289 676246 400317
rect 673898 400277 673904 400289
rect 676240 400277 676246 400289
rect 676298 400277 676304 400329
rect 48112 400203 48118 400255
rect 48170 400243 48176 400255
rect 58768 400243 58774 400255
rect 48170 400215 58774 400243
rect 48170 400203 48176 400215
rect 58768 400203 58774 400215
rect 58826 400203 58832 400255
rect 47920 400129 47926 400181
rect 47978 400169 47984 400181
rect 59728 400169 59734 400181
rect 47978 400141 59734 400169
rect 47978 400129 47984 400141
rect 59728 400129 59734 400141
rect 59786 400129 59792 400181
rect 670960 399019 670966 399071
rect 671018 399059 671024 399071
rect 676048 399059 676054 399071
rect 671018 399031 676054 399059
rect 671018 399019 671024 399031
rect 676048 399019 676054 399031
rect 676106 399019 676112 399071
rect 42064 394505 42070 394557
rect 42122 394545 42128 394557
rect 57616 394545 57622 394557
rect 42122 394517 57622 394545
rect 42122 394505 42128 394517
rect 57616 394505 57622 394517
rect 57674 394505 57680 394557
rect 675184 392507 675190 392559
rect 675242 392547 675248 392559
rect 676240 392547 676246 392559
rect 675242 392519 676246 392547
rect 675242 392507 675248 392519
rect 676240 392507 676246 392519
rect 676298 392507 676304 392559
rect 674992 391693 674998 391745
rect 675050 391733 675056 391745
rect 676240 391733 676246 391745
rect 675050 391705 676246 391733
rect 675050 391693 675056 391705
rect 676240 391693 676246 391705
rect 676298 391693 676304 391745
rect 650128 388807 650134 388859
rect 650186 388847 650192 388859
rect 679792 388847 679798 388859
rect 650186 388819 679798 388847
rect 650186 388807 650192 388819
rect 679792 388807 679798 388819
rect 679850 388807 679856 388859
rect 41584 385921 41590 385973
rect 41642 385961 41648 385973
rect 48016 385961 48022 385973
rect 41642 385933 48022 385961
rect 41642 385921 41648 385933
rect 48016 385921 48022 385933
rect 48074 385921 48080 385973
rect 675088 385921 675094 385973
rect 675146 385961 675152 385973
rect 675376 385961 675382 385973
rect 675146 385933 675382 385961
rect 675146 385921 675152 385933
rect 675376 385921 675382 385933
rect 675434 385921 675440 385973
rect 41584 385255 41590 385307
rect 41642 385295 41648 385307
rect 48208 385295 48214 385307
rect 41642 385267 48214 385295
rect 41642 385255 41648 385267
rect 48208 385255 48214 385267
rect 48266 385255 48272 385307
rect 41872 384959 41878 385011
rect 41930 384999 41936 385011
rect 48112 384999 48118 385011
rect 41930 384971 48118 384999
rect 41930 384959 41936 384971
rect 48112 384959 48118 384971
rect 48170 384959 48176 385011
rect 41584 384737 41590 384789
rect 41642 384777 41648 384789
rect 43216 384777 43222 384789
rect 41642 384749 43222 384777
rect 41642 384737 41648 384749
rect 43216 384737 43222 384749
rect 43274 384737 43280 384789
rect 41584 383775 41590 383827
rect 41642 383815 41648 383827
rect 43312 383815 43318 383827
rect 41642 383787 43318 383815
rect 41642 383775 41648 383787
rect 43312 383775 43318 383787
rect 43370 383775 43376 383827
rect 41584 382295 41590 382347
rect 41642 382335 41648 382347
rect 43216 382335 43222 382347
rect 41642 382307 43222 382335
rect 41642 382295 41648 382307
rect 43216 382295 43222 382307
rect 43274 382295 43280 382347
rect 656560 381555 656566 381607
rect 656618 381595 656624 381607
rect 675088 381595 675094 381607
rect 656618 381567 675094 381595
rect 656618 381555 656624 381567
rect 675088 381555 675094 381567
rect 675146 381555 675152 381607
rect 41776 379483 41782 379535
rect 41834 379523 41840 379535
rect 42928 379523 42934 379535
rect 41834 379495 42934 379523
rect 41834 379483 41840 379495
rect 42928 379483 42934 379495
rect 42986 379483 42992 379535
rect 41584 377263 41590 377315
rect 41642 377303 41648 377315
rect 42832 377303 42838 377315
rect 41642 377275 42838 377303
rect 41642 377263 41648 377275
rect 42832 377263 42838 377275
rect 42890 377263 42896 377315
rect 41488 374303 41494 374355
rect 41546 374343 41552 374355
rect 42736 374343 42742 374355
rect 41546 374315 42742 374343
rect 41546 374303 41552 374315
rect 42736 374303 42742 374315
rect 42794 374303 42800 374355
rect 41776 374007 41782 374059
rect 41834 374047 41840 374059
rect 43024 374047 43030 374059
rect 41834 374019 43030 374047
rect 41834 374007 41840 374019
rect 43024 374007 43030 374019
rect 43082 374007 43088 374059
rect 37360 373859 37366 373911
rect 37418 373899 37424 373911
rect 41776 373899 41782 373911
rect 37418 373871 41782 373899
rect 37418 373859 37424 373871
rect 41776 373859 41782 373871
rect 41834 373859 41840 373911
rect 41584 373415 41590 373467
rect 41642 373455 41648 373467
rect 42544 373455 42550 373467
rect 41642 373427 42550 373455
rect 41642 373415 41648 373427
rect 42544 373415 42550 373427
rect 42602 373415 42608 373467
rect 41584 373267 41590 373319
rect 41642 373307 41648 373319
rect 47920 373307 47926 373319
rect 41642 373279 47926 373307
rect 41642 373267 41648 373279
rect 47920 373267 47926 373279
rect 47978 373267 47984 373319
rect 39952 372453 39958 372505
rect 40010 372493 40016 372505
rect 42256 372493 42262 372505
rect 40010 372465 42262 372493
rect 40010 372453 40016 372465
rect 42256 372453 42262 372465
rect 42314 372453 42320 372505
rect 41680 371935 41686 371987
rect 41738 371975 41744 371987
rect 42640 371975 42646 371987
rect 41738 371947 42646 371975
rect 41738 371935 41744 371947
rect 42640 371935 42646 371947
rect 42698 371935 42704 371987
rect 41776 370159 41782 370211
rect 41834 370159 41840 370211
rect 41794 369989 41822 370159
rect 41776 369937 41782 369989
rect 41834 369937 41840 369989
rect 42160 366533 42166 366585
rect 42218 366573 42224 366585
rect 42448 366573 42454 366585
rect 42218 366545 42454 366573
rect 42218 366533 42224 366545
rect 42448 366533 42454 366545
rect 42506 366533 42512 366585
rect 42256 364979 42262 365031
rect 42314 365019 42320 365031
rect 42544 365019 42550 365031
rect 42314 364991 42550 365019
rect 42314 364979 42320 364991
rect 42544 364979 42550 364991
rect 42602 364979 42608 365031
rect 42256 364461 42262 364513
rect 42314 364501 42320 364513
rect 42736 364501 42742 364513
rect 42314 364473 42742 364501
rect 42314 364461 42320 364473
rect 42736 364461 42742 364473
rect 42794 364461 42800 364513
rect 42160 363795 42166 363847
rect 42218 363835 42224 363847
rect 42640 363835 42646 363847
rect 42218 363807 42646 363835
rect 42218 363795 42224 363807
rect 42640 363795 42646 363807
rect 42698 363795 42704 363847
rect 42256 363721 42262 363773
rect 42314 363761 42320 363773
rect 43024 363761 43030 363773
rect 42314 363733 43030 363761
rect 42314 363721 42320 363733
rect 43024 363721 43030 363733
rect 43082 363721 43088 363773
rect 42064 362907 42070 362959
rect 42122 362947 42128 362959
rect 42928 362947 42934 362959
rect 42122 362919 42934 362947
rect 42122 362907 42128 362919
rect 42928 362907 42934 362919
rect 42986 362907 42992 362959
rect 42448 362833 42454 362885
rect 42506 362873 42512 362885
rect 58480 362873 58486 362885
rect 42506 362845 58486 362873
rect 42506 362833 42512 362845
rect 58480 362833 58486 362845
rect 58538 362833 58544 362885
rect 42352 359947 42358 359999
rect 42410 359987 42416 359999
rect 59152 359987 59158 359999
rect 42410 359959 59158 359987
rect 42410 359947 42416 359959
rect 59152 359947 59158 359959
rect 59210 359947 59216 359999
rect 655312 357283 655318 357335
rect 655370 357323 655376 357335
rect 676144 357323 676150 357335
rect 655370 357295 676150 357323
rect 655370 357283 655376 357295
rect 676144 357283 676150 357295
rect 676202 357283 676208 357335
rect 655216 357209 655222 357261
rect 655274 357249 655280 357261
rect 676240 357249 676246 357261
rect 655274 357221 676246 357249
rect 655274 357209 655280 357221
rect 676240 357209 676246 357221
rect 676298 357209 676304 357261
rect 655120 357135 655126 357187
rect 655178 357175 655184 357187
rect 676048 357175 676054 357187
rect 655178 357147 676054 357175
rect 655178 357135 655184 357147
rect 676048 357135 676054 357147
rect 676106 357135 676112 357187
rect 48016 357061 48022 357113
rect 48074 357101 48080 357113
rect 58192 357101 58198 357113
rect 48074 357073 58198 357101
rect 48074 357061 48080 357073
rect 58192 357061 58198 357073
rect 58250 357061 58256 357113
rect 48112 356987 48118 357039
rect 48170 357027 48176 357039
rect 59632 357027 59638 357039
rect 48170 356999 59638 357027
rect 48170 356987 48176 356999
rect 59632 356987 59638 356999
rect 59690 356987 59696 357039
rect 48208 356913 48214 356965
rect 48266 356953 48272 356965
rect 58576 356953 58582 356965
rect 48266 356925 58582 356953
rect 48266 356913 48272 356925
rect 58576 356913 58582 356925
rect 58634 356913 58640 356965
rect 673744 356765 673750 356817
rect 673802 356805 673808 356817
rect 676048 356805 676054 356817
rect 673802 356777 676054 356805
rect 673802 356765 673808 356777
rect 676048 356765 676054 356777
rect 676106 356765 676112 356817
rect 674512 352399 674518 352451
rect 674570 352439 674576 352451
rect 676048 352439 676054 352451
rect 674570 352411 676054 352439
rect 674570 352399 674576 352411
rect 676048 352399 676054 352411
rect 676106 352399 676112 352451
rect 674800 351363 674806 351415
rect 674858 351403 674864 351415
rect 676048 351403 676054 351415
rect 674858 351375 676054 351403
rect 674858 351363 674864 351375
rect 676048 351363 676054 351375
rect 676106 351363 676112 351415
rect 42160 351289 42166 351341
rect 42218 351329 42224 351341
rect 57616 351329 57622 351341
rect 42218 351301 57622 351329
rect 42218 351289 42224 351301
rect 57616 351289 57622 351301
rect 57674 351289 57680 351341
rect 674128 348551 674134 348603
rect 674186 348591 674192 348603
rect 676240 348591 676246 348603
rect 674186 348563 676246 348591
rect 674186 348551 674192 348563
rect 676240 348551 676246 348563
rect 676298 348551 676304 348603
rect 675184 348477 675190 348529
rect 675242 348517 675248 348529
rect 676048 348517 676054 348529
rect 675242 348489 676054 348517
rect 675242 348477 675248 348489
rect 676048 348477 676054 348489
rect 676106 348477 676112 348529
rect 650224 345813 650230 345865
rect 650282 345853 650288 345865
rect 679888 345853 679894 345865
rect 650282 345825 679894 345853
rect 650282 345813 650288 345825
rect 679888 345813 679894 345825
rect 679946 345813 679952 345865
rect 674896 345739 674902 345791
rect 674954 345779 674960 345791
rect 675952 345779 675958 345791
rect 674954 345751 675958 345779
rect 674954 345739 674960 345751
rect 675952 345739 675958 345751
rect 676010 345739 676016 345791
rect 674992 345665 674998 345717
rect 675050 345705 675056 345717
rect 676048 345705 676054 345717
rect 675050 345677 676054 345705
rect 675050 345665 675056 345677
rect 676048 345665 676054 345677
rect 676106 345665 676112 345717
rect 675088 345591 675094 345643
rect 675146 345631 675152 345643
rect 676240 345631 676246 345643
rect 675146 345603 676246 345631
rect 675146 345591 675152 345603
rect 676240 345591 676246 345603
rect 676298 345591 676304 345643
rect 41776 342779 41782 342831
rect 41834 342819 41840 342831
rect 48016 342819 48022 342831
rect 41834 342791 48022 342819
rect 41834 342779 41840 342791
rect 48016 342779 48022 342791
rect 48074 342779 48080 342831
rect 41776 342261 41782 342313
rect 41834 342301 41840 342313
rect 48112 342301 48118 342313
rect 41834 342273 48118 342301
rect 41834 342261 41840 342273
rect 48112 342261 48118 342273
rect 48170 342261 48176 342313
rect 41776 341743 41782 341795
rect 41834 341783 41840 341795
rect 48208 341783 48214 341795
rect 41834 341755 48214 341783
rect 41834 341743 41840 341755
rect 48208 341743 48214 341755
rect 48266 341743 48272 341795
rect 41776 341373 41782 341425
rect 41834 341413 41840 341425
rect 43312 341413 43318 341425
rect 41834 341385 43318 341413
rect 41834 341373 41840 341385
rect 43312 341373 43318 341385
rect 43370 341373 43376 341425
rect 675760 341373 675766 341425
rect 675818 341373 675824 341425
rect 675778 340759 675806 341373
rect 675760 340707 675766 340759
rect 675818 340707 675824 340759
rect 667792 340633 667798 340685
rect 667850 340673 667856 340685
rect 675472 340673 675478 340685
rect 667850 340645 675478 340673
rect 667850 340633 667856 340645
rect 675472 340633 675478 340645
rect 675530 340633 675536 340685
rect 41584 340559 41590 340611
rect 41642 340599 41648 340611
rect 43504 340599 43510 340611
rect 41642 340571 43510 340599
rect 41642 340559 41648 340571
rect 43504 340559 43510 340571
rect 43562 340559 43568 340611
rect 41776 340263 41782 340315
rect 41834 340303 41840 340315
rect 43408 340303 43414 340315
rect 41834 340275 43414 340303
rect 41834 340263 41840 340275
rect 43408 340263 43414 340275
rect 43466 340263 43472 340315
rect 674800 339745 674806 339797
rect 674858 339785 674864 339797
rect 675280 339785 675286 339797
rect 674858 339757 675286 339785
rect 674858 339745 674864 339757
rect 675280 339745 675286 339757
rect 675338 339745 675344 339797
rect 674512 339523 674518 339575
rect 674570 339563 674576 339575
rect 675376 339563 675382 339575
rect 674570 339535 675382 339563
rect 674570 339523 674576 339535
rect 675376 339523 675382 339535
rect 675434 339523 675440 339575
rect 41584 339079 41590 339131
rect 41642 339119 41648 339131
rect 43312 339119 43318 339131
rect 41642 339091 43318 339119
rect 41642 339079 41648 339091
rect 43312 339079 43318 339091
rect 43370 339079 43376 339131
rect 674128 336563 674134 336615
rect 674186 336603 674192 336615
rect 675376 336603 675382 336615
rect 674186 336575 675382 336603
rect 674186 336563 674192 336575
rect 675376 336563 675382 336575
rect 675434 336563 675440 336615
rect 41584 334195 41590 334247
rect 41642 334235 41648 334247
rect 42928 334235 42934 334247
rect 41642 334207 42934 334235
rect 41642 334195 41648 334207
rect 42928 334195 42934 334207
rect 42986 334195 42992 334247
rect 41872 334121 41878 334173
rect 41930 334161 41936 334173
rect 43024 334161 43030 334173
rect 41930 334133 43030 334161
rect 41930 334121 41936 334133
rect 43024 334121 43030 334133
rect 43082 334121 43088 334173
rect 41488 331087 41494 331139
rect 41546 331127 41552 331139
rect 42736 331127 42742 331139
rect 41546 331099 42742 331127
rect 41546 331087 41552 331099
rect 42736 331087 42742 331099
rect 42794 331087 42800 331139
rect 41392 331013 41398 331065
rect 41450 331053 41456 331065
rect 42832 331053 42838 331065
rect 41450 331025 42838 331053
rect 41450 331013 41456 331025
rect 42832 331013 42838 331025
rect 42890 331013 42896 331065
rect 39760 330643 39766 330695
rect 39818 330683 39824 330695
rect 42256 330683 42262 330695
rect 39818 330655 42262 330683
rect 39818 330643 39824 330655
rect 42256 330643 42262 330655
rect 42314 330643 42320 330695
rect 41872 330347 41878 330399
rect 41930 330387 41936 330399
rect 45232 330387 45238 330399
rect 41930 330359 45238 330387
rect 41930 330347 41936 330359
rect 45232 330347 45238 330359
rect 45290 330347 45296 330399
rect 41584 328571 41590 328623
rect 41642 328611 41648 328623
rect 42544 328611 42550 328623
rect 41642 328583 42550 328611
rect 41642 328571 41648 328583
rect 42544 328571 42550 328583
rect 42602 328571 42608 328623
rect 41680 328497 41686 328549
rect 41738 328537 41744 328549
rect 42640 328537 42646 328549
rect 41738 328509 42646 328537
rect 41738 328497 41744 328509
rect 42640 328497 42646 328509
rect 42698 328497 42704 328549
rect 654160 328275 654166 328327
rect 654218 328315 654224 328327
rect 667792 328315 667798 328327
rect 654218 328287 667798 328315
rect 654218 328275 654224 328287
rect 667792 328275 667798 328287
rect 667850 328275 667856 328327
rect 41776 327017 41782 327069
rect 41834 327017 41840 327069
rect 41794 326773 41822 327017
rect 41776 326721 41782 326773
rect 41834 326721 41840 326773
rect 42064 323317 42070 323369
rect 42122 323357 42128 323369
rect 42448 323357 42454 323369
rect 42122 323329 42454 323357
rect 42122 323317 42128 323329
rect 42448 323317 42454 323329
rect 42506 323317 42512 323369
rect 42256 321763 42262 321815
rect 42314 321803 42320 321815
rect 42544 321803 42550 321815
rect 42314 321775 42550 321803
rect 42314 321763 42320 321775
rect 42544 321763 42550 321775
rect 42602 321763 42608 321815
rect 42256 321245 42262 321297
rect 42314 321285 42320 321297
rect 42640 321285 42646 321297
rect 42314 321257 42646 321285
rect 42314 321245 42320 321257
rect 42640 321245 42646 321257
rect 42698 321245 42704 321297
rect 42160 321023 42166 321075
rect 42218 321063 42224 321075
rect 42736 321063 42742 321075
rect 42218 321035 42742 321063
rect 42218 321023 42224 321035
rect 42736 321023 42742 321035
rect 42794 321023 42800 321075
rect 42256 319913 42262 319965
rect 42314 319953 42320 319965
rect 42928 319953 42934 319965
rect 42314 319925 42934 319953
rect 42314 319913 42320 319925
rect 42928 319913 42934 319925
rect 42986 319913 42992 319965
rect 42448 319617 42454 319669
rect 42506 319657 42512 319669
rect 58480 319657 58486 319669
rect 42506 319629 58486 319657
rect 42506 319617 42512 319629
rect 58480 319617 58486 319629
rect 58538 319617 58544 319669
rect 42448 319395 42454 319447
rect 42506 319435 42512 319447
rect 42832 319435 42838 319447
rect 42506 319407 42838 319435
rect 42506 319395 42512 319407
rect 42832 319395 42838 319407
rect 42890 319395 42896 319447
rect 42448 316879 42454 316931
rect 42506 316919 42512 316931
rect 43024 316919 43030 316931
rect 42506 316891 43030 316919
rect 42506 316879 42512 316891
rect 43024 316879 43030 316891
rect 43082 316879 43088 316931
rect 42544 316731 42550 316783
rect 42602 316771 42608 316783
rect 59152 316771 59158 316783
rect 42602 316743 59158 316771
rect 42602 316731 42608 316743
rect 59152 316731 59158 316743
rect 59210 316731 59216 316783
rect 48208 313845 48214 313897
rect 48266 313885 48272 313897
rect 59632 313885 59638 313897
rect 48266 313857 59638 313885
rect 48266 313845 48272 313857
rect 59632 313845 59638 313857
rect 59690 313845 59696 313897
rect 48016 313771 48022 313823
rect 48074 313811 48080 313823
rect 58864 313811 58870 313823
rect 48074 313783 58870 313811
rect 48074 313771 48080 313783
rect 58864 313771 58870 313783
rect 58922 313771 58928 313823
rect 48112 313697 48118 313749
rect 48170 313737 48176 313749
rect 59632 313737 59638 313749
rect 48170 313709 59638 313737
rect 48170 313697 48176 313709
rect 59632 313697 59638 313709
rect 59690 313697 59696 313749
rect 654256 311181 654262 311233
rect 654314 311221 654320 311233
rect 676240 311221 676246 311233
rect 654314 311193 676246 311221
rect 654314 311181 654320 311193
rect 676240 311181 676246 311193
rect 676298 311181 676304 311233
rect 654160 311107 654166 311159
rect 654218 311147 654224 311159
rect 676144 311147 676150 311159
rect 654218 311119 676150 311147
rect 654218 311107 654224 311119
rect 676144 311107 676150 311119
rect 676202 311107 676208 311159
rect 654064 311033 654070 311085
rect 654122 311073 654128 311085
rect 676336 311073 676342 311085
rect 654122 311045 676342 311073
rect 654122 311033 654128 311045
rect 676336 311033 676342 311045
rect 676394 311033 676400 311085
rect 42160 308073 42166 308125
rect 42218 308113 42224 308125
rect 59152 308113 59158 308125
rect 42218 308085 59158 308113
rect 42218 308073 42224 308085
rect 59152 308073 59158 308085
rect 59210 308073 59216 308125
rect 674128 305261 674134 305313
rect 674186 305301 674192 305313
rect 676240 305301 676246 305313
rect 674186 305273 676246 305301
rect 674186 305261 674192 305273
rect 676240 305261 676246 305273
rect 676298 305261 676304 305313
rect 673936 302523 673942 302575
rect 673994 302563 674000 302575
rect 675952 302563 675958 302575
rect 673994 302535 675958 302563
rect 673994 302523 674000 302535
rect 675952 302523 675958 302535
rect 676010 302523 676016 302575
rect 674032 302449 674038 302501
rect 674090 302489 674096 302501
rect 676048 302489 676054 302501
rect 674090 302461 676054 302489
rect 674090 302449 674096 302461
rect 676048 302449 676054 302461
rect 676106 302449 676112 302501
rect 674224 302375 674230 302427
rect 674282 302415 674288 302427
rect 676240 302415 676246 302427
rect 674282 302387 676246 302415
rect 674282 302375 674288 302387
rect 676240 302375 676246 302387
rect 676298 302375 676304 302427
rect 43408 300895 43414 300947
rect 43466 300935 43472 300947
rect 63280 300935 63286 300947
rect 43466 300907 63286 300935
rect 43466 300895 43472 300907
rect 63280 300895 63286 300907
rect 63338 300895 63344 300947
rect 39760 299637 39766 299689
rect 39818 299677 39824 299689
rect 43408 299677 43414 299689
rect 39818 299649 43414 299677
rect 39818 299637 39824 299649
rect 43408 299637 43414 299649
rect 43466 299637 43472 299689
rect 41776 299563 41782 299615
rect 41834 299603 41840 299615
rect 43120 299603 43126 299615
rect 41834 299575 43126 299603
rect 41834 299563 41840 299575
rect 43120 299563 43126 299575
rect 43178 299563 43184 299615
rect 650320 299563 650326 299615
rect 650378 299603 650384 299615
rect 679984 299603 679990 299615
rect 650378 299575 679990 299603
rect 650378 299563 650384 299575
rect 679984 299563 679990 299575
rect 680042 299563 680048 299615
rect 41776 299119 41782 299171
rect 41834 299159 41840 299171
rect 51472 299159 51478 299171
rect 41834 299131 51478 299159
rect 41834 299119 41840 299131
rect 51472 299119 51478 299131
rect 51530 299119 51536 299171
rect 41776 298157 41782 298209
rect 41834 298197 41840 298209
rect 43504 298197 43510 298209
rect 41834 298169 43510 298197
rect 41834 298157 41840 298169
rect 43504 298157 43510 298169
rect 43562 298157 43568 298209
rect 43216 298083 43222 298135
rect 43274 298123 43280 298135
rect 61648 298123 61654 298135
rect 43274 298095 61654 298123
rect 43274 298083 43280 298095
rect 61648 298083 61654 298095
rect 61706 298083 61712 298135
rect 41776 297565 41782 297617
rect 41834 297605 41840 297617
rect 43408 297605 43414 297617
rect 41834 297577 43414 297605
rect 41834 297565 41840 297577
rect 43408 297565 43414 297577
rect 43466 297565 43472 297617
rect 41776 297047 41782 297099
rect 41834 297087 41840 297099
rect 43312 297087 43318 297099
rect 41834 297059 43318 297087
rect 41834 297047 41840 297059
rect 43312 297047 43318 297059
rect 43370 297047 43376 297099
rect 39952 296677 39958 296729
rect 40010 296717 40016 296729
rect 43216 296717 43222 296729
rect 40010 296689 43222 296717
rect 40010 296677 40016 296689
rect 43216 296677 43222 296689
rect 43274 296677 43280 296729
rect 674128 295937 674134 295989
rect 674186 295977 674192 295989
rect 675280 295977 675286 295989
rect 674186 295949 675286 295977
rect 674186 295937 674192 295949
rect 675280 295937 675286 295949
rect 675338 295937 675344 295989
rect 41584 295863 41590 295915
rect 41642 295903 41648 295915
rect 43216 295903 43222 295915
rect 41642 295875 43222 295903
rect 41642 295863 41648 295875
rect 43216 295863 43222 295875
rect 43274 295863 43280 295915
rect 674224 295715 674230 295767
rect 674282 295755 674288 295767
rect 675184 295755 675190 295767
rect 674282 295727 675190 295755
rect 674282 295715 674288 295727
rect 675184 295715 675190 295727
rect 675242 295715 675248 295767
rect 674032 294235 674038 294287
rect 674090 294275 674096 294287
rect 675184 294275 675190 294287
rect 674090 294247 675190 294275
rect 674090 294235 674096 294247
rect 675184 294235 675190 294247
rect 675242 294235 675248 294287
rect 39664 293717 39670 293769
rect 39722 293757 39728 293769
rect 58192 293757 58198 293769
rect 39722 293729 58198 293757
rect 39722 293717 39728 293729
rect 58192 293717 58198 293729
rect 58250 293717 58256 293769
rect 673936 291719 673942 291771
rect 673994 291759 674000 291771
rect 675184 291759 675190 291771
rect 673994 291731 675190 291759
rect 673994 291719 674000 291731
rect 675184 291719 675190 291731
rect 675242 291719 675248 291771
rect 43120 291571 43126 291623
rect 43178 291611 43184 291623
rect 59632 291611 59638 291623
rect 43178 291583 59638 291611
rect 43178 291571 43184 291583
rect 59632 291571 59638 291583
rect 59690 291571 59696 291623
rect 41584 291423 41590 291475
rect 41642 291463 41648 291475
rect 43120 291463 43126 291475
rect 41642 291435 43126 291463
rect 41642 291423 41648 291435
rect 43120 291423 43126 291435
rect 43178 291423 43184 291475
rect 41584 290905 41590 290957
rect 41642 290945 41648 290957
rect 42928 290945 42934 290957
rect 41642 290917 42934 290945
rect 41642 290905 41648 290917
rect 42928 290905 42934 290917
rect 42986 290905 42992 290957
rect 53296 290905 53302 290957
rect 53354 290945 53360 290957
rect 59440 290945 59446 290957
rect 53354 290917 59446 290945
rect 53354 290905 53360 290917
rect 59440 290905 59446 290917
rect 59498 290905 59504 290957
rect 656560 290831 656566 290883
rect 656618 290871 656624 290883
rect 675088 290871 675094 290883
rect 656618 290843 675094 290871
rect 656618 290831 656624 290843
rect 675088 290831 675094 290843
rect 675146 290831 675152 290883
rect 51472 288315 51478 288367
rect 51530 288355 51536 288367
rect 58864 288355 58870 288367
rect 51530 288327 58870 288355
rect 51530 288315 51536 288327
rect 58864 288315 58870 288327
rect 58922 288315 58928 288367
rect 48016 288019 48022 288071
rect 48074 288059 48080 288071
rect 59152 288059 59158 288071
rect 48074 288031 59158 288059
rect 48074 288019 48080 288031
rect 59152 288019 59158 288031
rect 59210 288019 59216 288071
rect 40240 287945 40246 287997
rect 40298 287985 40304 287997
rect 42640 287985 42646 287997
rect 40298 287957 42646 287985
rect 40298 287945 40304 287957
rect 42640 287945 42646 287957
rect 42698 287945 42704 287997
rect 41488 287871 41494 287923
rect 41546 287911 41552 287923
rect 42736 287911 42742 287923
rect 41546 287883 42742 287911
rect 41546 287871 41552 287883
rect 42736 287871 42742 287883
rect 42794 287871 42800 287923
rect 41872 287131 41878 287183
rect 41930 287171 41936 287183
rect 45520 287171 45526 287183
rect 41930 287143 45526 287171
rect 41930 287131 41936 287143
rect 45520 287131 45526 287143
rect 45578 287131 45584 287183
rect 41584 285207 41590 285259
rect 41642 285247 41648 285259
rect 42448 285247 42454 285259
rect 41642 285219 42454 285247
rect 41642 285207 41648 285219
rect 42448 285207 42454 285219
rect 42506 285207 42512 285259
rect 53200 285133 53206 285185
rect 53258 285173 53264 285185
rect 59248 285173 59254 285185
rect 53258 285145 59254 285173
rect 53258 285133 53264 285145
rect 59248 285133 59254 285145
rect 59306 285133 59312 285185
rect 653776 284245 653782 284297
rect 653834 284285 653840 284297
rect 658000 284285 658006 284297
rect 653834 284257 658006 284285
rect 653834 284245 653840 284257
rect 658000 284245 658006 284257
rect 658058 284245 658064 284297
rect 41776 283801 41782 283853
rect 41834 283801 41840 283853
rect 41794 283557 41822 283801
rect 41776 283505 41782 283557
rect 41834 283505 41840 283557
rect 50320 282321 50326 282373
rect 50378 282361 50384 282373
rect 58864 282361 58870 282373
rect 50378 282333 58870 282361
rect 50378 282321 50384 282333
rect 58864 282321 58870 282333
rect 58922 282321 58928 282373
rect 56176 282247 56182 282299
rect 56234 282287 56240 282299
rect 57616 282287 57622 282299
rect 56234 282259 57622 282287
rect 56234 282247 56240 282259
rect 57616 282247 57622 282259
rect 57674 282247 57680 282299
rect 42160 281729 42166 281781
rect 42218 281769 42224 281781
rect 42640 281769 42646 281781
rect 42218 281741 42646 281769
rect 42218 281729 42224 281741
rect 42640 281729 42646 281741
rect 42698 281729 42704 281781
rect 42064 280101 42070 280153
rect 42122 280141 42128 280153
rect 42832 280141 42838 280153
rect 42122 280113 42838 280141
rect 42122 280101 42128 280113
rect 42832 280101 42838 280113
rect 42890 280101 42896 280153
rect 42160 279879 42166 279931
rect 42218 279919 42224 279931
rect 42352 279919 42358 279931
rect 42218 279891 42358 279919
rect 42218 279879 42224 279891
rect 42352 279879 42358 279891
rect 42410 279879 42416 279931
rect 45328 279435 45334 279487
rect 45386 279475 45392 279487
rect 59536 279475 59542 279487
rect 45386 279447 59542 279475
rect 45386 279435 45392 279447
rect 59536 279435 59542 279447
rect 59594 279435 59600 279487
rect 654160 279435 654166 279487
rect 654218 279475 654224 279487
rect 663760 279475 663766 279487
rect 654218 279447 663766 279475
rect 654218 279435 654224 279447
rect 663760 279435 663766 279447
rect 663818 279435 663824 279487
rect 45424 279361 45430 279413
rect 45482 279401 45488 279413
rect 59248 279401 59254 279413
rect 45482 279373 59254 279401
rect 45482 279361 45488 279373
rect 59248 279361 59254 279373
rect 59306 279361 59312 279413
rect 42160 278473 42166 278525
rect 42218 278513 42224 278525
rect 43024 278513 43030 278525
rect 42218 278485 43030 278513
rect 42218 278473 42224 278485
rect 43024 278473 43030 278485
rect 43082 278473 43088 278525
rect 314896 278251 314902 278303
rect 314954 278291 314960 278303
rect 408304 278291 408310 278303
rect 314954 278263 408310 278291
rect 314954 278251 314960 278263
rect 408304 278251 408310 278263
rect 408362 278251 408368 278303
rect 316624 278177 316630 278229
rect 316682 278217 316688 278229
rect 411856 278217 411862 278229
rect 316682 278189 411862 278217
rect 316682 278177 316688 278189
rect 411856 278177 411862 278189
rect 411914 278177 411920 278229
rect 319504 278103 319510 278155
rect 319562 278143 319568 278155
rect 418960 278143 418966 278155
rect 319562 278115 418966 278143
rect 319562 278103 319568 278115
rect 418960 278103 418966 278115
rect 419018 278103 419024 278155
rect 320944 278029 320950 278081
rect 321002 278069 321008 278081
rect 422512 278069 422518 278081
rect 321002 278041 422518 278069
rect 321002 278029 321008 278041
rect 422512 278029 422518 278041
rect 422570 278029 422576 278081
rect 392272 277955 392278 278007
rect 392330 277995 392336 278007
rect 599824 277995 599830 278007
rect 392330 277967 599830 277995
rect 392330 277955 392336 277967
rect 599824 277955 599830 277967
rect 599882 277955 599888 278007
rect 675088 277955 675094 278007
rect 675146 277995 675152 278007
rect 679792 277995 679798 278007
rect 675146 277967 679798 277995
rect 675146 277955 675152 277967
rect 679792 277955 679798 277967
rect 679850 277955 679856 278007
rect 323824 277881 323830 277933
rect 323882 277921 323888 277933
rect 429616 277921 429622 277933
rect 323882 277893 429622 277921
rect 323882 277881 323888 277893
rect 429616 277881 429622 277893
rect 429674 277881 429680 277933
rect 42160 277807 42166 277859
rect 42218 277847 42224 277859
rect 42544 277847 42550 277859
rect 42218 277819 42550 277847
rect 42218 277807 42224 277819
rect 42544 277807 42550 277819
rect 42602 277807 42608 277859
rect 322096 277807 322102 277859
rect 322154 277847 322160 277859
rect 426352 277847 426358 277859
rect 322154 277819 426358 277847
rect 322154 277807 322160 277819
rect 426352 277807 426358 277819
rect 426410 277807 426416 277859
rect 317872 277733 317878 277785
rect 317930 277773 317936 277785
rect 415696 277773 415702 277785
rect 317930 277745 415702 277773
rect 317930 277733 317936 277745
rect 415696 277733 415702 277745
rect 415754 277733 415760 277785
rect 329296 277659 329302 277711
rect 329354 277699 329360 277711
rect 444112 277699 444118 277711
rect 329354 277671 444118 277699
rect 329354 277659 329360 277671
rect 444112 277659 444118 277671
rect 444170 277659 444176 277711
rect 332368 277585 332374 277637
rect 332426 277625 332432 277637
rect 451216 277625 451222 277637
rect 332426 277597 451222 277625
rect 332426 277585 332432 277597
rect 451216 277585 451222 277597
rect 451274 277585 451280 277637
rect 334960 277511 334966 277563
rect 335018 277551 335024 277563
rect 458224 277551 458230 277563
rect 335018 277523 458230 277551
rect 335018 277511 335024 277523
rect 458224 277511 458230 277523
rect 458282 277511 458288 277563
rect 337840 277437 337846 277489
rect 337898 277477 337904 277489
rect 465328 277477 465334 277489
rect 337898 277449 465334 277477
rect 337898 277437 337904 277449
rect 465328 277437 465334 277449
rect 465386 277437 465392 277489
rect 341008 277363 341014 277415
rect 341066 277403 341072 277415
rect 472432 277403 472438 277415
rect 341066 277375 472438 277403
rect 341066 277363 341072 277375
rect 472432 277363 472438 277375
rect 472490 277363 472496 277415
rect 343888 277289 343894 277341
rect 343946 277329 343952 277341
rect 479536 277329 479542 277341
rect 343946 277301 479542 277329
rect 343946 277289 343952 277301
rect 479536 277289 479542 277301
rect 479594 277289 479600 277341
rect 373840 277215 373846 277267
rect 373898 277255 373904 277267
rect 554032 277255 554038 277267
rect 373898 277227 554038 277255
rect 373898 277215 373904 277227
rect 554032 277215 554038 277227
rect 554090 277215 554096 277267
rect 375088 277141 375094 277193
rect 375146 277181 375152 277193
rect 557584 277181 557590 277193
rect 375146 277153 557590 277181
rect 375146 277141 375152 277153
rect 557584 277141 557590 277153
rect 557642 277141 557648 277193
rect 376816 277067 376822 277119
rect 376874 277107 376880 277119
rect 561136 277107 561142 277119
rect 376874 277079 561142 277107
rect 376874 277067 376880 277079
rect 561136 277067 561142 277079
rect 561194 277067 561200 277119
rect 377968 276993 377974 277045
rect 378026 277033 378032 277045
rect 564688 277033 564694 277045
rect 378026 277005 564694 277033
rect 378026 276993 378032 277005
rect 564688 276993 564694 277005
rect 564746 276993 564752 277045
rect 379408 276919 379414 276971
rect 379466 276959 379472 276971
rect 568240 276959 568246 276971
rect 379466 276931 568246 276959
rect 379466 276919 379472 276931
rect 568240 276919 568246 276931
rect 568298 276919 568304 276971
rect 381040 276845 381046 276897
rect 381098 276885 381104 276897
rect 571696 276885 571702 276897
rect 381098 276857 571702 276885
rect 381098 276845 381104 276857
rect 571696 276845 571702 276857
rect 571754 276845 571760 276897
rect 42352 276771 42358 276823
rect 42410 276811 42416 276823
rect 43120 276811 43126 276823
rect 42410 276783 43126 276811
rect 42410 276771 42416 276783
rect 43120 276771 43126 276783
rect 43178 276771 43184 276823
rect 382288 276771 382294 276823
rect 382346 276811 382352 276823
rect 575248 276811 575254 276823
rect 382346 276783 575254 276811
rect 382346 276771 382352 276783
rect 575248 276771 575254 276783
rect 575306 276771 575312 276823
rect 42544 276697 42550 276749
rect 42602 276737 42608 276749
rect 42928 276737 42934 276749
rect 42602 276709 42934 276737
rect 42602 276697 42608 276709
rect 42928 276697 42934 276709
rect 42986 276697 42992 276749
rect 383632 276697 383638 276749
rect 383690 276737 383696 276749
rect 578800 276737 578806 276749
rect 383690 276709 578806 276737
rect 383690 276697 383696 276709
rect 578800 276697 578806 276709
rect 578858 276697 578864 276749
rect 386512 276623 386518 276675
rect 386570 276663 386576 276675
rect 585904 276663 585910 276675
rect 386570 276635 585910 276663
rect 386570 276623 386576 276635
rect 585904 276623 585910 276635
rect 585962 276623 585968 276675
rect 385360 276549 385366 276601
rect 385418 276589 385424 276601
rect 582352 276589 582358 276601
rect 385418 276561 582358 276589
rect 385418 276549 385424 276561
rect 582352 276549 582358 276561
rect 582410 276549 582416 276601
rect 326416 276475 326422 276527
rect 326474 276515 326480 276527
rect 437008 276515 437014 276527
rect 326474 276487 437014 276515
rect 326474 276475 326480 276487
rect 437008 276475 437014 276487
rect 437066 276475 437072 276527
rect 42832 276401 42838 276453
rect 42890 276441 42896 276453
rect 59344 276441 59350 276453
rect 42890 276413 59350 276441
rect 42890 276401 42896 276413
rect 59344 276401 59350 276413
rect 59402 276401 59408 276453
rect 286096 276401 286102 276453
rect 286154 276441 286160 276453
rect 336496 276441 336502 276453
rect 286154 276413 336502 276441
rect 286154 276401 286160 276413
rect 336496 276401 336502 276413
rect 336554 276401 336560 276453
rect 359152 276401 359158 276453
rect 359210 276441 359216 276453
rect 517360 276441 517366 276453
rect 359210 276413 517366 276441
rect 359210 276401 359216 276413
rect 517360 276401 517366 276413
rect 517418 276401 517424 276453
rect 288688 276327 288694 276379
rect 288746 276367 288752 276379
rect 343600 276367 343606 276379
rect 288746 276339 343606 276367
rect 288746 276327 288752 276339
rect 343600 276327 343606 276339
rect 343658 276327 343664 276379
rect 361744 276327 361750 276379
rect 361802 276367 361808 276379
rect 524464 276367 524470 276379
rect 361802 276339 524470 276367
rect 361802 276327 361808 276339
rect 524464 276327 524470 276339
rect 524522 276327 524528 276379
rect 287344 276253 287350 276305
rect 287402 276293 287408 276305
rect 340048 276293 340054 276305
rect 287402 276265 340054 276293
rect 287402 276253 287408 276265
rect 340048 276253 340054 276265
rect 340106 276253 340112 276305
rect 364624 276253 364630 276305
rect 364682 276293 364688 276305
rect 531568 276293 531574 276305
rect 364682 276265 531574 276293
rect 364682 276253 364688 276265
rect 531568 276253 531574 276265
rect 531626 276253 531632 276305
rect 291856 276179 291862 276231
rect 291914 276219 291920 276231
rect 350704 276219 350710 276231
rect 291914 276191 350710 276219
rect 291914 276179 291920 276191
rect 350704 276179 350710 276191
rect 350762 276179 350768 276231
rect 367696 276179 367702 276231
rect 367754 276219 367760 276231
rect 538672 276219 538678 276231
rect 367754 276191 538678 276219
rect 367754 276179 367760 276191
rect 538672 276179 538678 276191
rect 538730 276179 538736 276231
rect 290320 276105 290326 276157
rect 290378 276145 290384 276157
rect 347152 276145 347158 276157
rect 290378 276117 347158 276145
rect 290378 276105 290384 276117
rect 347152 276105 347158 276117
rect 347210 276105 347216 276157
rect 370288 276105 370294 276157
rect 370346 276145 370352 276157
rect 545776 276145 545782 276157
rect 370346 276117 545782 276145
rect 370346 276105 370352 276117
rect 545776 276105 545782 276117
rect 545834 276105 545840 276157
rect 293008 276031 293014 276083
rect 293066 276071 293072 276083
rect 354256 276071 354262 276083
rect 293066 276043 354262 276071
rect 293066 276031 293072 276043
rect 354256 276031 354262 276043
rect 354314 276031 354320 276083
rect 371056 276031 371062 276083
rect 371114 276071 371120 276083
rect 546928 276071 546934 276083
rect 371114 276043 546934 276071
rect 371114 276031 371120 276043
rect 546928 276031 546934 276043
rect 546986 276031 546992 276083
rect 294640 275957 294646 276009
rect 294698 275997 294704 276009
rect 357808 275997 357814 276009
rect 294698 275969 357814 275997
rect 294698 275957 294704 275969
rect 357808 275957 357814 275969
rect 357866 275957 357872 276009
rect 371920 275957 371926 276009
rect 371978 275997 371984 276009
rect 549328 275997 549334 276009
rect 371978 275969 549334 275997
rect 371978 275957 371984 275969
rect 549328 275957 549334 275969
rect 549386 275957 549392 276009
rect 297328 275883 297334 275935
rect 297386 275923 297392 275935
rect 364912 275923 364918 275935
rect 297386 275895 364918 275923
rect 297386 275883 297392 275895
rect 364912 275883 364918 275895
rect 364970 275883 364976 275935
rect 373456 275883 373462 275935
rect 373514 275923 373520 275935
rect 552784 275923 552790 275935
rect 373514 275895 552790 275923
rect 373514 275883 373520 275895
rect 552784 275883 552790 275895
rect 552842 275883 552848 275935
rect 295888 275809 295894 275861
rect 295946 275849 295952 275861
rect 361360 275849 361366 275861
rect 295946 275821 361366 275849
rect 295946 275809 295952 275821
rect 361360 275809 361366 275821
rect 361418 275809 361424 275861
rect 374608 275809 374614 275861
rect 374666 275849 374672 275861
rect 556336 275849 556342 275861
rect 374666 275821 556342 275849
rect 374666 275809 374672 275821
rect 556336 275809 556342 275821
rect 556394 275809 556400 275861
rect 296464 275735 296470 275787
rect 296522 275775 296528 275787
rect 362512 275775 362518 275787
rect 296522 275747 362518 275775
rect 296522 275735 296528 275747
rect 362512 275735 362518 275747
rect 362570 275735 362576 275787
rect 377488 275735 377494 275787
rect 377546 275775 377552 275787
rect 563440 275775 563446 275787
rect 377546 275747 563446 275775
rect 377546 275735 377552 275747
rect 563440 275735 563446 275747
rect 563498 275735 563504 275787
rect 298960 275661 298966 275713
rect 299018 275701 299024 275713
rect 368464 275701 368470 275713
rect 299018 275673 368470 275701
rect 299018 275661 299024 275673
rect 368464 275661 368470 275673
rect 368522 275661 368528 275713
rect 376240 275661 376246 275713
rect 376298 275701 376304 275713
rect 559888 275701 559894 275713
rect 376298 275673 559894 275701
rect 376298 275661 376304 275673
rect 559888 275661 559894 275673
rect 559946 275661 559952 275713
rect 297808 275587 297814 275639
rect 297866 275627 297872 275639
rect 366064 275627 366070 275639
rect 297866 275599 366070 275627
rect 297866 275587 297872 275599
rect 366064 275587 366070 275599
rect 366122 275587 366128 275639
rect 380560 275587 380566 275639
rect 380618 275627 380624 275639
rect 570544 275627 570550 275639
rect 380618 275599 570550 275627
rect 380618 275587 380624 275599
rect 570544 275587 570550 275599
rect 570602 275587 570608 275639
rect 300208 275513 300214 275565
rect 300266 275553 300272 275565
rect 372016 275553 372022 275565
rect 300266 275525 372022 275553
rect 300266 275513 300272 275525
rect 372016 275513 372022 275525
rect 372074 275513 372080 275565
rect 381808 275513 381814 275565
rect 381866 275553 381872 275565
rect 574096 275553 574102 275565
rect 381866 275525 574102 275553
rect 381866 275513 381872 275525
rect 574096 275513 574102 275525
rect 574154 275513 574160 275565
rect 299152 275439 299158 275491
rect 299210 275479 299216 275491
rect 369616 275479 369622 275491
rect 299210 275451 369622 275479
rect 299210 275439 299216 275451
rect 369616 275439 369622 275451
rect 369674 275439 369680 275491
rect 388912 275439 388918 275491
rect 388970 275479 388976 275491
rect 591856 275479 591862 275491
rect 388970 275451 591862 275479
rect 388970 275439 388976 275451
rect 591856 275439 591862 275451
rect 591914 275439 591920 275491
rect 303280 275365 303286 275417
rect 303338 275405 303344 275417
rect 379120 275405 379126 275417
rect 303338 275377 379126 275405
rect 303338 275365 303344 275377
rect 379120 275365 379126 275377
rect 379178 275365 379184 275417
rect 389584 275365 389590 275417
rect 389642 275405 389648 275417
rect 593008 275405 593014 275417
rect 389642 275377 593014 275405
rect 389642 275365 389648 275377
rect 593008 275365 593014 275377
rect 593066 275365 593072 275417
rect 304432 275291 304438 275343
rect 304490 275331 304496 275343
rect 382576 275331 382582 275343
rect 304490 275303 382582 275331
rect 304490 275291 304496 275303
rect 382576 275291 382582 275303
rect 382634 275291 382640 275343
rect 391984 275291 391990 275343
rect 392042 275331 392048 275343
rect 598960 275331 598966 275343
rect 392042 275303 598966 275331
rect 392042 275291 392048 275303
rect 598960 275291 598966 275303
rect 599018 275291 599024 275343
rect 307312 275217 307318 275269
rect 307370 275257 307376 275269
rect 389680 275257 389686 275269
rect 307370 275229 389686 275257
rect 307370 275217 307376 275229
rect 389680 275217 389686 275229
rect 389738 275217 389744 275269
rect 396304 275217 396310 275269
rect 396362 275257 396368 275269
rect 609520 275257 609526 275269
rect 396362 275229 609526 275257
rect 396362 275217 396368 275229
rect 609520 275217 609526 275229
rect 609578 275217 609584 275269
rect 310384 275143 310390 275195
rect 310442 275183 310448 275195
rect 396784 275183 396790 275195
rect 310442 275155 396790 275183
rect 310442 275143 310448 275155
rect 396784 275143 396790 275155
rect 396842 275143 396848 275195
rect 404944 275143 404950 275195
rect 405002 275183 405008 275195
rect 405002 275155 407678 275183
rect 405002 275143 405008 275155
rect 314704 275069 314710 275121
rect 314762 275109 314768 275121
rect 407440 275109 407446 275121
rect 314762 275081 407446 275109
rect 314762 275069 314768 275081
rect 407440 275069 407446 275081
rect 407498 275069 407504 275121
rect 311632 274995 311638 275047
rect 311690 275035 311696 275047
rect 400336 275035 400342 275047
rect 311690 275007 400342 275035
rect 311690 274995 311696 275007
rect 400336 274995 400342 275007
rect 400394 274995 400400 275047
rect 407650 275035 407678 275155
rect 407728 275143 407734 275195
rect 407786 275183 407792 275195
rect 623728 275183 623734 275195
rect 407786 275155 623734 275183
rect 407786 275143 407792 275155
rect 623728 275143 623734 275155
rect 623786 275143 623792 275195
rect 408400 275069 408406 275121
rect 408458 275109 408464 275121
rect 635536 275109 635542 275121
rect 408458 275081 635542 275109
rect 408458 275069 408464 275081
rect 635536 275069 635542 275081
rect 635594 275069 635600 275121
rect 630832 275035 630838 275047
rect 407650 275007 630838 275035
rect 630832 274995 630838 275007
rect 630890 274995 630896 275047
rect 284464 274921 284470 274973
rect 284522 274961 284528 274973
rect 332944 274961 332950 274973
rect 284522 274933 332950 274961
rect 284522 274921 284528 274933
rect 332944 274921 332950 274933
rect 333002 274921 333008 274973
rect 356176 274921 356182 274973
rect 356234 274961 356240 274973
rect 510256 274961 510262 274973
rect 356234 274933 510262 274961
rect 356234 274921 356240 274933
rect 510256 274921 510262 274933
rect 510314 274921 510320 274973
rect 283024 274847 283030 274899
rect 283082 274887 283088 274899
rect 329392 274887 329398 274899
rect 283082 274859 329398 274887
rect 283082 274847 283088 274859
rect 329392 274847 329398 274859
rect 329450 274847 329456 274899
rect 344560 274847 344566 274899
rect 344618 274887 344624 274899
rect 481936 274887 481942 274899
rect 344618 274859 481942 274887
rect 344618 274847 344624 274859
rect 481936 274847 481942 274859
rect 481994 274847 482000 274899
rect 281776 274773 281782 274825
rect 281834 274813 281840 274825
rect 325840 274813 325846 274825
rect 281834 274785 325846 274813
rect 281834 274773 281840 274785
rect 325840 274773 325846 274785
rect 325898 274773 325904 274825
rect 339088 274773 339094 274825
rect 339146 274813 339152 274825
rect 467728 274813 467734 274825
rect 339146 274785 467734 274813
rect 339146 274773 339152 274785
rect 467728 274773 467734 274785
rect 467786 274773 467792 274825
rect 336016 274699 336022 274751
rect 336074 274739 336080 274751
rect 460624 274739 460630 274751
rect 336074 274711 460630 274739
rect 336074 274699 336080 274711
rect 460624 274699 460630 274711
rect 460682 274699 460688 274751
rect 333136 274625 333142 274677
rect 333194 274665 333200 274677
rect 453520 274665 453526 274677
rect 333194 274637 453526 274665
rect 333194 274625 333200 274637
rect 453520 274625 453526 274637
rect 453578 274625 453584 274677
rect 330448 274551 330454 274603
rect 330506 274591 330512 274603
rect 446416 274591 446422 274603
rect 330506 274563 446422 274591
rect 330506 274551 330512 274563
rect 446416 274551 446422 274563
rect 446474 274551 446480 274603
rect 328816 274477 328822 274529
rect 328874 274517 328880 274529
rect 442864 274517 442870 274529
rect 328874 274489 442870 274517
rect 328874 274477 328880 274489
rect 442864 274477 442870 274489
rect 442922 274477 442928 274529
rect 325936 274403 325942 274455
rect 325994 274443 326000 274455
rect 435856 274443 435862 274455
rect 325994 274415 435862 274443
rect 325994 274403 326000 274415
rect 435856 274403 435862 274415
rect 435914 274403 435920 274455
rect 323344 274329 323350 274381
rect 323402 274369 323408 274381
rect 428752 274369 428758 274381
rect 323402 274341 428758 274369
rect 323402 274329 323408 274341
rect 428752 274329 428758 274341
rect 428810 274329 428816 274381
rect 320176 274255 320182 274307
rect 320234 274295 320240 274307
rect 421648 274295 421654 274307
rect 320234 274267 421654 274295
rect 320234 274255 320240 274267
rect 421648 274255 421654 274267
rect 421706 274255 421712 274307
rect 315952 274181 315958 274233
rect 316010 274221 316016 274233
rect 410992 274221 410998 274233
rect 316010 274193 410998 274221
rect 316010 274181 316016 274193
rect 410992 274181 410998 274193
rect 411050 274181 411056 274233
rect 317296 274107 317302 274159
rect 317354 274147 317360 274159
rect 414544 274147 414550 274159
rect 317354 274119 414550 274147
rect 317354 274107 317360 274119
rect 414544 274107 414550 274119
rect 414602 274107 414608 274159
rect 348496 274033 348502 274085
rect 348554 274073 348560 274085
rect 401488 274073 401494 274085
rect 348554 274045 401494 274073
rect 348554 274033 348560 274045
rect 401488 274033 401494 274045
rect 401546 274033 401552 274085
rect 401776 274033 401782 274085
rect 401834 274073 401840 274085
rect 407728 274073 407734 274085
rect 401834 274045 407734 274073
rect 401834 274033 401840 274045
rect 407728 274033 407734 274045
rect 407786 274033 407792 274085
rect 326800 273959 326806 274011
rect 326858 273999 326864 274011
rect 373168 273999 373174 274011
rect 326858 273971 373174 273999
rect 326858 273959 326864 273971
rect 373168 273959 373174 273971
rect 373226 273959 373232 274011
rect 342160 273885 342166 273937
rect 342218 273925 342224 273937
rect 387376 273925 387382 273937
rect 342218 273897 387382 273925
rect 342218 273885 342224 273897
rect 387376 273885 387382 273897
rect 387434 273885 387440 273937
rect 334288 273811 334294 273863
rect 334346 273851 334352 273863
rect 380272 273851 380278 273863
rect 334346 273823 380278 273851
rect 334346 273811 334352 273823
rect 380272 273811 380278 273823
rect 380330 273811 380336 273863
rect 347056 273737 347062 273789
rect 347114 273777 347120 273789
rect 394480 273777 394486 273789
rect 347114 273749 394486 273777
rect 347114 273737 347120 273749
rect 394480 273737 394486 273749
rect 394538 273737 394544 273789
rect 331216 273663 331222 273715
rect 331274 273703 331280 273715
rect 376720 273703 376726 273715
rect 331274 273675 376726 273703
rect 331274 273663 331280 273675
rect 376720 273663 376726 273675
rect 376778 273663 376784 273715
rect 43024 273515 43030 273567
rect 43082 273555 43088 273567
rect 59152 273555 59158 273567
rect 43082 273527 59158 273555
rect 43082 273515 43088 273527
rect 59152 273515 59158 273527
rect 59210 273515 59216 273567
rect 160432 273515 160438 273567
rect 160490 273555 160496 273567
rect 207472 273555 207478 273567
rect 160490 273527 207478 273555
rect 160490 273515 160496 273527
rect 207472 273515 207478 273527
rect 207530 273515 207536 273567
rect 228976 273515 228982 273567
rect 229034 273555 229040 273567
rect 242416 273555 242422 273567
rect 229034 273527 242422 273555
rect 229034 273515 229040 273527
rect 242416 273515 242422 273527
rect 242474 273515 242480 273567
rect 271024 273515 271030 273567
rect 271082 273555 271088 273567
rect 299920 273555 299926 273567
rect 271082 273527 299926 273555
rect 271082 273515 271088 273527
rect 299920 273515 299926 273527
rect 299978 273515 299984 273567
rect 308368 273515 308374 273567
rect 308426 273555 308432 273567
rect 344752 273555 344758 273567
rect 308426 273527 344758 273555
rect 308426 273515 308432 273527
rect 344752 273515 344758 273527
rect 344810 273515 344816 273567
rect 350032 273515 350038 273567
rect 350090 273555 350096 273567
rect 494896 273555 494902 273567
rect 350090 273527 494902 273555
rect 350090 273515 350096 273527
rect 494896 273515 494902 273527
rect 494954 273515 494960 273567
rect 521296 273515 521302 273567
rect 521354 273555 521360 273567
rect 631984 273555 631990 273567
rect 521354 273527 631990 273555
rect 521354 273515 521360 273527
rect 631984 273515 631990 273527
rect 632042 273515 632048 273567
rect 130864 273441 130870 273493
rect 130922 273481 130928 273493
rect 190096 273481 190102 273493
rect 130922 273453 190102 273481
rect 130922 273441 130928 273453
rect 190096 273441 190102 273453
rect 190154 273441 190160 273493
rect 193552 273441 193558 273493
rect 193610 273481 193616 273493
rect 221488 273481 221494 273493
rect 193610 273453 221494 273481
rect 193610 273441 193616 273453
rect 221488 273441 221494 273453
rect 221546 273441 221552 273493
rect 277072 273441 277078 273493
rect 277130 273481 277136 273493
rect 314032 273481 314038 273493
rect 277130 273453 314038 273481
rect 277130 273441 277136 273453
rect 314032 273441 314038 273453
rect 314090 273441 314096 273493
rect 349456 273441 349462 273493
rect 349514 273481 349520 273493
rect 493744 273481 493750 273493
rect 349514 273453 493750 273481
rect 349514 273441 349520 273453
rect 493744 273441 493750 273453
rect 493802 273441 493808 273493
rect 529840 273441 529846 273493
rect 529898 273481 529904 273493
rect 624976 273481 624982 273493
rect 529898 273453 624982 273481
rect 529898 273441 529904 273453
rect 624976 273441 624982 273453
rect 625034 273441 625040 273493
rect 108400 273367 108406 273419
rect 108458 273407 108464 273419
rect 109360 273407 109366 273419
rect 108458 273379 109366 273407
rect 108458 273367 108464 273379
rect 109360 273367 109366 273379
rect 109418 273367 109424 273419
rect 122608 273367 122614 273419
rect 122666 273407 122672 273419
rect 123760 273407 123766 273419
rect 122666 273379 123766 273407
rect 122666 273367 122672 273379
rect 123760 273367 123766 273379
rect 123818 273367 123824 273419
rect 142672 273367 142678 273419
rect 142730 273407 142736 273419
rect 209584 273407 209590 273419
rect 142730 273379 209590 273407
rect 142730 273367 142736 273379
rect 209584 273367 209590 273379
rect 209642 273367 209648 273419
rect 277744 273367 277750 273419
rect 277802 273407 277808 273419
rect 316432 273407 316438 273419
rect 277802 273379 316438 273407
rect 277802 273367 277808 273379
rect 316432 273367 316438 273379
rect 316490 273367 316496 273419
rect 352432 273367 352438 273419
rect 352490 273407 352496 273419
rect 500848 273407 500854 273419
rect 352490 273379 500854 273407
rect 352490 273367 352496 273379
rect 500848 273367 500854 273379
rect 500906 273367 500912 273419
rect 135568 273293 135574 273345
rect 135626 273333 135632 273345
rect 209776 273333 209782 273345
rect 135626 273305 209782 273333
rect 135626 273293 135632 273305
rect 209776 273293 209782 273305
rect 209834 273293 209840 273345
rect 279664 273293 279670 273345
rect 279722 273333 279728 273345
rect 321136 273333 321142 273345
rect 279722 273305 321142 273333
rect 279722 273293 279728 273305
rect 321136 273293 321142 273305
rect 321194 273293 321200 273345
rect 352624 273293 352630 273345
rect 352682 273333 352688 273345
rect 502000 273333 502006 273345
rect 352682 273305 502006 273333
rect 352682 273293 352688 273305
rect 502000 273293 502006 273305
rect 502058 273293 502064 273345
rect 68272 273219 68278 273271
rect 68330 273259 68336 273271
rect 142480 273259 142486 273271
rect 68330 273231 142486 273259
rect 68330 273219 68336 273231
rect 142480 273219 142486 273231
rect 142538 273219 142544 273271
rect 153328 273219 153334 273271
rect 153386 273259 153392 273271
rect 207376 273259 207382 273271
rect 153386 273231 207382 273259
rect 153386 273219 153392 273231
rect 207376 273219 207382 273231
rect 207434 273219 207440 273271
rect 219568 273219 219574 273271
rect 219626 273259 219632 273271
rect 238672 273259 238678 273271
rect 219626 273231 238678 273259
rect 219626 273219 219632 273231
rect 238672 273219 238678 273231
rect 238730 273219 238736 273271
rect 278224 273219 278230 273271
rect 278282 273259 278288 273271
rect 317584 273259 317590 273271
rect 278282 273231 317590 273259
rect 278282 273219 278288 273231
rect 317584 273219 317590 273231
rect 317642 273219 317648 273271
rect 355504 273219 355510 273271
rect 355562 273259 355568 273271
rect 509104 273259 509110 273271
rect 355562 273231 509110 273259
rect 355562 273219 355568 273231
rect 509104 273219 509110 273231
rect 509162 273219 509168 273271
rect 509200 273219 509206 273271
rect 509258 273259 509264 273271
rect 548080 273259 548086 273271
rect 509258 273231 548086 273259
rect 509258 273219 509264 273231
rect 548080 273219 548086 273231
rect 548138 273219 548144 273271
rect 132016 273145 132022 273197
rect 132074 273185 132080 273197
rect 209872 273185 209878 273197
rect 132074 273157 209878 273185
rect 132074 273145 132080 273157
rect 209872 273145 209878 273157
rect 209930 273145 209936 273197
rect 220720 273145 220726 273197
rect 220778 273185 220784 273197
rect 239152 273185 239158 273197
rect 220778 273157 239158 273185
rect 220778 273145 220784 273157
rect 239152 273145 239158 273157
rect 239210 273145 239216 273197
rect 285616 273145 285622 273197
rect 285674 273185 285680 273197
rect 335344 273185 335350 273197
rect 285674 273157 335350 273185
rect 285674 273145 285680 273157
rect 335344 273145 335350 273157
rect 335402 273145 335408 273197
rect 355024 273145 355030 273197
rect 355082 273185 355088 273197
rect 507952 273185 507958 273197
rect 355082 273157 507958 273185
rect 355082 273145 355088 273157
rect 507952 273145 507958 273157
rect 508010 273145 508016 273197
rect 508240 273145 508246 273197
rect 508298 273185 508304 273197
rect 639088 273185 639094 273197
rect 508298 273157 639094 273185
rect 508298 273145 508304 273157
rect 639088 273145 639094 273157
rect 639146 273145 639152 273197
rect 127312 273071 127318 273123
rect 127370 273111 127376 273123
rect 209968 273111 209974 273123
rect 127370 273083 209974 273111
rect 127370 273071 127376 273083
rect 209968 273071 209974 273083
rect 210026 273071 210032 273123
rect 218320 273071 218326 273123
rect 218378 273111 218384 273123
rect 238096 273111 238102 273123
rect 218378 273083 238102 273111
rect 218378 273071 218384 273083
rect 238096 273071 238102 273083
rect 238154 273071 238160 273123
rect 286768 273071 286774 273123
rect 286826 273111 286832 273123
rect 338896 273111 338902 273123
rect 286826 273083 338902 273111
rect 286826 273071 286832 273083
rect 338896 273071 338902 273083
rect 338954 273071 338960 273123
rect 358576 273071 358582 273123
rect 358634 273111 358640 273123
rect 358634 273083 374942 273111
rect 358634 273071 358640 273083
rect 125008 272997 125014 273049
rect 125066 273037 125072 273049
rect 207280 273037 207286 273049
rect 125066 273009 207286 273037
rect 125066 272997 125072 273009
rect 207280 272997 207286 273009
rect 207338 272997 207344 273049
rect 217168 272997 217174 273049
rect 217226 273037 217232 273049
rect 237616 273037 237622 273049
rect 217226 273009 237622 273037
rect 217226 272997 217232 273009
rect 237616 272997 237622 273009
rect 237674 272997 237680 273049
rect 284944 272997 284950 273049
rect 285002 273037 285008 273049
rect 334192 273037 334198 273049
rect 285002 273009 334198 273037
rect 285002 272997 285008 273009
rect 334192 272997 334198 273009
rect 334250 272997 334256 273049
rect 360976 272997 360982 273049
rect 361034 273037 361040 273049
rect 374800 273037 374806 273049
rect 361034 273009 374806 273037
rect 361034 272997 361040 273009
rect 374800 272997 374806 273009
rect 374858 272997 374864 273049
rect 374914 273037 374942 273083
rect 374992 273071 374998 273123
rect 375050 273111 375056 273123
rect 514960 273111 514966 273123
rect 375050 273083 514966 273111
rect 375050 273071 375056 273083
rect 514960 273071 514966 273083
rect 515018 273071 515024 273123
rect 516208 273037 516214 273049
rect 374914 273009 516214 273037
rect 516208 272997 516214 273009
rect 516266 272997 516272 273049
rect 516304 272997 516310 273049
rect 516362 273037 516368 273049
rect 580048 273037 580054 273049
rect 516362 273009 580054 273037
rect 516362 272997 516368 273009
rect 580048 272997 580054 273009
rect 580106 272997 580112 273049
rect 128464 272923 128470 272975
rect 128522 272963 128528 272975
rect 210160 272963 210166 272975
rect 128522 272935 210166 272963
rect 128522 272923 128528 272935
rect 210160 272923 210166 272935
rect 210218 272923 210224 272975
rect 216016 272923 216022 272975
rect 216074 272963 216080 272975
rect 236944 272963 236950 272975
rect 216074 272935 236950 272963
rect 216074 272923 216080 272935
rect 236944 272923 236950 272935
rect 237002 272923 237008 272975
rect 274192 272923 274198 272975
rect 274250 272963 274256 272975
rect 306928 272963 306934 272975
rect 274250 272935 306934 272963
rect 274250 272923 274256 272935
rect 306928 272923 306934 272935
rect 306986 272923 306992 272975
rect 307024 272923 307030 272975
rect 307082 272963 307088 272975
rect 358960 272963 358966 272975
rect 307082 272935 358966 272963
rect 307082 272923 307088 272935
rect 358960 272923 358966 272935
rect 359018 272923 359024 272975
rect 361264 272923 361270 272975
rect 361322 272963 361328 272975
rect 523312 272963 523318 272975
rect 361322 272935 523318 272963
rect 361322 272923 361328 272935
rect 523312 272923 523318 272935
rect 523370 272923 523376 272975
rect 123664 272849 123670 272901
rect 123722 272889 123728 272901
rect 209008 272889 209014 272901
rect 123722 272861 209014 272889
rect 123722 272849 123728 272861
rect 209008 272849 209014 272861
rect 209066 272849 209072 272901
rect 236464 272889 236470 272901
rect 215986 272861 236470 272889
rect 116656 272775 116662 272827
rect 116714 272815 116720 272827
rect 207088 272815 207094 272827
rect 116714 272787 207094 272815
rect 116714 272775 116720 272787
rect 207088 272775 207094 272787
rect 207146 272775 207152 272827
rect 214768 272775 214774 272827
rect 214826 272815 214832 272827
rect 215986 272815 216014 272861
rect 236464 272849 236470 272861
rect 236522 272849 236528 272901
rect 289936 272849 289942 272901
rect 289994 272889 290000 272901
rect 346000 272889 346006 272901
rect 289994 272861 346006 272889
rect 289994 272849 290000 272861
rect 346000 272849 346006 272861
rect 346058 272849 346064 272901
rect 363568 272849 363574 272901
rect 363626 272889 363632 272901
rect 363626 272861 374750 272889
rect 363626 272849 363632 272861
rect 236272 272815 236278 272827
rect 214826 272787 216014 272815
rect 226210 272787 236278 272815
rect 214826 272775 214832 272787
rect 120208 272701 120214 272753
rect 120266 272741 120272 272753
rect 207856 272741 207862 272753
rect 120266 272713 207862 272741
rect 120266 272701 120272 272713
rect 207856 272701 207862 272713
rect 207914 272701 207920 272753
rect 212464 272701 212470 272753
rect 212522 272741 212528 272753
rect 225904 272741 225910 272753
rect 212522 272713 225910 272741
rect 212522 272701 212528 272713
rect 225904 272701 225910 272713
rect 225962 272701 225968 272753
rect 113104 272627 113110 272679
rect 113162 272667 113168 272679
rect 206032 272667 206038 272679
rect 113162 272639 206038 272667
rect 113162 272627 113168 272639
rect 206032 272627 206038 272639
rect 206090 272627 206096 272679
rect 213616 272627 213622 272679
rect 213674 272667 213680 272679
rect 226210 272667 226238 272787
rect 236272 272775 236278 272787
rect 236330 272775 236336 272827
rect 292240 272775 292246 272827
rect 292298 272815 292304 272827
rect 351856 272815 351862 272827
rect 292298 272787 351862 272815
rect 292298 272775 292304 272787
rect 351856 272775 351862 272787
rect 351914 272775 351920 272827
rect 364144 272775 364150 272827
rect 364202 272815 364208 272827
rect 374722 272815 374750 272861
rect 374800 272849 374806 272901
rect 374858 272889 374864 272901
rect 522064 272889 522070 272901
rect 374858 272861 522070 272889
rect 374858 272849 374864 272861
rect 522064 272849 522070 272861
rect 522122 272849 522128 272901
rect 523024 272849 523030 272901
rect 523082 272889 523088 272901
rect 583600 272889 583606 272901
rect 523082 272861 583606 272889
rect 523082 272849 523088 272861
rect 583600 272849 583606 272861
rect 583658 272849 583664 272901
rect 529168 272815 529174 272827
rect 364202 272787 374654 272815
rect 374722 272787 529174 272815
rect 364202 272775 364208 272787
rect 233680 272701 233686 272753
rect 233738 272741 233744 272753
rect 244048 272741 244054 272753
rect 233738 272713 244054 272741
rect 233738 272701 233744 272713
rect 244048 272701 244054 272713
rect 244106 272701 244112 272753
rect 292720 272701 292726 272753
rect 292778 272741 292784 272753
rect 353104 272741 353110 272753
rect 292778 272713 353110 272741
rect 292778 272701 292784 272713
rect 353104 272701 353110 272713
rect 353162 272701 353168 272753
rect 366544 272701 366550 272753
rect 366602 272741 366608 272753
rect 374512 272741 374518 272753
rect 366602 272713 374518 272741
rect 366602 272701 366608 272713
rect 374512 272701 374518 272713
rect 374570 272701 374576 272753
rect 374626 272741 374654 272787
rect 529168 272775 529174 272787
rect 529226 272775 529232 272827
rect 530416 272741 530422 272753
rect 374626 272713 530422 272741
rect 530416 272701 530422 272713
rect 530474 272701 530480 272753
rect 213674 272639 226238 272667
rect 213674 272627 213680 272639
rect 295408 272627 295414 272679
rect 295466 272667 295472 272679
rect 360208 272667 360214 272679
rect 295466 272639 360214 272667
rect 295466 272627 295472 272639
rect 360208 272627 360214 272639
rect 360266 272627 360272 272679
rect 367120 272627 367126 272679
rect 367178 272667 367184 272679
rect 537424 272667 537430 272679
rect 367178 272639 537430 272667
rect 367178 272627 367184 272639
rect 537424 272627 537430 272639
rect 537482 272627 537488 272679
rect 96592 272553 96598 272605
rect 96650 272593 96656 272605
rect 106672 272593 106678 272605
rect 96650 272565 106678 272593
rect 96650 272553 96656 272565
rect 106672 272553 106678 272565
rect 106730 272553 106736 272605
rect 110800 272553 110806 272605
rect 110858 272593 110864 272605
rect 205744 272593 205750 272605
rect 110858 272565 205750 272593
rect 110858 272553 110864 272565
rect 205744 272553 205750 272565
rect 205802 272553 205808 272605
rect 211216 272553 211222 272605
rect 211274 272593 211280 272605
rect 235024 272593 235030 272605
rect 211274 272565 235030 272593
rect 211274 272553 211280 272565
rect 235024 272553 235030 272565
rect 235082 272553 235088 272605
rect 270256 272553 270262 272605
rect 270314 272593 270320 272605
rect 297520 272593 297526 272605
rect 270314 272565 297526 272593
rect 270314 272553 270320 272565
rect 297520 272553 297526 272565
rect 297578 272553 297584 272605
rect 298288 272553 298294 272605
rect 298346 272593 298352 272605
rect 367216 272593 367222 272605
rect 298346 272565 367222 272593
rect 298346 272553 298352 272565
rect 367216 272553 367222 272565
rect 367274 272553 367280 272605
rect 372688 272553 372694 272605
rect 372746 272593 372752 272605
rect 372746 272565 374462 272593
rect 372746 272553 372752 272565
rect 106096 272479 106102 272531
rect 106154 272519 106160 272531
rect 204016 272519 204022 272531
rect 106154 272491 204022 272519
rect 106154 272479 106160 272491
rect 204016 272479 204022 272491
rect 204074 272479 204080 272531
rect 210064 272479 210070 272531
rect 210122 272519 210128 272531
rect 234544 272519 234550 272531
rect 210122 272491 234550 272519
rect 210122 272479 210128 272491
rect 234544 272479 234550 272491
rect 234602 272479 234608 272531
rect 270544 272479 270550 272531
rect 270602 272519 270608 272531
rect 298672 272519 298678 272531
rect 270602 272491 298678 272519
rect 270602 272479 270608 272491
rect 298672 272479 298678 272491
rect 298730 272479 298736 272531
rect 301360 272479 301366 272531
rect 301418 272519 301424 272531
rect 374320 272519 374326 272531
rect 301418 272491 374326 272519
rect 301418 272479 301424 272491
rect 374320 272479 374326 272491
rect 374378 272479 374384 272531
rect 374434 272519 374462 272565
rect 374512 272553 374518 272605
rect 374570 272593 374576 272605
rect 536272 272593 536278 272605
rect 374570 272565 536278 272593
rect 374570 272553 374576 272565
rect 536272 272553 536278 272565
rect 536330 272553 536336 272605
rect 551632 272519 551638 272531
rect 374434 272491 551638 272519
rect 551632 272479 551638 272491
rect 551690 272479 551696 272531
rect 103696 272405 103702 272457
rect 103754 272445 103760 272457
rect 203536 272445 203542 272457
rect 103754 272417 203542 272445
rect 103754 272405 103760 272417
rect 203536 272405 203542 272417
rect 203594 272405 203600 272457
rect 208912 272405 208918 272457
rect 208970 272445 208976 272457
rect 234352 272445 234358 272457
rect 208970 272417 234358 272445
rect 208970 272405 208976 272417
rect 234352 272405 234358 272417
rect 234410 272405 234416 272457
rect 234928 272405 234934 272457
rect 234986 272445 234992 272457
rect 244816 272445 244822 272457
rect 234986 272417 244822 272445
rect 234986 272405 234992 272417
rect 244816 272405 244822 272417
rect 244874 272405 244880 272457
rect 272752 272405 272758 272457
rect 272810 272445 272816 272457
rect 303472 272445 303478 272457
rect 272810 272417 303478 272445
rect 272810 272405 272816 272417
rect 303472 272405 303478 272417
rect 303530 272405 303536 272457
rect 303952 272405 303958 272457
rect 304010 272445 304016 272457
rect 381424 272445 381430 272457
rect 304010 272417 381430 272445
rect 304010 272405 304016 272417
rect 381424 272405 381430 272417
rect 381482 272405 381488 272457
rect 381520 272405 381526 272457
rect 381578 272445 381584 272457
rect 572944 272445 572950 272457
rect 381578 272417 572950 272445
rect 381578 272405 381584 272417
rect 572944 272405 572950 272417
rect 573002 272405 573008 272457
rect 98992 272331 98998 272383
rect 99050 272371 99056 272383
rect 199120 272371 199126 272383
rect 99050 272343 199126 272371
rect 99050 272331 99056 272343
rect 199120 272331 199126 272343
rect 199178 272331 199184 272383
rect 232528 272331 232534 272383
rect 232586 272371 232592 272383
rect 243664 272371 243670 272383
rect 232586 272343 243670 272371
rect 232586 272331 232592 272343
rect 243664 272331 243670 272343
rect 243722 272331 243728 272383
rect 273424 272331 273430 272383
rect 273482 272371 273488 272383
rect 305776 272371 305782 272383
rect 273482 272343 305782 272371
rect 273482 272331 273488 272343
rect 305776 272331 305782 272343
rect 305834 272331 305840 272383
rect 306832 272331 306838 272383
rect 306890 272371 306896 272383
rect 388528 272371 388534 272383
rect 306890 272343 388534 272371
rect 306890 272331 306896 272343
rect 388528 272331 388534 272343
rect 388586 272331 388592 272383
rect 407440 272331 407446 272383
rect 407498 272371 407504 272383
rect 587152 272371 587158 272383
rect 407498 272343 587158 272371
rect 407498 272331 407504 272343
rect 587152 272331 587158 272343
rect 587210 272331 587216 272383
rect 76528 272257 76534 272309
rect 76586 272297 76592 272309
rect 76586 272269 106622 272297
rect 76586 272257 76592 272269
rect 84784 272183 84790 272235
rect 84842 272223 84848 272235
rect 86320 272223 86326 272235
rect 84842 272195 86326 272223
rect 84842 272183 84848 272195
rect 86320 272183 86326 272195
rect 86378 272183 86384 272235
rect 104848 272183 104854 272235
rect 104906 272223 104912 272235
rect 106480 272223 106486 272235
rect 104906 272195 106486 272223
rect 104906 272183 104912 272195
rect 106480 272183 106486 272195
rect 106538 272183 106544 272235
rect 106594 272223 106622 272269
rect 106672 272257 106678 272309
rect 106730 272297 106736 272309
rect 201616 272297 201622 272309
rect 106730 272269 201622 272297
rect 106730 272257 106736 272269
rect 201616 272257 201622 272269
rect 201674 272257 201680 272309
rect 207664 272257 207670 272309
rect 207722 272297 207728 272309
rect 233872 272297 233878 272309
rect 207722 272269 233878 272297
rect 207722 272257 207728 272269
rect 233872 272257 233878 272269
rect 233930 272257 233936 272309
rect 236080 272257 236086 272309
rect 236138 272297 236144 272309
rect 245296 272297 245302 272309
rect 236138 272269 245302 272297
rect 236138 272257 236144 272269
rect 245296 272257 245302 272269
rect 245354 272257 245360 272309
rect 275344 272257 275350 272309
rect 275402 272297 275408 272309
rect 310480 272297 310486 272309
rect 275402 272269 310486 272297
rect 275402 272257 275408 272269
rect 310480 272257 310486 272269
rect 310538 272257 310544 272309
rect 395632 272297 395638 272309
rect 310594 272269 395638 272297
rect 195664 272223 195670 272235
rect 106594 272195 195670 272223
rect 195664 272183 195670 272195
rect 195722 272183 195728 272235
rect 198256 272183 198262 272235
rect 198314 272223 198320 272235
rect 224368 272223 224374 272235
rect 198314 272195 224374 272223
rect 198314 272183 198320 272195
rect 224368 272183 224374 272195
rect 224426 272183 224432 272235
rect 225904 272183 225910 272235
rect 225962 272223 225968 272235
rect 235696 272223 235702 272235
rect 225962 272195 235702 272223
rect 225962 272183 225968 272195
rect 235696 272183 235702 272195
rect 235754 272183 235760 272235
rect 275152 272183 275158 272235
rect 275210 272223 275216 272235
rect 309328 272223 309334 272235
rect 275210 272195 309334 272223
rect 275210 272183 275216 272195
rect 309328 272183 309334 272195
rect 309386 272183 309392 272235
rect 309904 272183 309910 272235
rect 309962 272223 309968 272235
rect 310594 272223 310622 272269
rect 395632 272257 395638 272269
rect 395690 272257 395696 272309
rect 395920 272257 395926 272309
rect 395978 272297 395984 272309
rect 608368 272297 608374 272309
rect 395978 272269 608374 272297
rect 395978 272257 395984 272269
rect 608368 272257 608374 272269
rect 608426 272257 608432 272309
rect 309962 272195 310622 272223
rect 309962 272183 309968 272195
rect 312784 272183 312790 272235
rect 312842 272223 312848 272235
rect 402736 272223 402742 272235
rect 312842 272195 402742 272223
rect 312842 272183 312848 272195
rect 402736 272183 402742 272195
rect 402794 272183 402800 272235
rect 402928 272183 402934 272235
rect 402986 272223 402992 272235
rect 622576 272223 622582 272235
rect 402986 272195 622582 272223
rect 402986 272183 402992 272195
rect 622576 272183 622582 272195
rect 622634 272183 622640 272235
rect 194704 272109 194710 272161
rect 194762 272149 194768 272161
rect 224464 272149 224470 272161
rect 194762 272121 224470 272149
rect 194762 272109 194768 272121
rect 224464 272109 224470 272121
rect 224522 272109 224528 272161
rect 227824 272109 227830 272161
rect 227882 272149 227888 272161
rect 242128 272149 242134 272161
rect 227882 272121 242134 272149
rect 227882 272109 227888 272121
rect 242128 272109 242134 272121
rect 242186 272109 242192 272161
rect 276304 272109 276310 272161
rect 276362 272149 276368 272161
rect 312880 272149 312886 272161
rect 276362 272121 312886 272149
rect 276362 272109 276368 272121
rect 312880 272109 312886 272121
rect 312938 272109 312944 272161
rect 315472 272109 315478 272161
rect 315530 272149 315536 272161
rect 409840 272149 409846 272161
rect 315530 272121 409846 272149
rect 315530 272109 315536 272121
rect 409840 272109 409846 272121
rect 409898 272109 409904 272161
rect 413680 272109 413686 272161
rect 413738 272149 413744 272161
rect 643888 272149 643894 272161
rect 413738 272121 643894 272149
rect 413738 272109 413744 272121
rect 643888 272109 643894 272121
rect 643946 272109 643952 272161
rect 119056 272035 119062 272087
rect 119114 272075 119120 272087
rect 120880 272075 120886 272087
rect 119114 272047 120886 272075
rect 119114 272035 119120 272047
rect 120880 272035 120886 272047
rect 120938 272035 120944 272087
rect 165136 272035 165142 272087
rect 165194 272075 165200 272087
rect 166960 272075 166966 272087
rect 165194 272047 166966 272075
rect 165194 272035 165200 272047
rect 166960 272035 166966 272047
rect 167018 272035 167024 272087
rect 167536 272035 167542 272087
rect 167594 272075 167600 272087
rect 210640 272075 210646 272087
rect 167594 272047 210646 272075
rect 167594 272035 167600 272047
rect 210640 272035 210646 272047
rect 210698 272035 210704 272087
rect 230128 272035 230134 272087
rect 230186 272075 230192 272087
rect 242896 272075 242902 272087
rect 230186 272047 242902 272075
rect 230186 272035 230192 272047
rect 242896 272035 242902 272047
rect 242954 272035 242960 272087
rect 299440 272035 299446 272087
rect 299498 272075 299504 272087
rect 299498 272047 302078 272075
rect 299498 272035 299504 272047
rect 174640 271961 174646 272013
rect 174698 272001 174704 272013
rect 210544 272001 210550 272013
rect 174698 271973 210550 272001
rect 174698 271961 174704 271973
rect 210544 271961 210550 271973
rect 210602 271961 210608 272013
rect 231376 271961 231382 272013
rect 231434 272001 231440 272013
rect 243088 272001 243094 272013
rect 231434 271973 243094 272001
rect 231434 271961 231440 271973
rect 243088 271961 243094 271973
rect 243146 271961 243152 272013
rect 301936 272001 301942 272013
rect 296626 271973 301942 272001
rect 159280 271887 159286 271939
rect 159338 271927 159344 271939
rect 192976 271927 192982 271939
rect 159338 271899 192982 271927
rect 159338 271887 159344 271899
rect 192976 271887 192982 271899
rect 193034 271887 193040 271939
rect 195856 271887 195862 271939
rect 195914 271927 195920 271939
rect 221680 271927 221686 271939
rect 195914 271899 221686 271927
rect 195914 271887 195920 271899
rect 221680 271887 221686 271899
rect 221738 271887 221744 271939
rect 272272 271887 272278 271939
rect 272330 271927 272336 271939
rect 296626 271927 296654 271973
rect 301936 271961 301942 271973
rect 301994 271961 302000 272013
rect 302050 272001 302078 272047
rect 306640 272035 306646 272087
rect 306698 272075 306704 272087
rect 328240 272075 328246 272087
rect 306698 272047 328246 272075
rect 306698 272035 306704 272047
rect 328240 272035 328246 272047
rect 328298 272035 328304 272087
rect 346960 272035 346966 272087
rect 347018 272075 347024 272087
rect 487792 272075 487798 272087
rect 347018 272047 487798 272075
rect 347018 272035 347024 272047
rect 487792 272035 487798 272047
rect 487850 272035 487856 272087
rect 327088 272001 327094 272013
rect 302050 271973 327094 272001
rect 327088 271961 327094 271973
rect 327146 271961 327152 272013
rect 346480 271961 346486 272013
rect 346538 272001 346544 272013
rect 486640 272001 486646 272013
rect 346538 271973 486646 272001
rect 346538 271961 346544 271973
rect 486640 271961 486646 271973
rect 486698 271961 486704 272013
rect 272330 271899 296654 271927
rect 272330 271887 272336 271899
rect 301072 271887 301078 271939
rect 301130 271927 301136 271939
rect 324688 271927 324694 271939
rect 301130 271899 324694 271927
rect 301130 271887 301136 271899
rect 324688 271887 324694 271899
rect 324746 271887 324752 271939
rect 344080 271887 344086 271939
rect 344138 271927 344144 271939
rect 480688 271927 480694 271939
rect 344138 271899 480694 271927
rect 344138 271887 344144 271899
rect 480688 271887 480694 271899
rect 480746 271887 480752 271939
rect 191152 271813 191158 271865
rect 191210 271853 191216 271865
rect 227152 271853 227158 271865
rect 191210 271825 227158 271853
rect 191210 271813 191216 271825
rect 227152 271813 227158 271825
rect 227210 271813 227216 271865
rect 299344 271813 299350 271865
rect 299402 271853 299408 271865
rect 306640 271853 306646 271865
rect 299402 271825 306646 271853
rect 299402 271813 299408 271825
rect 306640 271813 306646 271825
rect 306698 271813 306704 271865
rect 341488 271813 341494 271865
rect 341546 271853 341552 271865
rect 473680 271853 473686 271865
rect 341546 271825 473686 271853
rect 341546 271813 341552 271825
rect 473680 271813 473686 271825
rect 473738 271813 473744 271865
rect 147376 271739 147382 271791
rect 147434 271779 147440 271791
rect 149680 271779 149686 271791
rect 147434 271751 149686 271779
rect 147434 271739 147440 271751
rect 149680 271739 149686 271751
rect 149738 271739 149744 271791
rect 192304 271739 192310 271791
rect 192362 271779 192368 271791
rect 224560 271779 224566 271791
rect 192362 271751 224566 271779
rect 192362 271739 192368 271751
rect 224560 271739 224566 271751
rect 224618 271739 224624 271791
rect 338608 271739 338614 271791
rect 338666 271779 338672 271791
rect 466576 271779 466582 271791
rect 338666 271751 466582 271779
rect 338666 271739 338672 271751
rect 466576 271739 466582 271751
rect 466634 271739 466640 271791
rect 166288 271665 166294 271717
rect 166346 271705 166352 271717
rect 198640 271705 198646 271717
rect 166346 271677 198646 271705
rect 166346 271665 166352 271677
rect 198640 271665 198646 271677
rect 198698 271665 198704 271717
rect 199408 271665 199414 271717
rect 199466 271705 199472 271717
rect 221584 271705 221590 271717
rect 199466 271677 221590 271705
rect 199466 271665 199472 271677
rect 221584 271665 221590 271677
rect 221642 271665 221648 271717
rect 335440 271665 335446 271717
rect 335498 271705 335504 271717
rect 459472 271705 459478 271717
rect 335498 271677 459478 271705
rect 335498 271665 335504 271677
rect 459472 271665 459478 271677
rect 459530 271665 459536 271717
rect 75280 271591 75286 271643
rect 75338 271631 75344 271643
rect 77680 271631 77686 271643
rect 75338 271603 77686 271631
rect 75338 271591 75344 271603
rect 77680 271591 77686 271603
rect 77738 271591 77744 271643
rect 129712 271591 129718 271643
rect 129770 271631 129776 271643
rect 132400 271631 132406 271643
rect 129770 271603 132406 271631
rect 129770 271591 129776 271603
rect 132400 271591 132406 271603
rect 132458 271591 132464 271643
rect 181744 271591 181750 271643
rect 181802 271631 181808 271643
rect 210448 271631 210454 271643
rect 181802 271603 210454 271631
rect 181802 271591 181808 271603
rect 210448 271591 210454 271603
rect 210506 271591 210512 271643
rect 332560 271591 332566 271643
rect 332618 271631 332624 271643
rect 452368 271631 452374 271643
rect 332618 271603 452374 271631
rect 332618 271591 332624 271603
rect 452368 271591 452374 271603
rect 452426 271591 452432 271643
rect 89488 271517 89494 271569
rect 89546 271557 89552 271569
rect 92080 271557 92086 271569
rect 89546 271529 92086 271557
rect 89546 271517 89552 271529
rect 92080 271517 92086 271529
rect 92138 271517 92144 271569
rect 150928 271517 150934 271569
rect 150986 271557 150992 271569
rect 152368 271557 152374 271569
rect 150986 271529 152374 271557
rect 150986 271517 150992 271529
rect 152368 271517 152374 271529
rect 152426 271517 152432 271569
rect 180496 271517 180502 271569
rect 180554 271557 180560 271569
rect 205168 271557 205174 271569
rect 180554 271529 205174 271557
rect 180554 271517 180560 271529
rect 205168 271517 205174 271529
rect 205226 271517 205232 271569
rect 329968 271517 329974 271569
rect 330026 271557 330032 271569
rect 445264 271557 445270 271569
rect 330026 271529 445270 271557
rect 330026 271517 330032 271529
rect 445264 271517 445270 271529
rect 445322 271517 445328 271569
rect 185200 271443 185206 271495
rect 185258 271483 185264 271495
rect 210352 271483 210358 271495
rect 185258 271455 210358 271483
rect 185258 271443 185264 271455
rect 210352 271443 210358 271455
rect 210410 271443 210416 271495
rect 326896 271443 326902 271495
rect 326954 271483 326960 271495
rect 438160 271483 438166 271495
rect 326954 271455 438166 271483
rect 326954 271443 326960 271455
rect 438160 271443 438166 271455
rect 438218 271443 438224 271495
rect 173392 271369 173398 271421
rect 173450 271409 173456 271421
rect 200464 271409 200470 271421
rect 173450 271381 200470 271409
rect 173450 271369 173456 271381
rect 200464 271369 200470 271381
rect 200522 271369 200528 271421
rect 201808 271369 201814 271421
rect 201866 271409 201872 271421
rect 223696 271409 223702 271421
rect 201866 271381 223702 271409
rect 201866 271369 201872 271381
rect 223696 271369 223702 271381
rect 223754 271369 223760 271421
rect 324016 271369 324022 271421
rect 324074 271409 324080 271421
rect 431056 271409 431062 271421
rect 324074 271381 431062 271409
rect 324074 271369 324080 271381
rect 431056 271369 431062 271381
rect 431114 271369 431120 271421
rect 184048 271295 184054 271347
rect 184106 271335 184112 271347
rect 205936 271335 205942 271347
rect 184106 271307 205942 271335
rect 184106 271295 184112 271307
rect 205936 271295 205942 271307
rect 205994 271295 206000 271347
rect 321424 271295 321430 271347
rect 321482 271335 321488 271347
rect 423952 271335 423958 271347
rect 321482 271307 423958 271335
rect 321482 271295 321488 271307
rect 423952 271295 423958 271307
rect 424010 271295 424016 271347
rect 161584 271221 161590 271273
rect 161642 271261 161648 271273
rect 163888 271261 163894 271273
rect 161642 271233 163894 271261
rect 161642 271221 161648 271233
rect 163888 271221 163894 271233
rect 163946 271221 163952 271273
rect 188752 271221 188758 271273
rect 188810 271261 188816 271273
rect 210256 271261 210262 271273
rect 188810 271233 210262 271261
rect 188810 271221 188816 271233
rect 210256 271221 210262 271233
rect 210314 271221 210320 271273
rect 237232 271221 237238 271273
rect 237290 271261 237296 271273
rect 245584 271261 245590 271273
rect 237290 271233 245590 271261
rect 237290 271221 237296 271233
rect 245584 271221 245590 271233
rect 245642 271221 245648 271273
rect 318352 271221 318358 271273
rect 318410 271261 318416 271273
rect 416944 271261 416950 271273
rect 318410 271233 416950 271261
rect 318410 271221 318416 271233
rect 416944 271221 416950 271233
rect 417002 271221 417008 271273
rect 175792 271147 175798 271199
rect 175850 271187 175856 271199
rect 178288 271187 178294 271199
rect 175850 271159 178294 271187
rect 175850 271147 175856 271159
rect 178288 271147 178294 271159
rect 178346 271147 178352 271199
rect 187600 271147 187606 271199
rect 187658 271187 187664 271199
rect 205840 271187 205846 271199
rect 187658 271159 205846 271187
rect 187658 271147 187664 271159
rect 205840 271147 205846 271159
rect 205898 271147 205904 271199
rect 238480 271147 238486 271199
rect 238538 271187 238544 271199
rect 246064 271187 246070 271199
rect 238538 271159 246070 271187
rect 238538 271147 238544 271159
rect 246064 271147 246070 271159
rect 246122 271147 246128 271199
rect 357904 271147 357910 271199
rect 357962 271187 357968 271199
rect 374992 271187 374998 271199
rect 357962 271159 374998 271187
rect 357962 271147 357968 271159
rect 374992 271147 374998 271159
rect 375050 271147 375056 271199
rect 387280 271147 387286 271199
rect 387338 271187 387344 271199
rect 407440 271187 407446 271199
rect 387338 271159 407446 271187
rect 387338 271147 387344 271159
rect 407440 271147 407446 271159
rect 407498 271147 407504 271199
rect 85936 271073 85942 271125
rect 85994 271113 86000 271125
rect 198544 271113 198550 271125
rect 85994 271085 198550 271113
rect 85994 271073 86000 271085
rect 198544 271073 198550 271085
rect 198602 271073 198608 271125
rect 205360 271073 205366 271125
rect 205418 271113 205424 271125
rect 232624 271113 232630 271125
rect 205418 271085 232630 271113
rect 205418 271073 205424 271085
rect 232624 271073 232630 271085
rect 232682 271073 232688 271125
rect 240784 271073 240790 271125
rect 240842 271113 240848 271125
rect 247216 271113 247222 271125
rect 240842 271085 247222 271113
rect 240842 271073 240848 271085
rect 247216 271073 247222 271085
rect 247274 271073 247280 271125
rect 221872 270999 221878 271051
rect 221930 271039 221936 271051
rect 239344 271039 239350 271051
rect 221930 271011 239350 271039
rect 221930 270999 221936 271011
rect 239344 270999 239350 271011
rect 239402 270999 239408 271051
rect 239536 270999 239542 271051
rect 239594 271039 239600 271051
rect 241264 271039 241270 271051
rect 239594 271011 241270 271039
rect 239594 270999 239600 271011
rect 241264 270999 241270 271011
rect 241322 270999 241328 271051
rect 241936 270999 241942 271051
rect 241994 271039 242000 271051
rect 247696 271039 247702 271051
rect 241994 271011 247702 271039
rect 241994 270999 242000 271011
rect 247696 270999 247702 271011
rect 247754 270999 247760 271051
rect 223024 270925 223030 270977
rect 223082 270965 223088 270977
rect 240016 270965 240022 270977
rect 223082 270937 240022 270965
rect 223082 270925 223088 270937
rect 240016 270925 240022 270937
rect 240074 270925 240080 270977
rect 243184 270925 243190 270977
rect 243242 270965 243248 270977
rect 247984 270965 247990 270977
rect 243242 270937 247990 270965
rect 243242 270925 243248 270937
rect 247984 270925 247990 270937
rect 248042 270925 248048 270977
rect 342736 270925 342742 270977
rect 342794 270965 342800 270977
rect 348304 270965 348310 270977
rect 342794 270937 348310 270965
rect 342794 270925 342800 270937
rect 348304 270925 348310 270937
rect 348362 270925 348368 270977
rect 224272 270851 224278 270903
rect 224330 270891 224336 270903
rect 240496 270891 240502 270903
rect 224330 270863 240502 270891
rect 224330 270851 224336 270863
rect 240496 270851 240502 270863
rect 240554 270851 240560 270903
rect 244336 270851 244342 270903
rect 244394 270891 244400 270903
rect 248656 270891 248662 270903
rect 244394 270863 248662 270891
rect 244394 270851 244400 270863
rect 248656 270851 248662 270863
rect 248714 270851 248720 270903
rect 334096 270851 334102 270903
rect 334154 270891 334160 270903
rect 337744 270891 337750 270903
rect 334154 270863 337750 270891
rect 334154 270851 334160 270863
rect 337744 270851 337750 270863
rect 337802 270851 337808 270903
rect 225424 270777 225430 270829
rect 225482 270817 225488 270829
rect 241072 270817 241078 270829
rect 225482 270789 241078 270817
rect 225482 270777 225488 270789
rect 241072 270777 241078 270789
rect 241130 270777 241136 270829
rect 245488 270777 245494 270829
rect 245546 270817 245552 270829
rect 249136 270817 249142 270829
rect 245546 270789 249142 270817
rect 245546 270777 245552 270789
rect 249136 270777 249142 270789
rect 249194 270777 249200 270829
rect 351376 270777 351382 270829
rect 351434 270817 351440 270829
rect 355408 270817 355414 270829
rect 351434 270789 355414 270817
rect 351434 270777 351440 270789
rect 355408 270777 355414 270789
rect 355466 270777 355472 270829
rect 94192 270703 94198 270755
rect 94250 270743 94256 270755
rect 94960 270743 94966 270755
rect 94250 270715 94966 270743
rect 94250 270703 94256 270715
rect 94960 270703 94966 270715
rect 95018 270703 95024 270755
rect 101296 270703 101302 270755
rect 101354 270743 101360 270755
rect 103600 270743 103606 270755
rect 101354 270715 103606 270743
rect 101354 270703 101360 270715
rect 103600 270703 103606 270715
rect 103658 270703 103664 270755
rect 115504 270703 115510 270755
rect 115562 270743 115568 270755
rect 118000 270743 118006 270755
rect 115562 270715 118006 270743
rect 115562 270703 115568 270715
rect 118000 270703 118006 270715
rect 118058 270703 118064 270755
rect 133264 270703 133270 270755
rect 133322 270743 133328 270755
rect 135280 270743 135286 270755
rect 133322 270715 135286 270743
rect 133322 270703 133328 270715
rect 135280 270703 135286 270715
rect 135338 270703 135344 270755
rect 136816 270703 136822 270755
rect 136874 270743 136880 270755
rect 138160 270743 138166 270755
rect 136874 270715 138166 270743
rect 136874 270703 136880 270715
rect 138160 270703 138166 270715
rect 138218 270703 138224 270755
rect 154480 270703 154486 270755
rect 154538 270743 154544 270755
rect 155440 270743 155446 270755
rect 154538 270715 155446 270743
rect 154538 270703 154544 270715
rect 155440 270703 155446 270715
rect 155498 270703 155504 270755
rect 168688 270703 168694 270755
rect 168746 270743 168752 270755
rect 169840 270743 169846 270755
rect 168746 270715 169846 270743
rect 168746 270703 168752 270715
rect 169840 270703 169846 270715
rect 169898 270703 169904 270755
rect 179344 270703 179350 270755
rect 179402 270743 179408 270755
rect 181360 270743 181366 270755
rect 179402 270715 181366 270743
rect 179402 270703 179408 270715
rect 181360 270703 181366 270715
rect 181418 270703 181424 270755
rect 182896 270703 182902 270755
rect 182954 270743 182960 270755
rect 184240 270743 184246 270755
rect 182954 270715 184246 270743
rect 182954 270703 182960 270715
rect 184240 270703 184246 270715
rect 184298 270703 184304 270755
rect 185488 270703 185494 270755
rect 185546 270743 185552 270755
rect 186448 270743 186454 270755
rect 185546 270715 186454 270743
rect 185546 270703 185552 270715
rect 186448 270703 186454 270715
rect 186506 270703 186512 270755
rect 226576 270703 226582 270755
rect 226634 270743 226640 270755
rect 239536 270743 239542 270755
rect 226634 270715 239542 270743
rect 226634 270703 226640 270715
rect 239536 270703 239542 270715
rect 239594 270703 239600 270755
rect 239632 270703 239638 270755
rect 239690 270743 239696 270755
rect 246448 270743 246454 270755
rect 239690 270715 246454 270743
rect 239690 270703 239696 270715
rect 246448 270703 246454 270715
rect 246506 270703 246512 270755
rect 246736 270703 246742 270755
rect 246794 270743 246800 270755
rect 249616 270743 249622 270755
rect 246794 270715 249622 270743
rect 246794 270703 246800 270715
rect 249616 270703 249622 270715
rect 249674 270703 249680 270755
rect 337936 270703 337942 270755
rect 337994 270743 338000 270755
rect 341296 270743 341302 270755
rect 337994 270715 341302 270743
rect 337994 270703 338000 270715
rect 341296 270703 341302 270715
rect 341354 270703 341360 270755
rect 408976 270703 408982 270755
rect 409034 270743 409040 270755
rect 413392 270743 413398 270755
rect 409034 270715 413398 270743
rect 409034 270703 409040 270715
rect 413392 270703 413398 270715
rect 413450 270703 413456 270755
rect 146224 270629 146230 270681
rect 146282 270669 146288 270681
rect 214960 270669 214966 270681
rect 146282 270641 214966 270669
rect 146282 270629 146288 270641
rect 214960 270629 214966 270641
rect 215018 270629 215024 270681
rect 269680 270629 269686 270681
rect 269738 270669 269744 270681
rect 296368 270669 296374 270681
rect 269738 270641 296374 270669
rect 269738 270629 269744 270641
rect 296368 270629 296374 270641
rect 296426 270629 296432 270681
rect 356656 270669 356662 270681
rect 296482 270641 356662 270669
rect 141520 270555 141526 270607
rect 141578 270595 141584 270607
rect 213808 270595 213814 270607
rect 141578 270567 213814 270595
rect 141578 270555 141584 270567
rect 213808 270555 213814 270567
rect 213866 270555 213872 270607
rect 284368 270555 284374 270607
rect 284426 270595 284432 270607
rect 284656 270595 284662 270607
rect 284426 270567 284662 270595
rect 284426 270555 284432 270567
rect 284656 270555 284662 270567
rect 284714 270555 284720 270607
rect 284770 270567 288014 270595
rect 137968 270481 137974 270533
rect 138026 270521 138032 270533
rect 212656 270521 212662 270533
rect 138026 270493 212662 270521
rect 138026 270481 138032 270493
rect 212656 270481 212662 270493
rect 212714 270481 212720 270533
rect 262960 270481 262966 270533
rect 263018 270521 263024 270533
rect 279760 270521 279766 270533
rect 263018 270493 279766 270521
rect 263018 270481 263024 270493
rect 279760 270481 279766 270493
rect 279818 270481 279824 270533
rect 280144 270481 280150 270533
rect 280202 270521 280208 270533
rect 284770 270521 284798 270567
rect 280202 270493 284798 270521
rect 287986 270521 288014 270567
rect 293968 270555 293974 270607
rect 294026 270595 294032 270607
rect 296482 270595 296510 270641
rect 356656 270629 356662 270641
rect 356714 270629 356720 270681
rect 371248 270629 371254 270681
rect 371306 270669 371312 270681
rect 509200 270669 509206 270681
rect 371306 270641 509206 270669
rect 371306 270629 371312 270641
rect 509200 270629 509206 270641
rect 509258 270629 509264 270681
rect 294026 270567 296510 270595
rect 294026 270555 294032 270567
rect 296560 270555 296566 270607
rect 296618 270595 296624 270607
rect 315280 270595 315286 270607
rect 296618 270567 315286 270595
rect 296618 270555 296624 270567
rect 315280 270555 315286 270567
rect 315338 270555 315344 270607
rect 345424 270555 345430 270607
rect 345482 270595 345488 270607
rect 484240 270595 484246 270607
rect 345482 270567 484246 270595
rect 345482 270555 345488 270567
rect 484240 270555 484246 270567
rect 484298 270555 484304 270607
rect 322384 270521 322390 270533
rect 287986 270493 322390 270521
rect 280202 270481 280208 270493
rect 322384 270481 322390 270493
rect 322442 270481 322448 270533
rect 348400 270481 348406 270533
rect 348458 270521 348464 270533
rect 491344 270521 491350 270533
rect 348458 270493 491350 270521
rect 348458 270481 348464 270493
rect 491344 270481 491350 270493
rect 491402 270481 491408 270533
rect 134416 270407 134422 270459
rect 134474 270447 134480 270459
rect 211888 270447 211894 270459
rect 134474 270419 211894 270447
rect 134474 270407 134480 270419
rect 211888 270407 211894 270419
rect 211946 270407 211952 270459
rect 253936 270407 253942 270459
rect 253994 270447 254000 270459
rect 257296 270447 257302 270459
rect 253994 270419 257302 270447
rect 253994 270407 254000 270419
rect 257296 270407 257302 270419
rect 257354 270407 257360 270459
rect 262480 270407 262486 270459
rect 262538 270447 262544 270459
rect 278608 270447 278614 270459
rect 262538 270419 278614 270447
rect 262538 270407 262544 270419
rect 278608 270407 278614 270419
rect 278666 270407 278672 270459
rect 279280 270407 279286 270459
rect 279338 270447 279344 270459
rect 284272 270447 284278 270459
rect 279338 270419 284278 270447
rect 279338 270407 279344 270419
rect 284272 270407 284278 270419
rect 284330 270407 284336 270459
rect 284752 270407 284758 270459
rect 284810 270447 284816 270459
rect 318832 270447 318838 270459
rect 284810 270419 318838 270447
rect 284810 270407 284816 270419
rect 318832 270407 318838 270419
rect 318890 270407 318896 270459
rect 348112 270407 348118 270459
rect 348170 270447 348176 270459
rect 490192 270447 490198 270459
rect 348170 270419 490198 270447
rect 348170 270407 348176 270419
rect 490192 270407 490198 270419
rect 490250 270407 490256 270459
rect 121456 270333 121462 270385
rect 121514 270373 121520 270385
rect 208336 270373 208342 270385
rect 121514 270345 208342 270373
rect 121514 270333 121520 270345
rect 208336 270333 208342 270345
rect 208394 270333 208400 270385
rect 278896 270333 278902 270385
rect 278954 270373 278960 270385
rect 284368 270373 284374 270385
rect 278954 270345 284374 270373
rect 278954 270333 278960 270345
rect 284368 270333 284374 270345
rect 284426 270333 284432 270385
rect 284848 270333 284854 270385
rect 284906 270373 284912 270385
rect 323536 270373 323542 270385
rect 284906 270345 323542 270373
rect 284906 270333 284912 270345
rect 323536 270333 323542 270345
rect 323594 270333 323600 270385
rect 350704 270333 350710 270385
rect 350762 270373 350768 270385
rect 497296 270373 497302 270385
rect 350762 270345 497302 270373
rect 350762 270333 350768 270345
rect 497296 270333 497302 270345
rect 497354 270333 497360 270385
rect 117904 270259 117910 270311
rect 117962 270299 117968 270311
rect 207568 270299 207574 270311
rect 117962 270271 207574 270299
rect 117962 270259 117968 270271
rect 207568 270259 207574 270271
rect 207626 270259 207632 270311
rect 255280 270259 255286 270311
rect 255338 270299 255344 270311
rect 260848 270299 260854 270311
rect 255338 270271 260854 270299
rect 255338 270259 255344 270271
rect 260848 270259 260854 270271
rect 260906 270259 260912 270311
rect 262000 270259 262006 270311
rect 262058 270299 262064 270311
rect 277456 270299 277462 270311
rect 262058 270271 277462 270299
rect 262058 270259 262064 270271
rect 277456 270259 277462 270271
rect 277514 270259 277520 270311
rect 284560 270299 284566 270311
rect 277570 270271 284566 270299
rect 114352 270185 114358 270237
rect 114410 270225 114416 270237
rect 206416 270225 206422 270237
rect 114410 270197 206422 270225
rect 114410 270185 114416 270197
rect 206416 270185 206422 270197
rect 206474 270185 206480 270237
rect 210544 270185 210550 270237
rect 210602 270225 210608 270237
rect 222832 270225 222838 270237
rect 210602 270197 222838 270225
rect 210602 270185 210608 270197
rect 222832 270185 222838 270197
rect 222890 270185 222896 270237
rect 264880 270185 264886 270237
rect 264938 270225 264944 270237
rect 277570 270225 277598 270271
rect 284560 270259 284566 270271
rect 284618 270259 284624 270311
rect 284656 270259 284662 270311
rect 284714 270299 284720 270311
rect 319984 270299 319990 270311
rect 284714 270271 319990 270299
rect 284714 270259 284720 270271
rect 319984 270259 319990 270271
rect 320042 270259 320048 270311
rect 351280 270259 351286 270311
rect 351338 270299 351344 270311
rect 498448 270299 498454 270311
rect 351338 270271 498454 270299
rect 351338 270259 351344 270271
rect 498448 270259 498454 270271
rect 498506 270259 498512 270311
rect 264938 270197 277598 270225
rect 264938 270185 264944 270197
rect 283696 270185 283702 270237
rect 283754 270225 283760 270237
rect 330640 270225 330646 270237
rect 283754 270197 330646 270225
rect 283754 270185 283760 270197
rect 330640 270185 330646 270197
rect 330698 270185 330704 270237
rect 354064 270185 354070 270237
rect 354122 270225 354128 270237
rect 505552 270225 505558 270237
rect 354122 270197 505558 270225
rect 354122 270185 354128 270197
rect 505552 270185 505558 270197
rect 505610 270185 505616 270237
rect 109552 270111 109558 270163
rect 109610 270151 109616 270163
rect 205264 270151 205270 270163
rect 109610 270123 205270 270151
rect 109610 270111 109616 270123
rect 205264 270111 205270 270123
rect 205322 270111 205328 270163
rect 210352 270111 210358 270163
rect 210410 270151 210416 270163
rect 225520 270151 225526 270163
rect 210410 270123 225526 270151
rect 210410 270111 210416 270123
rect 225520 270111 225526 270123
rect 225578 270111 225584 270163
rect 264688 270111 264694 270163
rect 264746 270151 264752 270163
rect 283312 270151 283318 270163
rect 264746 270123 283318 270151
rect 264746 270111 264752 270123
rect 283312 270111 283318 270123
rect 283370 270111 283376 270163
rect 284176 270111 284182 270163
rect 284234 270151 284240 270163
rect 331792 270151 331798 270163
rect 284234 270123 331798 270151
rect 284234 270111 284240 270123
rect 331792 270111 331798 270123
rect 331850 270111 331856 270163
rect 353680 270111 353686 270163
rect 353738 270151 353744 270163
rect 504400 270151 504406 270163
rect 353738 270123 504406 270151
rect 353738 270111 353744 270123
rect 504400 270111 504406 270123
rect 504458 270111 504464 270163
rect 107248 270037 107254 270089
rect 107306 270077 107312 270089
rect 204688 270077 204694 270089
rect 107306 270049 204694 270077
rect 107306 270037 107312 270049
rect 204688 270037 204694 270049
rect 204746 270037 204752 270089
rect 210256 270037 210262 270089
rect 210314 270077 210320 270089
rect 226672 270077 226678 270089
rect 210314 270049 226678 270077
rect 210314 270037 210320 270049
rect 226672 270037 226678 270049
rect 226730 270037 226736 270089
rect 265360 270037 265366 270089
rect 265418 270077 265424 270089
rect 285712 270077 285718 270089
rect 265418 270049 285718 270077
rect 265418 270037 265424 270049
rect 285712 270037 285718 270049
rect 285770 270037 285776 270089
rect 286288 270037 286294 270089
rect 286346 270077 286352 270089
rect 334096 270077 334102 270089
rect 286346 270049 334102 270077
rect 286346 270037 286352 270049
rect 334096 270037 334102 270049
rect 334154 270037 334160 270089
rect 356752 270037 356758 270089
rect 356810 270077 356816 270089
rect 511504 270077 511510 270089
rect 356810 270049 511510 270077
rect 356810 270037 356816 270049
rect 511504 270037 511510 270049
rect 511562 270037 511568 270089
rect 102544 269963 102550 270015
rect 102602 270003 102608 270015
rect 203344 270003 203350 270015
rect 102602 269975 203350 270003
rect 102602 269963 102608 269975
rect 203344 269963 203350 269975
rect 203402 269963 203408 270015
rect 210448 269963 210454 270015
rect 210506 270003 210512 270015
rect 224752 270003 224758 270015
rect 210506 269975 224758 270003
rect 210506 269963 210512 269975
rect 224752 269963 224758 269975
rect 224810 269963 224816 270015
rect 267088 269963 267094 270015
rect 267146 270003 267152 270015
rect 289264 270003 289270 270015
rect 267146 269975 289270 270003
rect 267146 269963 267152 269975
rect 289264 269963 289270 269975
rect 289322 269963 289328 270015
rect 342448 270003 342454 270015
rect 289378 269975 342454 270003
rect 100144 269889 100150 269941
rect 100202 269929 100208 269941
rect 202864 269929 202870 269941
rect 100202 269901 202870 269929
rect 100202 269889 100208 269901
rect 202864 269889 202870 269901
rect 202922 269889 202928 269941
rect 205168 269889 205174 269941
rect 205226 269929 205232 269941
rect 224080 269929 224086 269941
rect 205226 269901 224086 269929
rect 205226 269889 205232 269901
rect 224080 269889 224086 269901
rect 224138 269889 224144 269941
rect 256240 269889 256246 269941
rect 256298 269929 256304 269941
rect 263248 269929 263254 269941
rect 256298 269901 263254 269929
rect 256298 269889 256304 269901
rect 263248 269889 263254 269901
rect 263306 269889 263312 269941
rect 266512 269889 266518 269941
rect 266570 269929 266576 269941
rect 266570 269901 277886 269929
rect 266570 269889 266576 269901
rect 95440 269815 95446 269867
rect 95498 269855 95504 269867
rect 185584 269855 185590 269867
rect 95498 269827 185590 269855
rect 95498 269815 95504 269827
rect 185584 269815 185590 269827
rect 185642 269815 185648 269867
rect 200944 269855 200950 269867
rect 185698 269827 200950 269855
rect 93040 269741 93046 269793
rect 93098 269781 93104 269793
rect 185698 269781 185726 269827
rect 200944 269815 200950 269827
rect 201002 269815 201008 269867
rect 205936 269815 205942 269867
rect 205994 269855 206000 269867
rect 225232 269855 225238 269867
rect 205994 269827 225238 269855
rect 205994 269815 206000 269827
rect 225232 269815 225238 269827
rect 225290 269815 225296 269867
rect 261808 269815 261814 269867
rect 261866 269855 261872 269867
rect 276208 269855 276214 269867
rect 261866 269827 276214 269855
rect 261866 269815 261872 269827
rect 276208 269815 276214 269827
rect 276266 269815 276272 269867
rect 277858 269855 277886 269901
rect 280624 269889 280630 269941
rect 280682 269929 280688 269941
rect 284848 269929 284854 269941
rect 280682 269901 284854 269929
rect 280682 269889 280688 269901
rect 284848 269889 284854 269901
rect 284906 269889 284912 269941
rect 288496 269889 288502 269941
rect 288554 269929 288560 269941
rect 289378 269929 289406 269975
rect 342448 269963 342454 269975
rect 342506 269963 342512 270015
rect 356944 269963 356950 270015
rect 357002 270003 357008 270015
rect 512656 270003 512662 270015
rect 357002 269975 512662 270003
rect 357002 269963 357008 269975
rect 512656 269963 512662 269975
rect 512714 269963 512720 270015
rect 337936 269929 337942 269941
rect 288554 269901 289406 269929
rect 290530 269901 337942 269929
rect 288554 269889 288560 269901
rect 288016 269855 288022 269867
rect 277858 269827 288022 269855
rect 288016 269815 288022 269827
rect 288074 269815 288080 269867
rect 199696 269781 199702 269793
rect 93098 269753 185726 269781
rect 185794 269753 199702 269781
rect 93098 269741 93104 269753
rect 90640 269667 90646 269719
rect 90698 269707 90704 269719
rect 185794 269707 185822 269753
rect 199696 269741 199702 269753
rect 199754 269741 199760 269793
rect 205840 269741 205846 269793
rect 205898 269781 205904 269793
rect 226000 269781 226006 269793
rect 205898 269753 226006 269781
rect 205898 269741 205904 269753
rect 226000 269741 226006 269753
rect 226058 269741 226064 269793
rect 255760 269741 255766 269793
rect 255818 269781 255824 269793
rect 262096 269781 262102 269793
rect 255818 269753 262102 269781
rect 255818 269741 255824 269753
rect 262096 269741 262102 269753
rect 262154 269741 262160 269793
rect 267280 269741 267286 269793
rect 267338 269781 267344 269793
rect 290416 269781 290422 269793
rect 267338 269753 290422 269781
rect 267338 269741 267344 269753
rect 290416 269741 290422 269753
rect 290474 269741 290480 269793
rect 198064 269707 198070 269719
rect 90698 269679 185822 269707
rect 195826 269679 198070 269707
rect 90698 269667 90704 269679
rect 83632 269593 83638 269645
rect 83690 269633 83696 269645
rect 195826 269633 195854 269679
rect 198064 269667 198070 269679
rect 198122 269667 198128 269719
rect 200464 269667 200470 269719
rect 200522 269707 200528 269719
rect 222352 269707 222358 269719
rect 200522 269679 222358 269707
rect 200522 269667 200528 269679
rect 222352 269667 222358 269679
rect 222410 269667 222416 269719
rect 287920 269667 287926 269719
rect 287978 269707 287984 269719
rect 290530 269707 290558 269901
rect 337936 269889 337942 269901
rect 337994 269889 338000 269941
rect 359824 269889 359830 269941
rect 359882 269929 359888 269941
rect 519760 269929 519766 269941
rect 359882 269901 519766 269929
rect 359882 269889 359888 269901
rect 519760 269889 519766 269901
rect 519818 269889 519824 269941
rect 290608 269815 290614 269867
rect 290666 269855 290672 269867
rect 342736 269855 342742 269867
rect 290666 269827 342742 269855
rect 290666 269815 290672 269827
rect 342736 269815 342742 269827
rect 342794 269815 342800 269867
rect 359344 269815 359350 269867
rect 359402 269855 359408 269867
rect 518512 269855 518518 269867
rect 359402 269827 518518 269855
rect 359402 269815 359408 269827
rect 518512 269815 518518 269827
rect 518570 269815 518576 269867
rect 291088 269741 291094 269793
rect 291146 269781 291152 269793
rect 349552 269781 349558 269793
rect 291146 269753 349558 269781
rect 291146 269741 291152 269753
rect 349552 269741 349558 269753
rect 349610 269741 349616 269793
rect 362800 269741 362806 269793
rect 362858 269781 362864 269793
rect 526864 269781 526870 269793
rect 362858 269753 526870 269781
rect 362858 269741 362864 269753
rect 526864 269741 526870 269753
rect 526922 269741 526928 269793
rect 287978 269679 290558 269707
rect 287978 269667 287984 269679
rect 362224 269667 362230 269719
rect 362282 269707 362288 269719
rect 525616 269707 525622 269719
rect 362282 269679 525622 269707
rect 362282 269667 362288 269679
rect 525616 269667 525622 269679
rect 525674 269667 525680 269719
rect 83690 269605 195854 269633
rect 83690 269593 83696 269605
rect 198640 269593 198646 269645
rect 198698 269633 198704 269645
rect 220528 269633 220534 269645
rect 198698 269605 220534 269633
rect 198698 269593 198704 269605
rect 220528 269593 220534 269605
rect 220586 269593 220592 269645
rect 249040 269593 249046 269645
rect 249098 269633 249104 269645
rect 250288 269633 250294 269645
rect 249098 269605 250294 269633
rect 249098 269593 249104 269605
rect 250288 269593 250294 269605
rect 250346 269593 250352 269645
rect 259888 269593 259894 269645
rect 259946 269633 259952 269645
rect 271504 269633 271510 269645
rect 259946 269605 271510 269633
rect 259946 269593 259952 269605
rect 271504 269593 271510 269605
rect 271562 269593 271568 269645
rect 276496 269593 276502 269645
rect 276554 269633 276560 269645
rect 291568 269633 291574 269645
rect 276554 269605 291574 269633
rect 276554 269593 276560 269605
rect 291568 269593 291574 269605
rect 291626 269593 291632 269645
rect 293488 269593 293494 269645
rect 293546 269633 293552 269645
rect 351376 269633 351382 269645
rect 293546 269605 351382 269633
rect 293546 269593 293552 269605
rect 351376 269593 351382 269605
rect 351434 269593 351440 269645
rect 365296 269593 365302 269645
rect 365354 269633 365360 269645
rect 532720 269633 532726 269645
rect 365354 269605 532726 269633
rect 365354 269593 365360 269605
rect 532720 269593 532726 269605
rect 532778 269593 532784 269645
rect 82384 269519 82390 269571
rect 82442 269559 82448 269571
rect 197392 269559 197398 269571
rect 82442 269531 197398 269559
rect 82442 269519 82448 269531
rect 197392 269519 197398 269531
rect 197450 269519 197456 269571
rect 206512 269519 206518 269571
rect 206570 269559 206576 269571
rect 233392 269559 233398 269571
rect 206570 269531 233398 269559
rect 206570 269519 206576 269531
rect 233392 269519 233398 269531
rect 233450 269519 233456 269571
rect 269200 269519 269206 269571
rect 269258 269559 269264 269571
rect 295120 269559 295126 269571
rect 269258 269531 295126 269559
rect 269258 269519 269264 269531
rect 295120 269519 295126 269531
rect 295178 269519 295184 269571
rect 297040 269519 297046 269571
rect 297098 269559 297104 269571
rect 363664 269559 363670 269571
rect 297098 269531 363670 269559
rect 297098 269519 297104 269531
rect 363664 269519 363670 269531
rect 363722 269519 363728 269571
rect 365680 269519 365686 269571
rect 365738 269559 365744 269571
rect 533872 269559 533878 269571
rect 365738 269531 533878 269559
rect 365738 269519 365744 269531
rect 533872 269519 533878 269531
rect 533930 269519 533936 269571
rect 87184 269445 87190 269497
rect 87242 269485 87248 269497
rect 199024 269485 199030 269497
rect 87242 269457 199030 269485
rect 87242 269445 87248 269457
rect 199024 269445 199030 269457
rect 199082 269445 199088 269497
rect 202960 269445 202966 269497
rect 203018 269485 203024 269497
rect 231952 269485 231958 269497
rect 203018 269457 231958 269485
rect 203018 269445 203024 269457
rect 231952 269445 231958 269457
rect 232010 269445 232016 269497
rect 268624 269445 268630 269497
rect 268682 269485 268688 269497
rect 293872 269485 293878 269497
rect 268682 269457 293878 269485
rect 268682 269445 268688 269457
rect 293872 269445 293878 269457
rect 293930 269445 293936 269497
rect 299632 269445 299638 269497
rect 299690 269485 299696 269497
rect 370768 269485 370774 269497
rect 299690 269457 370774 269485
rect 299690 269445 299696 269457
rect 370768 269445 370774 269457
rect 370826 269445 370832 269497
rect 379888 269445 379894 269497
rect 379946 269485 379952 269497
rect 569392 269485 569398 269497
rect 379946 269457 569398 269485
rect 379946 269445 379952 269457
rect 569392 269445 569398 269457
rect 569450 269445 569456 269497
rect 81232 269371 81238 269423
rect 81290 269411 81296 269423
rect 196816 269411 196822 269423
rect 81290 269383 196822 269411
rect 81290 269371 81296 269383
rect 196816 269371 196822 269383
rect 196874 269371 196880 269423
rect 204112 269371 204118 269423
rect 204170 269411 204176 269423
rect 232144 269411 232150 269423
rect 204170 269383 232150 269411
rect 204170 269371 204176 269383
rect 232144 269371 232150 269383
rect 232202 269371 232208 269423
rect 258640 269371 258646 269423
rect 258698 269411 258704 269423
rect 269104 269411 269110 269423
rect 258698 269383 269110 269411
rect 258698 269371 258704 269383
rect 269104 269371 269110 269383
rect 269162 269371 269168 269423
rect 272944 269371 272950 269423
rect 273002 269411 273008 269423
rect 304624 269411 304630 269423
rect 273002 269383 304630 269411
rect 273002 269371 273008 269383
rect 304624 269371 304630 269383
rect 304682 269371 304688 269423
rect 308272 269371 308278 269423
rect 308330 269411 308336 269423
rect 392080 269411 392086 269423
rect 308330 269383 392086 269411
rect 308330 269371 308336 269383
rect 392080 269371 392086 269383
rect 392138 269371 392144 269423
rect 394384 269371 394390 269423
rect 394442 269411 394448 269423
rect 604816 269411 604822 269423
rect 394442 269383 604822 269411
rect 394442 269371 394448 269383
rect 604816 269371 604822 269383
rect 604874 269371 604880 269423
rect 74128 269297 74134 269349
rect 74186 269337 74192 269349
rect 194992 269337 194998 269349
rect 74186 269309 194998 269337
rect 74186 269297 74192 269309
rect 194992 269297 194998 269309
rect 195050 269297 195056 269349
rect 200656 269297 200662 269349
rect 200714 269337 200720 269349
rect 230992 269337 230998 269349
rect 200714 269309 230998 269337
rect 200714 269297 200720 269309
rect 230992 269297 230998 269309
rect 231050 269297 231056 269349
rect 274672 269297 274678 269349
rect 274730 269337 274736 269349
rect 308176 269337 308182 269349
rect 274730 269309 308182 269337
rect 274730 269297 274736 269309
rect 308176 269297 308182 269309
rect 308234 269297 308240 269349
rect 311152 269297 311158 269349
rect 311210 269337 311216 269349
rect 399184 269337 399190 269349
rect 311210 269309 399190 269337
rect 311210 269297 311216 269309
rect 399184 269297 399190 269309
rect 399242 269297 399248 269349
rect 399952 269297 399958 269349
rect 400010 269337 400016 269349
rect 619024 269337 619030 269349
rect 400010 269309 619030 269337
rect 400010 269297 400016 269309
rect 619024 269297 619030 269309
rect 619082 269297 619088 269349
rect 67024 269223 67030 269275
rect 67082 269263 67088 269275
rect 192592 269263 192598 269275
rect 67082 269235 192598 269263
rect 67082 269223 67088 269235
rect 192592 269223 192598 269235
rect 192650 269223 192656 269275
rect 197104 269223 197110 269275
rect 197162 269263 197168 269275
rect 229552 269263 229558 269275
rect 197162 269235 229558 269263
rect 197162 269223 197168 269235
rect 229552 269223 229558 269235
rect 229610 269223 229616 269275
rect 260560 269223 260566 269275
rect 260618 269263 260624 269275
rect 273904 269263 273910 269275
rect 260618 269235 273910 269263
rect 260618 269223 260624 269235
rect 273904 269223 273910 269235
rect 273962 269223 273968 269275
rect 275824 269223 275830 269275
rect 275882 269263 275888 269275
rect 311728 269263 311734 269275
rect 275882 269235 311734 269263
rect 275882 269223 275888 269235
rect 311728 269223 311734 269235
rect 311786 269223 311792 269275
rect 314224 269223 314230 269275
rect 314282 269263 314288 269275
rect 406288 269263 406294 269275
rect 314282 269235 406294 269263
rect 314282 269223 314288 269235
rect 406288 269223 406294 269235
rect 406346 269223 406352 269275
rect 145072 269149 145078 269201
rect 145130 269189 145136 269201
rect 214480 269189 214486 269201
rect 145130 269161 214486 269189
rect 145130 269149 145136 269161
rect 214480 269149 214486 269161
rect 214538 269149 214544 269201
rect 286864 269189 286870 269201
rect 267826 269161 286870 269189
rect 149776 269075 149782 269127
rect 149834 269115 149840 269127
rect 216208 269115 216214 269127
rect 149834 269087 216214 269115
rect 149834 269075 149840 269087
rect 216208 269075 216214 269087
rect 216266 269075 216272 269127
rect 253360 269075 253366 269127
rect 253418 269115 253424 269127
rect 256144 269115 256150 269127
rect 253418 269087 256150 269115
rect 253418 269075 253424 269087
rect 256144 269075 256150 269087
rect 256202 269075 256208 269127
rect 257008 269075 257014 269127
rect 257066 269115 257072 269127
rect 264400 269115 264406 269127
rect 257066 269087 264406 269115
rect 257066 269075 257072 269087
rect 264400 269075 264406 269087
rect 264458 269075 264464 269127
rect 266032 269075 266038 269127
rect 266090 269115 266096 269127
rect 267826 269115 267854 269161
rect 286864 269149 286870 269161
rect 286922 269149 286928 269201
rect 286960 269149 286966 269201
rect 287018 269189 287024 269201
rect 292816 269189 292822 269201
rect 287018 269161 292822 269189
rect 287018 269149 287024 269161
rect 292816 269149 292822 269161
rect 292874 269149 292880 269201
rect 306352 269149 306358 269201
rect 306410 269189 306416 269201
rect 342160 269189 342166 269201
rect 306410 269161 342166 269189
rect 306410 269149 306416 269161
rect 342160 269149 342166 269161
rect 342218 269149 342224 269201
rect 345232 269149 345238 269201
rect 345290 269189 345296 269201
rect 483088 269189 483094 269201
rect 345290 269161 483094 269189
rect 345290 269149 345296 269161
rect 483088 269149 483094 269161
rect 483146 269149 483152 269201
rect 266090 269087 267854 269115
rect 266090 269075 266096 269087
rect 281296 269075 281302 269127
rect 281354 269115 281360 269127
rect 301072 269115 301078 269127
rect 281354 269087 301078 269115
rect 281354 269075 281360 269087
rect 301072 269075 301078 269087
rect 301130 269075 301136 269127
rect 303760 269075 303766 269127
rect 303818 269115 303824 269127
rect 334288 269115 334294 269127
rect 303818 269087 334294 269115
rect 303818 269075 303824 269087
rect 334288 269075 334294 269087
rect 334346 269075 334352 269127
rect 342640 269075 342646 269127
rect 342698 269115 342704 269127
rect 477136 269115 477142 269127
rect 342698 269087 477142 269115
rect 342698 269075 342704 269087
rect 477136 269075 477142 269087
rect 477194 269075 477200 269127
rect 148624 269001 148630 269053
rect 148682 269041 148688 269053
rect 215728 269041 215734 269053
rect 148682 269013 215734 269041
rect 148682 269001 148688 269013
rect 215728 269001 215734 269013
rect 215786 269001 215792 269053
rect 282064 269001 282070 269053
rect 282122 269041 282128 269053
rect 299440 269041 299446 269053
rect 282122 269013 299446 269041
rect 282122 269001 282128 269013
rect 299440 269001 299446 269013
rect 299498 269001 299504 269053
rect 305680 269001 305686 269053
rect 305738 269041 305744 269053
rect 384976 269041 384982 269053
rect 305738 269013 384982 269041
rect 305738 269001 305744 269013
rect 384976 269001 384982 269013
rect 385034 269001 385040 269053
rect 406576 269001 406582 269053
rect 406634 269041 406640 269053
rect 408400 269041 408406 269053
rect 406634 269013 408406 269041
rect 406634 269001 406640 269013
rect 408400 269001 408406 269013
rect 408458 269001 408464 269053
rect 152176 268927 152182 268979
rect 152234 268967 152240 268979
rect 216688 268967 216694 268979
rect 152234 268939 216694 268967
rect 152234 268927 152240 268939
rect 216688 268927 216694 268939
rect 216746 268927 216752 268979
rect 253168 268927 253174 268979
rect 253226 268967 253232 268979
rect 254992 268967 254998 268979
rect 253226 268939 254998 268967
rect 253226 268927 253232 268939
rect 254992 268927 254998 268939
rect 255050 268927 255056 268979
rect 259408 268927 259414 268979
rect 259466 268967 259472 268979
rect 270352 268967 270358 268979
rect 259466 268939 270358 268967
rect 259466 268927 259472 268939
rect 270352 268927 270358 268939
rect 270410 268927 270416 268979
rect 277552 268927 277558 268979
rect 277610 268967 277616 268979
rect 296560 268967 296566 268979
rect 277610 268939 296566 268967
rect 277610 268927 277616 268939
rect 296560 268927 296566 268939
rect 296618 268927 296624 268979
rect 302032 268927 302038 268979
rect 302090 268967 302096 268979
rect 331216 268967 331222 268979
rect 302090 268939 331222 268967
rect 302090 268927 302096 268939
rect 331216 268927 331222 268939
rect 331274 268927 331280 268979
rect 339760 268927 339766 268979
rect 339818 268967 339824 268979
rect 470128 268967 470134 268979
rect 339818 268939 470134 268967
rect 339818 268927 339824 268939
rect 470128 268927 470134 268939
rect 470186 268927 470192 268979
rect 156880 268853 156886 268905
rect 156938 268893 156944 268905
rect 218128 268893 218134 268905
rect 156938 268865 218134 268893
rect 156938 268853 156944 268865
rect 218128 268853 218134 268865
rect 218186 268853 218192 268905
rect 260080 268853 260086 268905
rect 260138 268893 260144 268905
rect 272656 268893 272662 268905
rect 260138 268865 272662 268893
rect 260138 268853 260144 268865
rect 272656 268853 272662 268865
rect 272714 268853 272720 268905
rect 300688 268853 300694 268905
rect 300746 268893 300752 268905
rect 326800 268893 326806 268905
rect 300746 268865 326806 268893
rect 300746 268853 300752 268865
rect 326800 268853 326806 268865
rect 326858 268853 326864 268905
rect 336880 268853 336886 268905
rect 336938 268893 336944 268905
rect 463024 268893 463030 268905
rect 336938 268865 463030 268893
rect 336938 268853 336944 268865
rect 463024 268853 463030 268865
rect 463082 268853 463088 268905
rect 163984 268779 163990 268831
rect 164042 268819 164048 268831
rect 219952 268819 219958 268831
rect 164042 268791 219958 268819
rect 164042 268779 164048 268791
rect 219952 268779 219958 268791
rect 220010 268779 220016 268831
rect 258160 268779 258166 268831
rect 258218 268819 258224 268831
rect 267952 268819 267958 268831
rect 258218 268791 267958 268819
rect 258218 268779 258224 268791
rect 267952 268779 267958 268791
rect 268010 268779 268016 268831
rect 268432 268779 268438 268831
rect 268490 268819 268496 268831
rect 286960 268819 286966 268831
rect 268490 268791 286966 268819
rect 268490 268779 268496 268791
rect 286960 268779 286966 268791
rect 287018 268779 287024 268831
rect 289168 268779 289174 268831
rect 289226 268819 289232 268831
rect 308368 268819 308374 268831
rect 289226 268791 308374 268819
rect 289226 268779 289232 268791
rect 308368 268779 308374 268791
rect 308426 268779 308432 268831
rect 334288 268779 334294 268831
rect 334346 268819 334352 268831
rect 455920 268819 455926 268831
rect 334346 268791 455926 268819
rect 334346 268779 334352 268791
rect 455920 268779 455926 268791
rect 455978 268779 455984 268831
rect 155728 268705 155734 268757
rect 155786 268745 155792 268757
rect 217360 268745 217366 268757
rect 155786 268717 217366 268745
rect 155786 268705 155792 268717
rect 217360 268705 217366 268717
rect 217418 268705 217424 268757
rect 257680 268705 257686 268757
rect 257738 268745 257744 268757
rect 266800 268745 266806 268757
rect 257738 268717 266806 268745
rect 257738 268705 257744 268717
rect 266800 268705 266806 268717
rect 266858 268705 266864 268757
rect 295216 268705 295222 268757
rect 295274 268745 295280 268757
rect 307024 268745 307030 268757
rect 295274 268717 307030 268745
rect 295274 268705 295280 268717
rect 307024 268705 307030 268717
rect 307082 268705 307088 268757
rect 331216 268705 331222 268757
rect 331274 268745 331280 268757
rect 448816 268745 448822 268757
rect 331274 268717 448822 268745
rect 331274 268705 331280 268717
rect 448816 268705 448822 268717
rect 448874 268705 448880 268757
rect 162832 268631 162838 268683
rect 162890 268671 162896 268683
rect 219280 268671 219286 268683
rect 162890 268643 219286 268671
rect 162890 268631 162896 268643
rect 219280 268631 219286 268643
rect 219338 268631 219344 268683
rect 254608 268631 254614 268683
rect 254666 268671 254672 268683
rect 258544 268671 258550 268683
rect 254666 268643 258550 268671
rect 254666 268631 254672 268643
rect 258544 268631 258550 268643
rect 258602 268631 258608 268683
rect 271504 268631 271510 268683
rect 271562 268671 271568 268683
rect 300976 268671 300982 268683
rect 271562 268643 300982 268671
rect 271562 268631 271568 268643
rect 300976 268631 300982 268643
rect 301034 268631 301040 268683
rect 328336 268631 328342 268683
rect 328394 268671 328400 268683
rect 441712 268671 441718 268683
rect 328394 268643 441718 268671
rect 328394 268631 328400 268643
rect 441712 268631 441718 268643
rect 441770 268631 441776 268683
rect 171088 268557 171094 268609
rect 171146 268597 171152 268609
rect 221776 268597 221782 268609
rect 171146 268569 221782 268597
rect 171146 268557 171152 268569
rect 221776 268557 221782 268569
rect 221834 268557 221840 268609
rect 325744 268557 325750 268609
rect 325802 268597 325808 268609
rect 434608 268597 434614 268609
rect 325802 268569 434614 268597
rect 325802 268557 325808 268569
rect 434608 268557 434614 268569
rect 434666 268557 434672 268609
rect 169744 268483 169750 268535
rect 169802 268523 169808 268535
rect 221200 268523 221206 268535
rect 169802 268495 221206 268523
rect 169802 268483 169808 268495
rect 221200 268483 221206 268495
rect 221258 268483 221264 268535
rect 261232 268483 261238 268535
rect 261290 268523 261296 268535
rect 275056 268523 275062 268535
rect 261290 268495 275062 268523
rect 261290 268483 261296 268495
rect 275056 268483 275062 268495
rect 275114 268483 275120 268535
rect 322576 268483 322582 268535
rect 322634 268523 322640 268535
rect 427504 268523 427510 268535
rect 322634 268495 427510 268523
rect 322634 268483 322640 268495
rect 427504 268483 427510 268495
rect 427562 268483 427568 268535
rect 176944 268409 176950 268461
rect 177002 268449 177008 268461
rect 223408 268449 223414 268461
rect 177002 268421 223414 268449
rect 177002 268409 177008 268421
rect 223408 268409 223414 268421
rect 223466 268409 223472 268461
rect 319696 268409 319702 268461
rect 319754 268449 319760 268461
rect 420496 268449 420502 268461
rect 319754 268421 420502 268449
rect 319754 268409 319760 268421
rect 420496 268409 420502 268421
rect 420554 268409 420560 268461
rect 178192 268335 178198 268387
rect 178250 268375 178256 268387
rect 223600 268375 223606 268387
rect 178250 268347 223606 268375
rect 178250 268335 178256 268347
rect 223600 268335 223606 268347
rect 223658 268335 223664 268387
rect 247888 268335 247894 268387
rect 247946 268375 247952 268387
rect 249808 268375 249814 268387
rect 247946 268347 249814 268375
rect 247946 268335 247952 268347
rect 249808 268335 249814 268347
rect 249866 268335 249872 268387
rect 255088 268335 255094 268387
rect 255146 268375 255152 268387
rect 259696 268375 259702 268387
rect 255146 268347 259702 268375
rect 255146 268335 255152 268347
rect 259696 268335 259702 268347
rect 259754 268335 259760 268387
rect 317104 268335 317110 268387
rect 317162 268375 317168 268387
rect 408976 268375 408982 268387
rect 317162 268347 408982 268375
rect 317162 268335 317168 268347
rect 408976 268335 408982 268347
rect 409034 268335 409040 268387
rect 185584 268261 185590 268313
rect 185642 268301 185648 268313
rect 201136 268301 201142 268313
rect 185642 268273 201142 268301
rect 185642 268261 185648 268273
rect 201136 268261 201142 268273
rect 201194 268261 201200 268313
rect 207472 268261 207478 268313
rect 207530 268301 207536 268313
rect 212464 268301 212470 268313
rect 207530 268273 212470 268301
rect 207530 268261 207536 268273
rect 212464 268261 212470 268273
rect 212522 268261 212528 268313
rect 221488 268261 221494 268313
rect 221546 268301 221552 268313
rect 227824 268301 227830 268313
rect 221546 268273 227830 268301
rect 221546 268261 221552 268273
rect 227824 268261 227830 268273
rect 227882 268261 227888 268313
rect 312304 268261 312310 268313
rect 312362 268301 312368 268313
rect 348496 268301 348502 268313
rect 312362 268273 348502 268301
rect 312362 268261 312368 268273
rect 348496 268261 348502 268273
rect 348554 268261 348560 268313
rect 192976 268187 192982 268239
rect 193034 268227 193040 268239
rect 218608 268227 218614 268239
rect 193034 268199 218614 268227
rect 193034 268187 193040 268199
rect 218608 268187 218614 268199
rect 218666 268187 218672 268239
rect 224368 268187 224374 268239
rect 224426 268227 224432 268239
rect 230032 268227 230038 268239
rect 224426 268199 230038 268227
rect 224426 268187 224432 268199
rect 230032 268187 230038 268199
rect 230090 268187 230096 268239
rect 257488 268187 257494 268239
rect 257546 268227 257552 268239
rect 265648 268227 265654 268239
rect 257546 268199 265654 268227
rect 257546 268187 257552 268199
rect 265648 268187 265654 268199
rect 265706 268187 265712 268239
rect 309232 268187 309238 268239
rect 309290 268227 309296 268239
rect 347056 268227 347062 268239
rect 309290 268199 347062 268227
rect 309290 268187 309296 268199
rect 347056 268187 347062 268199
rect 347114 268187 347120 268239
rect 408496 268187 408502 268239
rect 408554 268227 408560 268239
rect 640336 268227 640342 268239
rect 408554 268199 640342 268227
rect 408554 268187 408560 268199
rect 640336 268187 640342 268199
rect 640394 268187 640400 268239
rect 190096 268113 190102 268165
rect 190154 268153 190160 268165
rect 210736 268153 210742 268165
rect 190154 268125 210742 268153
rect 190154 268113 190160 268125
rect 210736 268113 210742 268125
rect 210794 268113 210800 268165
rect 223696 268113 223702 268165
rect 223754 268153 223760 268165
rect 231472 268153 231478 268165
rect 223754 268125 231478 268153
rect 223754 268113 223760 268125
rect 231472 268113 231478 268125
rect 231530 268113 231536 268165
rect 264112 268113 264118 268165
rect 264170 268153 264176 268165
rect 282160 268153 282166 268165
rect 264170 268125 282166 268153
rect 264170 268113 264176 268125
rect 282160 268113 282166 268125
rect 282218 268113 282224 268165
rect 302608 268113 302614 268165
rect 302666 268153 302672 268165
rect 377872 268153 377878 268165
rect 302666 268125 377878 268153
rect 302666 268113 302672 268125
rect 377872 268113 377878 268125
rect 377930 268113 377936 268165
rect 384112 268113 384118 268165
rect 384170 268153 384176 268165
rect 516304 268153 516310 268165
rect 384170 268125 516310 268153
rect 384170 268113 384176 268125
rect 516304 268113 516310 268125
rect 516362 268113 516368 268165
rect 207376 268039 207382 268091
rect 207434 268079 207440 268091
rect 216880 268079 216886 268091
rect 207434 268051 216886 268079
rect 207434 268039 207440 268051
rect 216880 268039 216886 268051
rect 216938 268039 216944 268091
rect 221584 268039 221590 268091
rect 221642 268079 221648 268091
rect 230512 268079 230518 268091
rect 221642 268051 230518 268079
rect 221642 268039 221648 268051
rect 230512 268039 230518 268051
rect 230570 268039 230576 268091
rect 252688 268039 252694 268091
rect 252746 268079 252752 268091
rect 253744 268079 253750 268091
rect 252746 268051 253750 268079
rect 252746 268039 252752 268051
rect 253744 268039 253750 268051
rect 253802 268039 253808 268091
rect 342160 268039 342166 268091
rect 342218 268079 342224 268091
rect 359440 268079 359446 268091
rect 342218 268051 359446 268079
rect 342218 268039 342224 268051
rect 359440 268039 359446 268051
rect 359498 268039 359504 268091
rect 209872 267965 209878 268017
rect 209930 268005 209936 268017
rect 211408 268005 211414 268017
rect 209930 267977 211414 268005
rect 209930 267965 209936 267977
rect 211408 267965 211414 267977
rect 211466 267965 211472 268017
rect 221680 267965 221686 268017
rect 221738 268005 221744 268017
rect 229072 268005 229078 268017
rect 221738 267977 229078 268005
rect 221738 267965 221744 267977
rect 229072 267965 229078 267977
rect 229130 267965 229136 268017
rect 333616 267965 333622 268017
rect 333674 268005 333680 268017
rect 351376 268005 351382 268017
rect 333674 267977 351382 268005
rect 333674 267965 333680 267977
rect 351376 267965 351382 267977
rect 351434 267965 351440 268017
rect 210640 267891 210646 267943
rect 210698 267931 210704 267943
rect 221008 267931 221014 267943
rect 210698 267903 221014 267931
rect 210698 267891 210704 267903
rect 221008 267891 221014 267903
rect 221066 267891 221072 267943
rect 224464 267891 224470 267943
rect 224522 267931 224528 267943
rect 228400 267931 228406 267943
rect 224522 267903 228406 267931
rect 224522 267891 224528 267903
rect 228400 267891 228406 267903
rect 228458 267891 228464 267943
rect 263632 267891 263638 267943
rect 263690 267931 263696 267943
rect 281008 267931 281014 267943
rect 263690 267903 281014 267931
rect 263690 267891 263696 267903
rect 281008 267891 281014 267903
rect 281066 267891 281072 267943
rect 282544 267891 282550 267943
rect 282602 267931 282608 267943
rect 299344 267931 299350 267943
rect 282602 267903 299350 267931
rect 282602 267891 282608 267903
rect 299344 267891 299350 267903
rect 299402 267891 299408 267943
rect 336688 267891 336694 267943
rect 336746 267931 336752 267943
rect 354256 267931 354262 267943
rect 336746 267903 354262 267931
rect 336746 267891 336752 267903
rect 354256 267891 354262 267903
rect 354314 267891 354320 267943
rect 199120 267817 199126 267869
rect 199178 267857 199184 267869
rect 202288 267857 202294 267869
rect 199178 267829 202294 267857
rect 199178 267817 199184 267829
rect 202288 267817 202294 267829
rect 202346 267817 202352 267869
rect 207280 267817 207286 267869
rect 207338 267857 207344 267869
rect 209488 267857 209494 267869
rect 207338 267829 209494 267857
rect 207338 267817 207344 267829
rect 209488 267817 209494 267829
rect 209546 267817 209552 267869
rect 209776 267817 209782 267869
rect 209834 267857 209840 267869
rect 212368 267857 212374 267869
rect 209834 267829 212374 267857
rect 209834 267817 209840 267829
rect 212368 267817 212374 267829
rect 212426 267817 212432 267869
rect 212464 267817 212470 267869
rect 212522 267857 212528 267869
rect 218896 267857 218902 267869
rect 212522 267829 218902 267857
rect 212522 267817 212528 267829
rect 218896 267817 218902 267829
rect 218954 267817 218960 267869
rect 224560 267817 224566 267869
rect 224618 267857 224624 267869
rect 227632 267857 227638 267869
rect 224618 267829 227638 267857
rect 224618 267817 224624 267829
rect 227632 267817 227638 267829
rect 227690 267817 227696 267869
rect 339280 267817 339286 267869
rect 339338 267857 339344 267869
rect 360400 267857 360406 267869
rect 339338 267829 360406 267857
rect 339338 267817 339344 267829
rect 360400 267817 360406 267829
rect 360458 267817 360464 267869
rect 401296 267817 401302 267869
rect 401354 267857 401360 267869
rect 402928 267857 402934 267869
rect 401354 267829 402934 267857
rect 401354 267817 401360 267829
rect 402928 267817 402934 267829
rect 402986 267817 402992 267869
rect 409936 267817 409942 267869
rect 409994 267857 410000 267869
rect 413680 267857 413686 267869
rect 409994 267829 413686 267857
rect 409994 267817 410000 267829
rect 413680 267817 413686 267829
rect 413738 267817 413744 267869
rect 351952 267743 351958 267795
rect 352010 267783 352016 267795
rect 499600 267783 499606 267795
rect 352010 267755 499606 267783
rect 352010 267743 352016 267755
rect 499600 267743 499606 267755
rect 499658 267743 499664 267795
rect 354832 267669 354838 267721
rect 354890 267709 354896 267721
rect 506704 267709 506710 267721
rect 354890 267681 506710 267709
rect 354890 267669 354896 267681
rect 506704 267669 506710 267681
rect 506762 267669 506768 267721
rect 357424 267595 357430 267647
rect 357482 267635 357488 267647
rect 513808 267635 513814 267647
rect 357482 267607 513814 267635
rect 357482 267595 357488 267607
rect 513808 267595 513814 267607
rect 513866 267595 513872 267647
rect 360304 267521 360310 267573
rect 360362 267561 360368 267573
rect 520912 267561 520918 267573
rect 360362 267533 520918 267561
rect 360362 267521 360368 267533
rect 520912 267521 520918 267533
rect 520970 267521 520976 267573
rect 363376 267447 363382 267499
rect 363434 267487 363440 267499
rect 528016 267487 528022 267499
rect 363434 267459 528022 267487
rect 363434 267447 363440 267459
rect 528016 267447 528022 267459
rect 528074 267447 528080 267499
rect 365968 267373 365974 267425
rect 366026 267413 366032 267425
rect 535120 267413 535126 267425
rect 366026 267385 535126 267413
rect 366026 267373 366032 267385
rect 535120 267373 535126 267385
rect 535178 267373 535184 267425
rect 368944 267299 368950 267351
rect 369002 267339 369008 267351
rect 542224 267339 542230 267351
rect 369002 267311 542230 267339
rect 369002 267299 369008 267311
rect 542224 267299 542230 267311
rect 542282 267299 542288 267351
rect 372496 267225 372502 267277
rect 372554 267265 372560 267277
rect 550480 267265 550486 267277
rect 372554 267237 550486 267265
rect 372554 267225 372560 267237
rect 550480 267225 550486 267237
rect 550538 267225 550544 267277
rect 384880 267151 384886 267203
rect 384938 267191 384944 267203
rect 581200 267191 581206 267203
rect 384938 267163 581206 267191
rect 384938 267151 384944 267163
rect 581200 267151 581206 267163
rect 581258 267151 581264 267203
rect 386032 267077 386038 267129
rect 386090 267117 386096 267129
rect 584752 267117 584758 267129
rect 386090 267089 584758 267117
rect 386090 267077 386096 267089
rect 584752 267077 584758 267089
rect 584810 267077 584816 267129
rect 387760 267003 387766 267055
rect 387818 267043 387824 267055
rect 588304 267043 588310 267055
rect 387818 267015 588310 267043
rect 387818 267003 387824 267015
rect 588304 267003 588310 267015
rect 588362 267003 588368 267055
rect 301840 266929 301846 266981
rect 301898 266969 301904 266981
rect 375280 266969 375286 266981
rect 301898 266941 375286 266969
rect 301898 266929 301904 266941
rect 375280 266929 375286 266941
rect 375338 266929 375344 266981
rect 394672 266929 394678 266981
rect 394730 266969 394736 266981
rect 606064 266969 606070 266981
rect 394730 266941 606070 266969
rect 394730 266929 394736 266941
rect 606064 266929 606070 266941
rect 606122 266929 606128 266981
rect 306160 266855 306166 266907
rect 306218 266895 306224 266907
rect 386128 266895 386134 266907
rect 306218 266867 386134 266895
rect 306218 266855 306224 266867
rect 386128 266855 386134 266867
rect 386186 266855 386192 266907
rect 393232 266855 393238 266907
rect 393290 266895 393296 266907
rect 602512 266895 602518 266907
rect 393290 266867 602518 266895
rect 393290 266855 393296 266867
rect 602512 266855 602518 266867
rect 602570 266855 602576 266907
rect 305008 266781 305014 266833
rect 305066 266821 305072 266833
rect 383824 266821 383830 266833
rect 305066 266793 383830 266821
rect 305066 266781 305072 266793
rect 383824 266781 383830 266793
rect 383882 266781 383888 266833
rect 397552 266781 397558 266833
rect 397610 266821 397616 266833
rect 613072 266821 613078 266833
rect 397610 266793 613078 266821
rect 397610 266781 397616 266793
rect 613072 266781 613078 266793
rect 613130 266781 613136 266833
rect 308752 266707 308758 266759
rect 308810 266747 308816 266759
rect 392944 266747 392950 266759
rect 308810 266719 392950 266747
rect 308810 266707 308816 266719
rect 392944 266707 392950 266719
rect 393002 266707 393008 266759
rect 398224 266707 398230 266759
rect 398282 266747 398288 266759
rect 614320 266747 614326 266759
rect 398282 266719 614326 266747
rect 398282 266707 398288 266719
rect 614320 266707 614326 266719
rect 614378 266707 614384 266759
rect 308080 266633 308086 266685
rect 308138 266673 308144 266685
rect 390928 266673 390934 266685
rect 308138 266645 390934 266673
rect 308138 266633 308144 266645
rect 390928 266633 390934 266645
rect 390986 266633 390992 266685
rect 400624 266633 400630 266685
rect 400682 266673 400688 266685
rect 620176 266673 620182 266685
rect 400682 266645 620182 266673
rect 400682 266633 400688 266645
rect 620176 266633 620182 266645
rect 620234 266633 620240 266685
rect 310672 266559 310678 266611
rect 310730 266599 310736 266611
rect 398032 266599 398038 266611
rect 310730 266571 398038 266599
rect 310730 266559 310736 266571
rect 398032 266559 398038 266571
rect 398090 266559 398096 266611
rect 403216 266559 403222 266611
rect 403274 266599 403280 266611
rect 627280 266599 627286 266611
rect 403274 266571 627286 266599
rect 403274 266559 403280 266571
rect 627280 266559 627286 266571
rect 627338 266559 627344 266611
rect 313552 266485 313558 266537
rect 313610 266525 313616 266537
rect 405040 266525 405046 266537
rect 313610 266497 405046 266525
rect 313610 266485 313616 266497
rect 405040 266485 405046 266497
rect 405098 266485 405104 266537
rect 406096 266485 406102 266537
rect 406154 266525 406160 266537
rect 634384 266525 634390 266537
rect 406154 266497 634390 266525
rect 406154 266485 406160 266497
rect 634384 266485 634390 266497
rect 634442 266485 634448 266537
rect 313072 266411 313078 266463
rect 313130 266451 313136 266463
rect 403888 266451 403894 266463
rect 313130 266423 403894 266451
rect 313130 266411 313136 266423
rect 403888 266411 403894 266423
rect 403946 266411 403952 266463
rect 409168 266411 409174 266463
rect 409226 266451 409232 266463
rect 641488 266451 641494 266463
rect 409226 266423 641494 266451
rect 409226 266411 409232 266423
rect 641488 266411 641494 266423
rect 641546 266411 641552 266463
rect 45040 266337 45046 266389
rect 45098 266377 45104 266389
rect 673744 266377 673750 266389
rect 45098 266349 673750 266377
rect 45098 266337 45104 266349
rect 673744 266337 673750 266349
rect 673802 266337 673808 266389
rect 348880 266263 348886 266315
rect 348938 266303 348944 266315
rect 492592 266303 492598 266315
rect 348938 266275 492598 266303
rect 348938 266263 348944 266275
rect 492592 266263 492598 266275
rect 492650 266263 492656 266315
rect 346000 266189 346006 266241
rect 346058 266229 346064 266241
rect 485488 266229 485494 266241
rect 346058 266201 485494 266229
rect 346058 266189 346064 266201
rect 485488 266189 485494 266201
rect 485546 266189 485552 266241
rect 343312 266115 343318 266167
rect 343370 266155 343376 266167
rect 478384 266155 478390 266167
rect 343370 266127 478390 266155
rect 343370 266115 343376 266127
rect 478384 266115 478390 266127
rect 478442 266115 478448 266167
rect 340240 266041 340246 266093
rect 340298 266081 340304 266093
rect 471280 266081 471286 266093
rect 340298 266053 471286 266081
rect 340298 266041 340304 266053
rect 471280 266041 471286 266053
rect 471338 266041 471344 266093
rect 337360 265967 337366 266019
rect 337418 266007 337424 266019
rect 464176 266007 464182 266019
rect 337418 265979 464182 266007
rect 337418 265967 337424 265979
rect 464176 265967 464182 265979
rect 464234 265967 464240 266019
rect 334768 265893 334774 265945
rect 334826 265933 334832 265945
rect 457072 265933 457078 265945
rect 334826 265905 457078 265933
rect 334826 265893 334832 265905
rect 457072 265893 457078 265905
rect 457130 265893 457136 265945
rect 331888 265819 331894 265871
rect 331946 265859 331952 265871
rect 449968 265859 449974 265871
rect 331946 265831 449974 265859
rect 331946 265819 331952 265831
rect 449968 265819 449974 265831
rect 450026 265819 450032 265871
rect 327568 265745 327574 265797
rect 327626 265785 327632 265797
rect 439312 265785 439318 265797
rect 327626 265757 439318 265785
rect 327626 265745 327632 265757
rect 439312 265745 439318 265757
rect 439370 265745 439376 265797
rect 324496 265671 324502 265723
rect 324554 265711 324560 265723
rect 432304 265711 432310 265723
rect 324554 265683 432310 265711
rect 324554 265671 324560 265683
rect 432304 265671 432310 265683
rect 432362 265671 432368 265723
rect 321616 265597 321622 265649
rect 321674 265637 321680 265649
rect 425200 265637 425206 265649
rect 321674 265609 425206 265637
rect 321674 265597 321680 265609
rect 425200 265597 425206 265609
rect 425258 265597 425264 265649
rect 408016 265523 408022 265575
rect 408074 265563 408080 265575
rect 508240 265563 508246 265575
rect 408074 265535 508246 265563
rect 408074 265523 408080 265535
rect 508240 265523 508246 265535
rect 508298 265523 508304 265575
rect 319024 265449 319030 265501
rect 319082 265489 319088 265501
rect 418096 265489 418102 265501
rect 319082 265461 418102 265489
rect 319082 265449 319088 265461
rect 418096 265449 418102 265461
rect 418154 265449 418160 265501
rect 656560 265375 656566 265427
rect 656618 265415 656624 265427
rect 676048 265415 676054 265427
rect 656618 265387 676054 265415
rect 656618 265375 656624 265387
rect 676048 265375 676054 265387
rect 676106 265375 676112 265427
rect 656272 265227 656278 265279
rect 656330 265267 656336 265279
rect 676240 265267 676246 265279
rect 656330 265239 676246 265267
rect 656330 265227 656336 265239
rect 676240 265227 676246 265239
rect 676298 265227 676304 265279
rect 656080 265079 656086 265131
rect 656138 265119 656144 265131
rect 676144 265119 676150 265131
rect 656138 265091 676150 265119
rect 656138 265079 656144 265091
rect 676144 265079 676150 265091
rect 676202 265079 676208 265131
rect 23056 265005 23062 265057
rect 23114 265045 23120 265057
rect 43504 265045 43510 265057
rect 23114 265017 43510 265045
rect 23114 265005 23120 265017
rect 43504 265005 43510 265017
rect 43562 265005 43568 265057
rect 673744 265005 673750 265057
rect 673802 265045 673808 265057
rect 676048 265045 676054 265057
rect 673802 265017 676054 265045
rect 673802 265005 673808 265017
rect 676048 265005 676054 265017
rect 676106 265005 676112 265057
rect 42160 264931 42166 264983
rect 42218 264971 42224 264983
rect 53296 264971 53302 264983
rect 42218 264943 53302 264971
rect 42218 264931 42224 264943
rect 53296 264931 53302 264943
rect 53354 264931 53360 264983
rect 669808 264971 669814 264983
rect 53506 264943 669814 264971
rect 45712 264783 45718 264835
rect 45770 264823 45776 264835
rect 53506 264823 53534 264943
rect 669808 264931 669814 264943
rect 669866 264931 669872 264983
rect 669616 264897 669622 264909
rect 45770 264795 53534 264823
rect 54706 264869 669622 264897
rect 45770 264783 45776 264795
rect 46000 264709 46006 264761
rect 46058 264749 46064 264761
rect 54706 264749 54734 264869
rect 669616 264857 669622 264869
rect 669674 264857 669680 264909
rect 359440 264783 359446 264835
rect 359498 264823 359504 264835
rect 475984 264823 475990 264835
rect 359498 264795 475990 264823
rect 359498 264783 359504 264795
rect 475984 264783 475990 264795
rect 476042 264783 476048 264835
rect 46058 264721 54734 264749
rect 46058 264709 46064 264721
rect 328048 264709 328054 264761
rect 328106 264749 328112 264761
rect 440560 264749 440566 264761
rect 328106 264721 440566 264749
rect 328106 264709 328112 264721
rect 440560 264709 440566 264721
rect 440618 264709 440624 264761
rect 331120 264635 331126 264687
rect 331178 264675 331184 264687
rect 447664 264675 447670 264687
rect 331178 264647 447670 264675
rect 331178 264635 331184 264647
rect 447664 264635 447670 264647
rect 447722 264635 447728 264687
rect 354256 264561 354262 264613
rect 354314 264601 354320 264613
rect 461776 264601 461782 264613
rect 354314 264573 461782 264601
rect 354314 264561 354320 264573
rect 461776 264561 461782 264573
rect 461834 264561 461840 264613
rect 360400 264487 360406 264539
rect 360458 264527 360464 264539
rect 468880 264527 468886 264539
rect 360458 264499 468886 264527
rect 360458 264487 360464 264499
rect 468880 264487 468886 264499
rect 468938 264487 468944 264539
rect 351376 264413 351382 264465
rect 351434 264453 351440 264465
rect 454768 264453 454774 264465
rect 351434 264425 454774 264453
rect 351434 264413 351440 264425
rect 454768 264413 454774 264425
rect 454826 264413 454832 264465
rect 399376 264117 399382 264169
rect 399434 264157 399440 264169
rect 410992 264157 410998 264169
rect 399434 264129 410998 264157
rect 399434 264117 399440 264129
rect 410992 264117 410998 264129
rect 411050 264117 411056 264169
rect 267712 264043 267718 264095
rect 267770 264083 267776 264095
rect 276496 264083 276502 264095
rect 267770 264055 276502 264083
rect 267770 264043 267776 264055
rect 276496 264043 276502 264055
rect 276554 264043 276560 264095
rect 324976 264043 324982 264095
rect 325034 264083 325040 264095
rect 433456 264083 433462 264095
rect 325034 264055 433462 264083
rect 325034 264043 325040 264055
rect 433456 264043 433462 264055
rect 433514 264043 433520 264095
rect 387952 263969 387958 264021
rect 388010 264009 388016 264021
rect 589456 264009 589462 264021
rect 388010 263981 589462 264009
rect 388010 263969 388016 263981
rect 589456 263969 589462 263981
rect 589514 263969 589520 264021
rect 390832 263895 390838 263947
rect 390890 263935 390896 263947
rect 596560 263935 596566 263947
rect 390890 263907 596566 263935
rect 390890 263895 390896 263907
rect 596560 263895 596566 263907
rect 596618 263895 596624 263947
rect 393904 263821 393910 263873
rect 393962 263861 393968 263873
rect 603664 263861 603670 263873
rect 393962 263833 603670 263861
rect 393962 263821 393968 263833
rect 603664 263821 603670 263833
rect 603722 263821 603728 263873
rect 396784 263747 396790 263799
rect 396842 263787 396848 263799
rect 610768 263787 610774 263799
rect 396842 263759 610774 263787
rect 396842 263747 396848 263759
rect 610768 263747 610774 263759
rect 610826 263747 610832 263799
rect 401104 263673 401110 263725
rect 401162 263713 401168 263725
rect 401162 263685 410750 263713
rect 401162 263673 401168 263685
rect 23344 263599 23350 263651
rect 23402 263639 23408 263651
rect 43312 263639 43318 263651
rect 23402 263611 43318 263639
rect 23402 263599 23408 263611
rect 43312 263599 43318 263611
rect 43370 263639 43376 263651
rect 46000 263639 46006 263651
rect 43370 263611 46006 263639
rect 43370 263599 43376 263611
rect 46000 263599 46006 263611
rect 46058 263599 46064 263651
rect 403984 263599 403990 263651
rect 404042 263639 404048 263651
rect 410722 263639 410750 263685
rect 410992 263673 410998 263725
rect 411050 263713 411056 263725
rect 617872 263713 617878 263725
rect 411050 263685 617878 263713
rect 411050 263673 411056 263685
rect 617872 263673 617878 263685
rect 617930 263673 617936 263725
rect 621424 263639 621430 263651
rect 404042 263611 410654 263639
rect 410722 263611 621430 263639
rect 404042 263599 404048 263611
rect 23248 263525 23254 263577
rect 23306 263565 23312 263577
rect 43216 263565 43222 263577
rect 23306 263537 43222 263565
rect 23306 263525 23312 263537
rect 43216 263525 43222 263537
rect 43274 263565 43280 263577
rect 45712 263565 45718 263577
rect 43274 263537 45718 263565
rect 43274 263525 43280 263537
rect 45712 263525 45718 263537
rect 45770 263525 45776 263577
rect 409648 263525 409654 263577
rect 409706 263525 409712 263577
rect 410626 263565 410654 263611
rect 621424 263599 621430 263611
rect 621482 263599 621488 263651
rect 628432 263565 628438 263577
rect 410626 263537 628438 263565
rect 628432 263525 628438 263537
rect 628490 263525 628496 263577
rect 409666 263491 409694 263525
rect 642640 263491 642646 263503
rect 409666 263463 642646 263491
rect 642640 263451 642646 263463
rect 642698 263451 642704 263503
rect 23152 262119 23158 262171
rect 23210 262159 23216 262171
rect 43312 262159 43318 262171
rect 23210 262131 43318 262159
rect 23210 262119 23216 262131
rect 43312 262119 43318 262131
rect 43370 262119 43376 262171
rect 420400 262119 420406 262171
rect 420458 262159 420464 262171
rect 606160 262159 606166 262171
rect 420458 262131 606166 262159
rect 420458 262119 420464 262131
rect 606160 262119 606166 262131
rect 606218 262119 606224 262171
rect 674800 262119 674806 262171
rect 674858 262159 674864 262171
rect 676240 262159 676246 262171
rect 674858 262131 676246 262159
rect 674858 262119 674864 262131
rect 676240 262119 676246 262131
rect 676298 262119 676304 262171
rect 187216 260639 187222 260691
rect 187274 260679 187280 260691
rect 189712 260679 189718 260691
rect 187274 260651 189718 260679
rect 187274 260639 187280 260651
rect 189712 260639 189718 260651
rect 189770 260639 189776 260691
rect 674608 259381 674614 259433
rect 674666 259421 674672 259433
rect 676048 259421 676054 259433
rect 674666 259393 676054 259421
rect 674666 259381 674672 259393
rect 676048 259381 676054 259393
rect 676106 259381 676112 259433
rect 420400 259233 420406 259285
rect 420458 259273 420464 259285
rect 606256 259273 606262 259285
rect 420458 259245 606262 259273
rect 420458 259233 420464 259245
rect 606256 259233 606262 259245
rect 606314 259233 606320 259285
rect 675184 259233 675190 259285
rect 675242 259273 675248 259285
rect 676048 259273 676054 259285
rect 675242 259245 676054 259273
rect 675242 259233 675248 259245
rect 676048 259233 676054 259245
rect 676106 259233 676112 259285
rect 674512 256939 674518 256991
rect 674570 256979 674576 256991
rect 676048 256979 676054 256991
rect 674570 256951 676054 256979
rect 674570 256939 674576 256951
rect 676048 256939 676054 256951
rect 676106 256939 676112 256991
rect 674704 256421 674710 256473
rect 674762 256461 674768 256473
rect 676048 256461 676054 256473
rect 674762 256433 676054 256461
rect 674762 256421 674768 256433
rect 676048 256421 676054 256433
rect 676106 256421 676112 256473
rect 40240 256347 40246 256399
rect 40298 256387 40304 256399
rect 59056 256387 59062 256399
rect 40298 256359 59062 256387
rect 40298 256347 40304 256359
rect 59056 256347 59062 256359
rect 59114 256347 59120 256399
rect 420400 256347 420406 256399
rect 420458 256387 420464 256399
rect 606352 256387 606358 256399
rect 420458 256359 606358 256387
rect 420458 256347 420464 256359
rect 606352 256347 606358 256359
rect 606410 256347 606416 256399
rect 674992 256347 674998 256399
rect 675050 256387 675056 256399
rect 676240 256387 676246 256399
rect 675050 256359 676246 256387
rect 675050 256347 675056 256359
rect 676240 256347 676246 256359
rect 676298 256347 676304 256399
rect 41776 255385 41782 255437
rect 41834 255425 41840 255437
rect 53200 255425 53206 255437
rect 41834 255397 53206 255425
rect 41834 255385 41840 255397
rect 53200 255385 53206 255397
rect 53258 255385 53264 255437
rect 47920 255089 47926 255141
rect 47978 255129 47984 255141
rect 186256 255129 186262 255141
rect 47978 255101 186262 255129
rect 47978 255089 47984 255101
rect 186256 255089 186262 255101
rect 186314 255089 186320 255141
rect 47728 255015 47734 255067
rect 47786 255055 47792 255067
rect 186064 255055 186070 255067
rect 47786 255027 186070 255055
rect 47786 255015 47792 255027
rect 186064 255015 186070 255027
rect 186122 255015 186128 255067
rect 41776 254941 41782 254993
rect 41834 254981 41840 254993
rect 43408 254981 43414 254993
rect 41834 254953 43414 254981
rect 41834 254941 41840 254953
rect 43408 254941 43414 254953
rect 43466 254941 43472 254993
rect 47824 254941 47830 254993
rect 47882 254981 47888 254993
rect 186448 254981 186454 254993
rect 47882 254953 186454 254981
rect 47882 254941 47888 254953
rect 186448 254941 186454 254953
rect 186506 254941 186512 254993
rect 44848 254867 44854 254919
rect 44906 254907 44912 254919
rect 185968 254907 185974 254919
rect 44906 254879 185974 254907
rect 44906 254867 44912 254879
rect 185968 254867 185974 254879
rect 186026 254867 186032 254919
rect 41776 254423 41782 254475
rect 41834 254463 41840 254475
rect 43216 254463 43222 254475
rect 41834 254435 43222 254463
rect 41834 254423 41840 254435
rect 43216 254423 43222 254435
rect 43274 254423 43280 254475
rect 41584 253609 41590 253661
rect 41642 253649 41648 253661
rect 56176 253649 56182 253661
rect 41642 253621 56182 253649
rect 41642 253609 41648 253621
rect 56176 253609 56182 253621
rect 56234 253609 56240 253661
rect 674896 253535 674902 253587
rect 674954 253575 674960 253587
rect 676048 253575 676054 253587
rect 674954 253547 676054 253575
rect 674954 253535 674960 253547
rect 676048 253535 676054 253547
rect 676106 253535 676112 253587
rect 44944 253461 44950 253513
rect 45002 253501 45008 253513
rect 58960 253501 58966 253513
rect 45002 253473 58966 253501
rect 45002 253461 45008 253473
rect 58960 253461 58966 253473
rect 59018 253461 59024 253513
rect 420400 253461 420406 253513
rect 420458 253501 420464 253513
rect 603280 253501 603286 253513
rect 420458 253473 603286 253501
rect 420458 253461 420464 253473
rect 603280 253461 603286 253473
rect 603338 253461 603344 253513
rect 646672 253461 646678 253513
rect 646730 253501 646736 253513
rect 679696 253501 679702 253513
rect 646730 253473 679702 253501
rect 646730 253461 646736 253473
rect 679696 253461 679702 253473
rect 679754 253461 679760 253513
rect 106480 252277 106486 252329
rect 106538 252317 106544 252329
rect 156880 252317 156886 252329
rect 106538 252289 156886 252317
rect 106538 252277 106544 252289
rect 156880 252277 156886 252289
rect 156938 252277 156944 252329
rect 92080 252203 92086 252255
rect 92138 252243 92144 252255
rect 145360 252243 145366 252255
rect 92138 252215 145366 252243
rect 92138 252203 92144 252215
rect 145360 252203 145366 252215
rect 145418 252203 145424 252255
rect 109360 252129 109366 252181
rect 109418 252169 109424 252181
rect 171280 252169 171286 252181
rect 109418 252141 171286 252169
rect 109418 252129 109424 252141
rect 171280 252129 171286 252141
rect 171338 252129 171344 252181
rect 97840 252055 97846 252107
rect 97898 252095 97904 252107
rect 182800 252095 182806 252107
rect 97898 252067 182806 252095
rect 97898 252055 97904 252067
rect 182800 252055 182806 252067
rect 182858 252055 182864 252107
rect 56080 251981 56086 252033
rect 56138 252021 56144 252033
rect 186640 252021 186646 252033
rect 56138 251993 186646 252021
rect 56138 251981 56144 251993
rect 186640 251981 186646 251993
rect 186698 251981 186704 252033
rect 665872 250649 665878 250701
rect 665930 250689 665936 250701
rect 675376 250689 675382 250701
rect 665930 250661 675382 250689
rect 665930 250649 665936 250661
rect 675376 250649 675382 250661
rect 675434 250649 675440 250701
rect 420400 250575 420406 250627
rect 420458 250615 420464 250627
rect 603376 250615 603382 250627
rect 420458 250587 603382 250615
rect 420458 250575 420464 250587
rect 603376 250575 603382 250587
rect 603434 250575 603440 250627
rect 674800 250205 674806 250257
rect 674858 250245 674864 250257
rect 675280 250245 675286 250257
rect 674858 250217 675286 250245
rect 674858 250205 674864 250217
rect 675280 250205 675286 250217
rect 675338 250205 675344 250257
rect 120880 249909 120886 249961
rect 120938 249949 120944 249961
rect 145648 249949 145654 249961
rect 120938 249921 145654 249949
rect 120938 249909 120944 249921
rect 145648 249909 145654 249921
rect 145706 249909 145712 249961
rect 132400 249835 132406 249887
rect 132458 249875 132464 249887
rect 159856 249875 159862 249887
rect 132458 249847 159862 249875
rect 132458 249835 132464 249847
rect 159856 249835 159862 249847
rect 159914 249835 159920 249887
rect 135280 249761 135286 249813
rect 135338 249801 135344 249813
rect 168496 249801 168502 249813
rect 135338 249773 168502 249801
rect 135338 249761 135344 249773
rect 168496 249761 168502 249773
rect 168554 249761 168560 249813
rect 138160 249687 138166 249739
rect 138218 249727 138224 249739
rect 171472 249727 171478 249739
rect 138218 249699 171478 249727
rect 138218 249687 138224 249699
rect 171472 249687 171478 249699
rect 171530 249687 171536 249739
rect 141040 249613 141046 249665
rect 141098 249653 141104 249665
rect 180016 249653 180022 249665
rect 141098 249625 180022 249653
rect 141098 249613 141104 249625
rect 180016 249613 180022 249625
rect 180074 249613 180080 249665
rect 123760 249539 123766 249591
rect 123818 249579 123824 249591
rect 165712 249579 165718 249591
rect 123818 249551 165718 249579
rect 123818 249539 123824 249551
rect 165712 249539 165718 249551
rect 165770 249539 165776 249591
rect 126640 249465 126646 249517
rect 126698 249505 126704 249517
rect 177040 249505 177046 249517
rect 126698 249477 177046 249505
rect 126698 249465 126704 249477
rect 177040 249465 177046 249477
rect 177098 249465 177104 249517
rect 94960 249391 94966 249443
rect 95018 249431 95024 249443
rect 154000 249431 154006 249443
rect 95018 249403 154006 249431
rect 95018 249391 95024 249403
rect 154000 249391 154006 249403
rect 154058 249391 154064 249443
rect 118000 249317 118006 249369
rect 118058 249357 118064 249369
rect 182896 249357 182902 249369
rect 118058 249329 182902 249357
rect 118058 249317 118064 249329
rect 182896 249317 182902 249329
rect 182954 249317 182960 249369
rect 77680 249243 77686 249295
rect 77738 249283 77744 249295
rect 145456 249283 145462 249295
rect 77738 249255 145462 249283
rect 77738 249243 77744 249255
rect 145456 249243 145462 249255
rect 145514 249243 145520 249295
rect 80560 249169 80566 249221
rect 80618 249209 80624 249221
rect 162640 249209 162646 249221
rect 80618 249181 162646 249209
rect 80618 249169 80624 249181
rect 162640 249169 162646 249181
rect 162698 249169 162704 249221
rect 86320 249095 86326 249147
rect 86378 249135 86384 249147
rect 174160 249135 174166 249147
rect 86378 249107 174166 249135
rect 86378 249095 86384 249107
rect 174160 249095 174166 249107
rect 174218 249095 174224 249147
rect 674608 249095 674614 249147
rect 674666 249135 674672 249147
rect 675280 249135 675286 249147
rect 674666 249107 675286 249135
rect 674666 249095 674672 249107
rect 675280 249095 675286 249107
rect 675338 249095 675344 249147
rect 41872 247837 41878 247889
rect 41930 247877 41936 247889
rect 42832 247877 42838 247889
rect 41930 247849 42838 247877
rect 41930 247837 41936 247849
rect 42832 247837 42838 247849
rect 42890 247837 42896 247889
rect 420304 247763 420310 247815
rect 420362 247803 420368 247815
rect 603472 247803 603478 247815
rect 420362 247775 603478 247803
rect 420362 247763 420368 247775
rect 603472 247763 603478 247775
rect 603530 247763 603536 247815
rect 420400 247689 420406 247741
rect 420458 247729 420464 247741
rect 629200 247729 629206 247741
rect 420458 247701 629206 247729
rect 420458 247689 420464 247701
rect 629200 247689 629206 247701
rect 629258 247689 629264 247741
rect 655888 247615 655894 247667
rect 655946 247655 655952 247667
rect 665872 247655 665878 247667
rect 655946 247627 665878 247655
rect 655946 247615 655952 247627
rect 665872 247615 665878 247627
rect 665930 247615 665936 247667
rect 674512 247467 674518 247519
rect 674570 247507 674576 247519
rect 675088 247507 675094 247519
rect 674570 247479 675094 247507
rect 674570 247467 674576 247479
rect 675088 247467 675094 247479
rect 675146 247467 675152 247519
rect 103600 246727 103606 246779
rect 103658 246767 103664 246779
rect 165520 246767 165526 246779
rect 103658 246739 165526 246767
rect 103658 246727 103664 246739
rect 165520 246727 165526 246739
rect 165578 246727 165584 246779
rect 112240 246653 112246 246705
rect 112298 246693 112304 246705
rect 185776 246693 185782 246705
rect 112298 246665 185782 246693
rect 112298 246653 112304 246665
rect 185776 246653 185782 246665
rect 185834 246653 185840 246705
rect 47536 246579 47542 246631
rect 47594 246619 47600 246631
rect 186352 246619 186358 246631
rect 47594 246591 186358 246619
rect 47594 246579 47600 246591
rect 186352 246579 186358 246591
rect 186410 246579 186416 246631
rect 47440 246505 47446 246557
rect 47498 246545 47504 246557
rect 186544 246545 186550 246557
rect 47498 246517 186550 246545
rect 47498 246505 47504 246517
rect 186544 246505 186550 246517
rect 186602 246505 186608 246557
rect 47632 246431 47638 246483
rect 47690 246471 47696 246483
rect 186736 246471 186742 246483
rect 47690 246443 186742 246471
rect 47690 246431 47696 246443
rect 186736 246431 186742 246443
rect 186794 246431 186800 246483
rect 45520 246357 45526 246409
rect 45578 246397 45584 246409
rect 186832 246397 186838 246409
rect 45578 246369 186838 246397
rect 45578 246357 45584 246369
rect 186832 246357 186838 246369
rect 186890 246357 186896 246409
rect 44560 246283 44566 246335
rect 44618 246323 44624 246335
rect 186160 246323 186166 246335
rect 44618 246295 186166 246323
rect 44618 246283 44624 246295
rect 186160 246283 186166 246295
rect 186218 246283 186224 246335
rect 45232 246209 45238 246261
rect 45290 246249 45296 246261
rect 187024 246249 187030 246261
rect 45290 246221 187030 246249
rect 45290 246209 45296 246221
rect 187024 246209 187030 246221
rect 187082 246209 187088 246261
rect 41584 245099 41590 245151
rect 41642 245139 41648 245151
rect 145744 245139 145750 245151
rect 41642 245111 145750 245139
rect 41642 245099 41648 245111
rect 145744 245099 145750 245111
rect 145802 245099 145808 245151
rect 41584 244951 41590 245003
rect 41642 244991 41648 245003
rect 145552 244991 145558 245003
rect 41642 244963 145558 244991
rect 41642 244951 41648 244963
rect 145552 244951 145558 244963
rect 145610 244951 145616 245003
rect 44752 244877 44758 244929
rect 44810 244917 44816 244929
rect 186928 244917 186934 244929
rect 44810 244889 186934 244917
rect 44810 244877 44816 244889
rect 186928 244877 186934 244889
rect 186986 244877 186992 244929
rect 420400 244803 420406 244855
rect 420458 244843 420464 244855
rect 629296 244843 629302 244855
rect 420458 244815 629302 244843
rect 420458 244803 420464 244815
rect 629296 244803 629302 244815
rect 629354 244803 629360 244855
rect 40240 244729 40246 244781
rect 40298 244769 40304 244781
rect 42448 244769 42454 244781
rect 40298 244741 42454 244769
rect 40298 244729 40304 244741
rect 42448 244729 42454 244741
rect 42506 244729 42512 244781
rect 41488 244655 41494 244707
rect 41546 244695 41552 244707
rect 42640 244695 42646 244707
rect 41546 244667 42646 244695
rect 41546 244655 41552 244667
rect 42640 244655 42646 244667
rect 42698 244655 42704 244707
rect 34480 243545 34486 243597
rect 34538 243585 34544 243597
rect 42352 243585 42358 243597
rect 34538 243557 42358 243585
rect 34538 243545 34544 243557
rect 42352 243545 42358 243557
rect 42410 243545 42416 243597
rect 41680 243175 41686 243227
rect 41738 243215 41744 243227
rect 42928 243215 42934 243227
rect 41738 243187 42934 243215
rect 41738 243175 41744 243187
rect 42928 243175 42934 243187
rect 42986 243175 42992 243227
rect 44656 242805 44662 242857
rect 44714 242845 44720 242857
rect 185584 242845 185590 242857
rect 44714 242817 185590 242845
rect 44714 242805 44720 242817
rect 185584 242805 185590 242817
rect 185642 242805 185648 242857
rect 44848 242731 44854 242783
rect 44906 242771 44912 242783
rect 185872 242771 185878 242783
rect 44906 242743 185878 242771
rect 44906 242731 44912 242743
rect 185872 242731 185878 242743
rect 185930 242731 185936 242783
rect 674704 242731 674710 242783
rect 674762 242771 674768 242783
rect 675376 242771 675382 242783
rect 674762 242743 675382 242771
rect 674762 242731 674768 242743
rect 675376 242731 675382 242743
rect 675434 242731 675440 242783
rect 44560 242657 44566 242709
rect 44618 242697 44624 242709
rect 185680 242697 185686 242709
rect 44618 242669 185686 242697
rect 44618 242657 44624 242669
rect 185680 242657 185686 242669
rect 185738 242657 185744 242709
rect 41584 242583 41590 242635
rect 41642 242623 41648 242635
rect 142576 242623 142582 242635
rect 41642 242595 142582 242623
rect 41642 242583 41648 242595
rect 142576 242583 142582 242595
rect 142634 242583 142640 242635
rect 41872 241917 41878 241969
rect 41930 241957 41936 241969
rect 43120 241957 43126 241969
rect 41930 241929 43126 241957
rect 41930 241917 41936 241929
rect 43120 241917 43126 241929
rect 43178 241917 43184 241969
rect 420400 241917 420406 241969
rect 420458 241957 420464 241969
rect 600400 241957 600406 241969
rect 420458 241929 600406 241957
rect 420458 241917 420464 241929
rect 600400 241917 600406 241929
rect 600458 241917 600464 241969
rect 41776 240585 41782 240637
rect 41834 240585 41840 240637
rect 41794 240415 41822 240585
rect 41776 240363 41782 240415
rect 41834 240363 41840 240415
rect 380848 239919 380854 239971
rect 380906 239959 380912 239971
rect 412048 239959 412054 239971
rect 380906 239931 412054 239959
rect 380906 239919 380912 239931
rect 412048 239919 412054 239931
rect 412106 239919 412112 239971
rect 409552 239845 409558 239897
rect 409610 239885 409616 239897
rect 412144 239885 412150 239897
rect 409610 239857 412150 239885
rect 409610 239845 409616 239857
rect 412144 239845 412150 239857
rect 412202 239845 412208 239897
rect 357136 239771 357142 239823
rect 357194 239811 357200 239823
rect 434608 239811 434614 239823
rect 357194 239783 434614 239811
rect 357194 239771 357200 239783
rect 434608 239771 434614 239783
rect 434666 239771 434672 239823
rect 377296 239697 377302 239749
rect 377354 239737 377360 239749
rect 446704 239737 446710 239749
rect 377354 239709 446710 239737
rect 377354 239697 377360 239709
rect 446704 239697 446710 239709
rect 446762 239697 446768 239749
rect 385360 239623 385366 239675
rect 385418 239663 385424 239675
rect 470896 239663 470902 239675
rect 385418 239635 470902 239663
rect 385418 239623 385424 239635
rect 470896 239623 470902 239635
rect 470954 239623 470960 239675
rect 374416 239549 374422 239601
rect 374474 239589 374480 239601
rect 488272 239589 488278 239601
rect 374474 239561 488278 239589
rect 374474 239549 374480 239561
rect 488272 239549 488278 239561
rect 488330 239549 488336 239601
rect 334288 239475 334294 239527
rect 334346 239515 334352 239527
rect 458800 239515 458806 239527
rect 334346 239487 458806 239515
rect 334346 239475 334352 239487
rect 458800 239475 458806 239487
rect 458858 239475 458864 239527
rect 394672 239401 394678 239453
rect 394730 239441 394736 239453
rect 532816 239441 532822 239453
rect 394730 239413 532822 239441
rect 394730 239401 394736 239413
rect 532816 239401 532822 239413
rect 532874 239401 532880 239453
rect 397936 239327 397942 239379
rect 397994 239367 398000 239379
rect 541456 239367 541462 239379
rect 397994 239339 541462 239367
rect 397994 239327 398000 239339
rect 541456 239327 541462 239339
rect 541514 239327 541520 239379
rect 406000 239253 406006 239305
rect 406058 239293 406064 239305
rect 550864 239293 550870 239305
rect 406058 239265 550870 239293
rect 406058 239253 406064 239265
rect 550864 239253 550870 239265
rect 550922 239253 550928 239305
rect 420400 239179 420406 239231
rect 420458 239219 420464 239231
rect 599152 239219 599158 239231
rect 420458 239191 599158 239219
rect 420458 239179 420464 239191
rect 599152 239179 599158 239191
rect 599210 239179 599216 239231
rect 350416 239105 350422 239157
rect 350474 239145 350480 239157
rect 508624 239145 508630 239157
rect 350474 239117 508630 239145
rect 350474 239105 350480 239117
rect 508624 239105 508630 239117
rect 508682 239105 508688 239157
rect 368560 239031 368566 239083
rect 368618 239071 368624 239083
rect 544816 239071 544822 239083
rect 368618 239043 544822 239071
rect 368618 239031 368624 239043
rect 544816 239031 544822 239043
rect 544874 239031 544880 239083
rect 324400 238957 324406 239009
rect 324458 238997 324464 239009
rect 455152 238997 455158 239009
rect 324458 238969 455158 238997
rect 324458 238957 324464 238969
rect 455152 238957 455158 238969
rect 455210 238957 455216 239009
rect 323920 238883 323926 238935
rect 323978 238923 323984 238935
rect 455056 238923 455062 238935
rect 323978 238895 455062 238923
rect 323978 238883 323984 238895
rect 455056 238883 455062 238895
rect 455114 238883 455120 238935
rect 326704 238809 326710 238861
rect 326762 238849 326768 238861
rect 462544 238849 462550 238861
rect 326762 238821 462550 238849
rect 326762 238809 326768 238821
rect 462544 238809 462550 238821
rect 462602 238809 462608 238861
rect 328912 238735 328918 238787
rect 328970 238775 328976 238787
rect 464752 238775 464758 238787
rect 328970 238747 464758 238775
rect 328970 238735 328976 238747
rect 464752 238735 464758 238747
rect 464810 238735 464816 238787
rect 329872 238661 329878 238713
rect 329930 238701 329936 238713
rect 468592 238701 468598 238713
rect 329930 238673 468598 238701
rect 329930 238661 329936 238673
rect 468592 238661 468598 238673
rect 468650 238661 468656 238713
rect 332656 238587 332662 238639
rect 332714 238627 332720 238639
rect 474640 238627 474646 238639
rect 332714 238599 474646 238627
rect 332714 238587 332720 238599
rect 474640 238587 474646 238599
rect 474698 238587 474704 238639
rect 42160 238513 42166 238565
rect 42218 238553 42224 238565
rect 42448 238553 42454 238565
rect 42218 238525 42454 238553
rect 42218 238513 42224 238525
rect 42448 238513 42454 238525
rect 42506 238513 42512 238565
rect 335728 238513 335734 238565
rect 335786 238553 335792 238565
rect 480688 238553 480694 238565
rect 335786 238525 480694 238553
rect 335786 238513 335792 238525
rect 480688 238513 480694 238525
rect 480746 238513 480752 238565
rect 336688 238439 336694 238491
rect 336746 238479 336752 238491
rect 478096 238479 478102 238491
rect 336746 238451 478102 238479
rect 336746 238439 336752 238451
rect 478096 238439 478102 238451
rect 478154 238439 478160 238491
rect 42544 238365 42550 238417
rect 42602 238365 42608 238417
rect 338992 238365 338998 238417
rect 339050 238405 339056 238417
rect 486736 238405 486742 238417
rect 339050 238377 486742 238405
rect 339050 238365 339056 238377
rect 486736 238365 486742 238377
rect 486794 238365 486800 238417
rect 42562 238121 42590 238365
rect 341776 238291 341782 238343
rect 341834 238331 341840 238343
rect 492784 238331 492790 238343
rect 341834 238303 492790 238331
rect 341834 238291 341840 238303
rect 492784 238291 492790 238303
rect 492842 238291 492848 238343
rect 345328 238217 345334 238269
rect 345386 238257 345392 238269
rect 500272 238257 500278 238269
rect 345386 238229 500278 238257
rect 345386 238217 345392 238229
rect 500272 238217 500278 238229
rect 500330 238217 500336 238269
rect 346672 238143 346678 238195
rect 346730 238183 346736 238195
rect 503344 238183 503350 238195
rect 346730 238155 503350 238183
rect 346730 238143 346736 238155
rect 503344 238143 503350 238155
rect 503402 238143 503408 238195
rect 42544 238069 42550 238121
rect 42602 238069 42608 238121
rect 349936 238069 349942 238121
rect 349994 238109 350000 238121
rect 509392 238109 509398 238121
rect 349994 238081 509398 238109
rect 349994 238069 350000 238081
rect 509392 238069 509398 238081
rect 509450 238069 509456 238121
rect 353488 237995 353494 238047
rect 353546 238035 353552 238047
rect 514672 238035 514678 238047
rect 353546 238007 514678 238035
rect 353546 237995 353552 238007
rect 514672 237995 514678 238007
rect 514730 237995 514736 238047
rect 352720 237921 352726 237973
rect 352778 237961 352784 237973
rect 512752 237961 512758 237973
rect 352778 237933 512758 237961
rect 352778 237921 352784 237933
rect 512752 237921 512758 237933
rect 512810 237921 512816 237973
rect 355696 237847 355702 237899
rect 355754 237887 355760 237899
rect 522160 237887 522166 237899
rect 355754 237859 522166 237887
rect 355754 237847 355760 237859
rect 522160 237847 522166 237859
rect 522218 237847 522224 237899
rect 363088 237773 363094 237825
rect 363146 237813 363152 237825
rect 535120 237813 535126 237825
rect 363146 237785 535126 237813
rect 363146 237773 363152 237785
rect 535120 237773 535126 237785
rect 535178 237773 535184 237825
rect 275344 237699 275350 237751
rect 275402 237739 275408 237751
rect 357520 237739 357526 237751
rect 275402 237711 357526 237739
rect 275402 237699 275408 237711
rect 357520 237699 357526 237711
rect 357578 237699 357584 237751
rect 361744 237699 361750 237751
rect 361802 237739 361808 237751
rect 533488 237739 533494 237751
rect 361802 237711 533494 237739
rect 361802 237699 361808 237711
rect 533488 237699 533494 237711
rect 533546 237699 533552 237751
rect 277072 237625 277078 237677
rect 277130 237665 277136 237677
rect 363664 237665 363670 237677
rect 277130 237637 363670 237665
rect 277130 237625 277136 237637
rect 363664 237625 363670 237637
rect 363722 237625 363728 237677
rect 364432 237625 364438 237677
rect 364490 237665 364496 237677
rect 535792 237665 535798 237677
rect 364490 237637 535798 237665
rect 364490 237625 364496 237637
rect 535792 237625 535798 237637
rect 535850 237625 535856 237677
rect 365872 237551 365878 237603
rect 365930 237591 365936 237603
rect 541072 237591 541078 237603
rect 365930 237563 541078 237591
rect 365930 237551 365936 237563
rect 541072 237551 541078 237563
rect 541130 237551 541136 237603
rect 320848 237477 320854 237529
rect 320906 237517 320912 237529
rect 450448 237517 450454 237529
rect 320906 237489 450454 237517
rect 320906 237477 320912 237489
rect 450448 237477 450454 237489
rect 450506 237477 450512 237529
rect 317584 237403 317590 237455
rect 317642 237443 317648 237455
rect 444496 237443 444502 237455
rect 317642 237415 444502 237443
rect 317642 237403 317648 237415
rect 444496 237403 444502 237415
rect 444554 237403 444560 237455
rect 317104 237329 317110 237381
rect 317162 237369 317168 237381
rect 440656 237369 440662 237381
rect 317162 237341 440662 237369
rect 317162 237329 317168 237341
rect 440656 237329 440662 237341
rect 440714 237329 440720 237381
rect 314800 237255 314806 237307
rect 314858 237295 314864 237307
rect 438352 237295 438358 237307
rect 314858 237267 438358 237295
rect 314858 237255 314864 237267
rect 438352 237255 438358 237267
rect 438410 237255 438416 237307
rect 311536 237181 311542 237233
rect 311594 237221 311600 237233
rect 432400 237221 432406 237233
rect 311594 237193 432406 237221
rect 311594 237181 311600 237193
rect 432400 237181 432406 237193
rect 432458 237181 432464 237233
rect 308560 237107 308566 237159
rect 308618 237147 308624 237159
rect 426352 237147 426358 237159
rect 308618 237119 426358 237147
rect 308618 237107 308624 237119
rect 426352 237107 426358 237119
rect 426410 237107 426416 237159
rect 310768 237033 310774 237085
rect 310826 237073 310832 237085
rect 428656 237073 428662 237085
rect 310826 237045 428662 237073
rect 310826 237033 310832 237045
rect 428656 237033 428662 237045
rect 428714 237033 428720 237085
rect 305776 236959 305782 237011
rect 305834 236999 305840 237011
rect 420304 236999 420310 237011
rect 305834 236971 420310 236999
rect 305834 236959 305840 236971
rect 420304 236959 420310 236971
rect 420362 236959 420368 237011
rect 298960 236885 298966 236937
rect 299018 236925 299024 236937
rect 404464 236925 404470 236937
rect 299018 236897 404470 236925
rect 299018 236885 299024 236897
rect 404464 236885 404470 236897
rect 404522 236885 404528 236937
rect 405904 236885 405910 236937
rect 405962 236925 405968 236937
rect 414448 236925 414454 236937
rect 405962 236897 414454 236925
rect 405962 236885 405968 236897
rect 414448 236885 414454 236897
rect 414506 236885 414512 236937
rect 279856 236811 279862 236863
rect 279914 236851 279920 236863
rect 370480 236851 370486 236863
rect 279914 236823 370486 236851
rect 279914 236811 279920 236823
rect 370480 236811 370486 236823
rect 370538 236811 370544 236863
rect 386992 236811 386998 236863
rect 387050 236851 387056 236863
rect 387568 236851 387574 236863
rect 387050 236823 387574 236851
rect 387050 236811 387056 236823
rect 387568 236811 387574 236823
rect 387626 236811 387632 236863
rect 397840 236811 397846 236863
rect 397898 236851 397904 236863
rect 413584 236851 413590 236863
rect 397898 236823 413590 236851
rect 397898 236811 397904 236823
rect 413584 236811 413590 236823
rect 413642 236811 413648 236863
rect 278416 236737 278422 236789
rect 278474 236777 278480 236789
rect 366736 236777 366742 236789
rect 278474 236749 366742 236777
rect 278474 236737 278480 236749
rect 366736 236737 366742 236749
rect 366794 236737 366800 236789
rect 382384 236737 382390 236789
rect 382442 236777 382448 236789
rect 398032 236777 398038 236789
rect 382442 236749 398038 236777
rect 382442 236737 382448 236749
rect 398032 236737 398038 236749
rect 398090 236737 398096 236789
rect 397072 236663 397078 236715
rect 397130 236703 397136 236715
rect 397744 236703 397750 236715
rect 397130 236675 397750 236703
rect 397130 236663 397136 236675
rect 397744 236663 397750 236675
rect 397802 236663 397808 236715
rect 397456 236589 397462 236641
rect 397514 236629 397520 236641
rect 413392 236629 413398 236641
rect 397514 236601 413398 236629
rect 397514 236589 397520 236601
rect 413392 236589 413398 236601
rect 413450 236589 413456 236641
rect 387184 236515 387190 236567
rect 387242 236555 387248 236567
rect 387856 236555 387862 236567
rect 387242 236527 387862 236555
rect 387242 236515 387248 236527
rect 387856 236515 387862 236527
rect 387914 236515 387920 236567
rect 397456 236441 397462 236493
rect 397514 236481 397520 236493
rect 397936 236481 397942 236493
rect 397514 236453 397942 236481
rect 397514 236441 397520 236453
rect 397936 236441 397942 236453
rect 397994 236441 398000 236493
rect 378160 236367 378166 236419
rect 378218 236407 378224 236419
rect 397360 236407 397366 236419
rect 378218 236379 397366 236407
rect 378218 236367 378224 236379
rect 397360 236367 397366 236379
rect 397418 236367 397424 236419
rect 410704 236367 410710 236419
rect 410762 236407 410768 236419
rect 442192 236407 442198 236419
rect 410762 236379 442198 236407
rect 410762 236367 410768 236379
rect 442192 236367 442198 236379
rect 442250 236367 442256 236419
rect 387088 236293 387094 236345
rect 387146 236333 387152 236345
rect 387472 236333 387478 236345
rect 387146 236305 387478 236333
rect 387146 236293 387152 236305
rect 387472 236293 387478 236305
rect 387530 236293 387536 236345
rect 390736 236293 390742 236345
rect 390794 236333 390800 236345
rect 492016 236333 492022 236345
rect 390794 236305 492022 236333
rect 390794 236293 390800 236305
rect 492016 236293 492022 236305
rect 492074 236293 492080 236345
rect 394576 236219 394582 236271
rect 394634 236259 394640 236271
rect 505648 236259 505654 236271
rect 394634 236231 505654 236259
rect 394634 236219 394640 236231
rect 505648 236219 505654 236231
rect 505706 236219 505712 236271
rect 400336 236145 400342 236197
rect 400394 236185 400400 236197
rect 523792 236185 523798 236197
rect 400394 236157 523798 236185
rect 400394 236145 400400 236157
rect 523792 236145 523798 236157
rect 523850 236145 523856 236197
rect 251056 236071 251062 236123
rect 251114 236111 251120 236123
rect 273616 236111 273622 236123
rect 251114 236083 273622 236111
rect 251114 236071 251120 236083
rect 273616 236071 273622 236083
rect 273674 236071 273680 236123
rect 277552 236071 277558 236123
rect 277610 236111 277616 236123
rect 313936 236111 313942 236123
rect 277610 236083 313942 236111
rect 277610 236071 277616 236083
rect 313936 236071 313942 236083
rect 313994 236071 314000 236123
rect 326128 236071 326134 236123
rect 326186 236111 326192 236123
rect 334288 236111 334294 236123
rect 326186 236083 334294 236111
rect 326186 236071 326192 236083
rect 334288 236071 334294 236083
rect 334346 236071 334352 236123
rect 341200 236071 341206 236123
rect 341258 236111 341264 236123
rect 374416 236111 374422 236123
rect 341258 236083 374422 236111
rect 341258 236071 341264 236083
rect 374416 236071 374422 236083
rect 374474 236071 374480 236123
rect 376336 236071 376342 236123
rect 376394 236111 376400 236123
rect 376394 236083 406142 236111
rect 376394 236071 376400 236083
rect 208432 235997 208438 236049
rect 208490 236037 208496 236049
rect 223216 236037 223222 236049
rect 208490 236009 223222 236037
rect 208490 235997 208496 236009
rect 223216 235997 223222 236009
rect 223274 235997 223280 236049
rect 247984 235997 247990 236049
rect 248042 236037 248048 236049
rect 248042 236009 271166 236037
rect 248042 235997 248048 236009
rect 209680 235923 209686 235975
rect 209738 235963 209744 235975
rect 226192 235963 226198 235975
rect 209738 235935 226198 235963
rect 209738 235923 209744 235935
rect 226192 235923 226198 235935
rect 226250 235923 226256 235975
rect 243280 235923 243286 235975
rect 243338 235963 243344 235975
rect 271024 235963 271030 235975
rect 243338 235935 271030 235963
rect 243338 235923 243344 235935
rect 271024 235923 271030 235935
rect 271082 235923 271088 235975
rect 271138 235963 271166 236009
rect 276112 235997 276118 236049
rect 276170 236037 276176 236049
rect 310192 236037 310198 236049
rect 276170 236009 310198 236037
rect 276170 235997 276176 236009
rect 310192 235997 310198 236009
rect 310250 235997 310256 236049
rect 313840 235997 313846 236049
rect 313898 236037 313904 236049
rect 357136 236037 357142 236049
rect 313898 236009 357142 236037
rect 313898 235997 313904 236009
rect 357136 235997 357142 236009
rect 357194 235997 357200 236049
rect 371824 235997 371830 236049
rect 371882 236037 371888 236049
rect 406000 236037 406006 236049
rect 371882 236009 406006 236037
rect 371882 235997 371888 236009
rect 406000 235997 406006 236009
rect 406058 235997 406064 236049
rect 276208 235963 276214 235975
rect 271138 235935 276214 235963
rect 276208 235923 276214 235935
rect 276266 235923 276272 235975
rect 280624 235923 280630 235975
rect 280682 235963 280688 235975
rect 322000 235963 322006 235975
rect 280682 235935 322006 235963
rect 280682 235923 280688 235935
rect 322000 235923 322006 235935
rect 322058 235923 322064 235975
rect 386704 235923 386710 235975
rect 386762 235963 386768 235975
rect 405616 235963 405622 235975
rect 386762 235935 405622 235963
rect 386762 235923 386768 235935
rect 405616 235923 405622 235935
rect 405674 235923 405680 235975
rect 406114 235963 406142 236083
rect 410032 236071 410038 236123
rect 410090 236111 410096 236123
rect 584560 236111 584566 236123
rect 410090 236083 584566 236111
rect 410090 236071 410096 236083
rect 584560 236071 584566 236083
rect 584618 236071 584624 236123
rect 406288 235997 406294 236049
rect 406346 236037 406352 236049
rect 415408 236037 415414 236049
rect 406346 236009 415414 236037
rect 406346 235997 406352 236009
rect 415408 235997 415414 236009
rect 415466 235997 415472 236049
rect 413872 235963 413878 235975
rect 406114 235935 413878 235963
rect 413872 235923 413878 235935
rect 413930 235923 413936 235975
rect 208912 235849 208918 235901
rect 208970 235889 208976 235901
rect 226960 235889 226966 235901
rect 208970 235861 226966 235889
rect 208970 235849 208976 235861
rect 226960 235849 226966 235861
rect 227018 235849 227024 235901
rect 234256 235849 234262 235901
rect 234314 235889 234320 235901
rect 264688 235889 264694 235901
rect 234314 235861 264694 235889
rect 234314 235849 234320 235861
rect 264688 235849 264694 235861
rect 264746 235849 264752 235901
rect 279280 235849 279286 235901
rect 279338 235889 279344 235901
rect 318256 235889 318262 235901
rect 279338 235861 318262 235889
rect 279338 235849 279344 235861
rect 318256 235849 318262 235861
rect 318314 235849 318320 235901
rect 326224 235849 326230 235901
rect 326282 235889 326288 235901
rect 460240 235889 460246 235901
rect 326282 235861 460246 235889
rect 326282 235849 326288 235861
rect 460240 235849 460246 235861
rect 460298 235849 460304 235901
rect 208816 235775 208822 235827
rect 208874 235815 208880 235827
rect 224752 235815 224758 235827
rect 208874 235787 224758 235815
rect 208874 235775 208880 235787
rect 224752 235775 224758 235787
rect 224810 235775 224816 235827
rect 237520 235775 237526 235827
rect 237578 235815 237584 235827
rect 268144 235815 268150 235827
rect 237578 235787 268150 235815
rect 237578 235775 237584 235787
rect 268144 235775 268150 235787
rect 268202 235775 268208 235827
rect 290320 235775 290326 235827
rect 290378 235815 290384 235827
rect 334096 235815 334102 235827
rect 290378 235787 334102 235815
rect 290378 235775 290384 235787
rect 334096 235775 334102 235787
rect 334154 235775 334160 235827
rect 343504 235775 343510 235827
rect 343562 235815 343568 235827
rect 495760 235815 495766 235827
rect 343562 235787 495766 235815
rect 343562 235775 343568 235787
rect 495760 235775 495766 235787
rect 495818 235775 495824 235827
rect 211216 235701 211222 235753
rect 211274 235741 211280 235753
rect 229264 235741 229270 235753
rect 211274 235713 229270 235741
rect 211274 235701 211280 235713
rect 229264 235701 229270 235713
rect 229322 235701 229328 235753
rect 231184 235701 231190 235753
rect 231242 235741 231248 235753
rect 259024 235741 259030 235753
rect 231242 235713 259030 235741
rect 231242 235701 231248 235713
rect 259024 235701 259030 235713
rect 259082 235701 259088 235753
rect 262864 235701 262870 235753
rect 262922 235741 262928 235753
rect 305008 235741 305014 235753
rect 262922 235713 305014 235741
rect 262922 235701 262928 235713
rect 305008 235701 305014 235713
rect 305066 235701 305072 235753
rect 317200 235701 317206 235753
rect 317258 235741 317264 235753
rect 410704 235741 410710 235753
rect 317258 235713 410710 235741
rect 317258 235701 317264 235713
rect 410704 235701 410710 235713
rect 410762 235701 410768 235753
rect 411856 235701 411862 235753
rect 411914 235741 411920 235753
rect 413680 235741 413686 235753
rect 411914 235713 413686 235741
rect 411914 235701 411920 235713
rect 413680 235701 413686 235713
rect 413738 235701 413744 235753
rect 210640 235627 210646 235679
rect 210698 235667 210704 235679
rect 230032 235667 230038 235679
rect 210698 235639 230038 235667
rect 210698 235627 210704 235639
rect 230032 235627 230038 235639
rect 230090 235627 230096 235679
rect 239344 235627 239350 235679
rect 239402 235667 239408 235679
rect 239402 235639 287006 235667
rect 239402 235627 239408 235639
rect 210064 235553 210070 235605
rect 210122 235593 210128 235605
rect 227824 235593 227830 235605
rect 210122 235565 227830 235593
rect 210122 235553 210128 235565
rect 227824 235553 227830 235565
rect 227882 235553 227888 235605
rect 236464 235553 236470 235605
rect 236522 235593 236528 235605
rect 282928 235593 282934 235605
rect 236522 235565 282934 235593
rect 236522 235553 236528 235565
rect 282928 235553 282934 235565
rect 282986 235553 282992 235605
rect 286978 235593 287006 235639
rect 287056 235627 287062 235679
rect 287114 235667 287120 235679
rect 318448 235667 318454 235679
rect 287114 235639 318454 235667
rect 287114 235627 287120 235639
rect 318448 235627 318454 235639
rect 318506 235627 318512 235679
rect 358000 235627 358006 235679
rect 358058 235667 358064 235679
rect 400336 235667 400342 235679
rect 358058 235639 400342 235667
rect 358058 235627 358064 235639
rect 400336 235627 400342 235639
rect 400394 235627 400400 235679
rect 408976 235667 408982 235679
rect 405538 235639 408982 235667
rect 287344 235593 287350 235605
rect 286978 235565 287350 235593
rect 287344 235553 287350 235565
rect 287402 235553 287408 235605
rect 311152 235553 311158 235605
rect 311210 235593 311216 235605
rect 405538 235593 405566 235639
rect 408976 235627 408982 235639
rect 409034 235627 409040 235679
rect 409168 235627 409174 235679
rect 409226 235667 409232 235679
rect 588880 235667 588886 235679
rect 409226 235639 588886 235667
rect 409226 235627 409232 235639
rect 588880 235627 588886 235639
rect 588938 235627 588944 235679
rect 311210 235565 405566 235593
rect 311210 235553 311216 235565
rect 405616 235553 405622 235605
rect 405674 235593 405680 235605
rect 411856 235593 411862 235605
rect 405674 235565 411862 235593
rect 405674 235553 405680 235565
rect 411856 235553 411862 235565
rect 411914 235553 411920 235605
rect 412144 235553 412150 235605
rect 412202 235593 412208 235605
rect 590512 235593 590518 235605
rect 412202 235565 590518 235593
rect 412202 235553 412208 235565
rect 590512 235553 590518 235565
rect 590570 235553 590576 235605
rect 212944 235479 212950 235531
rect 213002 235519 213008 235531
rect 232336 235519 232342 235531
rect 213002 235491 232342 235519
rect 213002 235479 213008 235491
rect 232336 235479 232342 235491
rect 232394 235479 232400 235531
rect 238000 235479 238006 235531
rect 238058 235519 238064 235531
rect 285904 235519 285910 235531
rect 238058 235491 285910 235519
rect 238058 235479 238064 235491
rect 285904 235479 285910 235491
rect 285962 235479 285968 235531
rect 299824 235479 299830 235531
rect 299882 235519 299888 235531
rect 354256 235519 354262 235531
rect 299882 235491 354262 235519
rect 299882 235479 299888 235491
rect 354256 235479 354262 235491
rect 354314 235479 354320 235531
rect 394960 235479 394966 235531
rect 395018 235519 395024 235531
rect 587344 235519 587350 235531
rect 395018 235491 587350 235519
rect 395018 235479 395024 235491
rect 587344 235479 587350 235491
rect 587402 235479 587408 235531
rect 42160 235405 42166 235457
rect 42218 235445 42224 235457
rect 42544 235445 42550 235457
rect 42218 235417 42550 235445
rect 42218 235405 42224 235417
rect 42544 235405 42550 235417
rect 42602 235405 42608 235457
rect 211984 235405 211990 235457
rect 212042 235445 212048 235457
rect 233008 235445 233014 235457
rect 212042 235417 233014 235445
rect 212042 235405 212048 235417
rect 233008 235405 233014 235417
rect 233066 235405 233072 235457
rect 242128 235405 242134 235457
rect 242186 235445 242192 235457
rect 293392 235445 293398 235457
rect 242186 235417 293398 235445
rect 242186 235405 242192 235417
rect 293392 235405 293398 235417
rect 293450 235405 293456 235457
rect 294832 235405 294838 235457
rect 294890 235445 294896 235457
rect 338896 235445 338902 235457
rect 294890 235417 338902 235445
rect 294890 235405 294896 235417
rect 338896 235405 338902 235417
rect 338954 235405 338960 235457
rect 339472 235405 339478 235457
rect 339530 235445 339536 235457
rect 395056 235445 395062 235457
rect 339530 235417 395062 235445
rect 339530 235405 339536 235417
rect 395056 235405 395062 235417
rect 395114 235405 395120 235457
rect 396784 235405 396790 235457
rect 396842 235445 396848 235457
rect 588400 235445 588406 235457
rect 396842 235417 588406 235445
rect 396842 235405 396848 235417
rect 588400 235405 588406 235417
rect 588458 235405 588464 235457
rect 214192 235331 214198 235383
rect 214250 235371 214256 235383
rect 220528 235371 220534 235383
rect 214250 235343 220534 235371
rect 214250 235331 214256 235343
rect 220528 235331 220534 235343
rect 220586 235331 220592 235383
rect 220624 235331 220630 235383
rect 220682 235371 220688 235383
rect 241840 235371 241846 235383
rect 220682 235343 241846 235371
rect 220682 235331 220688 235343
rect 241840 235331 241846 235343
rect 241898 235331 241904 235383
rect 249712 235331 249718 235383
rect 249770 235371 249776 235383
rect 302320 235371 302326 235383
rect 249770 235343 302326 235371
rect 249770 235331 249776 235343
rect 302320 235331 302326 235343
rect 302378 235331 302384 235383
rect 304816 235331 304822 235383
rect 304874 235371 304880 235383
rect 362320 235371 362326 235383
rect 304874 235343 362326 235371
rect 304874 235331 304880 235343
rect 362320 235331 362326 235343
rect 362378 235331 362384 235383
rect 393424 235331 393430 235383
rect 393482 235371 393488 235383
rect 587056 235371 587062 235383
rect 393482 235343 587062 235371
rect 393482 235331 393488 235343
rect 587056 235331 587062 235343
rect 587114 235331 587120 235383
rect 209296 235257 209302 235309
rect 209354 235297 209360 235309
rect 228496 235297 228502 235309
rect 209354 235269 228502 235297
rect 209354 235257 209360 235269
rect 228496 235257 228502 235269
rect 228554 235257 228560 235309
rect 229744 235257 229750 235309
rect 229802 235297 229808 235309
rect 253552 235297 253558 235309
rect 229802 235269 253558 235297
rect 229802 235257 229808 235269
rect 253552 235257 253558 235269
rect 253610 235257 253616 235309
rect 257488 235257 257494 235309
rect 257546 235297 257552 235309
rect 308176 235297 308182 235309
rect 257546 235269 308182 235297
rect 257546 235257 257552 235269
rect 308176 235257 308182 235269
rect 308234 235257 308240 235309
rect 334960 235257 334966 235309
rect 335018 235297 335024 235309
rect 391696 235297 391702 235309
rect 335018 235269 391702 235297
rect 335018 235257 335024 235269
rect 391696 235257 391702 235269
rect 391754 235257 391760 235309
rect 396304 235257 396310 235309
rect 396362 235297 396368 235309
rect 587632 235297 587638 235309
rect 396362 235269 587638 235297
rect 396362 235257 396368 235269
rect 587632 235257 587638 235269
rect 587690 235257 587696 235309
rect 42256 235183 42262 235235
rect 42314 235223 42320 235235
rect 42448 235223 42454 235235
rect 42314 235195 42454 235223
rect 42314 235183 42320 235195
rect 42448 235183 42454 235195
rect 42506 235183 42512 235235
rect 230704 235223 230710 235235
rect 215986 235195 230710 235223
rect 211600 235109 211606 235161
rect 211658 235149 211664 235161
rect 215986 235149 216014 235195
rect 230704 235183 230710 235195
rect 230762 235183 230768 235235
rect 232912 235183 232918 235235
rect 232970 235223 232976 235235
rect 232970 235195 247694 235223
rect 232970 235183 232976 235195
rect 211658 235121 216014 235149
rect 211658 235109 211664 235121
rect 223888 235109 223894 235161
rect 223946 235149 223952 235161
rect 244720 235149 244726 235161
rect 223946 235121 244726 235149
rect 223946 235109 223952 235121
rect 244720 235109 244726 235121
rect 244778 235109 244784 235161
rect 247666 235149 247694 235195
rect 288880 235183 288886 235235
rect 288938 235223 288944 235235
rect 345712 235223 345718 235235
rect 288938 235195 345718 235223
rect 288938 235183 288944 235195
rect 345712 235183 345718 235195
rect 345770 235183 345776 235235
rect 392176 235183 392182 235235
rect 392234 235223 392240 235235
rect 587248 235223 587254 235235
rect 392234 235195 587254 235223
rect 392234 235183 392240 235195
rect 587248 235183 587254 235195
rect 587306 235183 587312 235235
rect 262000 235149 262006 235161
rect 247666 235121 262006 235149
rect 262000 235109 262006 235121
rect 262058 235109 262064 235161
rect 266128 235109 266134 235161
rect 266186 235149 266192 235161
rect 324112 235149 324118 235161
rect 266186 235121 324118 235149
rect 266186 235109 266192 235121
rect 324112 235109 324118 235121
rect 324170 235109 324176 235161
rect 332176 235109 332182 235161
rect 332234 235149 332240 235161
rect 385360 235149 385366 235161
rect 332234 235121 385366 235149
rect 332234 235109 332240 235121
rect 385360 235109 385366 235121
rect 385418 235109 385424 235161
rect 387664 235109 387670 235161
rect 387722 235149 387728 235161
rect 583408 235149 583414 235161
rect 387722 235121 583414 235149
rect 387722 235109 387728 235121
rect 583408 235109 583414 235121
rect 583466 235109 583472 235161
rect 207472 235035 207478 235087
rect 207530 235075 207536 235087
rect 223984 235075 223990 235087
rect 207530 235047 223990 235075
rect 207530 235035 207536 235047
rect 223984 235035 223990 235047
rect 224042 235035 224048 235087
rect 246640 235035 246646 235087
rect 246698 235075 246704 235087
rect 299248 235075 299254 235087
rect 246698 235047 299254 235075
rect 246698 235035 246704 235047
rect 299248 235035 299254 235047
rect 299306 235035 299312 235087
rect 309328 235035 309334 235087
rect 309386 235075 309392 235087
rect 370576 235075 370582 235087
rect 309386 235047 370582 235075
rect 309386 235035 309392 235047
rect 370576 235035 370582 235047
rect 370634 235035 370640 235087
rect 394864 235035 394870 235087
rect 394922 235075 394928 235087
rect 596080 235075 596086 235087
rect 394922 235047 596086 235075
rect 394922 235035 394928 235047
rect 596080 235035 596086 235047
rect 596138 235035 596144 235087
rect 211024 234961 211030 235013
rect 211082 235001 211088 235013
rect 231568 235001 231574 235013
rect 211082 234973 231574 235001
rect 211082 234961 211088 234973
rect 231568 234961 231574 234973
rect 231626 234961 231632 235013
rect 243856 234961 243862 235013
rect 243914 235001 243920 235013
rect 296464 235001 296470 235013
rect 243914 234973 296470 235001
rect 243914 234961 243920 234973
rect 296464 234961 296470 234973
rect 296522 234961 296528 235013
rect 298000 234961 298006 235013
rect 298058 235001 298064 235013
rect 362416 235001 362422 235013
rect 298058 234973 362422 235001
rect 298058 234961 298064 234973
rect 362416 234961 362422 234973
rect 362474 234961 362480 235013
rect 362512 234961 362518 235013
rect 362570 235001 362576 235013
rect 394672 235001 394678 235013
rect 362570 234973 394678 235001
rect 362570 234961 362576 234973
rect 394672 234961 394678 234973
rect 394730 234961 394736 235013
rect 398992 234961 398998 235013
rect 399050 235001 399056 235013
rect 605968 235001 605974 235013
rect 399050 234973 605974 235001
rect 399050 234961 399056 234973
rect 605968 234961 605974 234973
rect 606026 234961 606032 235013
rect 213424 234887 213430 234939
rect 213482 234927 213488 234939
rect 213482 234899 216014 234927
rect 213482 234887 213488 234899
rect 204400 234813 204406 234865
rect 204458 234853 204464 234865
rect 210160 234853 210166 234865
rect 204458 234825 210166 234853
rect 204458 234813 204464 234825
rect 210160 234813 210166 234825
rect 210218 234813 210224 234865
rect 204784 234739 204790 234791
rect 204842 234779 204848 234791
rect 210448 234779 210454 234791
rect 204842 234751 210454 234779
rect 204842 234739 204848 234751
rect 210448 234739 210454 234751
rect 210506 234739 210512 234791
rect 215986 234779 216014 234899
rect 220528 234887 220534 234939
rect 220586 234927 220592 234939
rect 235312 234927 235318 234939
rect 220586 234899 235318 234927
rect 220586 234887 220592 234899
rect 235312 234887 235318 234899
rect 235370 234887 235376 234939
rect 235696 234887 235702 234939
rect 235754 234927 235760 234939
rect 265072 234927 265078 234939
rect 235754 234899 265078 234927
rect 235754 234887 235760 234899
rect 265072 234887 265078 234899
rect 265130 234887 265136 234939
rect 268912 234887 268918 234939
rect 268970 234927 268976 234939
rect 331408 234927 331414 234939
rect 268970 234899 331414 234927
rect 268970 234887 268976 234899
rect 331408 234887 331414 234899
rect 331466 234887 331472 234939
rect 333424 234887 333430 234939
rect 333482 234927 333488 234939
rect 394768 234927 394774 234939
rect 333482 234899 394774 234927
rect 333482 234887 333488 234899
rect 394768 234887 394774 234899
rect 394826 234887 394832 234939
rect 398608 234887 398614 234939
rect 398666 234927 398672 234939
rect 605296 234927 605302 234939
rect 398666 234899 605302 234927
rect 398666 234887 398672 234899
rect 605296 234887 605302 234899
rect 605354 234887 605360 234939
rect 225520 234813 225526 234865
rect 225578 234853 225584 234865
rect 260176 234853 260182 234865
rect 225578 234825 260182 234853
rect 225578 234813 225584 234825
rect 260176 234813 260182 234825
rect 260234 234813 260240 234865
rect 260272 234813 260278 234865
rect 260330 234853 260336 234865
rect 323152 234853 323158 234865
rect 260330 234825 323158 234853
rect 260330 234813 260336 234825
rect 323152 234813 323158 234825
rect 323210 234813 323216 234865
rect 327664 234813 327670 234865
rect 327722 234853 327728 234865
rect 392464 234853 392470 234865
rect 327722 234825 392470 234853
rect 327722 234813 327728 234825
rect 392464 234813 392470 234825
rect 392522 234813 392528 234865
rect 403600 234813 403606 234865
rect 403658 234853 403664 234865
rect 615856 234853 615862 234865
rect 403658 234825 615862 234853
rect 403658 234813 403664 234825
rect 615856 234813 615862 234825
rect 615914 234813 615920 234865
rect 236080 234779 236086 234791
rect 215986 234751 236086 234779
rect 236080 234739 236086 234751
rect 236138 234739 236144 234791
rect 254224 234739 254230 234791
rect 254282 234779 254288 234791
rect 306736 234779 306742 234791
rect 254282 234751 306742 234779
rect 254282 234739 254288 234751
rect 306736 234739 306742 234751
rect 306794 234739 306800 234791
rect 321616 234739 321622 234791
rect 321674 234779 321680 234791
rect 387280 234779 387286 234791
rect 321674 234751 387286 234779
rect 321674 234739 321680 234751
rect 387280 234739 387286 234751
rect 387338 234739 387344 234791
rect 406672 234739 406678 234791
rect 406730 234779 406736 234791
rect 621808 234779 621814 234791
rect 406730 234751 621814 234779
rect 406730 234739 406736 234751
rect 621808 234739 621814 234751
rect 621866 234739 621872 234791
rect 206512 234665 206518 234717
rect 206570 234705 206576 234717
rect 222448 234705 222454 234717
rect 206570 234677 222454 234705
rect 206570 234665 206576 234677
rect 222448 234665 222454 234677
rect 222506 234665 222512 234717
rect 225136 234665 225142 234717
rect 225194 234705 225200 234717
rect 247696 234705 247702 234717
rect 225194 234677 247702 234705
rect 225194 234665 225200 234677
rect 247696 234665 247702 234677
rect 247754 234665 247760 234717
rect 251152 234665 251158 234717
rect 251210 234705 251216 234717
rect 304144 234705 304150 234717
rect 251210 234677 304150 234705
rect 251210 234665 251216 234677
rect 304144 234665 304150 234677
rect 304202 234665 304208 234717
rect 315280 234665 315286 234717
rect 315338 234705 315344 234717
rect 394672 234705 394678 234717
rect 315338 234677 394678 234705
rect 315338 234665 315344 234677
rect 394672 234665 394678 234677
rect 394730 234665 394736 234717
rect 408112 234665 408118 234717
rect 408170 234705 408176 234717
rect 624880 234705 624886 234717
rect 408170 234677 624886 234705
rect 408170 234665 408176 234677
rect 624880 234665 624886 234677
rect 624938 234665 624944 234717
rect 202864 234591 202870 234643
rect 202922 234631 202928 234643
rect 214864 234631 214870 234643
rect 202922 234603 214870 234631
rect 202922 234591 202928 234603
rect 214864 234591 214870 234603
rect 214922 234591 214928 234643
rect 222256 234591 222262 234643
rect 222314 234631 222320 234643
rect 222314 234603 227534 234631
rect 222314 234591 222320 234603
rect 202000 234517 202006 234569
rect 202058 234557 202064 234569
rect 213424 234557 213430 234569
rect 202058 234529 213430 234557
rect 202058 234517 202064 234529
rect 213424 234517 213430 234529
rect 213482 234517 213488 234569
rect 227506 234557 227534 234603
rect 240208 234591 240214 234643
rect 240266 234631 240272 234643
rect 263824 234631 263830 234643
rect 240266 234603 263830 234631
rect 240266 234591 240272 234603
rect 263824 234591 263830 234603
rect 263882 234591 263888 234643
rect 267472 234591 267478 234643
rect 267530 234631 267536 234643
rect 282352 234631 282358 234643
rect 267530 234603 282358 234631
rect 267530 234591 267536 234603
rect 282352 234591 282358 234603
rect 282410 234591 282416 234643
rect 286672 234591 286678 234643
rect 286730 234631 286736 234643
rect 325744 234631 325750 234643
rect 286730 234603 325750 234631
rect 286730 234591 286736 234603
rect 325744 234591 325750 234603
rect 325802 234591 325808 234643
rect 329296 234591 329302 234643
rect 329354 234631 329360 234643
rect 449296 234631 449302 234643
rect 329354 234603 449302 234631
rect 329354 234591 329360 234603
rect 449296 234591 449302 234603
rect 449354 234591 449360 234643
rect 243952 234557 243958 234569
rect 227506 234529 243958 234557
rect 243952 234517 243958 234529
rect 244010 234517 244016 234569
rect 250576 234557 250582 234569
rect 247666 234529 250582 234557
rect 206128 234443 206134 234495
rect 206186 234483 206192 234495
rect 211984 234483 211990 234495
rect 206186 234455 211990 234483
rect 206186 234443 206192 234455
rect 211984 234443 211990 234455
rect 212042 234443 212048 234495
rect 235600 234443 235606 234495
rect 235658 234483 235664 234495
rect 247666 234483 247694 234529
rect 250576 234517 250582 234529
rect 250634 234517 250640 234569
rect 255280 234517 255286 234569
rect 255338 234557 255344 234569
rect 278032 234557 278038 234569
rect 255338 234529 278038 234557
rect 255338 234517 255344 234529
rect 278032 234517 278038 234529
rect 278090 234517 278096 234569
rect 283888 234517 283894 234569
rect 283946 234557 283952 234569
rect 322192 234557 322198 234569
rect 283946 234529 322198 234557
rect 283946 234517 283952 234529
rect 322192 234517 322198 234529
rect 322250 234517 322256 234569
rect 323536 234517 323542 234569
rect 323594 234557 323600 234569
rect 434896 234557 434902 234569
rect 323594 234529 434902 234557
rect 323594 234517 323600 234529
rect 434896 234517 434902 234529
rect 434954 234517 434960 234569
rect 235658 234455 247694 234483
rect 235658 234443 235664 234455
rect 250480 234443 250486 234495
rect 250538 234483 250544 234495
rect 267952 234483 267958 234495
rect 250538 234455 267958 234483
rect 250538 234443 250544 234455
rect 267952 234443 267958 234455
rect 268010 234443 268016 234495
rect 273040 234443 273046 234495
rect 273098 234483 273104 234495
rect 305104 234483 305110 234495
rect 273098 234455 305110 234483
rect 273098 234443 273104 234455
rect 305104 234443 305110 234455
rect 305162 234443 305168 234495
rect 314416 234443 314422 234495
rect 314474 234483 314480 234495
rect 426160 234483 426166 234495
rect 314474 234455 426166 234483
rect 314474 234443 314480 234455
rect 426160 234443 426166 234455
rect 426218 234443 426224 234495
rect 206992 234369 206998 234421
rect 207050 234409 207056 234421
rect 221776 234409 221782 234421
rect 207050 234381 221782 234409
rect 207050 234369 207056 234381
rect 221776 234369 221782 234381
rect 221834 234369 221840 234421
rect 237040 234369 237046 234421
rect 237098 234409 237104 234421
rect 258928 234409 258934 234421
rect 237098 234381 258934 234409
rect 237098 234369 237104 234381
rect 258928 234369 258934 234381
rect 258986 234369 258992 234421
rect 262480 234369 262486 234421
rect 262538 234409 262544 234421
rect 290896 234409 290902 234421
rect 262538 234381 290902 234409
rect 262538 234369 262544 234381
rect 290896 234369 290902 234381
rect 290954 234369 290960 234421
rect 292912 234369 292918 234421
rect 292970 234409 292976 234421
rect 311152 234409 311158 234421
rect 292970 234381 311158 234409
rect 292970 234369 292976 234381
rect 311152 234369 311158 234381
rect 311210 234369 311216 234421
rect 312688 234369 312694 234421
rect 312746 234409 312752 234421
rect 407440 234409 407446 234421
rect 312746 234381 407446 234409
rect 312746 234369 312752 234381
rect 407440 234369 407446 234381
rect 407498 234369 407504 234421
rect 203248 234295 203254 234347
rect 203306 234335 203312 234347
rect 206800 234335 206806 234347
rect 203306 234307 206806 234335
rect 203306 234295 203312 234307
rect 206800 234295 206806 234307
rect 206858 234295 206864 234347
rect 206896 234295 206902 234347
rect 206954 234335 206960 234347
rect 220240 234335 220246 234347
rect 206954 234307 220246 234335
rect 206954 234295 206960 234307
rect 220240 234295 220246 234307
rect 220298 234295 220304 234347
rect 239824 234295 239830 234347
rect 239882 234335 239888 234347
rect 260944 234335 260950 234347
rect 239882 234307 260950 234335
rect 239882 234295 239888 234307
rect 260944 234295 260950 234307
rect 261002 234295 261008 234347
rect 271600 234295 271606 234347
rect 271658 234335 271664 234347
rect 302128 234335 302134 234347
rect 271658 234307 302134 234335
rect 271658 234295 271664 234307
rect 302128 234295 302134 234307
rect 302186 234295 302192 234347
rect 308464 234295 308470 234347
rect 308522 234335 308528 234347
rect 414736 234335 414742 234347
rect 308522 234307 414742 234335
rect 308522 234295 308528 234307
rect 414736 234295 414742 234307
rect 414794 234295 414800 234347
rect 42256 234221 42262 234273
rect 42314 234261 42320 234273
rect 42928 234261 42934 234273
rect 42314 234233 42934 234261
rect 42314 234221 42320 234233
rect 42928 234221 42934 234233
rect 42986 234221 42992 234273
rect 201520 234221 201526 234273
rect 201578 234261 201584 234273
rect 211888 234261 211894 234273
rect 201578 234233 211894 234261
rect 201578 234221 201584 234233
rect 211888 234221 211894 234233
rect 211946 234221 211952 234273
rect 211984 234221 211990 234273
rect 212042 234261 212048 234273
rect 221008 234261 221014 234273
rect 212042 234233 221014 234261
rect 212042 234221 212048 234233
rect 221008 234221 221014 234233
rect 221066 234221 221072 234273
rect 242896 234221 242902 234273
rect 242954 234261 242960 234273
rect 261136 234261 261142 234273
rect 242954 234233 261142 234261
rect 242954 234221 242960 234233
rect 261136 234221 261142 234233
rect 261194 234221 261200 234273
rect 261232 234221 261238 234273
rect 261290 234261 261296 234273
rect 288016 234261 288022 234273
rect 261290 234233 288022 234261
rect 261290 234221 261296 234233
rect 288016 234221 288022 234233
rect 288074 234221 288080 234273
rect 295216 234221 295222 234273
rect 295274 234261 295280 234273
rect 348688 234261 348694 234273
rect 295274 234233 348694 234261
rect 295274 234221 295280 234233
rect 348688 234221 348694 234233
rect 348746 234221 348752 234273
rect 352144 234221 352150 234273
rect 352202 234261 352208 234273
rect 398128 234261 398134 234273
rect 352202 234233 398134 234261
rect 352202 234221 352208 234233
rect 398128 234221 398134 234233
rect 398186 234221 398192 234273
rect 398224 234221 398230 234273
rect 398282 234261 398288 234273
rect 406000 234261 406006 234273
rect 398282 234233 406006 234261
rect 398282 234221 398288 234233
rect 406000 234221 406006 234233
rect 406058 234221 406064 234273
rect 407248 234221 407254 234273
rect 407306 234261 407312 234273
rect 503920 234261 503926 234273
rect 407306 234233 503926 234261
rect 407306 234221 407312 234233
rect 503920 234221 503926 234233
rect 503978 234221 503984 234273
rect 200272 234147 200278 234199
rect 200330 234187 200336 234199
rect 210352 234187 210358 234199
rect 200330 234159 210358 234187
rect 200330 234147 200336 234159
rect 210352 234147 210358 234159
rect 210410 234147 210416 234199
rect 210448 234147 210454 234199
rect 210506 234187 210512 234199
rect 219376 234187 219382 234199
rect 210506 234159 219382 234187
rect 210506 234147 210512 234159
rect 219376 234147 219382 234159
rect 219434 234147 219440 234199
rect 256528 234147 256534 234199
rect 256586 234187 256592 234199
rect 279280 234187 279286 234199
rect 256586 234159 279286 234187
rect 256586 234147 256592 234159
rect 279280 234147 279286 234159
rect 279338 234147 279344 234199
rect 283984 234147 283990 234199
rect 284042 234187 284048 234199
rect 311344 234187 311350 234199
rect 284042 234159 311350 234187
rect 284042 234147 284048 234159
rect 311344 234147 311350 234159
rect 311402 234147 311408 234199
rect 318352 234147 318358 234199
rect 318410 234187 318416 234199
rect 371632 234187 371638 234199
rect 318410 234159 371638 234187
rect 318410 234147 318416 234159
rect 371632 234147 371638 234159
rect 371690 234147 371696 234199
rect 378544 234147 378550 234199
rect 378602 234187 378608 234199
rect 399184 234187 399190 234199
rect 378602 234159 399190 234187
rect 378602 234147 378608 234159
rect 399184 234147 399190 234159
rect 399242 234147 399248 234199
rect 403504 234147 403510 234199
rect 403562 234187 403568 234199
rect 495376 234187 495382 234199
rect 403562 234159 495382 234187
rect 403562 234147 403568 234159
rect 495376 234147 495382 234159
rect 495434 234147 495440 234199
rect 200176 234073 200182 234125
rect 200234 234113 200240 234125
rect 208816 234113 208822 234125
rect 200234 234085 208822 234113
rect 200234 234073 200240 234085
rect 208816 234073 208822 234085
rect 208874 234073 208880 234125
rect 225520 234113 225526 234125
rect 211906 234085 225526 234113
rect 198736 233999 198742 234051
rect 198794 234039 198800 234051
rect 207376 234039 207382 234051
rect 198794 234011 207382 234039
rect 198794 233999 198800 234011
rect 207376 233999 207382 234011
rect 207434 233999 207440 234051
rect 207856 233999 207862 234051
rect 207914 234039 207920 234051
rect 211906 234039 211934 234085
rect 225520 234073 225526 234085
rect 225578 234073 225584 234125
rect 244336 234073 244342 234125
rect 244394 234113 244400 234125
rect 264880 234113 264886 234125
rect 244394 234085 264886 234113
rect 244394 234073 244400 234085
rect 264880 234073 264886 234085
rect 264938 234073 264944 234125
rect 268528 234073 268534 234125
rect 268586 234113 268592 234125
rect 293776 234113 293782 234125
rect 268586 234085 293782 234113
rect 268586 234073 268592 234085
rect 293776 234073 293782 234085
rect 293834 234073 293840 234125
rect 295696 234073 295702 234125
rect 295754 234113 295760 234125
rect 341200 234113 341206 234125
rect 295754 234085 341206 234113
rect 295754 234073 295760 234085
rect 341200 234073 341206 234085
rect 341258 234073 341264 234125
rect 345904 234073 345910 234125
rect 345962 234113 345968 234125
rect 400144 234113 400150 234125
rect 345962 234085 400150 234113
rect 345962 234073 345968 234085
rect 400144 234073 400150 234085
rect 400202 234073 400208 234125
rect 401776 234073 401782 234125
rect 401834 234113 401840 234125
rect 484624 234113 484630 234125
rect 401834 234085 484630 234113
rect 401834 234073 401840 234085
rect 484624 234073 484630 234085
rect 484682 234073 484688 234125
rect 207914 234011 211934 234039
rect 207914 233999 207920 234011
rect 247408 233999 247414 234051
rect 247466 234039 247472 234051
rect 266320 234039 266326 234051
rect 247466 234011 266326 234039
rect 247466 233999 247472 234011
rect 266320 233999 266326 234011
rect 266378 233999 266384 234051
rect 267088 233999 267094 234051
rect 267146 234039 267152 234051
rect 290992 234039 290998 234051
rect 267146 234011 290998 234039
rect 267146 233999 267152 234011
rect 290992 233999 290998 234011
rect 291050 233999 291056 234051
rect 301648 233999 301654 234051
rect 301706 234039 301712 234051
rect 344080 234039 344086 234051
rect 301706 234011 344086 234039
rect 301706 233999 301712 234011
rect 344080 233999 344086 234011
rect 344138 233999 344144 234051
rect 344368 233999 344374 234051
rect 344426 234039 344432 234051
rect 394864 234039 394870 234051
rect 344426 234011 394870 234039
rect 344426 233999 344432 234011
rect 394864 233999 394870 234011
rect 394922 233999 394928 234051
rect 396688 233999 396694 234051
rect 396746 234039 396752 234051
rect 475216 234039 475222 234051
rect 396746 234011 475222 234039
rect 396746 233999 396752 234011
rect 475216 233999 475222 234011
rect 475274 233999 475280 234051
rect 198352 233925 198358 233977
rect 198410 233965 198416 233977
rect 205936 233965 205942 233977
rect 198410 233937 205942 233965
rect 198410 233925 198416 233937
rect 205936 233925 205942 233937
rect 205994 233925 206000 233977
rect 206800 233925 206806 233977
rect 206858 233965 206864 233977
rect 216496 233965 216502 233977
rect 206858 233937 216502 233965
rect 206858 233925 206864 233937
rect 216496 233925 216502 233937
rect 216554 233925 216560 233977
rect 259792 233925 259798 233977
rect 259850 233965 259856 233977
rect 281200 233965 281206 233977
rect 259850 233937 281206 233965
rect 259850 233925 259856 233937
rect 281200 233925 281206 233937
rect 281258 233925 281264 233977
rect 305200 233925 305206 233977
rect 305258 233965 305264 233977
rect 351376 233965 351382 233977
rect 305258 233937 351382 233965
rect 305258 233925 305264 233937
rect 351376 233925 351382 233937
rect 351434 233925 351440 233977
rect 361264 233925 361270 233977
rect 361322 233965 361328 233977
rect 432016 233965 432022 233977
rect 361322 233937 432022 233965
rect 361322 233925 361328 233937
rect 432016 233925 432022 233937
rect 432074 233925 432080 233977
rect 197488 233851 197494 233903
rect 197546 233891 197552 233903
rect 204304 233891 204310 233903
rect 197546 233863 204310 233891
rect 197546 233851 197552 233863
rect 204304 233851 204310 233863
rect 204362 233851 204368 233903
rect 205168 233851 205174 233903
rect 205226 233891 205232 233903
rect 217168 233891 217174 233903
rect 205226 233863 217174 233891
rect 205226 233851 205232 233863
rect 217168 233851 217174 233863
rect 217226 233851 217232 233903
rect 258352 233851 258358 233903
rect 258410 233891 258416 233903
rect 279184 233891 279190 233903
rect 258410 233863 279190 233891
rect 258410 233851 258416 233863
rect 279184 233851 279190 233863
rect 279242 233851 279248 233903
rect 296080 233851 296086 233903
rect 296138 233891 296144 233903
rect 339088 233891 339094 233903
rect 296138 233863 339094 233891
rect 296138 233851 296144 233863
rect 339088 233851 339094 233863
rect 339146 233851 339152 233903
rect 370288 233851 370294 233903
rect 370346 233891 370352 233903
rect 427888 233891 427894 233903
rect 370346 233863 427894 233891
rect 370346 233851 370352 233863
rect 427888 233851 427894 233863
rect 427946 233851 427952 233903
rect 196912 233777 196918 233829
rect 196970 233817 196976 233829
rect 202864 233817 202870 233829
rect 196970 233789 202870 233817
rect 196970 233777 196976 233789
rect 202864 233777 202870 233789
rect 202922 233777 202928 233829
rect 204208 233777 204214 233829
rect 204266 233817 204272 233829
rect 215536 233817 215542 233829
rect 204266 233789 215542 233817
rect 204266 233777 204272 233789
rect 215536 233777 215542 233789
rect 215594 233777 215600 233829
rect 253456 233777 253462 233829
rect 253514 233817 253520 233829
rect 270832 233817 270838 233829
rect 253514 233789 270838 233817
rect 253514 233777 253520 233789
rect 270832 233777 270838 233789
rect 270890 233777 270896 233829
rect 285136 233777 285142 233829
rect 285194 233817 285200 233829
rect 325360 233817 325366 233829
rect 285194 233789 325366 233817
rect 285194 233777 285200 233789
rect 325360 233777 325366 233789
rect 325418 233777 325424 233829
rect 354928 233777 354934 233829
rect 354986 233817 354992 233829
rect 407344 233817 407350 233829
rect 354986 233789 407350 233817
rect 354986 233777 354992 233789
rect 407344 233777 407350 233789
rect 407402 233777 407408 233829
rect 407440 233777 407446 233829
rect 407498 233817 407504 233829
rect 423280 233817 423286 233829
rect 407498 233789 423286 233817
rect 407498 233777 407504 233789
rect 423280 233777 423286 233789
rect 423338 233777 423344 233829
rect 196528 233703 196534 233755
rect 196586 233743 196592 233755
rect 200560 233743 200566 233755
rect 196586 233715 200566 233743
rect 196586 233703 196592 233715
rect 200560 233703 200566 233715
rect 200618 233703 200624 233755
rect 201040 233703 201046 233755
rect 201098 233743 201104 233755
rect 209680 233743 209686 233755
rect 201098 233715 209686 233743
rect 201098 233703 201104 233715
rect 209680 233703 209686 233715
rect 209738 233703 209744 233755
rect 210160 233703 210166 233755
rect 210218 233743 210224 233755
rect 217936 233743 217942 233755
rect 210218 233715 217942 233743
rect 210218 233703 210224 233715
rect 217936 233703 217942 233715
rect 217994 233703 218000 233755
rect 294448 233703 294454 233755
rect 294506 233743 294512 233755
rect 331216 233743 331222 233755
rect 294506 233715 331222 233743
rect 294506 233703 294512 233715
rect 331216 233703 331222 233715
rect 331274 233703 331280 233755
rect 338032 233703 338038 233755
rect 338090 233743 338096 233755
rect 386128 233743 386134 233755
rect 338090 233715 386134 233743
rect 338090 233703 338096 233715
rect 386128 233703 386134 233715
rect 386186 233703 386192 233755
rect 398128 233703 398134 233755
rect 398186 233743 398192 233755
rect 403024 233743 403030 233755
rect 398186 233715 403030 233743
rect 398186 233703 398192 233715
rect 403024 233703 403030 233715
rect 403082 233703 403088 233755
rect 408976 233703 408982 233755
rect 409034 233743 409040 233755
rect 410608 233743 410614 233755
rect 409034 233715 410614 233743
rect 409034 233703 409040 233715
rect 410608 233703 410614 233715
rect 410666 233703 410672 233755
rect 195664 233629 195670 233681
rect 195722 233669 195728 233681
rect 201328 233669 201334 233681
rect 195722 233641 201334 233669
rect 195722 233629 195728 233641
rect 201328 233629 201334 233641
rect 201386 233629 201392 233681
rect 202480 233629 202486 233681
rect 202538 233669 202544 233681
rect 212560 233669 212566 233681
rect 202538 233641 212566 233669
rect 202538 233629 202544 233641
rect 212560 233629 212566 233641
rect 212618 233629 212624 233681
rect 306256 233629 306262 233681
rect 306314 233669 306320 233681
rect 344464 233669 344470 233681
rect 306314 233641 344470 233669
rect 306314 233629 306320 233641
rect 344464 233629 344470 233641
rect 344522 233629 344528 233681
rect 363472 233629 363478 233681
rect 363530 233669 363536 233681
rect 363760 233669 363766 233681
rect 363530 233641 363766 233669
rect 363530 233629 363536 233641
rect 363760 233629 363766 233641
rect 363818 233629 363824 233681
rect 383632 233629 383638 233681
rect 383690 233669 383696 233681
rect 408112 233669 408118 233681
rect 383690 233641 408118 233669
rect 383690 233629 383696 233641
rect 408112 233629 408118 233641
rect 408170 233629 408176 233681
rect 194224 233555 194230 233607
rect 194282 233595 194288 233607
rect 198352 233595 198358 233607
rect 194282 233567 198358 233595
rect 194282 233555 194288 233567
rect 198352 233555 198358 233567
rect 198410 233555 198416 233607
rect 199120 233555 199126 233607
rect 199178 233595 199184 233607
rect 205072 233595 205078 233607
rect 199178 233567 205078 233595
rect 199178 233555 199184 233567
rect 205072 233555 205078 233567
rect 205130 233555 205136 233607
rect 205552 233555 205558 233607
rect 205610 233595 205616 233607
rect 205610 233567 210782 233595
rect 205610 233555 205616 233567
rect 192880 233481 192886 233533
rect 192938 233521 192944 233533
rect 195280 233521 195286 233533
rect 192938 233493 195286 233521
rect 192938 233481 192944 233493
rect 195280 233481 195286 233493
rect 195338 233481 195344 233533
rect 195568 233481 195574 233533
rect 195626 233521 195632 233533
rect 199792 233521 199798 233533
rect 195626 233493 199798 233521
rect 195626 233481 195632 233493
rect 199792 233481 199798 233493
rect 199850 233481 199856 233533
rect 200656 233481 200662 233533
rect 200714 233521 200720 233533
rect 208144 233521 208150 233533
rect 200714 233493 208150 233521
rect 200714 233481 200720 233493
rect 208144 233481 208150 233493
rect 208202 233481 208208 233533
rect 210754 233521 210782 233567
rect 228400 233555 228406 233607
rect 228458 233595 228464 233607
rect 238096 233595 238102 233607
rect 228458 233567 238102 233595
rect 228458 233555 228464 233567
rect 238096 233555 238102 233567
rect 238154 233555 238160 233607
rect 259888 233555 259894 233607
rect 259946 233595 259952 233607
rect 267760 233595 267766 233607
rect 259946 233567 267766 233595
rect 259946 233555 259952 233567
rect 267760 233555 267766 233567
rect 267818 233555 267824 233607
rect 302896 233555 302902 233607
rect 302954 233595 302960 233607
rect 337360 233595 337366 233607
rect 302954 233567 337366 233595
rect 302954 233555 302960 233567
rect 337360 233555 337366 233567
rect 337418 233555 337424 233607
rect 348880 233555 348886 233607
rect 348938 233595 348944 233607
rect 394576 233595 394582 233607
rect 348938 233567 394582 233595
rect 348938 233555 348944 233567
rect 394576 233555 394582 233567
rect 394634 233555 394640 233607
rect 218704 233521 218710 233533
rect 210754 233493 218710 233521
rect 218704 233481 218710 233493
rect 218762 233481 218768 233533
rect 240592 233481 240598 233533
rect 240650 233521 240656 233533
rect 290416 233521 290422 233533
rect 240650 233493 290422 233521
rect 240650 233481 240656 233493
rect 290416 233481 290422 233493
rect 290474 233481 290480 233533
rect 297232 233481 297238 233533
rect 297290 233521 297296 233533
rect 328336 233521 328342 233533
rect 297290 233493 328342 233521
rect 297290 233481 297296 233493
rect 328336 233481 328342 233493
rect 328394 233481 328400 233533
rect 338608 233481 338614 233533
rect 338666 233521 338672 233533
rect 466480 233521 466486 233533
rect 338666 233493 466486 233521
rect 338666 233481 338672 233493
rect 466480 233481 466486 233493
rect 466538 233481 466544 233533
rect 42448 233407 42454 233459
rect 42506 233447 42512 233459
rect 43120 233447 43126 233459
rect 42506 233419 43126 233447
rect 42506 233407 42512 233419
rect 43120 233407 43126 233419
rect 43178 233407 43184 233459
rect 193840 233407 193846 233459
rect 193898 233447 193904 233459
rect 196816 233447 196822 233459
rect 193898 233419 196822 233447
rect 193898 233407 193904 233419
rect 196816 233407 196822 233419
rect 196874 233407 196880 233459
rect 197968 233407 197974 233459
rect 198026 233447 198032 233459
rect 203632 233447 203638 233459
rect 198026 233419 203638 233447
rect 198026 233407 198032 233419
rect 203632 233407 203638 233419
rect 203690 233407 203696 233459
rect 203920 233407 203926 233459
rect 203978 233447 203984 233459
rect 214192 233447 214198 233459
rect 203978 233419 214198 233447
rect 203978 233407 203984 233419
rect 214192 233407 214198 233419
rect 214250 233407 214256 233459
rect 264400 233407 264406 233459
rect 264458 233447 264464 233459
rect 271792 233447 271798 233459
rect 264458 233419 271798 233447
rect 264458 233407 264464 233419
rect 271792 233407 271798 233419
rect 271850 233407 271856 233459
rect 287440 233407 287446 233459
rect 287498 233447 287504 233459
rect 311248 233447 311254 233459
rect 287498 233419 311254 233447
rect 287498 233407 287504 233419
rect 311248 233407 311254 233419
rect 311306 233407 311312 233459
rect 320272 233407 320278 233459
rect 320330 233447 320336 233459
rect 448240 233447 448246 233459
rect 320330 233419 448246 233447
rect 320330 233407 320336 233419
rect 448240 233407 448246 233419
rect 448298 233407 448304 233459
rect 193264 233333 193270 233385
rect 193322 233373 193328 233385
rect 194608 233373 194614 233385
rect 193322 233345 194614 233373
rect 193322 233333 193328 233345
rect 194608 233333 194614 233345
rect 194666 233333 194672 233385
rect 195184 233333 195190 233385
rect 195242 233373 195248 233385
rect 197488 233373 197494 233385
rect 195242 233345 197494 233373
rect 195242 233333 195248 233345
rect 197488 233333 197494 233345
rect 197546 233333 197552 233385
rect 197872 233333 197878 233385
rect 197930 233373 197936 233385
rect 202096 233373 202102 233385
rect 197930 233345 202102 233373
rect 197930 233333 197936 233345
rect 202096 233333 202102 233345
rect 202154 233333 202160 233385
rect 202384 233333 202390 233385
rect 202442 233373 202448 233385
rect 211120 233373 211126 233385
rect 202442 233345 211126 233373
rect 202442 233333 202448 233345
rect 211120 233333 211126 233345
rect 211178 233333 211184 233385
rect 226672 233333 226678 233385
rect 226730 233373 226736 233385
rect 238960 233373 238966 233385
rect 226730 233345 238966 233373
rect 226730 233333 226736 233345
rect 238960 233333 238966 233345
rect 239018 233333 239024 233385
rect 261616 233333 261622 233385
rect 261674 233373 261680 233385
rect 269008 233373 269014 233385
rect 261674 233345 269014 233373
rect 261674 233333 261680 233345
rect 269008 233333 269014 233345
rect 269066 233333 269072 233385
rect 270448 233333 270454 233385
rect 270506 233373 270512 233385
rect 275056 233373 275062 233385
rect 270506 233345 275062 233373
rect 270506 233333 270512 233345
rect 275056 233333 275062 233345
rect 275114 233333 275120 233385
rect 288400 233333 288406 233385
rect 288458 233373 288464 233385
rect 311056 233373 311062 233385
rect 288458 233345 311062 233373
rect 288458 233333 288464 233345
rect 311056 233333 311062 233345
rect 311114 233333 311120 233385
rect 324784 233333 324790 233385
rect 324842 233373 324848 233385
rect 327280 233373 327286 233385
rect 324842 233345 327286 233373
rect 324842 233333 324848 233345
rect 327280 233333 327286 233345
rect 327338 233333 327344 233385
rect 335344 233333 335350 233385
rect 335402 233373 335408 233385
rect 463600 233373 463606 233385
rect 335402 233345 463606 233373
rect 335402 233333 335408 233345
rect 463600 233333 463606 233345
rect 463658 233333 463664 233385
rect 192400 233259 192406 233311
rect 192458 233299 192464 233311
rect 193744 233299 193750 233311
rect 192458 233271 193750 233299
rect 192458 233259 192464 233271
rect 193744 233259 193750 233271
rect 193802 233259 193808 233311
rect 194704 233259 194710 233311
rect 194762 233299 194768 233311
rect 196048 233299 196054 233311
rect 194762 233271 196054 233299
rect 194762 233259 194768 233271
rect 196048 233259 196054 233271
rect 196106 233259 196112 233311
rect 196144 233259 196150 233311
rect 196202 233299 196208 233311
rect 199120 233299 199126 233311
rect 196202 233271 199126 233299
rect 196202 233259 196208 233271
rect 199120 233259 199126 233271
rect 199178 233259 199184 233311
rect 199696 233259 199702 233311
rect 199754 233299 199760 233311
rect 206608 233299 206614 233311
rect 199754 233271 206614 233299
rect 199754 233259 199760 233271
rect 206608 233259 206614 233271
rect 206666 233259 206672 233311
rect 253840 233259 253846 233311
rect 253898 233299 253904 233311
rect 256240 233299 256246 233311
rect 253898 233271 256246 233299
rect 253898 233259 253904 233271
rect 256240 233259 256246 233271
rect 256298 233259 256304 233311
rect 257968 233259 257974 233311
rect 258026 233299 258032 233311
rect 269104 233299 269110 233311
rect 258026 233271 269110 233299
rect 258026 233259 258032 233271
rect 269104 233259 269110 233271
rect 269162 233259 269168 233311
rect 270256 233259 270262 233311
rect 270314 233299 270320 233311
rect 273520 233299 273526 233311
rect 270314 233271 273526 233299
rect 270314 233259 270320 233271
rect 273520 233259 273526 233271
rect 273578 233259 273584 233311
rect 297136 233259 297142 233311
rect 297194 233299 297200 233311
rect 317872 233299 317878 233311
rect 297194 233271 317878 233299
rect 297194 233259 297200 233271
rect 317872 233259 317878 233271
rect 317930 233259 317936 233311
rect 319888 233259 319894 233311
rect 319946 233299 319952 233311
rect 377296 233299 377302 233311
rect 319946 233271 377302 233299
rect 319946 233259 319952 233271
rect 377296 233259 377302 233271
rect 377354 233259 377360 233311
rect 380464 233259 380470 233311
rect 380522 233299 380528 233311
rect 382960 233299 382966 233311
rect 380522 233271 382966 233299
rect 380522 233259 380528 233271
rect 382960 233259 382966 233271
rect 383018 233259 383024 233311
rect 395920 233259 395926 233311
rect 395978 233299 395984 233311
rect 400240 233299 400246 233311
rect 395978 233271 400246 233299
rect 395978 233259 395984 233271
rect 400240 233259 400246 233271
rect 400298 233259 400304 233311
rect 401200 233259 401206 233311
rect 401258 233299 401264 233311
rect 408880 233299 408886 233311
rect 401258 233271 408886 233299
rect 401258 233259 401264 233271
rect 408880 233259 408886 233271
rect 408938 233259 408944 233311
rect 258736 233185 258742 233237
rect 258794 233225 258800 233237
rect 326704 233225 326710 233237
rect 258794 233197 326710 233225
rect 258794 233185 258800 233197
rect 326704 233185 326710 233197
rect 326762 233185 326768 233237
rect 340816 233185 340822 233237
rect 340874 233225 340880 233237
rect 491248 233225 491254 233237
rect 340874 233197 491254 233225
rect 340874 233185 340880 233197
rect 491248 233185 491254 233197
rect 491306 233185 491312 233237
rect 495376 233185 495382 233237
rect 495434 233225 495440 233237
rect 614992 233225 614998 233237
rect 495434 233197 614998 233225
rect 495434 233185 495440 233197
rect 614992 233185 614998 233197
rect 615050 233185 615056 233237
rect 260656 233111 260662 233163
rect 260714 233151 260720 233163
rect 331312 233151 331318 233163
rect 260714 233123 331318 233151
rect 260714 233111 260720 233123
rect 331312 233111 331318 233123
rect 331370 233111 331376 233163
rect 347056 233111 347062 233163
rect 347114 233151 347120 233163
rect 501040 233151 501046 233163
rect 347114 233123 501046 233151
rect 347114 233111 347120 233123
rect 501040 233111 501046 233123
rect 501098 233111 501104 233163
rect 262096 233037 262102 233089
rect 262154 233077 262160 233089
rect 334192 233077 334198 233089
rect 262154 233049 334198 233077
rect 262154 233037 262160 233049
rect 334192 233037 334198 233049
rect 334250 233037 334256 233089
rect 350320 233037 350326 233089
rect 350378 233077 350384 233089
rect 507088 233077 507094 233089
rect 350378 233049 507094 233077
rect 350378 233037 350384 233049
rect 507088 233037 507094 233049
rect 507146 233037 507152 233089
rect 265744 232963 265750 233015
rect 265802 233003 265808 233015
rect 338032 233003 338038 233015
rect 265802 232975 338038 233003
rect 265802 232963 265808 232975
rect 338032 232963 338038 232975
rect 338090 232963 338096 233015
rect 353104 232963 353110 233015
rect 353162 233003 353168 233015
rect 513136 233003 513142 233015
rect 353162 232975 513142 233003
rect 353162 232963 353168 232975
rect 513136 232963 513142 232975
rect 513194 232963 513200 233015
rect 281296 232889 281302 232941
rect 281354 232929 281360 232941
rect 288976 232929 288982 232941
rect 281354 232901 288982 232929
rect 281354 232889 281360 232901
rect 288976 232889 288982 232901
rect 289034 232889 289040 232941
rect 289936 232889 289942 232941
rect 289994 232929 290000 232941
rect 382768 232929 382774 232941
rect 289994 232901 382774 232929
rect 289994 232889 290000 232901
rect 382768 232889 382774 232901
rect 382826 232889 382832 232941
rect 410032 232889 410038 232941
rect 410090 232929 410096 232941
rect 572080 232929 572086 232941
rect 410090 232901 572086 232929
rect 410090 232889 410096 232901
rect 572080 232889 572086 232901
rect 572138 232889 572144 232941
rect 263920 232815 263926 232867
rect 263978 232855 263984 232867
rect 337264 232855 337270 232867
rect 263978 232827 337270 232855
rect 263978 232815 263984 232827
rect 337264 232815 337270 232827
rect 337322 232815 337328 232867
rect 356272 232815 356278 232867
rect 356330 232855 356336 232867
rect 519184 232855 519190 232867
rect 356330 232827 519190 232855
rect 356330 232815 356336 232827
rect 519184 232815 519190 232827
rect 519242 232815 519248 232867
rect 216592 232741 216598 232793
rect 216650 232781 216656 232793
rect 242128 232781 242134 232793
rect 216650 232753 242134 232781
rect 216650 232741 216656 232753
rect 242128 232741 242134 232753
rect 242186 232741 242192 232793
rect 265168 232741 265174 232793
rect 265226 232781 265232 232793
rect 340240 232781 340246 232793
rect 265226 232753 340246 232781
rect 265226 232741 265232 232753
rect 340240 232741 340246 232753
rect 340298 232741 340304 232793
rect 359056 232741 359062 232793
rect 359114 232781 359120 232793
rect 525232 232781 525238 232793
rect 359114 232753 525238 232781
rect 359114 232741 359120 232753
rect 525232 232741 525238 232753
rect 525290 232741 525296 232793
rect 237616 232667 237622 232719
rect 237674 232707 237680 232719
rect 284368 232707 284374 232719
rect 237674 232679 284374 232707
rect 237674 232667 237680 232679
rect 284368 232667 284374 232679
rect 284426 232667 284432 232719
rect 295312 232667 295318 232719
rect 295370 232707 295376 232719
rect 397360 232707 397366 232719
rect 295370 232679 397366 232707
rect 295370 232667 295376 232679
rect 397360 232667 397366 232679
rect 397418 232667 397424 232719
rect 399184 232667 399190 232719
rect 399242 232707 399248 232719
rect 566704 232707 566710 232719
rect 399242 232679 566710 232707
rect 399242 232667 399248 232679
rect 566704 232667 566710 232679
rect 566762 232667 566768 232719
rect 219760 232593 219766 232645
rect 219818 232633 219824 232645
rect 248080 232633 248086 232645
rect 219818 232605 248086 232633
rect 219818 232593 219824 232605
rect 248080 232593 248086 232605
rect 248138 232593 248144 232645
rect 266608 232593 266614 232645
rect 266666 232633 266672 232645
rect 343216 232633 343222 232645
rect 266666 232605 343222 232633
rect 266666 232593 266672 232605
rect 343216 232593 343222 232605
rect 343274 232593 343280 232645
rect 362128 232593 362134 232645
rect 362186 232633 362192 232645
rect 531280 232633 531286 232645
rect 362186 232605 531286 232633
rect 362186 232593 362192 232605
rect 531280 232593 531286 232605
rect 531338 232593 531344 232645
rect 218032 232519 218038 232571
rect 218090 232559 218096 232571
rect 245104 232559 245110 232571
rect 218090 232531 245110 232559
rect 218090 232519 218096 232531
rect 245104 232519 245110 232531
rect 245162 232519 245168 232571
rect 268432 232519 268438 232571
rect 268490 232559 268496 232571
rect 346288 232559 346294 232571
rect 268490 232531 346294 232559
rect 268490 232519 268496 232531
rect 346288 232519 346294 232531
rect 346346 232519 346352 232571
rect 346768 232519 346774 232571
rect 346826 232559 346832 232571
rect 356080 232559 356086 232571
rect 346826 232531 356086 232559
rect 346826 232519 346832 232531
rect 356080 232519 356086 232531
rect 356138 232519 356144 232571
rect 365392 232519 365398 232571
rect 365450 232559 365456 232571
rect 537232 232559 537238 232571
rect 365450 232531 537238 232559
rect 365450 232519 365456 232531
rect 537232 232519 537238 232531
rect 537290 232519 537296 232571
rect 221104 232445 221110 232497
rect 221162 232485 221168 232497
rect 251152 232485 251158 232497
rect 221162 232457 251158 232485
rect 221162 232445 221168 232457
rect 251152 232445 251158 232457
rect 251210 232445 251216 232497
rect 269680 232445 269686 232497
rect 269738 232485 269744 232497
rect 349360 232485 349366 232497
rect 269738 232457 349366 232485
rect 269738 232445 269744 232457
rect 349360 232445 349366 232457
rect 349418 232445 349424 232497
rect 365008 232445 365014 232497
rect 365066 232485 365072 232497
rect 539536 232485 539542 232497
rect 365066 232457 539542 232485
rect 365066 232445 365072 232457
rect 539536 232445 539542 232457
rect 539594 232445 539600 232497
rect 222544 232371 222550 232423
rect 222602 232411 222608 232423
rect 254224 232411 254230 232423
rect 222602 232383 254230 232411
rect 222602 232371 222608 232383
rect 254224 232371 254230 232383
rect 254282 232371 254288 232423
rect 271216 232371 271222 232423
rect 271274 232411 271280 232423
rect 271274 232383 346910 232411
rect 271274 232371 271280 232383
rect 222928 232297 222934 232349
rect 222986 232337 222992 232349
rect 255664 232337 255670 232349
rect 222986 232309 255670 232337
rect 222986 232297 222992 232309
rect 255664 232297 255670 232309
rect 255722 232297 255728 232349
rect 274864 232297 274870 232349
rect 274922 232337 274928 232349
rect 346768 232337 346774 232349
rect 274922 232309 346774 232337
rect 274922 232297 274928 232309
rect 346768 232297 346774 232309
rect 346826 232297 346832 232349
rect 346882 232337 346910 232383
rect 346960 232371 346966 232423
rect 347018 232411 347024 232423
rect 361360 232411 361366 232423
rect 347018 232383 361366 232411
rect 347018 232371 347024 232383
rect 361360 232371 361366 232383
rect 361418 232371 361424 232423
rect 368176 232371 368182 232423
rect 368234 232411 368240 232423
rect 543376 232411 543382 232423
rect 368234 232383 543382 232411
rect 368234 232371 368240 232383
rect 543376 232371 543382 232383
rect 543434 232371 543440 232423
rect 352336 232337 352342 232349
rect 346882 232309 352342 232337
rect 352336 232297 352342 232309
rect 352394 232297 352400 232349
rect 366256 232297 366262 232349
rect 366314 232337 366320 232349
rect 542608 232337 542614 232349
rect 366314 232309 542614 232337
rect 366314 232297 366320 232309
rect 542608 232297 542614 232309
rect 542666 232297 542672 232349
rect 224272 232223 224278 232275
rect 224330 232263 224336 232275
rect 257200 232263 257206 232275
rect 224330 232235 257206 232263
rect 224330 232223 224336 232235
rect 257200 232223 257206 232235
rect 257258 232223 257264 232275
rect 274192 232223 274198 232275
rect 274250 232263 274256 232275
rect 358288 232263 358294 232275
rect 274250 232235 358294 232263
rect 274250 232223 274256 232235
rect 358288 232223 358294 232235
rect 358346 232223 358352 232275
rect 369520 232223 369526 232275
rect 369578 232263 369584 232275
rect 548560 232263 548566 232275
rect 369578 232235 548566 232263
rect 369578 232223 369584 232235
rect 548560 232223 548566 232235
rect 548618 232223 548624 232275
rect 147856 232149 147862 232201
rect 147914 232189 147920 232201
rect 154096 232189 154102 232201
rect 147914 232161 154102 232189
rect 147914 232149 147920 232161
rect 154096 232149 154102 232161
rect 154154 232149 154160 232201
rect 226288 232149 226294 232201
rect 226346 232189 226352 232201
rect 261712 232189 261718 232201
rect 226346 232161 261718 232189
rect 226346 232149 226352 232161
rect 261712 232149 261718 232161
rect 261770 232149 261776 232201
rect 272944 232149 272950 232201
rect 273002 232189 273008 232201
rect 355312 232189 355318 232201
rect 273002 232161 355318 232189
rect 273002 232149 273008 232161
rect 355312 232149 355318 232161
rect 355370 232149 355376 232201
rect 372688 232149 372694 232201
rect 372746 232189 372752 232201
rect 552400 232189 552406 232201
rect 372746 232161 552406 232189
rect 372746 232149 372752 232161
rect 552400 232149 552406 232161
rect 552458 232149 552464 232201
rect 227056 232075 227062 232127
rect 227114 232115 227120 232127
rect 263248 232115 263254 232127
rect 227114 232087 263254 232115
rect 227114 232075 227120 232087
rect 263248 232075 263254 232087
rect 263306 232075 263312 232127
rect 277456 232075 277462 232127
rect 277514 232115 277520 232127
rect 364432 232115 364438 232127
rect 277514 232087 364438 232115
rect 277514 232075 277520 232087
rect 364432 232075 364438 232087
rect 364490 232075 364496 232127
rect 368080 232075 368086 232127
rect 368138 232115 368144 232127
rect 545584 232115 545590 232127
rect 368138 232087 545590 232115
rect 368138 232075 368144 232087
rect 545584 232075 545590 232087
rect 545642 232075 545648 232127
rect 233872 232001 233878 232053
rect 233930 232041 233936 232053
rect 274480 232041 274486 232053
rect 233930 232013 274486 232041
rect 233930 232001 233936 232013
rect 274480 232001 274486 232013
rect 274538 232001 274544 232053
rect 275728 232001 275734 232053
rect 275786 232041 275792 232053
rect 346960 232041 346966 232053
rect 275786 232013 346966 232041
rect 275786 232001 275792 232013
rect 346960 232001 346966 232013
rect 347018 232001 347024 232053
rect 354256 232001 354262 232053
rect 354314 232041 354320 232053
rect 367120 232041 367126 232053
rect 354314 232013 367126 232041
rect 354314 232001 354320 232013
rect 367120 232001 367126 232013
rect 367178 232001 367184 232053
rect 372304 232001 372310 232053
rect 372362 232041 372368 232053
rect 554704 232041 554710 232053
rect 372362 232013 554710 232041
rect 372362 232001 372368 232013
rect 554704 232001 554710 232013
rect 554762 232001 554768 232053
rect 234832 231927 234838 231979
rect 234890 231967 234896 231979
rect 278320 231967 278326 231979
rect 234890 231939 278326 231967
rect 234890 231927 234896 231939
rect 278320 231927 278326 231939
rect 278378 231927 278384 231979
rect 280240 231927 280246 231979
rect 280298 231967 280304 231979
rect 370384 231967 370390 231979
rect 280298 231939 370390 231967
rect 280298 231927 280304 231939
rect 370384 231927 370390 231939
rect 370442 231927 370448 231979
rect 374512 231927 374518 231979
rect 374570 231967 374576 231979
rect 557008 231967 557014 231979
rect 374570 231939 557014 231967
rect 374570 231927 374576 231939
rect 557008 231927 557014 231939
rect 557066 231927 557072 231979
rect 233200 231853 233206 231905
rect 233258 231893 233264 231905
rect 275344 231893 275350 231905
rect 233258 231865 275350 231893
rect 233258 231853 233264 231865
rect 275344 231853 275350 231865
rect 275402 231853 275408 231905
rect 278992 231853 278998 231905
rect 279050 231893 279056 231905
rect 367408 231893 367414 231905
rect 279050 231865 367414 231893
rect 279050 231853 279056 231865
rect 367408 231853 367414 231865
rect 367466 231853 367472 231905
rect 375760 231853 375766 231905
rect 375818 231893 375824 231905
rect 558352 231893 558358 231905
rect 375818 231865 558358 231893
rect 375818 231853 375824 231865
rect 558352 231853 558358 231865
rect 558410 231853 558416 231905
rect 235984 231779 235990 231831
rect 236042 231819 236048 231831
rect 281296 231819 281302 231831
rect 236042 231791 281302 231819
rect 236042 231779 236048 231791
rect 281296 231779 281302 231791
rect 281354 231779 281360 231831
rect 281968 231779 281974 231831
rect 282026 231819 282032 231831
rect 373456 231819 373462 231831
rect 282026 231791 373462 231819
rect 282026 231779 282032 231791
rect 373456 231779 373462 231791
rect 373514 231779 373520 231831
rect 378928 231779 378934 231831
rect 378986 231819 378992 231831
rect 564496 231819 564502 231831
rect 378986 231791 564502 231819
rect 378986 231779 378992 231791
rect 564496 231779 564502 231791
rect 564554 231779 564560 231831
rect 259120 231705 259126 231757
rect 259178 231745 259184 231757
rect 328144 231745 328150 231757
rect 259178 231717 328150 231745
rect 259178 231705 259184 231717
rect 328144 231705 328150 231717
rect 328202 231705 328208 231757
rect 337552 231705 337558 231757
rect 337610 231745 337616 231757
rect 485200 231745 485206 231757
rect 337610 231717 485206 231745
rect 337610 231705 337616 231717
rect 485200 231705 485206 231717
rect 485258 231705 485264 231757
rect 257584 231631 257590 231683
rect 257642 231671 257648 231683
rect 325168 231671 325174 231683
rect 257642 231643 325174 231671
rect 257642 231631 257648 231643
rect 325168 231631 325174 231643
rect 325226 231631 325232 231683
rect 334864 231631 334870 231683
rect 334922 231671 334928 231683
rect 479152 231671 479158 231683
rect 334922 231643 479158 231671
rect 334922 231631 334928 231643
rect 479152 231631 479158 231643
rect 479210 231631 479216 231683
rect 255760 231557 255766 231609
rect 255818 231597 255824 231609
rect 320656 231597 320662 231609
rect 255818 231569 320662 231597
rect 255818 231557 255824 231569
rect 320656 231557 320662 231569
rect 320714 231557 320720 231609
rect 327088 231557 327094 231609
rect 327146 231597 327152 231609
rect 464080 231597 464086 231609
rect 327146 231569 464086 231597
rect 327146 231557 327152 231569
rect 464080 231557 464086 231569
rect 464138 231557 464144 231609
rect 248368 231483 248374 231535
rect 248426 231523 248432 231535
rect 305488 231523 305494 231535
rect 248426 231495 305494 231523
rect 248426 231483 248432 231495
rect 305488 231483 305494 231495
rect 305546 231483 305552 231535
rect 312208 231483 312214 231535
rect 312266 231523 312272 231535
rect 433840 231523 433846 231535
rect 312266 231495 433846 231523
rect 312266 231483 312272 231495
rect 433840 231483 433846 231495
rect 433898 231483 433904 231535
rect 290800 231409 290806 231461
rect 290858 231449 290864 231461
rect 374608 231449 374614 231461
rect 290858 231421 374614 231449
rect 290858 231409 290864 231421
rect 374608 231409 374614 231421
rect 374666 231409 374672 231461
rect 403120 231409 403126 231461
rect 403178 231449 403184 231461
rect 520720 231449 520726 231461
rect 403178 231421 520726 231449
rect 403178 231409 403184 231421
rect 520720 231409 520726 231421
rect 520778 231409 520784 231461
rect 292528 231335 292534 231387
rect 292586 231375 292592 231387
rect 379984 231375 379990 231387
rect 292586 231347 379990 231375
rect 292586 231335 292592 231347
rect 379984 231335 379990 231347
rect 380042 231335 380048 231387
rect 400144 231335 400150 231387
rect 400202 231375 400208 231387
rect 499600 231375 499606 231387
rect 400202 231347 499606 231375
rect 400202 231335 400208 231347
rect 499600 231335 499606 231347
rect 499658 231335 499664 231387
rect 245200 231261 245206 231313
rect 245258 231301 245264 231313
rect 299440 231301 299446 231313
rect 245258 231273 299446 231301
rect 245258 231261 245264 231273
rect 299440 231261 299446 231273
rect 299498 231261 299504 231313
rect 300208 231261 300214 231313
rect 300266 231301 300272 231313
rect 385840 231301 385846 231313
rect 300266 231273 385846 231301
rect 300266 231261 300272 231273
rect 385840 231261 385846 231273
rect 385898 231261 385904 231313
rect 395056 231261 395062 231313
rect 395114 231301 395120 231313
rect 485968 231301 485974 231313
rect 395114 231273 485974 231301
rect 395114 231261 395120 231273
rect 485968 231261 485974 231273
rect 486026 231261 486032 231313
rect 293488 231187 293494 231239
rect 293546 231227 293552 231239
rect 365584 231227 365590 231239
rect 293546 231199 365590 231227
rect 293546 231187 293552 231199
rect 365584 231187 365590 231199
rect 365642 231187 365648 231239
rect 394768 231187 394774 231239
rect 394826 231227 394832 231239
rect 473872 231227 473878 231239
rect 394826 231199 473878 231227
rect 394826 231187 394832 231199
rect 473872 231187 473878 231199
rect 473930 231187 473936 231239
rect 256144 231113 256150 231165
rect 256202 231153 256208 231165
rect 322096 231153 322102 231165
rect 256202 231125 322102 231153
rect 256202 231113 256208 231125
rect 322096 231113 322102 231125
rect 322154 231113 322160 231165
rect 337360 231113 337366 231165
rect 337418 231153 337424 231165
rect 337418 231125 414686 231153
rect 337418 231113 337424 231125
rect 252976 231039 252982 231091
rect 253034 231079 253040 231091
rect 314512 231079 314518 231091
rect 253034 231051 314518 231079
rect 253034 231039 253040 231051
rect 314512 231039 314518 231051
rect 314570 231039 314576 231091
rect 344464 231039 344470 231091
rect 344522 231079 344528 231091
rect 344522 231051 407534 231079
rect 344522 231039 344528 231051
rect 308176 230965 308182 231017
rect 308234 231005 308240 231017
rect 323632 231005 323638 231017
rect 308234 230977 323638 231005
rect 308234 230965 308240 230977
rect 323632 230965 323638 230977
rect 323690 230965 323696 231017
rect 328336 230965 328342 231017
rect 328394 231005 328400 231017
rect 401392 231005 401398 231017
rect 328394 230977 401398 231005
rect 328394 230965 328400 230977
rect 401392 230965 401398 230977
rect 401450 230965 401456 231017
rect 323152 230891 323158 230943
rect 323210 230931 323216 230943
rect 329584 230931 329590 230943
rect 323210 230903 329590 230931
rect 323210 230891 323216 230903
rect 329584 230891 329590 230903
rect 329642 230891 329648 230943
rect 331216 230891 331222 230943
rect 331274 230931 331280 230943
rect 395344 230931 395350 230943
rect 331274 230903 395350 230931
rect 331274 230891 331280 230903
rect 395344 230891 395350 230903
rect 395402 230891 395408 230943
rect 407506 230931 407534 231051
rect 414658 231005 414686 231125
rect 414736 231113 414742 231165
rect 414794 231153 414800 231165
rect 424048 231153 424054 231165
rect 414794 231125 424054 231153
rect 414794 231113 414800 231125
rect 424048 231113 424054 231125
rect 424106 231113 424112 231165
rect 415696 231005 415702 231017
rect 414658 230977 415702 231005
rect 415696 230965 415702 230977
rect 415754 230965 415760 231017
rect 419536 230931 419542 230943
rect 407506 230903 419542 230931
rect 419536 230891 419542 230903
rect 419594 230891 419600 230943
rect 325744 230817 325750 230869
rect 325802 230857 325808 230869
rect 380272 230857 380278 230869
rect 325802 230829 380278 230857
rect 325802 230817 325808 230829
rect 380272 230817 380278 230829
rect 380330 230817 380336 230869
rect 387280 230817 387286 230869
rect 387338 230857 387344 230869
rect 449680 230857 449686 230869
rect 387338 230829 449686 230857
rect 387338 230817 387344 230829
rect 449680 230817 449686 230829
rect 449738 230817 449744 230869
rect 290704 230743 290710 230795
rect 290762 230783 290768 230795
rect 297328 230783 297334 230795
rect 290762 230755 297334 230783
rect 290762 230743 290768 230755
rect 297328 230743 297334 230755
rect 297386 230743 297392 230795
rect 313936 230743 313942 230795
rect 313994 230783 314000 230795
rect 362128 230783 362134 230795
rect 313994 230755 362134 230783
rect 313994 230743 314000 230755
rect 362128 230743 362134 230755
rect 362186 230743 362192 230795
rect 362320 230743 362326 230795
rect 362378 230783 362384 230795
rect 416464 230783 416470 230795
rect 362378 230755 416470 230783
rect 362378 230743 362384 230755
rect 416464 230743 416470 230755
rect 416522 230743 416528 230795
rect 318256 230669 318262 230721
rect 318314 230709 318320 230721
rect 365104 230709 365110 230721
rect 318314 230681 365110 230709
rect 318314 230669 318320 230681
rect 365104 230669 365110 230681
rect 365162 230669 365168 230721
rect 367120 230669 367126 230721
rect 367178 230709 367184 230721
rect 409648 230709 409654 230721
rect 367178 230681 409654 230709
rect 367178 230669 367184 230681
rect 409648 230669 409654 230681
rect 409706 230669 409712 230721
rect 302320 230595 302326 230647
rect 302378 230635 302384 230647
rect 308560 230635 308566 230647
rect 302378 230607 308566 230635
rect 302378 230595 302384 230607
rect 308560 230595 308566 230607
rect 308618 230595 308624 230647
rect 322192 230595 322198 230647
rect 322250 230635 322256 230647
rect 374128 230635 374134 230647
rect 322250 230607 374134 230635
rect 322250 230595 322256 230607
rect 374128 230595 374134 230607
rect 374186 230595 374192 230647
rect 306736 230521 306742 230573
rect 306794 230561 306800 230573
rect 317584 230561 317590 230573
rect 306794 230533 317590 230561
rect 306794 230521 306800 230533
rect 317584 230521 317590 230533
rect 317642 230521 317648 230573
rect 325360 230521 325366 230573
rect 325418 230561 325424 230573
rect 377104 230561 377110 230573
rect 325418 230533 377110 230561
rect 325418 230521 325424 230533
rect 377104 230521 377110 230533
rect 377162 230521 377168 230573
rect 149392 230447 149398 230499
rect 149450 230487 149456 230499
rect 156976 230487 156982 230499
rect 149450 230459 156982 230487
rect 149450 230447 149456 230459
rect 156976 230447 156982 230459
rect 157034 230447 157040 230499
rect 299248 230447 299254 230499
rect 299306 230487 299312 230499
rect 302512 230487 302518 230499
rect 299306 230459 302518 230487
rect 299306 230447 299312 230459
rect 302512 230447 302518 230459
rect 302570 230447 302576 230499
rect 304144 230447 304150 230499
rect 304202 230487 304208 230499
rect 311632 230487 311638 230499
rect 304202 230459 311638 230487
rect 304202 230447 304208 230459
rect 311632 230447 311638 230459
rect 311690 230447 311696 230499
rect 322000 230447 322006 230499
rect 322058 230487 322064 230499
rect 368176 230487 368182 230499
rect 322058 230459 368182 230487
rect 322058 230447 322064 230459
rect 368176 230447 368182 230459
rect 368234 230447 368240 230499
rect 426160 230447 426166 230499
rect 426218 230487 426224 230499
rect 436144 230487 436150 230499
rect 426218 230459 436150 230487
rect 426218 230447 426224 230459
rect 436144 230447 436150 230459
rect 436202 230447 436208 230499
rect 246160 230373 246166 230425
rect 246218 230413 246224 230425
rect 298672 230413 298678 230425
rect 246218 230385 298678 230413
rect 246218 230373 246224 230385
rect 298672 230373 298678 230385
rect 298730 230373 298736 230425
rect 324016 230373 324022 230425
rect 324074 230413 324080 230425
rect 346960 230413 346966 230425
rect 324074 230385 346966 230413
rect 324074 230373 324080 230385
rect 346960 230373 346966 230385
rect 347018 230373 347024 230425
rect 369904 230373 369910 230425
rect 369962 230413 369968 230425
rect 387280 230413 387286 230425
rect 369962 230385 387286 230413
rect 369962 230373 369968 230385
rect 387280 230373 387286 230385
rect 387338 230373 387344 230425
rect 434896 230373 434902 230425
rect 434954 230413 434960 230425
rect 454288 230413 454294 230425
rect 434954 230385 454294 230413
rect 434954 230373 434960 230385
rect 454288 230373 454294 230385
rect 454346 230373 454352 230425
rect 245776 230299 245782 230351
rect 245834 230339 245840 230351
rect 300976 230339 300982 230351
rect 245834 230311 300982 230339
rect 245834 230299 245840 230311
rect 300976 230299 300982 230311
rect 301034 230299 301040 230351
rect 314896 230299 314902 230351
rect 314954 230339 314960 230351
rect 439984 230339 439990 230351
rect 314954 230311 439990 230339
rect 314954 230299 314960 230311
rect 439984 230299 439990 230311
rect 440042 230299 440048 230351
rect 248944 230225 248950 230277
rect 249002 230265 249008 230277
rect 304816 230265 304822 230277
rect 249002 230237 304822 230265
rect 249002 230225 249008 230237
rect 304816 230225 304822 230237
rect 304874 230225 304880 230277
rect 317968 230225 317974 230277
rect 318026 230265 318032 230277
rect 445936 230265 445942 230277
rect 318026 230237 445942 230265
rect 318026 230225 318032 230237
rect 445936 230225 445942 230237
rect 445994 230225 446000 230277
rect 247024 230151 247030 230203
rect 247082 230191 247088 230203
rect 303952 230191 303958 230203
rect 247082 230163 303958 230191
rect 247082 230151 247088 230163
rect 303952 230151 303958 230163
rect 304010 230151 304016 230203
rect 313456 230151 313462 230203
rect 313514 230191 313520 230203
rect 436912 230191 436918 230203
rect 313514 230163 436918 230191
rect 313514 230151 313520 230163
rect 436912 230151 436918 230163
rect 436970 230151 436976 230203
rect 449296 230151 449302 230203
rect 449354 230191 449360 230203
rect 466384 230191 466390 230203
rect 449354 230163 466390 230191
rect 449354 230151 449360 230163
rect 466384 230151 466390 230163
rect 466442 230151 466448 230203
rect 248752 230077 248758 230129
rect 248810 230117 248816 230129
rect 307024 230117 307030 230129
rect 248810 230089 307030 230117
rect 248810 230077 248816 230089
rect 307024 230077 307030 230089
rect 307082 230077 307088 230129
rect 325840 230077 325846 230129
rect 325898 230117 325904 230129
rect 461008 230117 461014 230129
rect 325898 230089 461014 230117
rect 325898 230077 325904 230089
rect 461008 230077 461014 230089
rect 461066 230077 461072 230129
rect 463600 230077 463606 230129
rect 463658 230117 463664 230129
rect 478384 230117 478390 230129
rect 463658 230089 478390 230117
rect 463658 230077 463664 230089
rect 478384 230077 478390 230089
rect 478442 230077 478448 230129
rect 251920 230003 251926 230055
rect 251978 230043 251984 230055
rect 310768 230043 310774 230055
rect 251978 230015 310774 230043
rect 251978 230003 251984 230015
rect 310768 230003 310774 230015
rect 310826 230003 310832 230055
rect 328528 230003 328534 230055
rect 328586 230043 328592 230055
rect 328586 230015 341534 230043
rect 328586 230003 328592 230015
rect 251536 229929 251542 229981
rect 251594 229969 251600 229981
rect 313072 229969 313078 229981
rect 251594 229941 313078 229969
rect 251594 229929 251600 229941
rect 313072 229929 313078 229941
rect 313130 229929 313136 229981
rect 331600 229929 331606 229981
rect 331658 229969 331664 229981
rect 341506 229969 341534 230015
rect 346960 230003 346966 230055
rect 347018 230043 347024 230055
rect 458032 230043 458038 230055
rect 347018 230015 458038 230043
rect 347018 230003 347024 230015
rect 458032 230003 458038 230015
rect 458090 230003 458096 230055
rect 466480 230003 466486 230055
rect 466538 230043 466544 230055
rect 484432 230043 484438 230055
rect 466538 230015 484438 230043
rect 466538 230003 466544 230015
rect 484432 230003 484438 230015
rect 484490 230003 484496 230055
rect 503920 230003 503926 230055
rect 503978 230043 503984 230055
rect 622672 230043 622678 230055
rect 503978 230015 622678 230043
rect 503978 230003 503984 230015
rect 622672 230003 622678 230015
rect 622730 230003 622736 230055
rect 467056 229969 467062 229981
rect 331658 229941 336974 229969
rect 341506 229941 467062 229969
rect 331658 229929 331664 229941
rect 227440 229855 227446 229907
rect 227498 229895 227504 229907
rect 264784 229895 264790 229907
rect 227498 229867 264790 229895
rect 227498 229855 227504 229867
rect 264784 229855 264790 229867
rect 264842 229855 264848 229907
rect 290896 229855 290902 229907
rect 290954 229895 290960 229907
rect 331888 229895 331894 229907
rect 290954 229867 331894 229895
rect 290954 229855 290960 229867
rect 331888 229855 331894 229867
rect 331946 229855 331952 229907
rect 336946 229895 336974 229941
rect 467056 229929 467062 229941
rect 467114 229929 467120 229981
rect 475216 229929 475222 229981
rect 475274 229969 475280 229981
rect 601456 229969 601462 229981
rect 475274 229941 601462 229969
rect 475274 229929 475280 229941
rect 601456 229929 601462 229941
rect 601514 229929 601520 229981
rect 473104 229895 473110 229907
rect 336946 229867 473110 229895
rect 473104 229855 473110 229867
rect 473162 229855 473168 229907
rect 480880 229855 480886 229907
rect 480938 229895 480944 229907
rect 609040 229895 609046 229907
rect 480938 229867 609046 229895
rect 480938 229855 480944 229867
rect 609040 229855 609046 229867
rect 609098 229855 609104 229907
rect 254800 229781 254806 229833
rect 254858 229821 254864 229833
rect 319120 229821 319126 229833
rect 254858 229793 319126 229821
rect 254858 229781 254864 229793
rect 319120 229781 319126 229793
rect 319178 229781 319184 229833
rect 336304 229781 336310 229833
rect 336362 229821 336368 229833
rect 482128 229821 482134 229833
rect 336362 229793 482134 229821
rect 336362 229781 336368 229793
rect 482128 229781 482134 229793
rect 482186 229781 482192 229833
rect 484624 229781 484630 229833
rect 484682 229821 484688 229833
rect 612112 229821 612118 229833
rect 484682 229793 612118 229821
rect 484682 229781 484688 229793
rect 612112 229781 612118 229793
rect 612170 229781 612176 229833
rect 220144 229707 220150 229759
rect 220202 229747 220208 229759
rect 249712 229747 249718 229759
rect 220202 229719 249718 229747
rect 220202 229707 220208 229719
rect 249712 229707 249718 229719
rect 249770 229707 249776 229759
rect 253072 229707 253078 229759
rect 253130 229747 253136 229759
rect 316144 229747 316150 229759
rect 253130 229719 316150 229747
rect 253130 229707 253136 229719
rect 316144 229707 316150 229719
rect 316202 229707 316208 229759
rect 348496 229707 348502 229759
rect 348554 229747 348560 229759
rect 504016 229747 504022 229759
rect 348554 229719 504022 229747
rect 348554 229707 348560 229719
rect 504016 229707 504022 229719
rect 504074 229707 504080 229759
rect 244240 229633 244246 229685
rect 244298 229673 244304 229685
rect 298000 229673 298006 229685
rect 244298 229645 298006 229673
rect 244298 229633 244304 229645
rect 298000 229633 298006 229645
rect 298058 229633 298064 229685
rect 298576 229633 298582 229685
rect 298634 229673 298640 229685
rect 406768 229673 406774 229685
rect 298634 229645 406774 229673
rect 298634 229633 298640 229645
rect 406768 229633 406774 229645
rect 406826 229633 406832 229685
rect 409840 229633 409846 229685
rect 409898 229673 409904 229685
rect 565936 229673 565942 229685
rect 409898 229645 565942 229673
rect 409898 229633 409904 229645
rect 565936 229633 565942 229645
rect 565994 229633 566000 229685
rect 221584 229559 221590 229611
rect 221642 229599 221648 229611
rect 252592 229599 252598 229611
rect 221642 229571 252598 229599
rect 221642 229559 221648 229571
rect 252592 229559 252598 229571
rect 252650 229559 252656 229611
rect 255184 229559 255190 229611
rect 255242 229599 255248 229611
rect 316816 229599 316822 229611
rect 255242 229571 316822 229599
rect 255242 229559 255248 229571
rect 316816 229559 316822 229571
rect 316874 229559 316880 229611
rect 351760 229559 351766 229611
rect 351818 229599 351824 229611
rect 510160 229599 510166 229611
rect 351818 229571 510166 229599
rect 351818 229559 351824 229571
rect 510160 229559 510166 229571
rect 510218 229559 510224 229611
rect 264304 229485 264310 229537
rect 264362 229525 264368 229537
rect 334960 229525 334966 229537
rect 264362 229497 334966 229525
rect 264362 229485 264368 229497
rect 334960 229485 334966 229497
rect 335018 229485 335024 229537
rect 354832 229485 354838 229537
rect 354890 229525 354896 229537
rect 516112 229525 516118 229537
rect 354890 229497 516118 229525
rect 354890 229485 354896 229497
rect 516112 229485 516118 229497
rect 516170 229485 516176 229537
rect 228880 229411 228886 229463
rect 228938 229451 228944 229463
rect 267856 229451 267862 229463
rect 228938 229423 267862 229451
rect 228938 229411 228944 229423
rect 267856 229411 267862 229423
rect 267914 229411 267920 229463
rect 283504 229411 283510 229463
rect 283562 229451 283568 229463
rect 368848 229451 368854 229463
rect 283562 229423 368854 229451
rect 283562 229411 283568 229423
rect 368848 229411 368854 229423
rect 368906 229411 368912 229463
rect 380080 229411 380086 229463
rect 380138 229451 380144 229463
rect 538864 229451 538870 229463
rect 380138 229423 538870 229451
rect 380138 229411 380144 229423
rect 538864 229411 538870 229423
rect 538922 229411 538928 229463
rect 230320 229337 230326 229389
rect 230378 229377 230384 229389
rect 269296 229377 269302 229389
rect 230378 229349 269302 229377
rect 230378 229337 230384 229349
rect 269296 229337 269302 229349
rect 269354 229337 269360 229389
rect 273520 229337 273526 229389
rect 273578 229377 273584 229389
rect 347056 229377 347062 229389
rect 273578 229349 347062 229377
rect 273578 229337 273584 229349
rect 347056 229337 347062 229349
rect 347114 229337 347120 229389
rect 357616 229337 357622 229389
rect 357674 229377 357680 229389
rect 522160 229377 522166 229389
rect 357674 229349 522166 229377
rect 357674 229337 357680 229349
rect 522160 229337 522166 229349
rect 522218 229337 522224 229389
rect 233488 229263 233494 229315
rect 233546 229303 233552 229315
rect 276784 229303 276790 229315
rect 233546 229275 276790 229303
rect 233546 229263 233552 229275
rect 276784 229263 276790 229275
rect 276842 229263 276848 229315
rect 284752 229263 284758 229315
rect 284810 229303 284816 229315
rect 284810 229275 294110 229303
rect 284810 229263 284816 229275
rect 146896 229189 146902 229241
rect 146954 229229 146960 229241
rect 151312 229229 151318 229241
rect 146954 229201 151318 229229
rect 146954 229189 146960 229201
rect 151312 229189 151318 229201
rect 151370 229189 151376 229241
rect 231952 229189 231958 229241
rect 232010 229229 232016 229241
rect 273808 229229 273814 229241
rect 232010 229201 273814 229229
rect 232010 229189 232016 229201
rect 273808 229189 273814 229201
rect 273866 229189 273872 229241
rect 286288 229189 286294 229241
rect 286346 229229 286352 229241
rect 293968 229229 293974 229241
rect 286346 229201 293974 229229
rect 286346 229189 286352 229201
rect 293968 229189 293974 229201
rect 294026 229189 294032 229241
rect 294082 229229 294110 229275
rect 294160 229263 294166 229315
rect 294218 229303 294224 229315
rect 371248 229303 371254 229315
rect 294218 229275 371254 229303
rect 294218 229263 294224 229275
rect 371248 229263 371254 229275
rect 371306 229263 371312 229315
rect 374224 229263 374230 229315
rect 374282 229303 374288 229315
rect 374282 229275 377294 229303
rect 374282 229263 374288 229275
rect 371536 229229 371542 229241
rect 294082 229201 371542 229229
rect 371536 229189 371542 229201
rect 371594 229189 371600 229241
rect 377266 229229 377294 229275
rect 387280 229263 387286 229315
rect 387338 229303 387344 229315
rect 546352 229303 546358 229315
rect 387338 229275 546358 229303
rect 387338 229263 387344 229275
rect 546352 229263 546358 229275
rect 546410 229263 546416 229315
rect 555280 229229 555286 229241
rect 377266 229201 555286 229229
rect 555280 229189 555286 229201
rect 555338 229189 555344 229241
rect 235216 229115 235222 229167
rect 235274 229155 235280 229167
rect 279856 229155 279862 229167
rect 235274 229127 279862 229155
rect 235274 229115 235280 229127
rect 279856 229115 279862 229127
rect 279914 229115 279920 229167
rect 287920 229115 287926 229167
rect 287978 229155 287984 229167
rect 374416 229155 374422 229167
rect 287978 229127 374422 229155
rect 287978 229115 287984 229127
rect 374416 229115 374422 229127
rect 374474 229115 374480 229167
rect 377200 229115 377206 229167
rect 377258 229155 377264 229167
rect 561424 229155 561430 229167
rect 377258 229127 561430 229155
rect 377258 229115 377264 229127
rect 561424 229115 561430 229127
rect 561482 229115 561488 229167
rect 238384 229041 238390 229093
rect 238442 229081 238448 229093
rect 283600 229081 283606 229093
rect 238442 229053 283606 229081
rect 238442 229041 238448 229053
rect 283600 229041 283606 229053
rect 283658 229041 283664 229093
rect 291184 229041 291190 229093
rect 291242 229081 291248 229093
rect 291242 229053 293918 229081
rect 291242 229041 291248 229053
rect 215248 228967 215254 229019
rect 215306 229007 215312 229019
rect 239056 229007 239062 229019
rect 215306 228979 239062 229007
rect 215306 228967 215312 228979
rect 239056 228967 239062 228979
rect 239114 228967 239120 229019
rect 241072 228967 241078 229019
rect 241130 229007 241136 229019
rect 291952 229007 291958 229019
rect 241130 228979 291958 229007
rect 241130 228967 241136 228979
rect 291952 228967 291958 228979
rect 292010 228967 292016 229019
rect 293890 229007 293918 229053
rect 293968 229041 293974 229093
rect 294026 229081 294032 229093
rect 374512 229081 374518 229093
rect 294026 229053 374518 229081
rect 294026 229041 294032 229053
rect 374512 229041 374518 229053
rect 374570 229041 374576 229093
rect 376816 229041 376822 229093
rect 376874 229081 376880 229093
rect 563632 229081 563638 229093
rect 376874 229053 563638 229081
rect 376874 229041 376880 229053
rect 563632 229041 563638 229053
rect 563690 229041 563696 229093
rect 382864 229007 382870 229019
rect 293890 228979 382870 229007
rect 382864 228967 382870 228979
rect 382922 228967 382928 229019
rect 382960 228967 382966 229019
rect 383018 229007 383024 229019
rect 567376 229007 567382 229019
rect 383018 228979 567382 229007
rect 383018 228967 383024 228979
rect 567376 228967 567382 228979
rect 567434 228967 567440 229019
rect 242512 228893 242518 228945
rect 242570 228933 242576 228945
rect 294928 228933 294934 228945
rect 242570 228905 294934 228933
rect 242570 228893 242576 228905
rect 294928 228893 294934 228905
rect 294986 228893 294992 228945
rect 308944 228893 308950 228945
rect 309002 228933 309008 228945
rect 427792 228933 427798 228945
rect 309002 228905 427798 228933
rect 309002 228893 309008 228905
rect 427792 228893 427798 228905
rect 427850 228893 427856 228945
rect 427888 228893 427894 228945
rect 427946 228933 427952 228945
rect 547888 228933 547894 228945
rect 427946 228905 547894 228933
rect 427946 228893 427952 228905
rect 547888 228893 547894 228905
rect 547946 228893 547952 228945
rect 239728 228819 239734 228871
rect 239786 228859 239792 228871
rect 288880 228859 288886 228871
rect 239786 228831 288886 228859
rect 239786 228819 239792 228831
rect 288880 228819 288886 228831
rect 288938 228819 288944 228871
rect 294160 228859 294166 228871
rect 289282 228831 294166 228859
rect 241648 228745 241654 228797
rect 241706 228785 241712 228797
rect 241706 228757 276494 228785
rect 241706 228745 241712 228757
rect 231856 228671 231862 228723
rect 231914 228711 231920 228723
rect 272272 228711 272278 228723
rect 231914 228683 272278 228711
rect 231914 228671 231920 228683
rect 272272 228671 272278 228683
rect 272330 228671 272336 228723
rect 230608 228597 230614 228649
rect 230666 228637 230672 228649
rect 270736 228637 270742 228649
rect 230666 228609 270742 228637
rect 230666 228597 230672 228609
rect 270736 228597 270742 228609
rect 270794 228597 270800 228649
rect 276466 228637 276494 228757
rect 282160 228671 282166 228723
rect 282218 228711 282224 228723
rect 289282 228711 289310 228831
rect 294160 228819 294166 228831
rect 294218 228819 294224 228871
rect 310672 228819 310678 228871
rect 310730 228859 310736 228871
rect 430864 228859 430870 228871
rect 310730 228831 430870 228859
rect 310730 228819 310736 228831
rect 430864 228819 430870 228831
rect 430922 228819 430928 228871
rect 432016 228819 432022 228871
rect 432074 228859 432080 228871
rect 529744 228859 529750 228871
rect 432074 228831 529750 228859
rect 432074 228819 432080 228831
rect 529744 228819 529750 228831
rect 529802 228819 529808 228871
rect 304432 228745 304438 228797
rect 304490 228785 304496 228797
rect 418768 228785 418774 228797
rect 304490 228757 418774 228785
rect 304490 228745 304496 228757
rect 418768 228745 418774 228757
rect 418826 228745 418832 228797
rect 282218 228683 289310 228711
rect 282218 228671 282224 228683
rect 289360 228671 289366 228723
rect 289418 228711 289424 228723
rect 289418 228683 296654 228711
rect 289418 228671 289424 228683
rect 289744 228637 289750 228649
rect 276466 228609 289750 228637
rect 289744 228597 289750 228609
rect 289802 228597 289808 228649
rect 293872 228597 293878 228649
rect 293930 228637 293936 228649
rect 295792 228637 295798 228649
rect 293930 228609 295798 228637
rect 293930 228597 293936 228609
rect 295792 228597 295798 228609
rect 295850 228597 295856 228649
rect 296626 228637 296654 228683
rect 306160 228671 306166 228723
rect 306218 228711 306224 228723
rect 421840 228711 421846 228723
rect 306218 228683 421846 228711
rect 306218 228671 306224 228683
rect 421840 228671 421846 228683
rect 421898 228671 421904 228723
rect 380080 228637 380086 228649
rect 296626 228609 380086 228637
rect 380080 228597 380086 228609
rect 380138 228597 380144 228649
rect 407344 228597 407350 228649
rect 407402 228637 407408 228649
rect 517648 228637 517654 228649
rect 407402 228609 517654 228637
rect 407402 228597 407408 228609
rect 517648 228597 517654 228609
rect 517706 228597 517712 228649
rect 190192 228523 190198 228575
rect 190250 228563 190256 228575
rect 192304 228563 192310 228575
rect 190250 228535 192310 228563
rect 190250 228523 190256 228535
rect 192304 228523 192310 228535
rect 192362 228523 192368 228575
rect 228784 228523 228790 228575
rect 228842 228563 228848 228575
rect 266224 228563 266230 228575
rect 228842 228535 266230 228563
rect 228842 228523 228848 228535
rect 266224 228523 266230 228535
rect 266282 228523 266288 228575
rect 266320 228523 266326 228575
rect 266378 228563 266384 228575
rect 301744 228563 301750 228575
rect 266378 228535 301750 228563
rect 266378 228523 266384 228535
rect 301744 228523 301750 228535
rect 301802 228523 301808 228575
rect 303472 228523 303478 228575
rect 303530 228563 303536 228575
rect 413488 228563 413494 228575
rect 303530 228535 413494 228563
rect 303530 228523 303536 228535
rect 413488 228523 413494 228535
rect 413546 228523 413552 228575
rect 455056 228523 455062 228575
rect 455114 228563 455120 228575
rect 456496 228563 456502 228575
rect 455114 228535 456502 228563
rect 455114 228523 455120 228535
rect 456496 228523 456502 228535
rect 456554 228523 456560 228575
rect 535792 228523 535798 228575
rect 535850 228563 535856 228575
rect 538000 228563 538006 228575
rect 535850 228535 538006 228563
rect 535850 228523 535856 228535
rect 538000 228523 538006 228535
rect 538058 228523 538064 228575
rect 544336 228523 544342 228575
rect 544394 228563 544400 228575
rect 547120 228563 547126 228575
rect 544394 228535 547126 228563
rect 544394 228523 544400 228535
rect 547120 228523 547126 228535
rect 547178 228523 547184 228575
rect 556144 228523 556150 228575
rect 556202 228563 556208 228575
rect 558448 228563 558454 228575
rect 556202 228535 558454 228563
rect 556202 228523 556208 228535
rect 558448 228523 558454 228535
rect 558506 228523 558512 228575
rect 224368 228449 224374 228501
rect 224426 228489 224432 228501
rect 258736 228489 258742 228501
rect 224426 228461 258742 228489
rect 224426 228449 224432 228461
rect 258736 228449 258742 228461
rect 258794 228449 258800 228501
rect 270832 228449 270838 228501
rect 270890 228489 270896 228501
rect 313840 228489 313846 228501
rect 270890 228461 313846 228489
rect 270890 228449 270896 228461
rect 313840 228449 313846 228461
rect 313898 228449 313904 228501
rect 317872 228449 317878 228501
rect 317930 228489 317936 228501
rect 403696 228489 403702 228501
rect 317930 228461 403702 228489
rect 317930 228449 317936 228461
rect 403696 228449 403702 228461
rect 403754 228449 403760 228501
rect 405328 228449 405334 228501
rect 405386 228489 405392 228501
rect 502576 228489 502582 228501
rect 405386 228461 502582 228489
rect 405386 228449 405392 228461
rect 502576 228449 502582 228461
rect 502634 228449 502640 228501
rect 264880 228375 264886 228427
rect 264938 228415 264944 228427
rect 295696 228415 295702 228427
rect 264938 228387 295702 228415
rect 264938 228375 264944 228387
rect 295696 228375 295702 228387
rect 295754 228375 295760 228427
rect 295792 228375 295798 228427
rect 295850 228415 295856 228427
rect 382960 228415 382966 228427
rect 295850 228387 382966 228415
rect 295850 228375 295856 228387
rect 382960 228375 382966 228387
rect 383018 228375 383024 228427
rect 391696 228375 391702 228427
rect 391754 228415 391760 228427
rect 476944 228415 476950 228427
rect 391754 228387 476950 228415
rect 391754 228375 391760 228387
rect 476944 228375 476950 228387
rect 477002 228375 477008 228427
rect 535792 228375 535798 228427
rect 535850 228415 535856 228427
rect 537904 228415 537910 228427
rect 535850 228387 537910 228415
rect 535850 228375 535856 228387
rect 537904 228375 537910 228387
rect 537962 228375 537968 228427
rect 267952 228301 267958 228353
rect 268010 228341 268016 228353
rect 307696 228341 307702 228353
rect 268010 228313 307702 228341
rect 268010 228301 268016 228313
rect 307696 228301 307702 228313
rect 307754 228301 307760 228353
rect 311152 228301 311158 228353
rect 311210 228341 311216 228353
rect 392368 228341 392374 228353
rect 311210 228313 392374 228341
rect 311210 228301 311216 228313
rect 392368 228301 392374 228313
rect 392426 228301 392432 228353
rect 392464 228301 392470 228353
rect 392522 228341 392528 228353
rect 461872 228341 461878 228353
rect 392522 228313 461878 228341
rect 392522 228301 392528 228313
rect 461872 228301 461878 228313
rect 461930 228301 461936 228353
rect 261136 228227 261142 228279
rect 261194 228267 261200 228279
rect 292624 228267 292630 228279
rect 261194 228239 292630 228267
rect 261194 228227 261200 228239
rect 292624 228227 292630 228239
rect 292682 228227 292688 228279
rect 311056 228227 311062 228279
rect 311114 228267 311120 228279
rect 383248 228267 383254 228279
rect 311114 228239 383254 228267
rect 311114 228227 311120 228239
rect 383248 228227 383254 228239
rect 383306 228227 383312 228279
rect 394672 228227 394678 228279
rect 394730 228267 394736 228279
rect 437680 228267 437686 228279
rect 394730 228239 437686 228267
rect 394730 228227 394736 228239
rect 437680 228227 437686 228239
rect 437738 228227 437744 228279
rect 269104 228153 269110 228205
rect 269162 228193 269168 228205
rect 322960 228193 322966 228205
rect 269162 228165 322966 228193
rect 269162 228153 269168 228165
rect 322960 228153 322966 228165
rect 323018 228153 323024 228205
rect 344080 228153 344086 228205
rect 344138 228193 344144 228205
rect 412720 228193 412726 228205
rect 344138 228165 412726 228193
rect 344138 228153 344144 228165
rect 412720 228153 412726 228165
rect 412778 228153 412784 228205
rect 250576 228079 250582 228131
rect 250634 228119 250640 228131
rect 277552 228119 277558 228131
rect 250634 228091 277558 228119
rect 250634 228079 250640 228091
rect 277552 228079 277558 228091
rect 277610 228079 277616 228131
rect 290992 228079 290998 228131
rect 291050 228119 291056 228131
rect 341008 228119 341014 228131
rect 291050 228091 341014 228119
rect 291050 228079 291056 228091
rect 341008 228079 341014 228091
rect 341066 228079 341072 228131
rect 341200 228079 341206 228131
rect 341258 228119 341264 228131
rect 398320 228119 398326 228131
rect 341258 228091 398326 228119
rect 341258 228079 341264 228091
rect 398320 228079 398326 228091
rect 398378 228079 398384 228131
rect 260944 228005 260950 228057
rect 261002 228045 261008 228057
rect 286672 228045 286678 228057
rect 261002 228017 286678 228045
rect 261002 228005 261008 228017
rect 286672 228005 286678 228017
rect 286730 228005 286736 228057
rect 305104 228005 305110 228057
rect 305162 228045 305168 228057
rect 310096 228045 310102 228057
rect 305162 228017 310102 228045
rect 305162 228005 305168 228017
rect 310096 228005 310102 228017
rect 310154 228005 310160 228057
rect 310192 228005 310198 228057
rect 310250 228045 310256 228057
rect 310250 228017 357134 228045
rect 310250 228005 310256 228017
rect 258928 227931 258934 227983
rect 258986 227971 258992 227983
rect 280624 227971 280630 227983
rect 258986 227943 280630 227971
rect 258986 227931 258992 227943
rect 280624 227931 280630 227943
rect 280682 227931 280688 227983
rect 293776 227931 293782 227983
rect 293834 227971 293840 227983
rect 343984 227971 343990 227983
rect 293834 227943 343990 227971
rect 293834 227931 293840 227943
rect 343984 227931 343990 227943
rect 344042 227931 344048 227983
rect 357106 227971 357134 228017
rect 357520 228005 357526 228057
rect 357578 228045 357584 228057
rect 359920 228045 359926 228057
rect 357578 228017 359926 228045
rect 357578 228005 357584 228017
rect 359920 228005 359926 228017
rect 359978 228005 359984 228057
rect 368944 228005 368950 228057
rect 369002 228045 369008 228057
rect 370480 228045 370486 228057
rect 369002 228017 370486 228045
rect 369002 228005 369008 228017
rect 370480 228005 370486 228017
rect 370538 228005 370544 228057
rect 370576 228005 370582 228057
rect 370634 228045 370640 228057
rect 425584 228045 425590 228057
rect 370634 228017 425590 228045
rect 370634 228005 370640 228017
rect 425584 228005 425590 228017
rect 425642 228005 425648 228057
rect 359152 227971 359158 227983
rect 357106 227943 359158 227971
rect 359152 227931 359158 227943
rect 359210 227931 359216 227983
rect 302128 227857 302134 227909
rect 302186 227897 302192 227909
rect 350032 227897 350038 227909
rect 302186 227869 350038 227897
rect 302186 227857 302192 227869
rect 350032 227857 350038 227869
rect 350090 227857 350096 227909
rect 250192 227783 250198 227835
rect 250250 227823 250256 227835
rect 310000 227823 310006 227835
rect 250250 227795 310006 227823
rect 250250 227783 250256 227795
rect 310000 227783 310006 227795
rect 310058 227783 310064 227835
rect 310096 227783 310102 227835
rect 310154 227823 310160 227835
rect 353104 227823 353110 227835
rect 310154 227795 353110 227823
rect 310154 227783 310160 227795
rect 353104 227783 353110 227795
rect 353162 227783 353168 227835
rect 281200 227709 281206 227761
rect 281258 227749 281264 227761
rect 325840 227749 325846 227761
rect 281258 227721 325846 227749
rect 281258 227709 281264 227721
rect 325840 227709 325846 227721
rect 325898 227709 325904 227761
rect 279280 227635 279286 227687
rect 279338 227675 279344 227687
rect 319888 227675 319894 227687
rect 279338 227647 319894 227675
rect 279338 227635 279344 227647
rect 319888 227635 319894 227647
rect 319946 227635 319952 227687
rect 321232 227635 321238 227687
rect 321290 227675 321296 227687
rect 451984 227675 451990 227687
rect 321290 227647 451990 227675
rect 321290 227635 321296 227647
rect 451984 227635 451990 227647
rect 452042 227635 452048 227687
rect 149392 227561 149398 227613
rect 149450 227601 149456 227613
rect 174256 227601 174262 227613
rect 149450 227573 174262 227601
rect 149450 227561 149456 227573
rect 174256 227561 174262 227573
rect 174314 227561 174320 227613
rect 288016 227561 288022 227613
rect 288074 227601 288080 227613
rect 328912 227601 328918 227613
rect 288074 227573 328918 227601
rect 288074 227561 288080 227573
rect 328912 227561 328918 227573
rect 328970 227561 328976 227613
rect 387760 227561 387766 227613
rect 387818 227601 387824 227613
rect 396400 227601 396406 227613
rect 387818 227573 396406 227601
rect 387818 227561 387824 227573
rect 396400 227561 396406 227573
rect 396458 227561 396464 227613
rect 423280 227561 423286 227613
rect 423338 227601 423344 227613
rect 433168 227601 433174 227613
rect 423338 227573 433174 227601
rect 423338 227561 423344 227573
rect 433168 227561 433174 227573
rect 433226 227561 433232 227613
rect 187120 227487 187126 227539
rect 187178 227527 187184 227539
rect 190768 227527 190774 227539
rect 187178 227499 190774 227527
rect 187178 227487 187184 227499
rect 190768 227487 190774 227499
rect 190826 227487 190832 227539
rect 217456 227487 217462 227539
rect 217514 227527 217520 227539
rect 241264 227527 241270 227539
rect 217514 227499 241270 227527
rect 217514 227487 217520 227499
rect 241264 227487 241270 227499
rect 241322 227487 241328 227539
rect 244720 227487 244726 227539
rect 244778 227527 244784 227539
rect 254896 227527 254902 227539
rect 244778 227499 254902 227527
rect 244778 227487 244784 227499
rect 254896 227487 254902 227499
rect 254954 227487 254960 227539
rect 306256 227527 306262 227539
rect 255106 227499 306262 227527
rect 215728 227413 215734 227465
rect 215786 227453 215792 227465
rect 238384 227453 238390 227465
rect 215786 227425 238390 227453
rect 215786 227413 215792 227425
rect 238384 227413 238390 227425
rect 238442 227413 238448 227465
rect 217072 227339 217078 227391
rect 217130 227379 217136 227391
rect 243568 227379 243574 227391
rect 217130 227351 243574 227379
rect 217130 227339 217136 227351
rect 243568 227339 243574 227351
rect 243626 227339 243632 227391
rect 249328 227339 249334 227391
rect 249386 227379 249392 227391
rect 255106 227379 255134 227499
rect 306256 227487 306262 227499
rect 306314 227487 306320 227539
rect 311344 227487 311350 227539
rect 311402 227527 311408 227539
rect 375760 227527 375766 227539
rect 311402 227499 375766 227527
rect 311402 227487 311408 227499
rect 375760 227487 375766 227499
rect 375818 227487 375824 227539
rect 388912 227487 388918 227539
rect 388970 227527 388976 227539
rect 586384 227527 586390 227539
rect 388970 227499 586390 227527
rect 388970 227487 388976 227499
rect 586384 227487 586390 227499
rect 586442 227487 586448 227539
rect 591472 227487 591478 227539
rect 591530 227527 591536 227539
rect 594640 227527 594646 227539
rect 591530 227499 594646 227527
rect 591530 227487 591536 227499
rect 594640 227487 594646 227499
rect 594698 227487 594704 227539
rect 606256 227487 606262 227539
rect 606314 227527 606320 227539
rect 606314 227499 619214 227527
rect 606314 227487 606320 227499
rect 256240 227413 256246 227465
rect 256298 227453 256304 227465
rect 315376 227453 315382 227465
rect 256298 227425 315382 227453
rect 256298 227413 256304 227425
rect 315376 227413 315382 227425
rect 315434 227413 315440 227465
rect 318448 227413 318454 227465
rect 318506 227453 318512 227465
rect 381808 227453 381814 227465
rect 318506 227425 381814 227453
rect 318506 227413 318512 227425
rect 381808 227413 381814 227425
rect 381866 227413 381872 227465
rect 388528 227413 388534 227465
rect 388586 227453 388592 227465
rect 585616 227453 585622 227465
rect 388586 227425 585622 227453
rect 388586 227413 388592 227425
rect 585616 227413 585622 227425
rect 585674 227413 585680 227465
rect 587632 227413 587638 227465
rect 587690 227453 587696 227465
rect 600784 227453 600790 227465
rect 587690 227425 600790 227453
rect 587690 227413 587696 227425
rect 600784 227413 600790 227425
rect 600842 227413 600848 227465
rect 619186 227453 619214 227499
rect 629296 227487 629302 227539
rect 629354 227527 629360 227539
rect 634000 227527 634006 227539
rect 629354 227499 634006 227527
rect 629354 227487 629360 227499
rect 634000 227487 634006 227499
rect 634058 227487 634064 227539
rect 639184 227453 639190 227465
rect 619186 227425 639190 227453
rect 639184 227413 639190 227425
rect 639242 227413 639248 227465
rect 249386 227351 255134 227379
rect 249386 227339 249392 227351
rect 278032 227339 278038 227391
rect 278090 227379 278096 227391
rect 279280 227379 279286 227391
rect 278090 227351 279286 227379
rect 278090 227339 278096 227351
rect 279280 227339 279286 227351
rect 279338 227339 279344 227391
rect 311248 227339 311254 227391
rect 311306 227379 311312 227391
rect 384016 227379 384022 227391
rect 311306 227351 384022 227379
rect 311306 227339 311312 227351
rect 384016 227339 384022 227351
rect 384074 227339 384080 227391
rect 390448 227339 390454 227391
rect 390506 227379 390512 227391
rect 589360 227379 589366 227391
rect 390506 227351 589366 227379
rect 390506 227339 390512 227351
rect 589360 227339 589366 227351
rect 589418 227339 589424 227391
rect 590416 227339 590422 227391
rect 590474 227379 590480 227391
rect 627856 227379 627862 227391
rect 590474 227351 627862 227379
rect 590474 227339 590480 227351
rect 627856 227339 627862 227351
rect 627914 227339 627920 227391
rect 219472 227265 219478 227317
rect 219530 227305 219536 227317
rect 245872 227305 245878 227317
rect 219530 227277 245878 227305
rect 219530 227265 219536 227277
rect 245872 227265 245878 227277
rect 245930 227265 245936 227317
rect 275056 227265 275062 227317
rect 275114 227305 275120 227317
rect 348592 227305 348598 227317
rect 275114 227277 348598 227305
rect 275114 227265 275120 227277
rect 348592 227265 348598 227277
rect 348650 227265 348656 227317
rect 390064 227265 390070 227317
rect 390122 227305 390128 227317
rect 390122 227277 395294 227305
rect 390122 227265 390128 227277
rect 217840 227191 217846 227243
rect 217898 227231 217904 227243
rect 242896 227231 242902 227243
rect 217898 227203 242902 227231
rect 217898 227191 217904 227203
rect 242896 227191 242902 227203
rect 242954 227191 242960 227243
rect 271984 227191 271990 227243
rect 272042 227231 272048 227243
rect 351568 227231 351574 227243
rect 272042 227203 351574 227231
rect 272042 227191 272048 227203
rect 351568 227191 351574 227203
rect 351626 227191 351632 227243
rect 365584 227191 365590 227243
rect 365642 227231 365648 227243
rect 367120 227231 367126 227243
rect 365642 227203 367126 227231
rect 365642 227191 365648 227203
rect 367120 227191 367126 227203
rect 367178 227191 367184 227243
rect 390832 227191 390838 227243
rect 390890 227231 390896 227243
rect 395266 227231 395294 227277
rect 396400 227265 396406 227317
rect 396458 227305 396464 227317
rect 407440 227305 407446 227317
rect 396458 227277 407446 227305
rect 396458 227265 396464 227277
rect 407440 227265 407446 227277
rect 407498 227265 407504 227317
rect 587440 227265 587446 227317
rect 587498 227305 587504 227317
rect 630160 227305 630166 227317
rect 587498 227277 630166 227305
rect 587498 227265 587504 227277
rect 630160 227265 630166 227277
rect 630218 227265 630224 227317
rect 588592 227231 588598 227243
rect 390890 227203 395198 227231
rect 395266 227203 588598 227231
rect 390890 227191 390896 227203
rect 220336 227117 220342 227169
rect 220394 227157 220400 227169
rect 247408 227157 247414 227169
rect 220394 227129 247414 227157
rect 220394 227117 220400 227129
rect 247408 227117 247414 227129
rect 247466 227117 247472 227169
rect 263824 227117 263830 227169
rect 263882 227157 263888 227169
rect 288112 227157 288118 227169
rect 263882 227129 288118 227157
rect 263882 227117 263888 227129
rect 288112 227117 288118 227129
rect 288170 227117 288176 227169
rect 288976 227117 288982 227169
rect 289034 227157 289040 227169
rect 369616 227157 369622 227169
rect 289034 227129 369622 227157
rect 289034 227117 289040 227129
rect 369616 227117 369622 227129
rect 369674 227117 369680 227169
rect 392656 227117 392662 227169
rect 392714 227157 392720 227169
rect 395170 227157 395198 227203
rect 588592 227191 588598 227203
rect 588650 227191 588656 227243
rect 588880 227191 588886 227243
rect 588938 227231 588944 227243
rect 626416 227231 626422 227243
rect 588938 227203 626422 227231
rect 588938 227191 588944 227203
rect 626416 227191 626422 227203
rect 626474 227191 626480 227243
rect 590128 227157 590134 227169
rect 392714 227129 395102 227157
rect 395170 227129 590134 227157
rect 392714 227117 392720 227129
rect 238768 227043 238774 227095
rect 238826 227083 238832 227095
rect 252112 227083 252118 227095
rect 238826 227055 252118 227083
rect 238826 227043 238832 227055
rect 252112 227043 252118 227055
rect 252170 227043 252176 227095
rect 275248 227043 275254 227095
rect 275306 227083 275312 227095
rect 275306 227055 357134 227083
rect 275306 227043 275312 227055
rect 213040 226969 213046 227021
rect 213098 227009 213104 227021
rect 233776 227009 233782 227021
rect 213098 226981 233782 227009
rect 213098 226969 213104 226981
rect 233776 226969 233782 226981
rect 233834 226969 233840 227021
rect 238096 226969 238102 227021
rect 238154 227009 238160 227021
rect 264016 227009 264022 227021
rect 238154 226981 264022 227009
rect 238154 226969 238160 226981
rect 264016 226969 264022 226981
rect 264074 226969 264080 227021
rect 276688 226969 276694 227021
rect 276746 227009 276752 227021
rect 357106 227009 357134 227055
rect 359824 227043 359830 227095
rect 359882 227083 359888 227095
rect 393136 227083 393142 227095
rect 359882 227055 393142 227083
rect 359882 227043 359888 227055
rect 393136 227043 393142 227055
rect 393194 227043 393200 227095
rect 357616 227009 357622 227021
rect 276746 226981 347006 227009
rect 357106 226981 357622 227009
rect 276746 226969 276752 226981
rect 221680 226895 221686 226947
rect 221738 226935 221744 226947
rect 250384 226935 250390 226947
rect 221738 226907 250390 226935
rect 221738 226895 221744 226907
rect 250384 226895 250390 226907
rect 250442 226895 250448 226947
rect 253552 226895 253558 226947
rect 253610 226935 253616 226947
rect 266992 226935 266998 226947
rect 253610 226907 266998 226935
rect 253610 226895 253616 226907
rect 266992 226895 266998 226907
rect 267050 226895 267056 226947
rect 273424 226895 273430 226947
rect 273482 226935 273488 226947
rect 346978 226935 347006 226981
rect 357616 226969 357622 226981
rect 357674 226969 357680 227021
rect 365680 226969 365686 227021
rect 365738 227009 365744 227021
rect 393808 227009 393814 227021
rect 365738 226981 393814 227009
rect 365738 226969 365744 226981
rect 393808 226969 393814 226981
rect 393866 226969 393872 227021
rect 395074 227009 395102 227129
rect 590128 227117 590134 227129
rect 590186 227117 590192 227169
rect 590896 227117 590902 227169
rect 590954 227157 590960 227169
rect 630928 227157 630934 227169
rect 590954 227129 630934 227157
rect 590954 227117 590960 227129
rect 630928 227117 630934 227129
rect 630986 227117 630992 227169
rect 397648 227043 397654 227095
rect 397706 227083 397712 227095
rect 407344 227083 407350 227095
rect 397706 227055 407350 227083
rect 397706 227043 397712 227055
rect 407344 227043 407350 227055
rect 407402 227043 407408 227095
rect 407440 227043 407446 227095
rect 407498 227083 407504 227095
rect 584080 227083 584086 227095
rect 407498 227055 584086 227083
rect 407498 227043 407504 227055
rect 584080 227043 584086 227055
rect 584138 227043 584144 227095
rect 590512 227043 590518 227095
rect 590570 227083 590576 227095
rect 632368 227083 632374 227095
rect 590570 227055 632374 227083
rect 590570 227043 590576 227055
rect 632368 227043 632374 227055
rect 632426 227043 632432 227095
rect 593968 227009 593974 227021
rect 395074 226981 593974 227009
rect 593968 226969 593974 226981
rect 594026 226969 594032 227021
rect 599152 226969 599158 227021
rect 599210 226969 599216 227021
rect 606352 226969 606358 227021
rect 606410 227009 606416 227021
rect 638512 227009 638518 227021
rect 606410 226981 638518 227009
rect 606410 226969 606416 226981
rect 638512 226969 638518 226981
rect 638570 226969 638576 227021
rect 360592 226935 360598 226947
rect 273482 226907 346910 226935
rect 346978 226907 360598 226935
rect 273482 226895 273488 226907
rect 224848 226821 224854 226873
rect 224906 226861 224912 226873
rect 256432 226861 256438 226873
rect 224906 226833 256438 226861
rect 224906 226821 224912 226833
rect 256432 226821 256438 226833
rect 256490 226821 256496 226873
rect 324112 226821 324118 226873
rect 324170 226861 324176 226873
rect 339472 226861 339478 226873
rect 324170 226833 339478 226861
rect 324170 226821 324176 226833
rect 339472 226821 339478 226833
rect 339530 226821 339536 226873
rect 346882 226861 346910 226907
rect 360592 226895 360598 226907
rect 360650 226895 360656 226947
rect 367024 226895 367030 226947
rect 367082 226935 367088 226947
rect 408208 226935 408214 226947
rect 367082 226907 408214 226935
rect 367082 226895 367088 226907
rect 408208 226895 408214 226907
rect 408266 226895 408272 226947
rect 587344 226895 587350 226947
rect 587402 226935 587408 226947
rect 598480 226935 598486 226947
rect 587402 226907 598486 226935
rect 587402 226895 587408 226907
rect 598480 226895 598486 226907
rect 598538 226895 598544 226947
rect 599170 226935 599198 226969
rect 633136 226935 633142 226947
rect 599170 226907 633142 226935
rect 633136 226895 633142 226907
rect 633194 226895 633200 226947
rect 354544 226861 354550 226873
rect 346882 226833 354550 226861
rect 354544 226821 354550 226833
rect 354602 226821 354608 226873
rect 355888 226821 355894 226873
rect 355946 226861 355952 226873
rect 366832 226861 366838 226873
rect 355946 226833 366838 226861
rect 355946 226821 355952 226833
rect 366832 226821 366838 226833
rect 366890 226821 366896 226873
rect 367120 226821 367126 226873
rect 367178 226861 367184 226873
rect 396112 226861 396118 226873
rect 367178 226833 396118 226861
rect 367178 226821 367184 226833
rect 396112 226821 396118 226833
rect 396170 226821 396176 226873
rect 599152 226861 599158 226873
rect 396514 226833 599158 226861
rect 223312 226747 223318 226799
rect 223370 226787 223376 226799
rect 253456 226787 253462 226799
rect 223370 226759 253462 226787
rect 223370 226747 223376 226759
rect 253456 226747 253462 226759
rect 253514 226747 253520 226799
rect 257104 226747 257110 226799
rect 257162 226787 257168 226799
rect 273232 226787 273238 226799
rect 257162 226759 273238 226787
rect 257162 226747 257168 226759
rect 273232 226747 273238 226759
rect 273290 226747 273296 226799
rect 279760 226747 279766 226799
rect 279818 226787 279824 226799
rect 366736 226787 366742 226799
rect 279818 226759 366742 226787
rect 279818 226747 279824 226759
rect 366736 226747 366742 226759
rect 366794 226747 366800 226799
rect 386608 226747 386614 226799
rect 386666 226787 386672 226799
rect 388720 226787 388726 226799
rect 386666 226759 388726 226787
rect 386666 226747 386672 226759
rect 388720 226747 388726 226759
rect 388778 226747 388784 226799
rect 395536 226747 395542 226799
rect 395594 226787 395600 226799
rect 396514 226787 396542 226833
rect 599152 226821 599158 226833
rect 599210 226821 599216 226873
rect 600400 226821 600406 226873
rect 600458 226861 600464 226873
rect 634672 226861 634678 226873
rect 600458 226833 634678 226861
rect 600458 226821 600464 226833
rect 634672 226821 634678 226833
rect 634730 226821 634736 226873
rect 395594 226759 396542 226787
rect 395594 226747 395600 226759
rect 397456 226747 397462 226799
rect 397514 226787 397520 226799
rect 400624 226787 400630 226799
rect 397514 226759 400630 226787
rect 397514 226747 397520 226759
rect 400624 226747 400630 226759
rect 400682 226747 400688 226799
rect 407344 226747 407350 226799
rect 407402 226787 407408 226799
rect 407402 226759 603230 226787
rect 407402 226747 407408 226759
rect 149392 226673 149398 226725
rect 149450 226713 149456 226725
rect 159760 226713 159766 226725
rect 149450 226685 159766 226713
rect 149450 226673 149456 226685
rect 159760 226673 159766 226685
rect 159818 226673 159824 226725
rect 227920 226673 227926 226725
rect 227978 226713 227984 226725
rect 262480 226713 262486 226725
rect 227978 226685 262486 226713
rect 227978 226673 227984 226685
rect 262480 226673 262486 226685
rect 262538 226673 262544 226725
rect 282544 226673 282550 226725
rect 282602 226713 282608 226725
rect 372688 226713 372694 226725
rect 282602 226685 372694 226713
rect 282602 226673 282608 226685
rect 372688 226673 372694 226685
rect 372746 226673 372752 226725
rect 374608 226673 374614 226725
rect 374666 226713 374672 226725
rect 391504 226713 391510 226725
rect 374666 226685 391510 226713
rect 374666 226673 374672 226685
rect 391504 226673 391510 226685
rect 391562 226673 391568 226725
rect 397168 226673 397174 226725
rect 397226 226713 397232 226725
rect 602992 226713 602998 226725
rect 397226 226685 602998 226713
rect 397226 226673 397232 226685
rect 602992 226673 602998 226685
rect 603050 226673 603056 226725
rect 226576 226599 226582 226651
rect 226634 226639 226640 226651
rect 259408 226639 259414 226651
rect 226634 226611 259414 226639
rect 226634 226599 226640 226611
rect 259408 226599 259414 226611
rect 259466 226599 259472 226651
rect 285712 226599 285718 226651
rect 285770 226639 285776 226651
rect 378736 226639 378742 226651
rect 285770 226611 378742 226639
rect 285770 226599 285776 226611
rect 378736 226599 378742 226611
rect 378794 226599 378800 226651
rect 382960 226599 382966 226651
rect 383018 226639 383024 226651
rect 397648 226639 397654 226651
rect 383018 226611 397654 226639
rect 383018 226599 383024 226611
rect 397648 226599 397654 226611
rect 397706 226599 397712 226651
rect 400816 226599 400822 226651
rect 400874 226639 400880 226651
rect 603202 226639 603230 226759
rect 603376 226747 603382 226799
rect 603434 226787 603440 226799
rect 636880 226787 636886 226799
rect 603434 226759 636886 226787
rect 603434 226747 603440 226759
rect 636880 226747 636886 226759
rect 636938 226747 636944 226799
rect 603280 226673 603286 226725
rect 603338 226713 603344 226725
rect 637744 226713 637750 226725
rect 603338 226685 637750 226713
rect 603338 226673 603344 226685
rect 637744 226673 637750 226685
rect 637802 226673 637808 226725
rect 603664 226639 603670 226651
rect 400874 226611 417614 226639
rect 603202 226611 603670 226639
rect 400874 226599 400880 226611
rect 229552 226525 229558 226577
rect 229610 226565 229616 226577
rect 265552 226565 265558 226577
rect 229610 226537 265558 226565
rect 229610 226525 229616 226537
rect 265552 226525 265558 226537
rect 265610 226525 265616 226577
rect 271024 226525 271030 226577
rect 271082 226565 271088 226577
rect 294256 226565 294262 226577
rect 271082 226537 294262 226565
rect 271082 226525 271088 226537
rect 294256 226525 294262 226537
rect 294314 226525 294320 226577
rect 297328 226525 297334 226577
rect 297386 226565 297392 226577
rect 390064 226565 390070 226577
rect 297386 226537 390070 226565
rect 297386 226525 297392 226537
rect 390064 226525 390070 226537
rect 390122 226525 390128 226577
rect 402352 226525 402358 226577
rect 402410 226565 402416 226577
rect 417586 226565 417614 226611
rect 603664 226599 603670 226611
rect 603722 226599 603728 226651
rect 606160 226599 606166 226651
rect 606218 226639 606224 226651
rect 639952 226639 639958 226651
rect 606218 226611 639958 226639
rect 606218 226599 606224 226611
rect 639952 226599 639958 226611
rect 640010 226599 640016 226651
rect 609808 226565 609814 226577
rect 402410 226537 417470 226565
rect 417586 226537 609814 226565
rect 402410 226525 402416 226537
rect 247696 226451 247702 226503
rect 247754 226491 247760 226503
rect 257968 226491 257974 226503
rect 247754 226463 257974 226491
rect 247754 226451 247760 226463
rect 257968 226451 257974 226463
rect 258026 226451 258032 226503
rect 268144 226451 268150 226503
rect 268202 226491 268208 226503
rect 282064 226491 282070 226503
rect 268202 226463 282070 226491
rect 268202 226451 268208 226463
rect 282064 226451 282070 226463
rect 282122 226451 282128 226503
rect 288496 226451 288502 226503
rect 288554 226491 288560 226503
rect 384784 226491 384790 226503
rect 288554 226463 384790 226491
rect 288554 226451 288560 226463
rect 384784 226451 384790 226463
rect 384842 226451 384848 226503
rect 385744 226451 385750 226503
rect 385802 226491 385808 226503
rect 394768 226491 394774 226503
rect 385802 226463 394774 226491
rect 385802 226451 385808 226463
rect 394768 226451 394774 226463
rect 394826 226451 394832 226503
rect 402640 226451 402646 226503
rect 402698 226491 402704 226503
rect 417442 226491 417470 226537
rect 609808 226525 609814 226537
rect 609866 226525 609872 226577
rect 612784 226491 612790 226503
rect 402698 226463 417374 226491
rect 417442 226463 612790 226491
rect 402698 226451 402704 226463
rect 232528 226377 232534 226429
rect 232586 226417 232592 226429
rect 271600 226417 271606 226429
rect 232586 226389 271606 226417
rect 232586 226377 232592 226389
rect 271600 226377 271606 226389
rect 271658 226377 271664 226429
rect 284656 226377 284662 226429
rect 284714 226417 284720 226429
rect 378064 226417 378070 226429
rect 284714 226389 378070 226417
rect 284714 226377 284720 226389
rect 378064 226377 378070 226389
rect 378122 226377 378128 226429
rect 382672 226377 382678 226429
rect 382730 226417 382736 226429
rect 386992 226417 386998 226429
rect 382730 226389 386998 226417
rect 382730 226377 382736 226389
rect 386992 226377 386998 226389
rect 387050 226377 387056 226429
rect 404944 226377 404950 226429
rect 405002 226417 405008 226429
rect 417346 226417 417374 226463
rect 612784 226451 612790 226463
rect 612842 226451 612848 226503
rect 613552 226417 613558 226429
rect 405002 226389 417278 226417
rect 417346 226389 613558 226417
rect 405002 226377 405008 226389
rect 147184 226303 147190 226355
rect 147242 226343 147248 226355
rect 151216 226343 151222 226355
rect 147242 226315 151222 226343
rect 147242 226303 147248 226315
rect 151216 226303 151222 226315
rect 151274 226303 151280 226355
rect 213808 226303 213814 226355
rect 213866 226343 213872 226355
rect 237520 226343 237526 226355
rect 213866 226315 237526 226343
rect 213866 226303 213872 226315
rect 237520 226303 237526 226315
rect 237578 226303 237584 226355
rect 241744 226303 241750 226355
rect 241802 226343 241808 226355
rect 241802 226315 252062 226343
rect 241802 226303 241808 226315
rect 216400 226229 216406 226281
rect 216458 226269 216464 226281
rect 239824 226269 239830 226281
rect 216458 226241 239830 226269
rect 216458 226229 216464 226241
rect 239824 226229 239830 226241
rect 239882 226229 239888 226281
rect 245008 226229 245014 226281
rect 245066 226269 245072 226281
rect 252034 226269 252062 226315
rect 252112 226303 252118 226355
rect 252170 226343 252176 226355
rect 285136 226343 285142 226355
rect 252170 226315 285142 226343
rect 252170 226303 252176 226315
rect 285136 226303 285142 226315
rect 285194 226303 285200 226355
rect 291568 226303 291574 226355
rect 291626 226343 291632 226355
rect 390832 226343 390838 226355
rect 291626 226315 390838 226343
rect 291626 226303 291632 226315
rect 390832 226303 390838 226315
rect 390890 226303 390896 226355
rect 407728 226303 407734 226355
rect 407786 226343 407792 226355
rect 417250 226343 417278 226389
rect 613552 226377 613558 226389
rect 613610 226377 613616 226429
rect 629200 226377 629206 226429
rect 629258 226417 629264 226429
rect 635440 226417 635446 226429
rect 629258 226389 635446 226417
rect 629258 226377 629264 226389
rect 635440 226377 635446 226389
rect 635498 226377 635504 226429
rect 618064 226343 618070 226355
rect 407786 226315 417182 226343
rect 417250 226315 618070 226343
rect 407786 226303 407792 226315
rect 291184 226269 291190 226281
rect 245066 226241 251966 226269
rect 252034 226241 291190 226269
rect 245066 226229 245072 226241
rect 215632 226155 215638 226207
rect 215690 226195 215696 226207
rect 240592 226195 240598 226207
rect 215690 226167 240598 226195
rect 215690 226155 215696 226167
rect 240592 226155 240598 226167
rect 240650 226155 240656 226207
rect 246544 226155 246550 226207
rect 246602 226195 246608 226207
rect 251938 226195 251966 226241
rect 291184 226229 291190 226241
rect 291242 226229 291248 226281
rect 297616 226229 297622 226281
rect 297674 226269 297680 226281
rect 402832 226269 402838 226281
rect 297674 226241 402838 226269
rect 297674 226229 297680 226241
rect 402832 226229 402838 226241
rect 402890 226229 402896 226281
rect 410416 226229 410422 226281
rect 410474 226269 410480 226281
rect 417154 226269 417182 226315
rect 618064 226303 618070 226315
rect 618122 226303 618128 226355
rect 624112 226269 624118 226281
rect 410474 226241 414014 226269
rect 417154 226241 624118 226269
rect 410474 226229 410480 226241
rect 297232 226195 297238 226207
rect 246602 226167 251870 226195
rect 251938 226167 297238 226195
rect 246602 226155 246608 226167
rect 151120 226081 151126 226133
rect 151178 226121 151184 226133
rect 187120 226121 187126 226133
rect 151178 226093 187126 226121
rect 151178 226081 151184 226093
rect 187120 226081 187126 226093
rect 187178 226081 187184 226133
rect 218320 226081 218326 226133
rect 218378 226121 218384 226133
rect 246640 226121 246646 226133
rect 218378 226093 246646 226121
rect 218378 226081 218384 226093
rect 246640 226081 246646 226093
rect 246698 226081 246704 226133
rect 251842 226121 251870 226167
rect 297232 226155 297238 226167
rect 297290 226155 297296 226207
rect 301264 226155 301270 226207
rect 301322 226195 301328 226207
rect 411280 226195 411286 226207
rect 301322 226167 411286 226195
rect 301322 226155 301328 226167
rect 411280 226155 411286 226167
rect 411338 226155 411344 226207
rect 413986 226195 414014 226241
rect 624112 226229 624118 226241
rect 624170 226229 624176 226281
rect 629392 226195 629398 226207
rect 413986 226167 629398 226195
rect 629392 226155 629398 226167
rect 629450 226155 629456 226207
rect 300208 226121 300214 226133
rect 251842 226093 300214 226121
rect 300208 226081 300214 226093
rect 300266 226081 300272 226133
rect 300688 226081 300694 226133
rect 300746 226121 300752 226133
rect 408976 226121 408982 226133
rect 300746 226093 408982 226121
rect 300746 226081 300752 226093
rect 408976 226081 408982 226093
rect 409034 226081 409040 226133
rect 411664 226081 411670 226133
rect 411722 226121 411728 226133
rect 631696 226121 631702 226133
rect 411722 226093 631702 226121
rect 411722 226081 411728 226093
rect 631696 226081 631702 226093
rect 631754 226081 631760 226133
rect 214576 226007 214582 226059
rect 214634 226047 214640 226059
rect 236848 226047 236854 226059
rect 214634 226019 236854 226047
rect 214634 226007 214640 226019
rect 236848 226007 236854 226019
rect 236906 226007 236912 226059
rect 238960 226007 238966 226059
rect 239018 226047 239024 226059
rect 261040 226047 261046 226059
rect 239018 226019 261046 226047
rect 239018 226007 239024 226019
rect 261040 226007 261046 226019
rect 261098 226007 261104 226059
rect 271792 226007 271798 226059
rect 271850 226047 271856 226059
rect 336400 226047 336406 226059
rect 271850 226019 336406 226047
rect 271850 226007 271856 226019
rect 336400 226007 336406 226019
rect 336458 226007 336464 226059
rect 379984 226007 379990 226059
rect 380042 226047 380048 226059
rect 394576 226047 394582 226059
rect 380042 226019 394582 226047
rect 380042 226007 380048 226019
rect 394576 226007 394582 226019
rect 394634 226007 394640 226059
rect 394672 226007 394678 226059
rect 394730 226047 394736 226059
rect 582640 226047 582646 226059
rect 394730 226019 582646 226047
rect 394730 226007 394736 226019
rect 582640 226007 582646 226019
rect 582698 226007 582704 226059
rect 584560 226007 584566 226059
rect 584618 226047 584624 226059
rect 584618 226019 584990 226047
rect 584618 226007 584624 226019
rect 212368 225933 212374 225985
rect 212426 225973 212432 225985
rect 234544 225973 234550 225985
rect 212426 225945 234550 225973
rect 212426 225933 212432 225945
rect 234544 225933 234550 225945
rect 234602 225933 234608 225985
rect 267760 225933 267766 225985
rect 267818 225973 267824 225985
rect 267818 225945 273182 225973
rect 267818 225933 267824 225945
rect 218800 225859 218806 225911
rect 218858 225899 218864 225911
rect 244336 225899 244342 225911
rect 218858 225871 244342 225899
rect 218858 225859 218864 225871
rect 244336 225859 244342 225871
rect 244394 225859 244400 225911
rect 262000 225859 262006 225911
rect 262058 225899 262064 225911
rect 273040 225899 273046 225911
rect 262058 225871 273046 225899
rect 262058 225859 262064 225871
rect 273040 225859 273046 225871
rect 273098 225859 273104 225911
rect 273154 225899 273182 225945
rect 273232 225933 273238 225985
rect 273290 225973 273296 225985
rect 321328 225973 321334 225985
rect 273290 225945 321334 225973
rect 273290 225933 273296 225945
rect 321328 225933 321334 225945
rect 321386 225933 321392 225985
rect 374320 225933 374326 225985
rect 374378 225973 374384 225985
rect 387760 225973 387766 225985
rect 374378 225945 387766 225973
rect 374378 225933 374384 225945
rect 387760 225933 387766 225945
rect 387818 225933 387824 225985
rect 388144 225933 388150 225985
rect 388202 225973 388208 225985
rect 584848 225973 584854 225985
rect 388202 225945 584854 225973
rect 388202 225933 388208 225945
rect 584848 225933 584854 225945
rect 584906 225933 584912 225985
rect 584962 225973 584990 226019
rect 587056 226007 587062 226059
rect 587114 226047 587120 226059
rect 595408 226047 595414 226059
rect 587114 226019 595414 226047
rect 587114 226007 587120 226019
rect 595408 226007 595414 226019
rect 595466 226007 595472 226059
rect 628624 226047 628630 226059
rect 599026 226019 628630 226047
rect 599026 225973 599054 226019
rect 628624 226007 628630 226019
rect 628682 226007 628688 226059
rect 584962 225945 599054 225973
rect 603472 225933 603478 225985
rect 603530 225973 603536 225985
rect 636208 225973 636214 225985
rect 603530 225945 636214 225973
rect 603530 225933 603536 225945
rect 636208 225933 636214 225945
rect 636266 225933 636272 225985
rect 327376 225899 327382 225911
rect 273154 225871 327382 225899
rect 327376 225859 327382 225871
rect 327434 225859 327440 225911
rect 331408 225859 331414 225911
rect 331466 225899 331472 225911
rect 345520 225899 345526 225911
rect 331466 225871 345526 225899
rect 331466 225859 331472 225871
rect 345520 225859 345526 225871
rect 345578 225859 345584 225911
rect 382672 225899 382678 225911
rect 368626 225871 382678 225899
rect 269008 225785 269014 225837
rect 269066 225825 269072 225837
rect 330448 225825 330454 225837
rect 269066 225797 330454 225825
rect 269066 225785 269072 225797
rect 330448 225785 330454 225797
rect 330506 225785 330512 225837
rect 345712 225785 345718 225837
rect 345770 225825 345776 225837
rect 368626 225825 368654 225871
rect 382672 225859 382678 225871
rect 382730 225859 382736 225911
rect 382864 225859 382870 225911
rect 382922 225899 382928 225911
rect 386416 225899 386422 225911
rect 382922 225871 386422 225899
rect 382922 225859 382928 225871
rect 386416 225859 386422 225871
rect 386474 225859 386480 225911
rect 387376 225859 387382 225911
rect 387434 225899 387440 225911
rect 394672 225899 394678 225911
rect 387434 225871 394678 225899
rect 387434 225859 387440 225871
rect 394672 225859 394678 225871
rect 394730 225859 394736 225911
rect 394768 225859 394774 225911
rect 394826 225899 394832 225911
rect 579568 225899 579574 225911
rect 394826 225871 579574 225899
rect 394826 225859 394832 225871
rect 579568 225859 579574 225871
rect 579626 225859 579632 225911
rect 345770 225797 368654 225825
rect 345770 225785 345776 225797
rect 374416 225785 374422 225837
rect 374474 225825 374480 225837
rect 385552 225825 385558 225837
rect 374474 225797 385558 225825
rect 374474 225785 374480 225797
rect 385552 225785 385558 225797
rect 385610 225785 385616 225837
rect 388816 225785 388822 225837
rect 388874 225825 388880 225837
rect 581104 225825 581110 225837
rect 388874 225797 581110 225825
rect 388874 225785 388880 225797
rect 581104 225785 581110 225797
rect 581162 225785 581168 225837
rect 588400 225785 588406 225837
rect 588458 225825 588464 225837
rect 602224 225825 602230 225837
rect 588458 225797 602230 225825
rect 588458 225785 588464 225797
rect 602224 225785 602230 225797
rect 602282 225785 602288 225837
rect 231088 225711 231094 225763
rect 231146 225751 231152 225763
rect 268528 225751 268534 225763
rect 231146 225723 268534 225751
rect 231146 225711 231152 225723
rect 268528 225711 268534 225723
rect 268586 225711 268592 225763
rect 279184 225711 279190 225763
rect 279242 225751 279248 225763
rect 324400 225751 324406 225763
rect 279242 225723 324406 225751
rect 279242 225711 279248 225723
rect 324400 225711 324406 225723
rect 324458 225711 324464 225763
rect 338896 225711 338902 225763
rect 338954 225751 338960 225763
rect 396880 225751 396886 225763
rect 338954 225723 396886 225751
rect 338954 225711 338960 225723
rect 396880 225711 396886 225723
rect 396938 225711 396944 225763
rect 408880 225711 408886 225763
rect 408938 225751 408944 225763
rect 610480 225751 610486 225763
rect 408938 225723 610486 225751
rect 408938 225711 408944 225723
rect 610480 225711 610486 225723
rect 610538 225711 610544 225763
rect 265072 225637 265078 225689
rect 265130 225677 265136 225689
rect 279088 225677 279094 225689
rect 265130 225649 279094 225677
rect 265130 225637 265136 225649
rect 279088 225637 279094 225649
rect 279146 225637 279152 225689
rect 279280 225637 279286 225689
rect 279338 225677 279344 225689
rect 318352 225677 318358 225689
rect 279338 225649 318358 225677
rect 279338 225637 279344 225649
rect 318352 225637 318358 225649
rect 318410 225637 318416 225689
rect 321712 225637 321718 225689
rect 321770 225677 321776 225689
rect 451216 225677 451222 225689
rect 321770 225649 451222 225677
rect 321770 225637 321776 225649
rect 451216 225637 451222 225649
rect 451274 225637 451280 225689
rect 587248 225637 587254 225689
rect 587306 225677 587312 225689
rect 592336 225677 592342 225689
rect 587306 225649 592342 225677
rect 587306 225637 587312 225649
rect 592336 225637 592342 225649
rect 592394 225637 592400 225689
rect 241840 225563 241846 225615
rect 241898 225603 241904 225615
rect 248848 225603 248854 225615
rect 241898 225575 248854 225603
rect 241898 225563 241904 225575
rect 248848 225563 248854 225575
rect 248906 225563 248912 225615
rect 309328 225603 309334 225615
rect 276610 225575 309334 225603
rect 42160 225415 42166 225467
rect 42218 225455 42224 225467
rect 48016 225455 48022 225467
rect 42218 225427 48022 225455
rect 42218 225415 42224 225427
rect 48016 225415 48022 225427
rect 48074 225415 48080 225467
rect 259024 225415 259030 225467
rect 259082 225455 259088 225467
rect 269968 225455 269974 225467
rect 259082 225427 269974 225455
rect 259082 225415 259088 225427
rect 269968 225415 269974 225427
rect 270026 225415 270032 225467
rect 273616 225415 273622 225467
rect 273674 225455 273680 225467
rect 276610 225455 276638 225575
rect 309328 225563 309334 225575
rect 309386 225563 309392 225615
rect 315760 225563 315766 225615
rect 315818 225603 315824 225615
rect 439120 225603 439126 225615
rect 315818 225575 439126 225603
rect 315818 225563 315824 225575
rect 439120 225563 439126 225575
rect 439178 225563 439184 225615
rect 309904 225489 309910 225541
rect 309962 225529 309968 225541
rect 427024 225529 427030 225541
rect 309962 225501 427030 225529
rect 309962 225489 309968 225501
rect 427024 225489 427030 225501
rect 427082 225489 427088 225541
rect 273674 225427 276638 225455
rect 273674 225415 273680 225427
rect 306640 225415 306646 225467
rect 306698 225455 306704 225467
rect 420976 225455 420982 225467
rect 306698 225427 420982 225455
rect 306698 225415 306704 225427
rect 420976 225415 420982 225427
rect 421034 225415 421040 225467
rect 264688 225341 264694 225393
rect 264746 225381 264752 225393
rect 276112 225381 276118 225393
rect 264746 225353 276118 225381
rect 264746 225341 264752 225353
rect 276112 225341 276118 225353
rect 276170 225341 276176 225393
rect 276208 225341 276214 225393
rect 276266 225381 276272 225393
rect 303184 225381 303190 225393
rect 276266 225353 303190 225381
rect 276266 225341 276272 225353
rect 303184 225341 303190 225353
rect 303242 225341 303248 225393
rect 303856 225341 303862 225393
rect 303914 225381 303920 225393
rect 415024 225381 415030 225393
rect 303914 225353 415030 225381
rect 303914 225341 303920 225353
rect 415024 225341 415030 225353
rect 415082 225341 415088 225393
rect 302224 225267 302230 225319
rect 302282 225307 302288 225319
rect 411952 225307 411958 225319
rect 302282 225279 411958 225307
rect 302282 225267 302288 225279
rect 411952 225267 411958 225279
rect 412010 225267 412016 225319
rect 282352 225193 282358 225245
rect 282410 225233 282416 225245
rect 342544 225233 342550 225245
rect 282410 225205 342550 225233
rect 282410 225193 282416 225205
rect 342544 225193 342550 225205
rect 342602 225193 342608 225245
rect 351376 225193 351382 225245
rect 351434 225233 351440 225245
rect 418000 225233 418006 225245
rect 351434 225205 418006 225233
rect 351434 225193 351440 225205
rect 418000 225193 418006 225205
rect 418058 225193 418064 225245
rect 243952 225119 243958 225171
rect 244010 225159 244016 225171
rect 251920 225159 251926 225171
rect 244010 225131 251926 225159
rect 244010 225119 244016 225131
rect 251920 225119 251926 225131
rect 251978 225119 251984 225171
rect 305008 225119 305014 225171
rect 305066 225159 305072 225171
rect 333520 225159 333526 225171
rect 305066 225131 333526 225159
rect 305066 225119 305072 225131
rect 333520 225119 333526 225131
rect 333578 225119 333584 225171
rect 339088 225119 339094 225171
rect 339146 225159 339152 225171
rect 399952 225159 399958 225171
rect 339146 225131 399958 225159
rect 339146 225119 339152 225131
rect 399952 225119 399958 225131
rect 400010 225119 400016 225171
rect 606736 225159 606742 225171
rect 417586 225131 606742 225159
rect 252688 225045 252694 225097
rect 252746 225085 252752 225097
rect 312304 225085 312310 225097
rect 252746 225057 312310 225085
rect 252746 225045 252752 225057
rect 312304 225045 312310 225057
rect 312362 225045 312368 225097
rect 348688 225045 348694 225097
rect 348746 225085 348752 225097
rect 399088 225085 399094 225097
rect 348746 225057 399094 225085
rect 348746 225045 348752 225057
rect 399088 225045 399094 225057
rect 399146 225045 399152 225097
rect 399376 225045 399382 225097
rect 399434 225085 399440 225097
rect 417586 225085 417614 225131
rect 606736 225119 606742 225131
rect 606794 225119 606800 225171
rect 399434 225057 417614 225085
rect 399434 225045 399440 225057
rect 368848 224971 368854 225023
rect 368906 225011 368912 225023
rect 376432 225011 376438 225023
rect 368906 224983 376438 225011
rect 368906 224971 368912 224983
rect 376432 224971 376438 224983
rect 376490 224971 376496 225023
rect 378640 224971 378646 225023
rect 378698 225011 378704 225023
rect 405136 225011 405142 225023
rect 378698 224983 405142 225011
rect 378698 224971 378704 224983
rect 405136 224971 405142 224983
rect 405194 224971 405200 225023
rect 362800 224897 362806 224949
rect 362858 224937 362864 224949
rect 402160 224937 402166 224949
rect 362858 224909 402166 224937
rect 362858 224897 362864 224909
rect 402160 224897 402166 224909
rect 402218 224897 402224 224949
rect 149392 224823 149398 224875
rect 149450 224863 149456 224875
rect 162736 224863 162742 224875
rect 149450 224835 162742 224863
rect 149450 224823 149456 224835
rect 162736 224823 162742 224835
rect 162794 224823 162800 224875
rect 277936 224823 277942 224875
rect 277994 224863 278000 224875
rect 363664 224863 363670 224875
rect 277994 224835 363670 224863
rect 277994 224823 278000 224835
rect 363664 224823 363670 224835
rect 363722 224823 363728 224875
rect 371536 224823 371542 224875
rect 371594 224863 371600 224875
rect 379504 224863 379510 224875
rect 371594 224835 379510 224863
rect 371594 224823 371600 224835
rect 379504 224823 379510 224835
rect 379562 224823 379568 224875
rect 380080 224823 380086 224875
rect 380138 224863 380144 224875
rect 388624 224863 388630 224875
rect 380138 224835 388630 224863
rect 380138 224823 380144 224835
rect 388624 224823 388630 224835
rect 388682 224823 388688 224875
rect 407440 224863 407446 224875
rect 388786 224835 407446 224863
rect 334096 224749 334102 224801
rect 334154 224789 334160 224801
rect 374320 224789 374326 224801
rect 334154 224761 374326 224789
rect 334154 224749 334160 224761
rect 374320 224749 374326 224761
rect 374378 224749 374384 224801
rect 374512 224749 374518 224801
rect 374570 224789 374576 224801
rect 382576 224789 382582 224801
rect 374570 224761 382582 224789
rect 374570 224749 374576 224761
rect 382576 224749 382582 224761
rect 382634 224749 382640 224801
rect 385840 224749 385846 224801
rect 385898 224789 385904 224801
rect 388786 224789 388814 224835
rect 407440 224823 407446 224835
rect 407498 224823 407504 224875
rect 385898 224761 388814 224789
rect 385898 224749 385904 224761
rect 392272 224749 392278 224801
rect 392330 224789 392336 224801
rect 593104 224789 593110 224801
rect 392330 224761 593110 224789
rect 392330 224749 392336 224761
rect 593104 224749 593110 224761
rect 593162 224749 593168 224801
rect 362416 224675 362422 224727
rect 362474 224715 362480 224727
rect 378640 224715 378646 224727
rect 362474 224687 378646 224715
rect 362474 224675 362480 224687
rect 378640 224675 378646 224687
rect 378698 224675 378704 224727
rect 382768 224675 382774 224727
rect 382826 224715 382832 224727
rect 386320 224715 386326 224727
rect 382826 224687 386326 224715
rect 382826 224675 382832 224687
rect 386320 224675 386326 224687
rect 386378 224675 386384 224727
rect 386416 224675 386422 224727
rect 386474 224715 386480 224727
rect 389296 224715 389302 224727
rect 386474 224687 389302 224715
rect 386474 224675 386480 224687
rect 389296 224675 389302 224687
rect 389354 224675 389360 224727
rect 389488 224675 389494 224727
rect 389546 224715 389552 224727
rect 587152 224715 587158 224727
rect 389546 224687 587158 224715
rect 389546 224675 389552 224687
rect 587152 224675 587158 224687
rect 587210 224675 587216 224727
rect 596080 224675 596086 224727
rect 596138 224715 596144 224727
rect 597712 224715 597718 224727
rect 596138 224687 597718 224715
rect 596138 224675 596144 224687
rect 597712 224675 597718 224687
rect 597770 224675 597776 224727
rect 316336 224601 316342 224653
rect 316394 224641 316400 224653
rect 441424 224641 441430 224653
rect 316394 224613 441430 224641
rect 316394 224601 316400 224613
rect 441424 224601 441430 224613
rect 441482 224601 441488 224653
rect 319408 224527 319414 224579
rect 319466 224567 319472 224579
rect 447472 224567 447478 224579
rect 319466 224539 447478 224567
rect 319466 224527 319472 224539
rect 447472 224527 447478 224539
rect 447530 224527 447536 224579
rect 323248 224453 323254 224505
rect 323306 224493 323312 224505
rect 452752 224493 452758 224505
rect 323306 224465 452758 224493
rect 323306 224453 323312 224465
rect 452752 224453 452758 224465
rect 452810 224453 452816 224505
rect 322288 224379 322294 224431
rect 322346 224419 322352 224431
rect 453424 224419 453430 224431
rect 322346 224391 453430 224419
rect 322346 224379 322352 224391
rect 453424 224379 453430 224391
rect 453482 224379 453488 224431
rect 325264 224305 325270 224357
rect 325322 224345 325328 224357
rect 459568 224345 459574 224357
rect 325322 224317 459574 224345
rect 325322 224305 325328 224317
rect 459568 224305 459574 224317
rect 459626 224305 459632 224357
rect 331504 224231 331510 224283
rect 331562 224271 331568 224283
rect 471568 224271 471574 224283
rect 331562 224243 471574 224271
rect 331562 224231 331568 224243
rect 471568 224231 471574 224243
rect 471626 224231 471632 224283
rect 330736 224157 330742 224209
rect 330794 224197 330800 224209
rect 467824 224197 467830 224209
rect 330794 224169 467830 224197
rect 330794 224157 330800 224169
rect 467824 224157 467830 224169
rect 467882 224157 467888 224209
rect 553264 224157 553270 224209
rect 553322 224197 553328 224209
rect 555376 224197 555382 224209
rect 553322 224169 555382 224197
rect 553322 224157 553328 224169
rect 555376 224157 555382 224169
rect 555434 224157 555440 224209
rect 328240 224083 328246 224135
rect 328298 224123 328304 224135
rect 465616 224123 465622 224135
rect 328298 224095 465622 224123
rect 328298 224083 328304 224095
rect 465616 224083 465622 224095
rect 465674 224083 465680 224135
rect 334480 224009 334486 224061
rect 334538 224049 334544 224061
rect 477616 224049 477622 224061
rect 334538 224021 477622 224049
rect 334538 224009 334544 224021
rect 477616 224009 477622 224021
rect 477674 224009 477680 224061
rect 337168 223935 337174 223987
rect 337226 223975 337232 223987
rect 483760 223975 483766 223987
rect 337226 223947 483766 223975
rect 337226 223935 337232 223947
rect 483760 223935 483766 223947
rect 483818 223935 483824 223987
rect 340432 223861 340438 223913
rect 340490 223901 340496 223913
rect 489712 223901 489718 223913
rect 340490 223873 489718 223901
rect 340490 223861 340496 223873
rect 489712 223861 489718 223873
rect 489770 223861 489776 223913
rect 343600 223787 343606 223839
rect 343658 223827 343664 223839
rect 497296 223827 497302 223839
rect 343658 223799 497302 223827
rect 343658 223787 343664 223799
rect 497296 223787 497302 223799
rect 497354 223787 497360 223839
rect 263536 223713 263542 223765
rect 263594 223753 263600 223765
rect 335728 223753 335734 223765
rect 263594 223725 335734 223753
rect 263594 223713 263600 223725
rect 335728 223713 335734 223725
rect 335786 223713 335792 223765
rect 346576 223713 346582 223765
rect 346634 223753 346640 223765
rect 501808 223753 501814 223765
rect 346634 223725 501814 223753
rect 346634 223713 346640 223725
rect 501808 223713 501814 223725
rect 501866 223713 501872 223765
rect 261904 223639 261910 223691
rect 261962 223679 261968 223691
rect 332656 223679 332662 223691
rect 261962 223651 332662 223679
rect 261962 223639 261968 223651
rect 332656 223639 332662 223651
rect 332714 223639 332720 223691
rect 349552 223639 349558 223691
rect 349610 223679 349616 223691
rect 507856 223679 507862 223691
rect 349610 223651 507862 223679
rect 349610 223639 349616 223651
rect 507856 223639 507862 223651
rect 507914 223639 507920 223691
rect 266416 223565 266422 223617
rect 266474 223605 266480 223617
rect 341776 223605 341782 223617
rect 266474 223577 341782 223605
rect 266474 223565 266480 223577
rect 341776 223565 341782 223577
rect 341834 223565 341840 223617
rect 348112 223565 348118 223617
rect 348170 223605 348176 223617
rect 506320 223605 506326 223617
rect 348170 223577 506326 223605
rect 348170 223565 348176 223577
rect 506320 223565 506326 223577
rect 506378 223565 506384 223617
rect 268048 223491 268054 223543
rect 268106 223531 268112 223543
rect 344848 223531 344854 223543
rect 268106 223503 344854 223531
rect 268106 223491 268112 223503
rect 344848 223491 344854 223503
rect 344906 223491 344912 223543
rect 348016 223491 348022 223543
rect 348074 223531 348080 223543
rect 504784 223531 504790 223543
rect 348074 223503 504790 223531
rect 348074 223491 348080 223503
rect 504784 223491 504790 223503
rect 504842 223491 504848 223543
rect 264592 223417 264598 223469
rect 264650 223457 264656 223469
rect 338704 223457 338710 223469
rect 264650 223429 338710 223457
rect 264650 223417 264656 223429
rect 338704 223417 338710 223429
rect 338762 223417 338768 223469
rect 352528 223417 352534 223469
rect 352586 223457 352592 223469
rect 513904 223457 513910 223469
rect 352586 223429 513910 223457
rect 352586 223417 352592 223429
rect 513904 223417 513910 223429
rect 513962 223417 513968 223469
rect 270928 223343 270934 223395
rect 270986 223383 270992 223395
rect 350800 223383 350806 223395
rect 270986 223355 350806 223383
rect 270986 223343 270992 223355
rect 350800 223343 350806 223355
rect 350858 223343 350864 223395
rect 351088 223343 351094 223395
rect 351146 223383 351152 223395
rect 510832 223383 510838 223395
rect 351146 223355 510838 223383
rect 351146 223343 351152 223355
rect 510832 223343 510838 223355
rect 510890 223343 510896 223395
rect 269392 223269 269398 223321
rect 269450 223309 269456 223321
rect 347728 223309 347734 223321
rect 269450 223281 347734 223309
rect 269450 223269 269456 223281
rect 347728 223269 347734 223281
rect 347786 223269 347792 223321
rect 351184 223269 351190 223321
rect 351242 223309 351248 223321
rect 512368 223309 512374 223321
rect 351242 223281 512374 223309
rect 351242 223269 351248 223281
rect 512368 223269 512374 223281
rect 512426 223269 512432 223321
rect 272560 223195 272566 223247
rect 272618 223235 272624 223247
rect 353872 223235 353878 223247
rect 272618 223207 353878 223235
rect 272618 223195 272624 223207
rect 353872 223195 353878 223207
rect 353930 223195 353936 223247
rect 353968 223195 353974 223247
rect 354026 223235 354032 223247
rect 516976 223235 516982 223247
rect 354026 223207 516982 223235
rect 354026 223195 354032 223207
rect 516976 223195 516982 223207
rect 517034 223195 517040 223247
rect 313360 223121 313366 223173
rect 313418 223161 313424 223173
rect 435376 223161 435382 223173
rect 313418 223133 435382 223161
rect 313418 223121 313424 223133
rect 435376 223121 435382 223133
rect 435434 223121 435440 223173
rect 310288 223047 310294 223099
rect 310346 223087 310352 223099
rect 429328 223087 429334 223099
rect 310346 223059 429334 223087
rect 310346 223047 310352 223059
rect 429328 223047 429334 223059
rect 429386 223047 429392 223099
rect 312592 222973 312598 223025
rect 312650 223013 312656 223025
rect 431536 223013 431542 223025
rect 312650 222985 431542 223013
rect 312650 222973 312656 222985
rect 431536 222973 431542 222985
rect 431594 222973 431600 223025
rect 307216 222899 307222 222951
rect 307274 222939 307280 222951
rect 423280 222939 423286 222951
rect 307274 222911 423286 222939
rect 307274 222899 307280 222911
rect 423280 222899 423286 222911
rect 423338 222899 423344 222951
rect 304240 222825 304246 222877
rect 304298 222865 304304 222877
rect 417232 222865 417238 222877
rect 304298 222837 417238 222865
rect 304298 222825 304304 222837
rect 417232 222825 417238 222837
rect 417290 222825 417296 222877
rect 307984 222751 307990 222803
rect 308042 222791 308048 222803
rect 422512 222791 422518 222803
rect 308042 222763 422518 222791
rect 308042 222751 308048 222763
rect 422512 222751 422518 222763
rect 422570 222751 422576 222803
rect 286192 222677 286198 222729
rect 286250 222717 286256 222729
rect 381040 222717 381046 222729
rect 286250 222689 381046 222717
rect 286250 222677 286256 222689
rect 381040 222677 381046 222689
rect 381098 222677 381104 222729
rect 403024 222677 403030 222729
rect 403082 222717 403088 222729
rect 511600 222717 511606 222729
rect 403082 222689 511606 222717
rect 403082 222677 403088 222689
rect 511600 222677 511606 222689
rect 511658 222677 511664 222729
rect 302800 222603 302806 222655
rect 302858 222643 302864 222655
rect 414256 222643 414262 222655
rect 302858 222615 414262 222643
rect 302858 222603 302864 222615
rect 414256 222603 414262 222615
rect 414314 222603 414320 222655
rect 302032 222529 302038 222581
rect 302090 222569 302096 222581
rect 410512 222569 410518 222581
rect 302090 222541 410518 222569
rect 302090 222529 302096 222541
rect 410512 222529 410518 222541
rect 410570 222529 410576 222581
rect 410608 222529 410614 222581
rect 410666 222569 410672 222581
rect 430096 222569 430102 222581
rect 410666 222541 430102 222569
rect 410666 222529 410672 222541
rect 430096 222529 430102 222541
rect 430154 222529 430160 222581
rect 283024 222455 283030 222507
rect 283082 222495 283088 222507
rect 374992 222495 374998 222507
rect 283082 222467 374998 222495
rect 283082 222455 283088 222467
rect 374992 222455 374998 222467
rect 375050 222455 375056 222507
rect 394864 222455 394870 222507
rect 394922 222495 394928 222507
rect 496528 222495 496534 222507
rect 394922 222467 496534 222495
rect 394922 222455 394928 222467
rect 496528 222455 496534 222467
rect 496586 222455 496592 222507
rect 281584 222381 281590 222433
rect 281642 222421 281648 222433
rect 371920 222421 371926 222433
rect 281642 222393 371926 222421
rect 281642 222381 281648 222393
rect 371920 222381 371926 222393
rect 371978 222381 371984 222433
rect 386128 222381 386134 222433
rect 386186 222421 386192 222433
rect 482896 222421 482902 222433
rect 386186 222393 482902 222421
rect 386186 222381 386192 222393
rect 482896 222381 482902 222393
rect 482954 222381 482960 222433
rect 274096 222307 274102 222359
rect 274154 222347 274160 222359
rect 356848 222347 356854 222359
rect 274154 222319 356854 222347
rect 274154 222307 274160 222319
rect 356848 222307 356854 222319
rect 356906 222307 356912 222359
rect 371632 222307 371638 222359
rect 371690 222347 371696 222359
rect 443728 222347 443734 222359
rect 371690 222319 443734 222347
rect 371690 222307 371696 222319
rect 443728 222307 443734 222319
rect 443786 222307 443792 222359
rect 149392 221863 149398 221915
rect 149450 221903 149456 221915
rect 168400 221903 168406 221915
rect 149450 221875 168406 221903
rect 149450 221863 149456 221875
rect 168400 221863 168406 221875
rect 168458 221863 168464 221915
rect 149488 221789 149494 221841
rect 149546 221829 149552 221841
rect 171376 221829 171382 221841
rect 149546 221801 171382 221829
rect 149546 221789 149552 221801
rect 171376 221789 171382 221801
rect 171434 221789 171440 221841
rect 656176 221789 656182 221841
rect 656234 221829 656240 221841
rect 676240 221829 676246 221841
rect 656234 221801 676246 221829
rect 656234 221789 656240 221801
rect 676240 221789 676246 221801
rect 676298 221789 676304 221841
rect 145744 221715 145750 221767
rect 145802 221755 145808 221767
rect 184336 221755 184342 221767
rect 145802 221727 184342 221755
rect 145802 221715 145808 221727
rect 184336 221715 184342 221727
rect 184394 221715 184400 221767
rect 478096 221715 478102 221767
rect 478154 221755 478160 221767
rect 479968 221755 479974 221767
rect 478154 221727 479974 221755
rect 478154 221715 478160 221727
rect 479968 221715 479974 221727
rect 480026 221715 480032 221767
rect 512752 221715 512758 221767
rect 512810 221755 512816 221767
rect 515392 221755 515398 221767
rect 512810 221727 515398 221755
rect 512810 221715 512816 221727
rect 515392 221715 515398 221727
rect 515450 221715 515456 221767
rect 146896 221419 146902 221471
rect 146954 221459 146960 221471
rect 151408 221459 151414 221471
rect 146954 221431 151414 221459
rect 146954 221419 146960 221431
rect 151408 221419 151414 221431
rect 151466 221419 151472 221471
rect 673840 219495 673846 219547
rect 673898 219535 673904 219547
rect 676048 219535 676054 219547
rect 673898 219507 676054 219535
rect 673898 219495 673904 219507
rect 676048 219495 676054 219507
rect 676106 219495 676112 219547
rect 655984 219199 655990 219251
rect 656042 219239 656048 219251
rect 676240 219239 676246 219251
rect 656042 219211 676246 219239
rect 656042 219199 656048 219211
rect 676240 219199 676246 219211
rect 676298 219199 676304 219251
rect 147664 219051 147670 219103
rect 147722 219091 147728 219103
rect 179920 219091 179926 219103
rect 147722 219063 179926 219091
rect 147722 219051 147728 219063
rect 179920 219051 179926 219063
rect 179978 219051 179984 219103
rect 655792 219051 655798 219103
rect 655850 219091 655856 219103
rect 676144 219091 676150 219103
rect 655850 219063 676150 219091
rect 655850 219051 655856 219063
rect 676144 219051 676150 219063
rect 676202 219051 676208 219103
rect 149392 218977 149398 219029
rect 149450 219017 149456 219029
rect 165616 219017 165622 219029
rect 149450 218989 165622 219017
rect 149450 218977 149456 218989
rect 165616 218977 165622 218989
rect 165674 218977 165680 219029
rect 143056 218829 143062 218881
rect 143114 218869 143120 218881
rect 184336 218869 184342 218881
rect 143114 218841 184342 218869
rect 143114 218829 143120 218841
rect 184336 218829 184342 218841
rect 184394 218829 184400 218881
rect 149488 216091 149494 216143
rect 149546 216131 149552 216143
rect 174352 216131 174358 216143
rect 149546 216103 174358 216131
rect 149546 216091 149552 216103
rect 174352 216091 174358 216103
rect 174410 216091 174416 216143
rect 149392 216017 149398 216069
rect 149450 216057 149456 216069
rect 177136 216057 177142 216069
rect 149450 216029 177142 216057
rect 149450 216017 149456 216029
rect 177136 216017 177142 216029
rect 177194 216017 177200 216069
rect 675088 216017 675094 216069
rect 675146 216057 675152 216069
rect 676048 216057 676054 216069
rect 675146 216029 676054 216057
rect 675146 216017 675152 216029
rect 676048 216017 676054 216029
rect 676106 216017 676112 216069
rect 149392 214389 149398 214441
rect 149450 214429 149456 214441
rect 159952 214429 159958 214441
rect 149450 214401 159958 214429
rect 149450 214389 149456 214401
rect 159952 214389 159958 214401
rect 160010 214389 160016 214441
rect 147088 214019 147094 214071
rect 147146 214059 147152 214071
rect 151696 214059 151702 214071
rect 147146 214031 151702 214059
rect 147146 214019 147152 214031
rect 151696 214019 151702 214031
rect 151754 214019 151760 214071
rect 41776 213279 41782 213331
rect 41834 213319 41840 213331
rect 45424 213319 45430 213331
rect 41834 213291 45430 213319
rect 41834 213279 41840 213291
rect 45424 213279 45430 213291
rect 45482 213279 45488 213331
rect 674704 213279 674710 213331
rect 674762 213319 674768 213331
rect 676240 213319 676246 213331
rect 674762 213291 676246 213319
rect 674762 213279 674768 213291
rect 676240 213279 676246 213291
rect 676298 213279 676304 213331
rect 674800 213205 674806 213257
rect 674858 213245 674864 213257
rect 675952 213245 675958 213257
rect 674858 213217 675958 213245
rect 674858 213205 674864 213217
rect 675952 213205 675958 213217
rect 676010 213205 676016 213257
rect 675280 213131 675286 213183
rect 675338 213171 675344 213183
rect 676048 213171 676054 213183
rect 675338 213143 676054 213171
rect 675338 213131 675344 213143
rect 676048 213131 676054 213143
rect 676106 213131 676112 213183
rect 41584 212909 41590 212961
rect 41642 212949 41648 212961
rect 45328 212949 45334 212961
rect 41642 212921 45334 212949
rect 41642 212909 41648 212921
rect 45328 212909 45334 212921
rect 45386 212909 45392 212961
rect 146896 212835 146902 212887
rect 146954 212875 146960 212887
rect 152080 212875 152086 212887
rect 146954 212847 152086 212875
rect 146954 212835 146960 212847
rect 152080 212835 152086 212847
rect 152138 212835 152144 212887
rect 41776 212169 41782 212221
rect 41834 212209 41840 212221
rect 44944 212209 44950 212221
rect 41834 212181 44950 212209
rect 41834 212169 41840 212181
rect 44944 212169 44950 212181
rect 45002 212169 45008 212221
rect 674512 212095 674518 212147
rect 674570 212135 674576 212147
rect 676048 212135 676054 212147
rect 674570 212107 676054 212135
rect 674570 212095 674576 212107
rect 676048 212095 676054 212107
rect 676106 212095 676112 212147
rect 41776 211725 41782 211777
rect 41834 211765 41840 211777
rect 43216 211765 43222 211777
rect 41834 211737 43222 211765
rect 41834 211725 41840 211737
rect 43216 211725 43222 211737
rect 43274 211725 43280 211777
rect 41584 211429 41590 211481
rect 41642 211469 41648 211481
rect 44848 211469 44854 211481
rect 41642 211441 44854 211469
rect 41642 211429 41648 211441
rect 44848 211429 44854 211441
rect 44906 211429 44912 211481
rect 41776 210689 41782 210741
rect 41834 210729 41840 210741
rect 50608 210729 50614 210741
rect 41834 210701 50614 210729
rect 41834 210689 41840 210701
rect 50608 210689 50614 210701
rect 50666 210689 50672 210741
rect 674608 210393 674614 210445
rect 674666 210433 674672 210445
rect 675952 210433 675958 210445
rect 674666 210405 675958 210433
rect 674666 210393 674672 210405
rect 675952 210393 675958 210405
rect 676010 210393 676016 210445
rect 147472 210319 147478 210371
rect 147530 210359 147536 210371
rect 151600 210359 151606 210371
rect 147530 210331 151606 210359
rect 147530 210319 147536 210331
rect 151600 210319 151606 210331
rect 151658 210319 151664 210371
rect 674896 210319 674902 210371
rect 674954 210359 674960 210371
rect 676240 210359 676246 210371
rect 674954 210331 676246 210359
rect 674954 210319 674960 210331
rect 676240 210319 676246 210331
rect 676298 210319 676304 210371
rect 147376 210245 147382 210297
rect 147434 210285 147440 210297
rect 151792 210285 151798 210297
rect 147434 210257 151798 210285
rect 147434 210245 147440 210257
rect 151792 210245 151798 210257
rect 151850 210245 151856 210297
rect 674992 210245 674998 210297
rect 675050 210285 675056 210297
rect 676048 210285 676054 210297
rect 675050 210257 676054 210285
rect 675050 210245 675056 210257
rect 676048 210245 676054 210257
rect 676106 210245 676112 210297
rect 41776 210171 41782 210223
rect 41834 210211 41840 210223
rect 43312 210211 43318 210223
rect 41834 210183 43318 210211
rect 41834 210171 41840 210183
rect 43312 210171 43318 210183
rect 43370 210171 43376 210223
rect 41584 209949 41590 210001
rect 41642 209989 41648 210001
rect 50416 209989 50422 210001
rect 41642 209961 50422 209989
rect 41642 209949 41648 209961
rect 50416 209949 50422 209961
rect 50474 209949 50480 210001
rect 41584 209357 41590 209409
rect 41642 209397 41648 209409
rect 43504 209397 43510 209409
rect 41642 209369 43510 209397
rect 41642 209357 41648 209369
rect 43504 209357 43510 209369
rect 43562 209357 43568 209409
rect 147184 207877 147190 207929
rect 147242 207917 147248 207929
rect 151504 207917 151510 207929
rect 147242 207889 151510 207917
rect 147242 207877 147248 207889
rect 151504 207877 151510 207889
rect 151562 207877 151568 207929
rect 41776 207507 41782 207559
rect 41834 207547 41840 207559
rect 42928 207547 42934 207559
rect 41834 207519 42934 207547
rect 41834 207507 41840 207519
rect 42928 207507 42934 207519
rect 42986 207507 42992 207559
rect 146896 207359 146902 207411
rect 146954 207399 146960 207411
rect 151888 207399 151894 207411
rect 146954 207371 151894 207399
rect 146954 207359 146960 207371
rect 151888 207359 151894 207371
rect 151946 207359 151952 207411
rect 646768 207359 646774 207411
rect 646826 207399 646832 207411
rect 679792 207399 679798 207411
rect 646826 207371 679798 207399
rect 646826 207359 646832 207371
rect 679792 207359 679798 207371
rect 679850 207359 679856 207411
rect 147280 206101 147286 206153
rect 147338 206141 147344 206153
rect 151984 206141 151990 206153
rect 147338 206113 151990 206141
rect 147338 206101 147344 206113
rect 151984 206101 151990 206113
rect 152042 206101 152048 206153
rect 675760 206101 675766 206153
rect 675818 206101 675824 206153
rect 675088 205657 675094 205709
rect 675146 205697 675152 205709
rect 675472 205697 675478 205709
rect 675146 205669 675478 205697
rect 675146 205657 675152 205669
rect 675472 205657 675478 205669
rect 675530 205657 675536 205709
rect 675778 205635 675806 206101
rect 675760 205583 675766 205635
rect 675818 205583 675824 205635
rect 149392 204473 149398 204525
rect 149450 204513 149456 204525
rect 182992 204513 182998 204525
rect 149450 204485 182998 204513
rect 149450 204473 149456 204485
rect 182992 204473 182998 204485
rect 183050 204473 183056 204525
rect 674800 202031 674806 202083
rect 674858 202071 674864 202083
rect 675184 202071 675190 202083
rect 674858 202043 675190 202071
rect 674858 202031 674864 202043
rect 675184 202031 675190 202043
rect 675242 202031 675248 202083
rect 41584 201735 41590 201787
rect 41642 201775 41648 201787
rect 42544 201775 42550 201787
rect 41642 201747 42550 201775
rect 41642 201735 41648 201747
rect 42544 201735 42550 201747
rect 42602 201735 42608 201787
rect 149392 201735 149398 201787
rect 149450 201775 149456 201787
rect 174448 201775 174454 201787
rect 149450 201747 174454 201775
rect 149450 201735 149456 201747
rect 174448 201735 174454 201747
rect 174506 201735 174512 201787
rect 41968 201661 41974 201713
rect 42026 201701 42032 201713
rect 44752 201701 44758 201713
rect 42026 201673 44758 201701
rect 42026 201661 42032 201673
rect 44752 201661 44758 201673
rect 44810 201661 44816 201713
rect 149488 201661 149494 201713
rect 149546 201701 149552 201713
rect 177232 201701 177238 201713
rect 149546 201673 177238 201701
rect 149546 201661 149552 201673
rect 177232 201661 177238 201673
rect 177290 201661 177296 201713
rect 41872 201587 41878 201639
rect 41930 201627 41936 201639
rect 42736 201627 42742 201639
rect 41930 201599 42742 201627
rect 41930 201587 41936 201599
rect 42736 201587 42742 201599
rect 42794 201587 42800 201639
rect 149296 201587 149302 201639
rect 149354 201627 149360 201639
rect 180112 201627 180118 201639
rect 149354 201599 180118 201627
rect 149354 201587 149360 201599
rect 180112 201587 180118 201599
rect 180170 201587 180176 201639
rect 41584 201513 41590 201565
rect 41642 201553 41648 201565
rect 44560 201553 44566 201565
rect 41642 201525 44566 201553
rect 41642 201513 41648 201525
rect 44560 201513 44566 201525
rect 44618 201513 44624 201565
rect 143056 201513 143062 201565
rect 143114 201553 143120 201565
rect 185968 201553 185974 201565
rect 143114 201525 185974 201553
rect 143114 201513 143120 201525
rect 185968 201513 185974 201525
rect 186026 201513 186032 201565
rect 655600 201513 655606 201565
rect 655658 201553 655664 201565
rect 675088 201553 675094 201565
rect 655658 201525 675094 201553
rect 655658 201513 655664 201525
rect 675088 201513 675094 201525
rect 675146 201513 675152 201565
rect 674704 201291 674710 201343
rect 674762 201331 674768 201343
rect 675376 201331 675382 201343
rect 674762 201303 675382 201331
rect 674762 201291 674768 201303
rect 675376 201291 675382 201303
rect 675434 201291 675440 201343
rect 41584 200921 41590 200973
rect 41642 200961 41648 200973
rect 44656 200961 44662 200973
rect 41642 200933 44662 200961
rect 41642 200921 41648 200933
rect 44656 200921 44662 200933
rect 44714 200921 44720 200973
rect 34480 200403 34486 200455
rect 34538 200443 34544 200455
rect 42640 200443 42646 200455
rect 34538 200415 42646 200443
rect 34538 200403 34544 200415
rect 42640 200403 42646 200415
rect 42698 200403 42704 200455
rect 34096 200329 34102 200381
rect 34154 200369 34160 200381
rect 42832 200369 42838 200381
rect 34154 200341 42838 200369
rect 34154 200329 34160 200341
rect 42832 200329 42838 200341
rect 42890 200329 42896 200381
rect 34192 200255 34198 200307
rect 34250 200295 34256 200307
rect 43024 200295 43030 200307
rect 34250 200267 43030 200295
rect 34250 200255 34256 200267
rect 43024 200255 43030 200267
rect 43082 200255 43088 200307
rect 34288 200181 34294 200233
rect 34346 200221 34352 200233
rect 42352 200221 42358 200233
rect 34346 200193 42358 200221
rect 34346 200181 34352 200193
rect 42352 200181 42358 200193
rect 42410 200181 42416 200233
rect 34384 200107 34390 200159
rect 34442 200147 34448 200159
rect 43120 200147 43126 200159
rect 34442 200119 43126 200147
rect 34442 200107 34448 200119
rect 43120 200107 43126 200119
rect 43178 200107 43184 200159
rect 147472 198775 147478 198827
rect 147530 198815 147536 198827
rect 154192 198815 154198 198827
rect 147530 198787 154198 198815
rect 147530 198775 147536 198787
rect 154192 198775 154198 198787
rect 154250 198775 154256 198827
rect 149392 198701 149398 198753
rect 149450 198741 149456 198753
rect 162832 198741 162838 198753
rect 149450 198713 162838 198741
rect 149450 198701 149456 198713
rect 162832 198701 162838 198713
rect 162890 198701 162896 198753
rect 181360 198593 181366 198605
rect 181321 198565 181366 198593
rect 181360 198553 181366 198565
rect 181418 198593 181424 198605
rect 185968 198593 185974 198605
rect 181418 198565 185974 198593
rect 181418 198553 181424 198565
rect 185968 198553 185974 198565
rect 186026 198553 186032 198605
rect 178288 198479 178294 198531
rect 178346 198519 178352 198531
rect 186064 198519 186070 198531
rect 178346 198491 186070 198519
rect 178346 198479 178352 198491
rect 186064 198479 186070 198491
rect 186122 198479 186128 198531
rect 674512 197147 674518 197199
rect 674570 197187 674576 197199
rect 675184 197187 675190 197199
rect 674570 197159 675190 197187
rect 674570 197147 674576 197159
rect 675184 197147 675190 197159
rect 675242 197147 675248 197199
rect 149392 195963 149398 196015
rect 149450 196003 149456 196015
rect 168592 196003 168598 196015
rect 149450 195975 168598 196003
rect 149450 195963 149456 195975
rect 168592 195963 168598 195975
rect 168650 195963 168656 196015
rect 149488 195889 149494 195941
rect 149546 195929 149552 195941
rect 171568 195929 171574 195941
rect 149546 195901 171574 195929
rect 149546 195889 149552 195901
rect 171568 195889 171574 195901
rect 171626 195889 171632 195941
rect 149392 195815 149398 195867
rect 149450 195855 149456 195867
rect 183088 195855 183094 195867
rect 149450 195827 183094 195855
rect 149450 195815 149456 195827
rect 183088 195815 183094 195827
rect 183146 195815 183152 195867
rect 166960 195741 166966 195793
rect 167018 195781 167024 195793
rect 184528 195781 184534 195793
rect 167018 195753 184534 195781
rect 167018 195741 167024 195753
rect 184528 195741 184534 195753
rect 184586 195741 184592 195793
rect 169840 195667 169846 195719
rect 169898 195707 169904 195719
rect 184432 195707 184438 195719
rect 169898 195679 184438 195707
rect 169898 195667 169904 195679
rect 184432 195667 184438 195679
rect 184490 195667 184496 195719
rect 172720 195593 172726 195645
rect 172778 195633 172784 195645
rect 184336 195633 184342 195645
rect 172778 195605 184342 195633
rect 172778 195593 172784 195605
rect 184336 195593 184342 195605
rect 184394 195593 184400 195645
rect 42256 194779 42262 194831
rect 42314 194819 42320 194831
rect 42928 194819 42934 194831
rect 42314 194791 42934 194819
rect 42314 194779 42320 194791
rect 42928 194779 42934 194791
rect 42986 194779 42992 194831
rect 149392 193151 149398 193203
rect 149450 193191 149456 193203
rect 160048 193191 160054 193203
rect 149450 193163 160054 193191
rect 149450 193151 149456 193163
rect 160048 193151 160054 193163
rect 160106 193151 160112 193203
rect 149488 193003 149494 193055
rect 149546 193043 149552 193055
rect 165808 193043 165814 193055
rect 149546 193015 165814 193043
rect 149546 193003 149552 193015
rect 165808 193003 165814 193015
rect 165866 193003 165872 193055
rect 152368 192929 152374 192981
rect 152426 192969 152432 192981
rect 184624 192969 184630 192981
rect 152426 192941 184630 192969
rect 152426 192929 152432 192941
rect 184624 192929 184630 192941
rect 184682 192929 184688 192981
rect 42352 192855 42358 192907
rect 42410 192895 42416 192907
rect 43120 192895 43126 192907
rect 42410 192867 43126 192895
rect 42410 192855 42416 192867
rect 43120 192855 43126 192867
rect 43178 192855 43184 192907
rect 155440 192855 155446 192907
rect 155498 192895 155504 192907
rect 184528 192895 184534 192907
rect 155498 192867 184534 192895
rect 155498 192855 155504 192867
rect 184528 192855 184534 192867
rect 184586 192855 184592 192907
rect 158128 192781 158134 192833
rect 158186 192821 158192 192833
rect 184336 192821 184342 192833
rect 158186 192793 184342 192821
rect 158186 192781 158192 192793
rect 184336 192781 184342 192793
rect 184394 192781 184400 192833
rect 163888 192707 163894 192759
rect 163946 192747 163952 192759
rect 184432 192747 184438 192759
rect 163946 192719 184438 192747
rect 163946 192707 163952 192719
rect 184432 192707 184438 192719
rect 184490 192707 184496 192759
rect 42640 191597 42646 191649
rect 42698 191637 42704 191649
rect 42928 191637 42934 191649
rect 42698 191609 42934 191637
rect 42698 191597 42704 191609
rect 42928 191597 42934 191609
rect 42986 191597 42992 191649
rect 147376 190191 147382 190243
rect 147434 190231 147440 190243
rect 154288 190231 154294 190243
rect 147434 190203 154294 190231
rect 147434 190191 147440 190203
rect 154288 190191 154294 190203
rect 154346 190191 154352 190243
rect 149392 190117 149398 190169
rect 149450 190157 149456 190169
rect 157072 190157 157078 190169
rect 149450 190129 157078 190157
rect 149450 190117 149456 190129
rect 157072 190117 157078 190129
rect 157130 190117 157136 190169
rect 143920 190043 143926 190095
rect 143978 190083 143984 190095
rect 184528 190083 184534 190095
rect 143978 190055 184534 190083
rect 143978 190043 143984 190055
rect 184528 190043 184534 190055
rect 184586 190043 184592 190095
rect 149680 189969 149686 190021
rect 149738 190009 149744 190021
rect 184336 190009 184342 190021
rect 149738 189981 184342 190009
rect 149738 189969 149744 189981
rect 184336 189969 184342 189981
rect 184394 189969 184400 190021
rect 171472 189895 171478 189947
rect 171530 189935 171536 189947
rect 184432 189935 184438 189947
rect 171530 189907 184438 189935
rect 171530 189895 171536 189907
rect 184432 189895 184438 189907
rect 184490 189895 184496 189947
rect 180016 189821 180022 189873
rect 180074 189861 180080 189873
rect 184336 189861 184342 189873
rect 180074 189833 184342 189861
rect 180074 189821 180080 189833
rect 184336 189821 184342 189833
rect 184394 189821 184400 189873
rect 159856 187157 159862 187209
rect 159914 187197 159920 187209
rect 184432 187197 184438 187209
rect 159914 187169 184438 187197
rect 159914 187157 159920 187169
rect 184432 187157 184438 187169
rect 184490 187157 184496 187209
rect 165712 187083 165718 187135
rect 165770 187123 165776 187135
rect 184528 187123 184534 187135
rect 165770 187095 184534 187123
rect 165770 187083 165776 187095
rect 184528 187083 184534 187095
rect 184586 187083 184592 187135
rect 168496 187009 168502 187061
rect 168554 187049 168560 187061
rect 184336 187049 184342 187061
rect 168554 187021 184342 187049
rect 168554 187009 168560 187021
rect 184336 187009 184342 187021
rect 184394 187009 184400 187061
rect 177040 186935 177046 186987
rect 177098 186975 177104 186987
rect 184624 186975 184630 186987
rect 177098 186947 184630 186975
rect 177098 186935 177104 186947
rect 184624 186935 184630 186947
rect 184682 186935 184688 186987
rect 149392 185751 149398 185803
rect 149450 185791 149456 185803
rect 186064 185791 186070 185803
rect 149450 185763 186070 185791
rect 149450 185751 149456 185763
rect 186064 185751 186070 185763
rect 186122 185751 186128 185803
rect 145648 184271 145654 184323
rect 145706 184311 145712 184323
rect 184336 184311 184342 184323
rect 145706 184283 184342 184311
rect 145706 184271 145712 184283
rect 184336 184271 184342 184283
rect 184394 184271 184400 184323
rect 171280 184197 171286 184249
rect 171338 184237 171344 184249
rect 184432 184237 184438 184249
rect 171338 184209 184438 184237
rect 171338 184197 171344 184209
rect 184432 184197 184438 184209
rect 184490 184197 184496 184249
rect 182896 184123 182902 184175
rect 182954 184163 182960 184175
rect 186736 184163 186742 184175
rect 182954 184135 186742 184163
rect 182954 184123 182960 184135
rect 186736 184123 186742 184135
rect 186794 184123 186800 184175
rect 645136 183087 645142 183139
rect 645194 183127 645200 183139
rect 649360 183127 649366 183139
rect 645194 183099 649366 183127
rect 645194 183087 645200 183099
rect 649360 183087 649366 183099
rect 649418 183087 649424 183139
rect 149488 182939 149494 182991
rect 149546 182979 149552 182991
rect 185968 182979 185974 182991
rect 149546 182951 185974 182979
rect 149546 182939 149552 182951
rect 185968 182939 185974 182951
rect 186026 182939 186032 182991
rect 149296 182865 149302 182917
rect 149354 182905 149360 182917
rect 186160 182905 186166 182917
rect 149354 182877 186166 182905
rect 149354 182865 149360 182877
rect 186160 182865 186166 182877
rect 186218 182865 186224 182917
rect 149392 181459 149398 181511
rect 149450 181499 149456 181511
rect 171472 181499 171478 181511
rect 149450 181471 171478 181499
rect 149450 181459 149456 181471
rect 171472 181459 171478 181471
rect 171530 181459 171536 181511
rect 182800 181385 182806 181437
rect 182858 181425 182864 181437
rect 184624 181425 184630 181437
rect 182858 181397 184630 181425
rect 182858 181385 182864 181397
rect 184624 181385 184630 181397
rect 184682 181385 184688 181437
rect 156880 181311 156886 181363
rect 156938 181351 156944 181363
rect 184336 181351 184342 181363
rect 156938 181323 184342 181351
rect 156938 181311 156944 181323
rect 184336 181311 184342 181323
rect 184394 181311 184400 181363
rect 165520 181237 165526 181289
rect 165578 181277 165584 181289
rect 184432 181277 184438 181289
rect 165578 181249 184438 181277
rect 165578 181237 165584 181249
rect 184432 181237 184438 181249
rect 184490 181237 184496 181289
rect 154000 181163 154006 181215
rect 154058 181203 154064 181215
rect 184528 181203 184534 181215
rect 154058 181175 184534 181203
rect 154058 181163 154064 181175
rect 184528 181163 184534 181175
rect 184586 181163 184592 181215
rect 149584 180053 149590 180105
rect 149642 180093 149648 180105
rect 185296 180093 185302 180105
rect 149642 180065 185302 180093
rect 149642 180053 149648 180065
rect 185296 180053 185302 180065
rect 185354 180053 185360 180105
rect 149200 179979 149206 180031
rect 149258 180019 149264 180031
rect 186448 180019 186454 180031
rect 149258 179991 186454 180019
rect 149258 179979 149264 179991
rect 186448 179979 186454 179991
rect 186506 179979 186512 180031
rect 645136 179387 645142 179439
rect 645194 179427 645200 179439
rect 649456 179427 649462 179439
rect 645194 179399 649462 179427
rect 645194 179387 645200 179399
rect 649456 179387 649462 179399
rect 649514 179387 649520 179439
rect 149392 178721 149398 178773
rect 149450 178761 149456 178773
rect 162928 178761 162934 178773
rect 149450 178733 162934 178761
rect 149450 178721 149456 178733
rect 162928 178721 162934 178733
rect 162986 178721 162992 178773
rect 149488 178647 149494 178699
rect 149546 178687 149552 178699
rect 165712 178687 165718 178699
rect 149546 178659 165718 178687
rect 149546 178647 149552 178659
rect 165712 178647 165718 178659
rect 165770 178647 165776 178699
rect 149296 178573 149302 178625
rect 149354 178613 149360 178625
rect 168496 178613 168502 178625
rect 149354 178585 168502 178613
rect 149354 178573 149360 178585
rect 168496 178573 168502 178585
rect 168554 178573 168560 178625
rect 42160 178499 42166 178551
rect 42218 178539 42224 178551
rect 50320 178539 50326 178551
rect 42218 178511 50326 178539
rect 42218 178499 42224 178511
rect 50320 178499 50326 178511
rect 50378 178499 50384 178551
rect 145360 178499 145366 178551
rect 145418 178539 145424 178551
rect 184432 178539 184438 178551
rect 145418 178511 184438 178539
rect 145418 178499 145424 178511
rect 184432 178499 184438 178511
rect 184490 178499 184496 178551
rect 162640 178425 162646 178477
rect 162698 178465 162704 178477
rect 184528 178465 184534 178477
rect 162698 178437 184534 178465
rect 162698 178425 162704 178437
rect 184528 178425 184534 178437
rect 184586 178425 184592 178477
rect 174160 178351 174166 178403
rect 174218 178391 174224 178403
rect 184336 178391 184342 178403
rect 174218 178363 184342 178391
rect 174218 178351 174224 178363
rect 184336 178351 184342 178363
rect 184394 178351 184400 178403
rect 149392 177241 149398 177293
rect 149450 177281 149456 177293
rect 156880 177281 156886 177293
rect 149450 177253 156886 177281
rect 149450 177241 149456 177253
rect 156880 177241 156886 177253
rect 156938 177241 156944 177293
rect 655696 176131 655702 176183
rect 655754 176171 655760 176183
rect 676144 176171 676150 176183
rect 655754 176143 676150 176171
rect 655754 176131 655760 176143
rect 676144 176131 676150 176143
rect 676202 176131 676208 176183
rect 147760 175983 147766 176035
rect 147818 176023 147824 176035
rect 154000 176023 154006 176035
rect 147818 175995 154006 176023
rect 147818 175983 147824 175995
rect 154000 175983 154006 175995
rect 154058 175983 154064 176035
rect 655504 175983 655510 176035
rect 655562 176023 655568 176035
rect 676240 176023 676246 176035
rect 655562 175995 676246 176023
rect 655562 175983 655568 175995
rect 676240 175983 676246 175995
rect 676298 175983 676304 176035
rect 655408 175835 655414 175887
rect 655466 175875 655472 175887
rect 676336 175875 676342 175887
rect 655466 175847 676342 175875
rect 655466 175835 655472 175847
rect 676336 175835 676342 175847
rect 676394 175835 676400 175887
rect 145552 175613 145558 175665
rect 145610 175653 145616 175665
rect 184432 175653 184438 175665
rect 145610 175625 184438 175653
rect 145610 175613 145616 175625
rect 184432 175613 184438 175625
rect 184490 175613 184496 175665
rect 145456 175539 145462 175591
rect 145514 175579 145520 175591
rect 184336 175579 184342 175591
rect 145514 175551 184342 175579
rect 145514 175539 145520 175551
rect 184336 175539 184342 175551
rect 184394 175539 184400 175591
rect 645136 174873 645142 174925
rect 645194 174913 645200 174925
rect 649552 174913 649558 174925
rect 645194 174885 649558 174913
rect 645194 174873 645200 174885
rect 649552 174873 649558 174885
rect 649610 174873 649616 174925
rect 148816 174281 148822 174333
rect 148874 174321 148880 174333
rect 149680 174321 149686 174333
rect 148874 174293 149686 174321
rect 148874 174281 148880 174293
rect 149680 174281 149686 174293
rect 149738 174281 149744 174333
rect 149200 174207 149206 174259
rect 149258 174247 149264 174259
rect 186256 174247 186262 174259
rect 149258 174219 186262 174247
rect 149258 174207 149264 174219
rect 186256 174207 186262 174219
rect 186314 174207 186320 174259
rect 149392 172801 149398 172853
rect 149450 172841 149456 172853
rect 182800 172841 182806 172853
rect 149450 172813 182806 172841
rect 149450 172801 149456 172813
rect 182800 172801 182806 172813
rect 182858 172801 182864 172853
rect 148336 172727 148342 172779
rect 148394 172767 148400 172779
rect 184624 172767 184630 172779
rect 148394 172739 184630 172767
rect 148394 172727 148400 172739
rect 184624 172727 184630 172739
rect 184682 172727 184688 172779
rect 148720 172653 148726 172705
rect 148778 172693 148784 172705
rect 184432 172693 184438 172705
rect 148778 172665 184438 172693
rect 148778 172653 148784 172665
rect 184432 172653 184438 172665
rect 184490 172653 184496 172705
rect 148528 172579 148534 172631
rect 148586 172619 148592 172631
rect 184336 172619 184342 172631
rect 148586 172591 184342 172619
rect 148586 172579 148592 172591
rect 184336 172579 184342 172591
rect 184394 172579 184400 172631
rect 149008 172505 149014 172557
rect 149066 172545 149072 172557
rect 184528 172545 184534 172557
rect 149066 172517 184534 172545
rect 149066 172505 149072 172517
rect 184528 172505 184534 172517
rect 184586 172505 184592 172557
rect 645136 171025 645142 171077
rect 645194 171065 645200 171077
rect 649648 171065 649654 171077
rect 645194 171037 649654 171065
rect 645194 171025 645200 171037
rect 649648 171025 649654 171037
rect 649706 171025 649712 171077
rect 675280 169915 675286 169967
rect 675338 169955 675344 169967
rect 676048 169955 676054 169967
rect 675338 169927 676054 169955
rect 675338 169915 675344 169927
rect 676048 169915 676054 169927
rect 676106 169915 676112 169967
rect 148240 169841 148246 169893
rect 148298 169881 148304 169893
rect 184432 169881 184438 169893
rect 148298 169853 184438 169881
rect 148298 169841 148304 169853
rect 184432 169841 184438 169853
rect 184490 169841 184496 169893
rect 148816 169767 148822 169819
rect 148874 169807 148880 169819
rect 184624 169807 184630 169819
rect 148874 169779 184630 169807
rect 148874 169767 148880 169779
rect 184624 169767 184630 169779
rect 184682 169767 184688 169819
rect 148624 169693 148630 169745
rect 148682 169733 148688 169745
rect 184336 169733 184342 169745
rect 148682 169705 184342 169733
rect 148682 169693 148688 169705
rect 184336 169693 184342 169705
rect 184394 169693 184400 169745
rect 149104 169619 149110 169671
rect 149162 169659 149168 169671
rect 184528 169659 184534 169671
rect 149162 169631 184534 169659
rect 149162 169619 149168 169631
rect 184528 169619 184534 169631
rect 184586 169619 184592 169671
rect 645136 168213 645142 168265
rect 645194 168253 645200 168265
rect 649840 168253 649846 168265
rect 645194 168225 649846 168253
rect 645194 168213 645200 168225
rect 649840 168213 649846 168225
rect 649898 168213 649904 168265
rect 674992 167103 674998 167155
rect 675050 167143 675056 167155
rect 676240 167143 676246 167155
rect 675050 167115 676246 167143
rect 675050 167103 675056 167115
rect 676240 167103 676246 167115
rect 676298 167103 676304 167155
rect 675184 167029 675190 167081
rect 675242 167069 675248 167081
rect 676048 167069 676054 167081
rect 675242 167041 676054 167069
rect 675242 167029 675248 167041
rect 676048 167029 676054 167041
rect 676106 167029 676112 167081
rect 148432 166955 148438 167007
rect 148490 166995 148496 167007
rect 184336 166995 184342 167007
rect 148490 166967 184342 166995
rect 148490 166955 148496 166967
rect 184336 166955 184342 166967
rect 184394 166955 184400 167007
rect 149680 166881 149686 166933
rect 149738 166921 149744 166933
rect 184432 166921 184438 166933
rect 149738 166893 184438 166921
rect 149738 166881 149744 166893
rect 184432 166881 184438 166893
rect 184490 166881 184496 166933
rect 154096 166807 154102 166859
rect 154154 166847 154160 166859
rect 184528 166847 184534 166859
rect 154154 166819 184534 166847
rect 154154 166807 154160 166819
rect 184528 166807 184534 166819
rect 184586 166807 184592 166859
rect 647056 164291 647062 164343
rect 647114 164331 647120 164343
rect 676240 164331 676246 164343
rect 647114 164303 676246 164331
rect 647114 164291 647120 164303
rect 676240 164291 676246 164303
rect 676298 164291 676304 164343
rect 646960 164217 646966 164269
rect 647018 164257 647024 164269
rect 676144 164257 676150 164269
rect 647018 164229 676150 164257
rect 647018 164217 647024 164229
rect 676144 164217 676150 164229
rect 676202 164217 676208 164269
rect 646864 164143 646870 164195
rect 646922 164183 646928 164195
rect 676048 164183 676054 164195
rect 646922 164155 676054 164183
rect 646922 164143 646928 164155
rect 676048 164143 676054 164155
rect 676106 164143 676112 164195
rect 151312 164069 151318 164121
rect 151370 164109 151376 164121
rect 184528 164109 184534 164121
rect 151370 164081 184534 164109
rect 151370 164069 151376 164081
rect 184528 164069 184534 164081
rect 184586 164069 184592 164121
rect 156976 163995 156982 164047
rect 157034 164035 157040 164047
rect 184336 164035 184342 164047
rect 157034 164007 184342 164035
rect 157034 163995 157040 164007
rect 184336 163995 184342 164007
rect 184394 163995 184400 164047
rect 159760 163921 159766 163973
rect 159818 163961 159824 163973
rect 184432 163961 184438 163973
rect 159818 163933 184438 163961
rect 159818 163921 159824 163933
rect 184432 163921 184438 163933
rect 184490 163921 184496 163973
rect 174256 163847 174262 163899
rect 174314 163887 174320 163899
rect 184336 163887 184342 163899
rect 174314 163859 184342 163887
rect 174314 163847 174320 163859
rect 184336 163847 184342 163859
rect 184394 163847 184400 163899
rect 645136 163329 645142 163381
rect 645194 163369 645200 163381
rect 649936 163369 649942 163381
rect 645194 163341 649942 163369
rect 645194 163329 645200 163341
rect 649936 163329 649942 163341
rect 649994 163329 650000 163381
rect 151216 161183 151222 161235
rect 151274 161223 151280 161235
rect 184432 161223 184438 161235
rect 151274 161195 184438 161223
rect 151274 161183 151280 161195
rect 184432 161183 184438 161195
rect 184490 161183 184496 161235
rect 162736 161109 162742 161161
rect 162794 161149 162800 161161
rect 184528 161149 184534 161161
rect 162794 161121 184534 161149
rect 162794 161109 162800 161121
rect 184528 161109 184534 161121
rect 184586 161109 184592 161161
rect 675664 161109 675670 161161
rect 675722 161109 675728 161161
rect 168400 161035 168406 161087
rect 168458 161075 168464 161087
rect 184624 161075 184630 161087
rect 168458 161047 184630 161075
rect 168458 161035 168464 161047
rect 184624 161035 184630 161047
rect 184682 161035 184688 161087
rect 171376 160961 171382 161013
rect 171434 161001 171440 161013
rect 184336 161001 184342 161013
rect 171434 160973 184342 161001
rect 171434 160961 171440 160973
rect 184336 160961 184342 160973
rect 184394 160961 184400 161013
rect 675682 160643 675710 161109
rect 675664 160591 675670 160643
rect 675722 160591 675728 160643
rect 670384 160443 670390 160495
rect 670442 160483 670448 160495
rect 675376 160483 675382 160495
rect 670442 160455 675382 160483
rect 670442 160443 670448 160455
rect 675376 160443 675382 160455
rect 675434 160443 675440 160495
rect 645136 159703 645142 159755
rect 645194 159743 645200 159755
rect 650032 159743 650038 159755
rect 645194 159715 650038 159743
rect 645194 159703 645200 159715
rect 650032 159703 650038 159715
rect 650090 159703 650096 159755
rect 147088 158445 147094 158497
rect 147146 158485 147152 158497
rect 151312 158485 151318 158497
rect 147146 158457 151318 158485
rect 147146 158445 147152 158457
rect 151312 158445 151318 158457
rect 151370 158445 151376 158497
rect 151408 158371 151414 158423
rect 151466 158411 151472 158423
rect 184336 158411 184342 158423
rect 151466 158383 184342 158411
rect 151466 158371 151472 158383
rect 184336 158371 184342 158383
rect 184394 158371 184400 158423
rect 165616 158297 165622 158349
rect 165674 158337 165680 158349
rect 184432 158337 184438 158349
rect 165674 158309 184438 158337
rect 165674 158297 165680 158309
rect 184432 158297 184438 158309
rect 184490 158297 184496 158349
rect 179920 158223 179926 158275
rect 179978 158263 179984 158275
rect 184528 158263 184534 158275
rect 179978 158235 184534 158263
rect 179978 158223 179984 158235
rect 184528 158223 184534 158235
rect 184586 158223 184592 158275
rect 177136 158149 177142 158201
rect 177194 158189 177200 158201
rect 184624 158189 184630 158201
rect 177194 158161 184630 158189
rect 177194 158149 177200 158161
rect 184624 158149 184630 158161
rect 184682 158149 184688 158201
rect 146896 156151 146902 156203
rect 146954 156191 146960 156203
rect 151216 156191 151222 156203
rect 146954 156163 151222 156191
rect 146954 156151 146960 156163
rect 151216 156151 151222 156163
rect 151274 156151 151280 156203
rect 645136 156003 645142 156055
rect 645194 156043 645200 156055
rect 650128 156043 650134 156055
rect 645194 156015 650134 156043
rect 645194 156003 645200 156015
rect 650128 156003 650134 156015
rect 650186 156003 650192 156055
rect 149680 155633 149686 155685
rect 149738 155673 149744 155685
rect 177040 155673 177046 155685
rect 149738 155645 177046 155673
rect 149738 155633 149744 155645
rect 177040 155633 177046 155645
rect 177098 155633 177104 155685
rect 148816 155559 148822 155611
rect 148874 155599 148880 155611
rect 180016 155599 180022 155611
rect 148874 155571 180022 155599
rect 148874 155559 148880 155571
rect 180016 155559 180022 155571
rect 180074 155559 180080 155611
rect 151696 155485 151702 155537
rect 151754 155525 151760 155537
rect 184528 155525 184534 155537
rect 151754 155497 184534 155525
rect 151754 155485 151760 155497
rect 184528 155485 184534 155497
rect 184586 155485 184592 155537
rect 658000 155485 658006 155537
rect 658058 155525 658064 155537
rect 670384 155525 670390 155537
rect 658058 155497 670390 155525
rect 658058 155485 658064 155497
rect 670384 155485 670390 155497
rect 670442 155485 670448 155537
rect 152080 155411 152086 155463
rect 152138 155451 152144 155463
rect 184624 155451 184630 155463
rect 152138 155423 184630 155451
rect 152138 155411 152144 155423
rect 184624 155411 184630 155423
rect 184682 155411 184688 155463
rect 159952 155337 159958 155389
rect 160010 155377 160016 155389
rect 184432 155377 184438 155389
rect 160010 155349 184438 155377
rect 160010 155337 160016 155349
rect 184432 155337 184438 155349
rect 184490 155337 184496 155389
rect 174352 155263 174358 155315
rect 174410 155303 174416 155315
rect 184336 155303 184342 155315
rect 174410 155275 184342 155303
rect 174410 155263 174416 155275
rect 184336 155263 184342 155275
rect 184394 155263 184400 155315
rect 148816 153191 148822 153243
rect 148874 153231 148880 153243
rect 149488 153231 149494 153243
rect 148874 153203 149494 153231
rect 148874 153191 148880 153203
rect 149488 153191 149494 153203
rect 149546 153191 149552 153243
rect 149488 152747 149494 152799
rect 149546 152787 149552 152799
rect 174160 152787 174166 152799
rect 149546 152759 174166 152787
rect 149546 152747 149552 152759
rect 174160 152747 174166 152759
rect 174218 152747 174224 152799
rect 149296 152673 149302 152725
rect 149354 152713 149360 152725
rect 182896 152713 182902 152725
rect 149354 152685 182902 152713
rect 149354 152673 149360 152685
rect 182896 152673 182902 152685
rect 182954 152673 182960 152725
rect 151888 152599 151894 152651
rect 151946 152639 151952 152651
rect 184528 152639 184534 152651
rect 151946 152611 184534 152639
rect 151946 152599 151952 152611
rect 184528 152599 184534 152611
rect 184586 152599 184592 152651
rect 151792 152525 151798 152577
rect 151850 152565 151856 152577
rect 184336 152565 184342 152577
rect 151850 152537 184342 152565
rect 151850 152525 151856 152537
rect 184336 152525 184342 152537
rect 184394 152525 184400 152577
rect 645136 152525 645142 152577
rect 645194 152565 645200 152577
rect 650224 152565 650230 152577
rect 645194 152537 650230 152565
rect 645194 152525 645200 152537
rect 650224 152525 650230 152537
rect 650282 152525 650288 152577
rect 151600 152451 151606 152503
rect 151658 152491 151664 152503
rect 184432 152491 184438 152503
rect 151658 152463 184438 152491
rect 151658 152451 151664 152463
rect 184432 152451 184438 152463
rect 184490 152451 184496 152503
rect 149296 149935 149302 149987
rect 149354 149975 149360 149987
rect 171376 149975 171382 149987
rect 149354 149947 171382 149975
rect 149354 149935 149360 149947
rect 171376 149935 171382 149947
rect 171434 149935 171440 149987
rect 149488 149861 149494 149913
rect 149546 149901 149552 149913
rect 174256 149901 174262 149913
rect 149546 149873 174262 149901
rect 149546 149861 149552 149873
rect 174256 149861 174262 149873
rect 174314 149861 174320 149913
rect 149680 149787 149686 149839
rect 149738 149827 149744 149839
rect 180208 149827 180214 149839
rect 149738 149799 180214 149827
rect 149738 149787 149744 149799
rect 180208 149787 180214 149799
rect 180266 149787 180272 149839
rect 182992 149713 182998 149765
rect 183050 149753 183056 149765
rect 186736 149753 186742 149765
rect 183050 149725 186742 149753
rect 183050 149713 183056 149725
rect 186736 149713 186742 149725
rect 186794 149713 186800 149765
rect 151984 149639 151990 149691
rect 152042 149679 152048 149691
rect 184432 149679 184438 149691
rect 152042 149651 184438 149679
rect 152042 149639 152048 149651
rect 184432 149639 184438 149651
rect 184490 149639 184496 149691
rect 180112 149565 180118 149617
rect 180170 149605 180176 149617
rect 184528 149605 184534 149617
rect 180170 149577 184534 149605
rect 180170 149565 180176 149577
rect 184528 149565 184534 149577
rect 184586 149565 184592 149617
rect 151504 149491 151510 149543
rect 151562 149531 151568 149543
rect 184336 149531 184342 149543
rect 151562 149503 184342 149531
rect 151562 149491 151568 149503
rect 184336 149491 184342 149503
rect 184394 149491 184400 149543
rect 645136 148159 645142 148211
rect 645194 148199 645200 148211
rect 650320 148199 650326 148211
rect 645194 148171 650326 148199
rect 645194 148159 645200 148171
rect 650320 148159 650326 148171
rect 650378 148159 650384 148211
rect 149488 146975 149494 147027
rect 149546 147015 149552 147027
rect 168400 147015 168406 147027
rect 149546 146987 168406 147015
rect 149546 146975 149552 146987
rect 168400 146975 168406 146987
rect 168458 146975 168464 147027
rect 149296 146901 149302 146953
rect 149354 146941 149360 146953
rect 177136 146941 177142 146953
rect 149354 146913 177142 146941
rect 149354 146901 149360 146913
rect 177136 146901 177142 146913
rect 177194 146901 177200 146953
rect 154192 146827 154198 146879
rect 154250 146867 154256 146879
rect 184528 146867 184534 146879
rect 154250 146839 184534 146867
rect 154250 146827 154256 146839
rect 184528 146827 184534 146839
rect 184586 146827 184592 146879
rect 162832 146753 162838 146805
rect 162890 146793 162896 146805
rect 184432 146793 184438 146805
rect 162890 146765 184438 146793
rect 162890 146753 162896 146765
rect 184432 146753 184438 146765
rect 184490 146753 184496 146805
rect 174448 146679 174454 146731
rect 174506 146719 174512 146731
rect 184336 146719 184342 146731
rect 174506 146691 184342 146719
rect 174506 146679 174512 146691
rect 184336 146679 184342 146691
rect 184394 146679 184400 146731
rect 177232 146605 177238 146657
rect 177290 146645 177296 146657
rect 184624 146645 184630 146657
rect 177290 146617 184630 146645
rect 177290 146605 177296 146617
rect 184624 146605 184630 146617
rect 184682 146605 184688 146657
rect 147664 145717 147670 145769
rect 147722 145757 147728 145769
rect 165520 145757 165526 145769
rect 147722 145729 165526 145757
rect 147722 145717 147728 145729
rect 165520 145717 165526 145729
rect 165578 145717 165584 145769
rect 147664 144015 147670 144067
rect 147722 144055 147728 144067
rect 162736 144055 162742 144067
rect 147722 144027 162742 144055
rect 147722 144015 147728 144027
rect 162736 144015 162742 144027
rect 162794 144015 162800 144067
rect 183088 143941 183094 143993
rect 183146 143981 183152 143993
rect 184624 143981 184630 143993
rect 183146 143953 184630 143981
rect 183146 143941 183152 143953
rect 184624 143941 184630 143953
rect 184682 143941 184688 143993
rect 168592 143867 168598 143919
rect 168650 143907 168656 143919
rect 184432 143907 184438 143919
rect 168650 143879 184438 143907
rect 168650 143867 168656 143879
rect 184432 143867 184438 143879
rect 184490 143867 184496 143919
rect 171568 143793 171574 143845
rect 171626 143833 171632 143845
rect 184336 143833 184342 143845
rect 171626 143805 184342 143833
rect 171626 143793 171632 143805
rect 184336 143793 184342 143805
rect 184394 143793 184400 143845
rect 165808 143719 165814 143771
rect 165866 143759 165872 143771
rect 184528 143759 184534 143771
rect 165866 143731 184534 143759
rect 165866 143719 165872 143731
rect 184528 143719 184534 143731
rect 184586 143719 184592 143771
rect 147280 142461 147286 142513
rect 147338 142501 147344 142513
rect 159856 142501 159862 142513
rect 147338 142473 159862 142501
rect 147338 142461 147344 142473
rect 159856 142461 159862 142473
rect 159914 142461 159920 142513
rect 147472 142165 147478 142217
rect 147530 142205 147536 142217
rect 156976 142205 156982 142217
rect 147530 142177 156982 142205
rect 147530 142165 147536 142177
rect 156976 142165 156982 142177
rect 157034 142165 157040 142217
rect 149680 141203 149686 141255
rect 149738 141243 149744 141255
rect 154096 141243 154102 141255
rect 149738 141215 154102 141243
rect 149738 141203 149744 141215
rect 154096 141203 154102 141215
rect 154154 141203 154160 141255
rect 154288 141055 154294 141107
rect 154346 141095 154352 141107
rect 184528 141095 184534 141107
rect 154346 141067 184534 141095
rect 154346 141055 154352 141067
rect 184528 141055 184534 141067
rect 184586 141055 184592 141107
rect 157072 140981 157078 141033
rect 157130 141021 157136 141033
rect 184432 141021 184438 141033
rect 157130 140993 184438 141021
rect 157130 140981 157136 140993
rect 184432 140981 184438 140993
rect 184490 140981 184496 141033
rect 160048 140907 160054 140959
rect 160106 140947 160112 140959
rect 184336 140947 184342 140959
rect 160106 140919 184342 140947
rect 160106 140907 160112 140919
rect 184336 140907 184342 140919
rect 184394 140907 184400 140959
rect 147472 140315 147478 140367
rect 147530 140355 147536 140367
rect 151120 140355 151126 140367
rect 147530 140327 151126 140355
rect 147530 140315 147536 140327
rect 151120 140315 151126 140327
rect 151178 140315 151184 140367
rect 147664 138243 147670 138295
rect 147722 138283 147728 138295
rect 159760 138283 159766 138295
rect 147722 138255 159766 138283
rect 147722 138243 147728 138255
rect 159760 138243 159766 138255
rect 159818 138243 159824 138295
rect 148624 136911 148630 136963
rect 148682 136911 148688 136963
rect 148336 136689 148342 136741
rect 148394 136729 148400 136741
rect 148642 136729 148670 136911
rect 149008 136837 149014 136889
rect 149066 136877 149072 136889
rect 149200 136877 149206 136889
rect 149066 136849 149206 136877
rect 149066 136837 149072 136849
rect 149200 136837 149206 136849
rect 149258 136837 149264 136889
rect 148816 136763 148822 136815
rect 148874 136763 148880 136815
rect 148394 136701 148670 136729
rect 148834 136729 148862 136763
rect 149200 136729 149206 136741
rect 148834 136701 149206 136729
rect 148394 136689 148400 136701
rect 149200 136689 149206 136701
rect 149258 136689 149264 136741
rect 149680 135431 149686 135483
rect 149738 135471 149744 135483
rect 171280 135471 171286 135483
rect 149738 135443 171286 135471
rect 149738 135431 149744 135443
rect 171280 135431 171286 135443
rect 171338 135431 171344 135483
rect 149584 135357 149590 135409
rect 149642 135397 149648 135409
rect 179920 135397 179926 135409
rect 149642 135369 179926 135397
rect 149642 135357 149648 135369
rect 179920 135357 179926 135369
rect 179978 135357 179984 135409
rect 168496 135283 168502 135335
rect 168554 135323 168560 135335
rect 184432 135323 184438 135335
rect 168554 135295 184438 135323
rect 168554 135283 168560 135295
rect 184432 135283 184438 135295
rect 184490 135283 184496 135335
rect 171472 135209 171478 135261
rect 171530 135249 171536 135261
rect 184336 135249 184342 135261
rect 171530 135221 184342 135249
rect 171530 135209 171536 135221
rect 184336 135209 184342 135221
rect 184394 135209 184400 135261
rect 177136 134321 177142 134373
rect 177194 134361 177200 134373
rect 184720 134361 184726 134373
rect 177194 134333 184726 134361
rect 177194 134321 177200 134333
rect 184720 134321 184726 134333
rect 184778 134321 184784 134373
rect 149680 132471 149686 132523
rect 149738 132511 149744 132523
rect 182992 132511 182998 132523
rect 149738 132483 182998 132511
rect 149738 132471 149744 132483
rect 182992 132471 182998 132483
rect 183050 132471 183056 132523
rect 154000 132397 154006 132449
rect 154058 132437 154064 132449
rect 184624 132437 184630 132449
rect 154058 132409 184630 132437
rect 154058 132397 154064 132409
rect 184624 132397 184630 132409
rect 184682 132397 184688 132449
rect 156880 132323 156886 132375
rect 156938 132363 156944 132375
rect 184528 132363 184534 132375
rect 156938 132335 184534 132363
rect 156938 132323 156944 132335
rect 184528 132323 184534 132335
rect 184586 132323 184592 132375
rect 162928 132249 162934 132301
rect 162986 132289 162992 132301
rect 184432 132289 184438 132301
rect 162986 132261 184438 132289
rect 162986 132249 162992 132261
rect 184432 132249 184438 132261
rect 184490 132249 184496 132301
rect 165712 132175 165718 132227
rect 165770 132215 165776 132227
rect 184336 132215 184342 132227
rect 165770 132187 184342 132215
rect 165770 132175 165776 132187
rect 184336 132175 184342 132187
rect 184394 132175 184400 132227
rect 655312 130103 655318 130155
rect 655370 130143 655376 130155
rect 676144 130143 676150 130155
rect 655370 130115 676150 130143
rect 655370 130103 655376 130115
rect 676144 130103 676150 130115
rect 676202 130103 676208 130155
rect 655216 129955 655222 130007
rect 655274 129995 655280 130007
rect 676240 129995 676246 130007
rect 655274 129967 676246 129995
rect 655274 129955 655280 129967
rect 676240 129955 676246 129967
rect 676298 129955 676304 130007
rect 655120 129807 655126 129859
rect 655178 129847 655184 129859
rect 676336 129847 676342 129859
rect 655178 129819 676342 129847
rect 655178 129807 655184 129819
rect 676336 129807 676342 129819
rect 676394 129807 676400 129859
rect 147472 129659 147478 129711
rect 147530 129699 147536 129711
rect 165616 129699 165622 129711
rect 147530 129671 165622 129699
rect 147530 129659 147536 129671
rect 165616 129659 165622 129671
rect 165674 129659 165680 129711
rect 149680 129585 149686 129637
rect 149738 129625 149744 129637
rect 168496 129625 168502 129637
rect 149738 129597 168502 129625
rect 149738 129585 149744 129597
rect 168496 129585 168502 129597
rect 168554 129585 168560 129637
rect 180208 129585 180214 129637
rect 180266 129625 180272 129637
rect 185680 129625 185686 129637
rect 180266 129597 185686 129625
rect 180266 129585 180272 129597
rect 185680 129585 185686 129597
rect 185738 129585 185744 129637
rect 645712 129585 645718 129637
rect 645770 129625 645776 129637
rect 676240 129625 676246 129637
rect 645770 129597 676246 129625
rect 645770 129585 645776 129597
rect 676240 129585 676246 129597
rect 676298 129585 676304 129637
rect 182800 129511 182806 129563
rect 182858 129551 182864 129563
rect 186736 129551 186742 129563
rect 182858 129523 186742 129551
rect 182858 129511 182864 129523
rect 186736 129511 186742 129523
rect 186794 129511 186800 129563
rect 149392 129437 149398 129489
rect 149450 129477 149456 129489
rect 184432 129477 184438 129489
rect 149450 129449 184438 129477
rect 149450 129437 149456 129449
rect 184432 129437 184438 129449
rect 184490 129437 184496 129489
rect 149488 129363 149494 129415
rect 149546 129403 149552 129415
rect 184528 129403 184534 129415
rect 149546 129375 184534 129403
rect 149546 129363 149552 129375
rect 184528 129363 184534 129375
rect 184586 129363 184592 129415
rect 149104 129289 149110 129341
rect 149162 129329 149168 129341
rect 184336 129329 184342 129341
rect 149162 129301 184342 129329
rect 149162 129289 149168 129301
rect 184336 129289 184342 129301
rect 184394 129289 184400 129341
rect 147664 127291 147670 127343
rect 147722 127331 147728 127343
rect 162640 127331 162646 127343
rect 147722 127303 162646 127331
rect 147722 127291 147728 127303
rect 162640 127291 162646 127303
rect 162698 127291 162704 127343
rect 646480 126847 646486 126899
rect 646538 126887 646544 126899
rect 676240 126887 676246 126899
rect 646538 126859 676246 126887
rect 646538 126847 646544 126859
rect 676240 126847 676246 126859
rect 676298 126847 676304 126899
rect 646576 126773 646582 126825
rect 646634 126813 646640 126825
rect 676144 126813 676150 126825
rect 646634 126785 676150 126813
rect 646634 126773 646640 126785
rect 676144 126773 676150 126785
rect 676202 126773 676208 126825
rect 674128 126699 674134 126751
rect 674186 126739 674192 126751
rect 676048 126739 676054 126751
rect 674186 126711 676054 126739
rect 674186 126699 674192 126711
rect 676048 126699 676054 126711
rect 676106 126699 676112 126751
rect 149008 126625 149014 126677
rect 149066 126665 149072 126677
rect 184432 126665 184438 126677
rect 149066 126637 184438 126665
rect 149066 126625 149072 126637
rect 184432 126625 184438 126637
rect 184490 126625 184496 126677
rect 148720 126551 148726 126603
rect 148778 126591 148784 126603
rect 184528 126591 184534 126603
rect 148778 126563 184534 126591
rect 148778 126551 148784 126563
rect 184528 126551 184534 126563
rect 184586 126551 184592 126603
rect 149200 126477 149206 126529
rect 149258 126517 149264 126529
rect 184336 126517 184342 126529
rect 149258 126489 184342 126517
rect 149258 126477 149264 126489
rect 184336 126477 184342 126489
rect 184394 126477 184400 126529
rect 674320 124627 674326 124679
rect 674378 124667 674384 124679
rect 676048 124667 676054 124679
rect 674378 124639 676054 124667
rect 674378 124627 674384 124639
rect 676048 124627 676054 124639
rect 676106 124627 676112 124679
rect 149392 124035 149398 124087
rect 149450 124075 149456 124087
rect 156880 124075 156886 124087
rect 149450 124047 156886 124075
rect 149450 124035 149456 124047
rect 156880 124035 156886 124047
rect 156938 124035 156944 124087
rect 674032 124035 674038 124087
rect 674090 124075 674096 124087
rect 675952 124075 675958 124087
rect 674090 124047 675958 124075
rect 674090 124035 674096 124047
rect 675952 124035 675958 124047
rect 676010 124035 676016 124087
rect 674416 123961 674422 124013
rect 674474 124001 674480 124013
rect 676048 124001 676054 124013
rect 674474 123973 676054 124001
rect 674474 123961 674480 123973
rect 676048 123961 676054 123973
rect 676106 123961 676112 124013
rect 675088 123887 675094 123939
rect 675146 123927 675152 123939
rect 676240 123927 676246 123939
rect 675146 123899 676246 123927
rect 675146 123887 675152 123899
rect 676240 123887 676246 123899
rect 676298 123887 676304 123939
rect 148432 123813 148438 123865
rect 148490 123853 148496 123865
rect 184528 123853 184534 123865
rect 148490 123825 184534 123853
rect 148490 123813 148496 123825
rect 184528 123813 184534 123825
rect 184586 123813 184592 123865
rect 148528 123739 148534 123791
rect 148586 123779 148592 123791
rect 184336 123779 184342 123791
rect 148586 123751 184342 123779
rect 148586 123739 148592 123751
rect 184336 123739 184342 123751
rect 184394 123739 184400 123791
rect 148240 123665 148246 123717
rect 148298 123705 148304 123717
rect 184432 123705 184438 123717
rect 148298 123677 184438 123705
rect 148298 123665 148304 123677
rect 184432 123665 184438 123677
rect 184490 123665 184496 123717
rect 148624 123591 148630 123643
rect 148682 123631 148688 123643
rect 184336 123631 184342 123643
rect 148682 123603 184342 123631
rect 148682 123591 148688 123603
rect 184336 123591 184342 123603
rect 184394 123591 184400 123643
rect 174256 122407 174262 122459
rect 174314 122447 174320 122459
rect 186160 122447 186166 122459
rect 174314 122419 186166 122447
rect 174314 122407 174320 122419
rect 186160 122407 186166 122419
rect 186218 122407 186224 122459
rect 674608 122111 674614 122163
rect 674666 122151 674672 122163
rect 676048 122151 676054 122163
rect 674666 122123 676054 122151
rect 674666 122111 674672 122123
rect 676048 122111 676054 122123
rect 676106 122111 676112 122163
rect 674512 121149 674518 121201
rect 674570 121189 674576 121201
rect 676048 121189 676054 121201
rect 674570 121161 676054 121189
rect 674570 121149 674576 121161
rect 676048 121149 676054 121161
rect 676106 121149 676112 121201
rect 674224 121075 674230 121127
rect 674282 121115 674288 121127
rect 676240 121115 676246 121127
rect 674282 121087 676246 121115
rect 674282 121075 674288 121087
rect 676240 121075 676246 121087
rect 676298 121075 676304 121127
rect 674800 121001 674806 121053
rect 674858 121041 674864 121053
rect 676048 121041 676054 121053
rect 674858 121013 676054 121041
rect 674858 121001 674864 121013
rect 676048 121001 676054 121013
rect 676106 121001 676112 121053
rect 148144 120927 148150 120979
rect 148202 120967 148208 120979
rect 184336 120967 184342 120979
rect 148202 120939 184342 120967
rect 148202 120927 148208 120939
rect 184336 120927 184342 120939
rect 184394 120927 184400 120979
rect 148336 120853 148342 120905
rect 148394 120893 148400 120905
rect 184432 120893 184438 120905
rect 148394 120865 184438 120893
rect 148394 120853 148400 120865
rect 184432 120853 184438 120865
rect 184490 120853 184496 120905
rect 171376 120779 171382 120831
rect 171434 120819 171440 120831
rect 184528 120819 184534 120831
rect 171434 120791 184534 120819
rect 171434 120779 171440 120791
rect 184528 120779 184534 120791
rect 184586 120779 184592 120831
rect 147472 119891 147478 119943
rect 147530 119931 147536 119943
rect 153136 119931 153142 119943
rect 147530 119903 153142 119931
rect 147530 119891 147536 119903
rect 153136 119891 153142 119903
rect 153194 119891 153200 119943
rect 647824 118337 647830 118389
rect 647882 118377 647888 118389
rect 676240 118377 676246 118389
rect 647882 118349 676246 118377
rect 647882 118337 647888 118349
rect 676240 118337 676246 118349
rect 676298 118337 676304 118389
rect 149392 118189 149398 118241
rect 149450 118229 149456 118241
rect 168592 118229 168598 118241
rect 149450 118201 168598 118229
rect 149450 118189 149456 118201
rect 168592 118189 168598 118201
rect 168650 118189 168656 118241
rect 647920 118189 647926 118241
rect 647978 118229 647984 118241
rect 676144 118229 676150 118241
rect 647978 118201 676150 118229
rect 647978 118189 647984 118201
rect 676144 118189 676150 118201
rect 676202 118189 676208 118241
rect 149488 118115 149494 118167
rect 149546 118155 149552 118167
rect 174256 118155 174262 118167
rect 149546 118127 174262 118155
rect 149546 118115 149552 118127
rect 174256 118115 174262 118127
rect 174314 118115 174320 118167
rect 645232 118115 645238 118167
rect 645290 118155 645296 118167
rect 676048 118155 676054 118167
rect 645290 118127 676054 118155
rect 645290 118115 645296 118127
rect 676048 118115 676054 118127
rect 676106 118115 676112 118167
rect 159856 118041 159862 118093
rect 159914 118081 159920 118093
rect 184624 118081 184630 118093
rect 159914 118053 184630 118081
rect 159914 118041 159920 118053
rect 184624 118041 184630 118053
rect 184682 118041 184688 118093
rect 162736 117967 162742 118019
rect 162794 118007 162800 118019
rect 184528 118007 184534 118019
rect 162794 117979 184534 118007
rect 162794 117967 162800 117979
rect 184528 117967 184534 117979
rect 184586 117967 184592 118019
rect 165520 117893 165526 117945
rect 165578 117933 165584 117945
rect 184432 117933 184438 117945
rect 165578 117905 184438 117933
rect 165578 117893 165584 117905
rect 184432 117893 184438 117905
rect 184490 117893 184496 117945
rect 168400 117819 168406 117871
rect 168458 117859 168464 117871
rect 184336 117859 184342 117871
rect 168458 117831 184342 117859
rect 168458 117819 168464 117831
rect 184336 117819 184342 117831
rect 184394 117819 184400 117871
rect 675088 115377 675094 115429
rect 675146 115417 675152 115429
rect 675280 115417 675286 115429
rect 675146 115389 675286 115417
rect 675146 115377 675152 115389
rect 675280 115377 675286 115389
rect 675338 115377 675344 115429
rect 149392 115303 149398 115355
rect 149450 115343 149456 115355
rect 162832 115343 162838 115355
rect 149450 115315 162838 115343
rect 149450 115303 149456 115315
rect 162832 115303 162838 115315
rect 162890 115303 162896 115355
rect 149488 115229 149494 115281
rect 149546 115269 149552 115281
rect 165712 115269 165718 115281
rect 149546 115241 165718 115269
rect 149546 115229 149552 115241
rect 165712 115229 165718 115241
rect 165770 115229 165776 115281
rect 647920 115229 647926 115281
rect 647978 115269 647984 115281
rect 665296 115269 665302 115281
rect 647978 115241 665302 115269
rect 647978 115229 647984 115241
rect 665296 115229 665302 115241
rect 665354 115229 665360 115281
rect 151312 115155 151318 115207
rect 151370 115195 151376 115207
rect 184528 115195 184534 115207
rect 151370 115167 184534 115195
rect 151370 115155 151376 115167
rect 184528 115155 184534 115167
rect 184586 115155 184592 115207
rect 663760 115155 663766 115207
rect 663818 115195 663824 115207
rect 665200 115195 665206 115207
rect 663818 115167 665206 115195
rect 663818 115155 663824 115167
rect 665200 115155 665206 115167
rect 665258 115155 665264 115207
rect 154096 115081 154102 115133
rect 154154 115121 154160 115133
rect 184432 115121 184438 115133
rect 154154 115093 184438 115121
rect 154154 115081 154160 115093
rect 184432 115081 184438 115093
rect 184490 115081 184496 115133
rect 156976 115007 156982 115059
rect 157034 115047 157040 115059
rect 184336 115047 184342 115059
rect 157034 115019 184342 115047
rect 157034 115007 157040 115019
rect 184336 115007 184342 115019
rect 184394 115007 184400 115059
rect 674416 114933 674422 114985
rect 674474 114973 674480 114985
rect 675184 114973 675190 114985
rect 674474 114945 675190 114973
rect 674474 114933 674480 114945
rect 675184 114933 675190 114945
rect 675242 114933 675248 114985
rect 674608 114563 674614 114615
rect 674666 114603 674672 114615
rect 674666 114575 675326 114603
rect 674666 114563 674672 114575
rect 675298 114393 675326 114575
rect 180016 114341 180022 114393
rect 180074 114381 180080 114393
rect 184624 114381 184630 114393
rect 180074 114353 184630 114381
rect 180074 114341 180080 114353
rect 184624 114341 184630 114353
rect 184682 114341 184688 114393
rect 675280 114341 675286 114393
rect 675338 114341 675344 114393
rect 674128 114119 674134 114171
rect 674186 114159 674192 114171
rect 675376 114159 675382 114171
rect 674186 114131 675382 114159
rect 674186 114119 674192 114131
rect 675376 114119 675382 114131
rect 675434 114119 675440 114171
rect 149488 113009 149494 113061
rect 149546 113049 149552 113061
rect 159856 113049 159862 113061
rect 149546 113021 159862 113049
rect 149546 113009 149552 113021
rect 159856 113009 159862 113021
rect 159914 113009 159920 113061
rect 674320 112491 674326 112543
rect 674378 112531 674384 112543
rect 675376 112531 675382 112543
rect 674378 112503 675382 112531
rect 674378 112491 674384 112503
rect 675376 112491 675382 112503
rect 675434 112491 675440 112543
rect 149392 112343 149398 112395
rect 149450 112383 149456 112395
rect 177136 112383 177142 112395
rect 149450 112355 177142 112383
rect 149450 112343 149456 112355
rect 177136 112343 177142 112355
rect 177194 112343 177200 112395
rect 151216 112269 151222 112321
rect 151274 112309 151280 112321
rect 184336 112309 184342 112321
rect 151274 112281 184342 112309
rect 151274 112269 151280 112281
rect 184336 112269 184342 112281
rect 184394 112269 184400 112321
rect 665200 112269 665206 112321
rect 665258 112309 665264 112321
rect 675088 112309 675094 112321
rect 665258 112281 675094 112309
rect 665258 112269 665264 112281
rect 675088 112269 675094 112281
rect 675146 112269 675152 112321
rect 182896 112195 182902 112247
rect 182954 112235 182960 112247
rect 184528 112235 184534 112247
rect 182954 112207 184534 112235
rect 182954 112195 182960 112207
rect 184528 112195 184534 112207
rect 184586 112195 184592 112247
rect 177040 112121 177046 112173
rect 177098 112161 177104 112173
rect 184432 112161 184438 112173
rect 177098 112133 184438 112161
rect 177098 112121 177104 112133
rect 184432 112121 184438 112133
rect 184490 112121 184496 112173
rect 674512 112121 674518 112173
rect 674570 112161 674576 112173
rect 675088 112161 675094 112173
rect 674570 112133 675094 112161
rect 674570 112121 674576 112133
rect 675088 112121 675094 112133
rect 675146 112121 675152 112173
rect 674032 111677 674038 111729
rect 674090 111717 674096 111729
rect 675376 111717 675382 111729
rect 674090 111689 675382 111717
rect 674090 111677 674096 111689
rect 675376 111677 675382 111689
rect 675434 111677 675440 111729
rect 149392 110789 149398 110841
rect 149450 110829 149456 110841
rect 156976 110829 156982 110841
rect 149450 110801 156982 110829
rect 149450 110789 149456 110801
rect 156976 110789 156982 110801
rect 157034 110789 157040 110841
rect 674224 110049 674230 110101
rect 674282 110089 674288 110101
rect 675088 110089 675094 110101
rect 674282 110061 675094 110089
rect 674282 110049 674288 110061
rect 675088 110049 675094 110061
rect 675146 110049 675152 110101
rect 148624 109531 148630 109583
rect 148682 109571 148688 109583
rect 154000 109571 154006 109583
rect 148682 109543 154006 109571
rect 148682 109531 148688 109543
rect 154000 109531 154006 109543
rect 154058 109531 154064 109583
rect 159760 109383 159766 109435
rect 159818 109423 159824 109435
rect 184432 109423 184438 109435
rect 159818 109395 184438 109423
rect 159818 109383 159824 109395
rect 184432 109383 184438 109395
rect 184490 109383 184496 109435
rect 174160 109309 174166 109361
rect 174218 109349 174224 109361
rect 184336 109349 184342 109361
rect 174218 109321 184342 109349
rect 174218 109309 174224 109321
rect 184336 109309 184342 109321
rect 184394 109309 184400 109361
rect 147184 108347 147190 108399
rect 147242 108387 147248 108399
rect 151120 108387 151126 108399
rect 147242 108359 151126 108387
rect 147242 108347 147248 108359
rect 151120 108347 151126 108359
rect 151178 108347 151184 108399
rect 182992 106497 182998 106549
rect 183050 106537 183056 106549
rect 184528 106537 184534 106549
rect 183050 106509 184534 106537
rect 183050 106497 183056 106509
rect 184528 106497 184534 106509
rect 184586 106497 184592 106549
rect 171280 106423 171286 106475
rect 171338 106463 171344 106475
rect 184336 106463 184342 106475
rect 171338 106435 184342 106463
rect 171338 106423 171344 106435
rect 184336 106423 184342 106435
rect 184394 106423 184400 106475
rect 179920 106349 179926 106401
rect 179978 106389 179984 106401
rect 185296 106389 185302 106401
rect 179978 106361 185302 106389
rect 179978 106349 179984 106361
rect 185296 106349 185302 106361
rect 185354 106349 185360 106401
rect 149008 106275 149014 106327
rect 149066 106315 149072 106327
rect 184432 106315 184438 106327
rect 149066 106287 184438 106315
rect 149066 106275 149072 106287
rect 184432 106275 184438 106287
rect 184490 106275 184496 106327
rect 153136 105091 153142 105143
rect 153194 105131 153200 105143
rect 184720 105131 184726 105143
rect 153194 105103 184726 105131
rect 153194 105091 153200 105103
rect 184720 105091 184726 105103
rect 184778 105091 184784 105143
rect 654064 104499 654070 104551
rect 654122 104539 654128 104551
rect 665200 104539 665206 104551
rect 654122 104511 665206 104539
rect 654122 104499 654128 104511
rect 665200 104499 665206 104511
rect 665258 104499 665264 104551
rect 647920 103907 647926 103959
rect 647978 103947 647984 103959
rect 661168 103947 661174 103959
rect 647978 103919 661174 103947
rect 647978 103907 647984 103919
rect 661168 103907 661174 103919
rect 661226 103907 661232 103959
rect 646096 103833 646102 103885
rect 646154 103873 646160 103885
rect 657520 103873 657526 103885
rect 646154 103845 657526 103873
rect 646154 103833 646160 103845
rect 657520 103833 657526 103845
rect 657578 103833 657584 103885
rect 643600 103685 643606 103737
rect 643658 103725 643664 103737
rect 665584 103725 665590 103737
rect 643658 103697 665590 103725
rect 643658 103685 643664 103697
rect 665584 103685 665590 103697
rect 665642 103685 665648 103737
rect 148816 103611 148822 103663
rect 148874 103651 148880 103663
rect 184432 103651 184438 103663
rect 148874 103623 184438 103651
rect 148874 103611 148880 103623
rect 184432 103611 184438 103623
rect 184490 103611 184496 103663
rect 149584 103537 149590 103589
rect 149642 103577 149648 103589
rect 184624 103577 184630 103589
rect 149642 103549 184630 103577
rect 149642 103537 149648 103549
rect 184624 103537 184630 103549
rect 184682 103537 184688 103589
rect 165616 103463 165622 103515
rect 165674 103503 165680 103515
rect 184528 103503 184534 103515
rect 165674 103475 184534 103503
rect 165674 103463 165680 103475
rect 184528 103463 184534 103475
rect 184586 103463 184592 103515
rect 168496 103389 168502 103441
rect 168554 103429 168560 103441
rect 184336 103429 184342 103441
rect 168554 103401 184342 103429
rect 168554 103389 168560 103401
rect 184336 103389 184342 103401
rect 184394 103389 184400 103441
rect 645136 102057 645142 102109
rect 645194 102097 645200 102109
rect 652432 102097 652438 102109
rect 645194 102069 652438 102097
rect 645194 102057 645200 102069
rect 652432 102057 652438 102069
rect 652490 102057 652496 102109
rect 149392 100799 149398 100851
rect 149450 100839 149456 100851
rect 171280 100839 171286 100851
rect 149450 100811 171286 100839
rect 149450 100799 149456 100811
rect 171280 100799 171286 100811
rect 171338 100799 171344 100851
rect 149296 100725 149302 100777
rect 149354 100765 149360 100777
rect 184432 100765 184438 100777
rect 149354 100737 184438 100765
rect 149354 100725 149360 100737
rect 184432 100725 184438 100737
rect 184490 100725 184496 100777
rect 149680 100651 149686 100703
rect 149738 100691 149744 100703
rect 184528 100691 184534 100703
rect 149738 100663 184534 100691
rect 149738 100651 149744 100663
rect 184528 100651 184534 100663
rect 184586 100651 184592 100703
rect 156880 100577 156886 100629
rect 156938 100617 156944 100629
rect 184624 100617 184630 100629
rect 156938 100589 184630 100617
rect 156938 100577 156944 100589
rect 184624 100577 184630 100589
rect 184682 100577 184688 100629
rect 162640 100503 162646 100555
rect 162698 100543 162704 100555
rect 184336 100543 184342 100555
rect 162698 100515 184342 100543
rect 162698 100503 162704 100515
rect 184336 100503 184342 100515
rect 184394 100503 184400 100555
rect 149392 97987 149398 98039
rect 149450 98027 149456 98039
rect 184240 98027 184246 98039
rect 149450 97999 184246 98027
rect 149450 97987 149456 97999
rect 184240 97987 184246 97999
rect 184298 97987 184304 98039
rect 149488 97913 149494 97965
rect 149546 97953 149552 97965
rect 186160 97953 186166 97965
rect 149546 97925 186166 97953
rect 149546 97913 149552 97925
rect 186160 97913 186166 97925
rect 186218 97913 186224 97965
rect 647920 97913 647926 97965
rect 647978 97953 647984 97965
rect 662512 97953 662518 97965
rect 647978 97925 662518 97953
rect 647978 97913 647984 97925
rect 662512 97913 662518 97925
rect 662570 97913 662576 97965
rect 148912 97839 148918 97891
rect 148970 97879 148976 97891
rect 184432 97879 184438 97891
rect 148970 97851 184438 97879
rect 148970 97839 148976 97851
rect 184432 97839 184438 97851
rect 184490 97839 184496 97891
rect 149200 97765 149206 97817
rect 149258 97805 149264 97817
rect 184336 97805 184342 97817
rect 149258 97777 184342 97805
rect 149258 97765 149264 97777
rect 184336 97765 184342 97777
rect 184394 97765 184400 97817
rect 645424 95915 645430 95967
rect 645482 95955 645488 95967
rect 653680 95955 653686 95967
rect 645482 95927 653686 95955
rect 645482 95915 645488 95927
rect 653680 95915 653686 95927
rect 653738 95915 653744 95967
rect 149488 95101 149494 95153
rect 149546 95141 149552 95153
rect 168208 95141 168214 95153
rect 149546 95113 168214 95141
rect 149546 95101 149552 95113
rect 168208 95101 168214 95113
rect 168266 95101 168272 95153
rect 149392 95027 149398 95079
rect 149450 95067 149456 95079
rect 179920 95067 179926 95079
rect 149450 95039 179926 95067
rect 149450 95027 149456 95039
rect 179920 95027 179926 95039
rect 179978 95027 179984 95079
rect 162832 94953 162838 95005
rect 162890 94993 162896 95005
rect 184624 94993 184630 95005
rect 162890 94965 184630 94993
rect 162890 94953 162896 94965
rect 184624 94953 184630 94965
rect 184682 94953 184688 95005
rect 165712 94879 165718 94931
rect 165770 94919 165776 94931
rect 184528 94919 184534 94931
rect 165770 94891 184534 94919
rect 165770 94879 165776 94891
rect 184528 94879 184534 94891
rect 184586 94879 184592 94931
rect 168592 94805 168598 94857
rect 168650 94845 168656 94857
rect 184432 94845 184438 94857
rect 168650 94817 184438 94845
rect 168650 94805 168656 94817
rect 184432 94805 184438 94817
rect 184490 94805 184496 94857
rect 174256 94731 174262 94783
rect 174314 94771 174320 94783
rect 184336 94771 184342 94783
rect 174314 94743 184342 94771
rect 174314 94731 174320 94743
rect 184336 94731 184342 94743
rect 184394 94731 184400 94783
rect 646768 92659 646774 92711
rect 646826 92699 646832 92711
rect 663088 92699 663094 92711
rect 646826 92671 663094 92699
rect 646826 92659 646832 92671
rect 663088 92659 663094 92671
rect 663146 92659 663152 92711
rect 646384 92363 646390 92415
rect 646442 92403 646448 92415
rect 660688 92403 660694 92415
rect 646442 92375 660694 92403
rect 646442 92363 646448 92375
rect 660688 92363 660694 92375
rect 660746 92363 660752 92415
rect 646672 92289 646678 92341
rect 646730 92329 646736 92341
rect 661744 92329 661750 92341
rect 646730 92301 661750 92329
rect 646730 92289 646736 92301
rect 661744 92289 661750 92301
rect 661802 92289 661808 92341
rect 149392 92215 149398 92267
rect 149450 92255 149456 92267
rect 162448 92255 162454 92267
rect 149450 92227 162454 92255
rect 149450 92215 149456 92227
rect 162448 92215 162454 92227
rect 162506 92215 162512 92267
rect 646864 92215 646870 92267
rect 646922 92255 646928 92267
rect 659824 92255 659830 92267
rect 646922 92227 659830 92255
rect 646922 92215 646928 92227
rect 659824 92215 659830 92227
rect 659882 92215 659888 92267
rect 149488 92141 149494 92193
rect 149546 92181 149552 92193
rect 165232 92181 165238 92193
rect 149546 92153 165238 92181
rect 149546 92141 149552 92153
rect 165232 92141 165238 92153
rect 165290 92141 165296 92193
rect 646960 92141 646966 92193
rect 647018 92181 647024 92193
rect 658864 92181 658870 92193
rect 647018 92153 658870 92181
rect 647018 92141 647024 92153
rect 658864 92141 658870 92153
rect 658922 92141 658928 92193
rect 148432 92067 148438 92119
rect 148490 92107 148496 92119
rect 184432 92107 184438 92119
rect 148490 92079 184438 92107
rect 148490 92067 148496 92079
rect 184432 92067 184438 92079
rect 184490 92067 184496 92119
rect 156976 91993 156982 92045
rect 157034 92033 157040 92045
rect 184528 92033 184534 92045
rect 157034 92005 184534 92033
rect 157034 91993 157040 92005
rect 184528 91993 184534 92005
rect 184586 91993 184592 92045
rect 159856 91919 159862 91971
rect 159914 91959 159920 91971
rect 184336 91959 184342 91971
rect 159914 91931 184342 91959
rect 159914 91919 159920 91931
rect 184336 91919 184342 91931
rect 184394 91919 184400 91971
rect 177136 91845 177142 91897
rect 177194 91885 177200 91897
rect 184624 91885 184630 91897
rect 177194 91857 184630 91885
rect 177194 91845 177200 91857
rect 184624 91845 184630 91857
rect 184682 91845 184688 91897
rect 149392 90069 149398 90121
rect 149450 90109 149456 90121
rect 159760 90109 159766 90121
rect 149450 90081 159766 90109
rect 149450 90069 149456 90081
rect 159760 90069 159766 90081
rect 159818 90069 159824 90121
rect 148336 89181 148342 89233
rect 148394 89221 148400 89233
rect 184528 89221 184534 89233
rect 148394 89193 184534 89221
rect 148394 89181 148400 89193
rect 184528 89181 184534 89193
rect 184586 89181 184592 89233
rect 148624 89107 148630 89159
rect 148682 89147 148688 89159
rect 184624 89147 184630 89159
rect 148682 89119 184630 89147
rect 148682 89107 148688 89119
rect 184624 89107 184630 89119
rect 184682 89107 184688 89159
rect 151120 89033 151126 89085
rect 151178 89073 151184 89085
rect 184432 89073 184438 89085
rect 151178 89045 184438 89073
rect 151178 89033 151184 89045
rect 184432 89033 184438 89045
rect 184490 89033 184496 89085
rect 154000 88959 154006 89011
rect 154058 88999 154064 89011
rect 184336 88999 184342 89011
rect 154058 88971 184342 88999
rect 154058 88959 154064 88971
rect 184336 88959 184342 88971
rect 184394 88959 184400 89011
rect 645904 87479 645910 87531
rect 645962 87519 645968 87531
rect 650896 87519 650902 87531
rect 645962 87491 650902 87519
rect 645962 87479 645968 87491
rect 650896 87479 650902 87491
rect 650954 87479 650960 87531
rect 647920 87257 647926 87309
rect 647978 87297 647984 87309
rect 658000 87297 658006 87309
rect 647978 87269 658006 87297
rect 647978 87257 647984 87269
rect 658000 87257 658006 87269
rect 658058 87257 658064 87309
rect 647152 87035 647158 87087
rect 647210 87075 647216 87087
rect 663280 87075 663286 87087
rect 647210 87047 663286 87075
rect 647210 87035 647216 87047
rect 663280 87035 663286 87047
rect 663338 87035 663344 87087
rect 149488 86739 149494 86791
rect 149546 86779 149552 86791
rect 156496 86779 156502 86791
rect 149546 86751 156502 86779
rect 149546 86739 149552 86751
rect 156496 86739 156502 86751
rect 156554 86739 156560 86791
rect 148624 86443 148630 86495
rect 148682 86483 148688 86495
rect 154096 86483 154102 86495
rect 148682 86455 154102 86483
rect 148682 86443 148688 86455
rect 154096 86443 154102 86455
rect 154154 86443 154160 86495
rect 148240 86369 148246 86421
rect 148298 86409 148304 86421
rect 184432 86409 184438 86421
rect 148298 86381 184438 86409
rect 148298 86369 148304 86381
rect 184432 86369 184438 86381
rect 184490 86369 184496 86421
rect 148528 86295 148534 86347
rect 148586 86335 148592 86347
rect 184528 86335 184534 86347
rect 148586 86307 184534 86335
rect 148586 86295 148592 86307
rect 184528 86295 184534 86307
rect 184586 86295 184592 86347
rect 148720 86221 148726 86273
rect 148778 86261 148784 86273
rect 184336 86261 184342 86273
rect 148778 86233 184342 86261
rect 148778 86221 148784 86233
rect 184336 86221 184342 86233
rect 184394 86221 184400 86273
rect 640720 84963 640726 85015
rect 640778 85003 640784 85015
rect 643600 85003 643606 85015
rect 640778 84975 643606 85003
rect 640778 84963 640784 84975
rect 643600 84963 643606 84975
rect 643658 84963 643664 85015
rect 645712 84149 645718 84201
rect 645770 84189 645776 84201
rect 657040 84189 657046 84201
rect 645770 84161 657046 84189
rect 645770 84149 645776 84161
rect 657040 84149 657046 84161
rect 657098 84149 657104 84201
rect 146992 83557 146998 83609
rect 147050 83597 147056 83609
rect 151120 83597 151126 83609
rect 147050 83569 151126 83597
rect 147050 83557 147056 83569
rect 151120 83557 151126 83569
rect 151178 83557 151184 83609
rect 646768 83557 646774 83609
rect 646826 83597 646832 83609
rect 653680 83597 653686 83609
rect 646826 83569 653686 83597
rect 646826 83557 646832 83569
rect 653680 83557 653686 83569
rect 653738 83557 653744 83609
rect 168208 83483 168214 83535
rect 168266 83523 168272 83535
rect 184432 83523 184438 83535
rect 168266 83495 184438 83523
rect 168266 83483 168272 83495
rect 184432 83483 184438 83495
rect 184490 83483 184496 83535
rect 171280 83409 171286 83461
rect 171338 83449 171344 83461
rect 184336 83449 184342 83461
rect 171338 83421 184342 83449
rect 171338 83409 171344 83421
rect 184336 83409 184342 83421
rect 184394 83409 184400 83461
rect 647920 81855 647926 81907
rect 647978 81895 647984 81907
rect 663280 81895 663286 81907
rect 647978 81867 663286 81895
rect 647978 81855 647984 81867
rect 663280 81855 663286 81867
rect 663338 81855 663344 81907
rect 647824 81781 647830 81833
rect 647882 81821 647888 81833
rect 663376 81821 663382 81833
rect 647882 81793 663382 81821
rect 647882 81781 647888 81793
rect 663376 81781 663382 81793
rect 663434 81781 663440 81833
rect 657040 81633 657046 81685
rect 657098 81673 657104 81685
rect 658576 81673 658582 81685
rect 657098 81645 658582 81673
rect 657098 81633 657104 81645
rect 658576 81633 658582 81645
rect 658634 81633 658640 81685
rect 647728 81559 647734 81611
rect 647786 81599 647792 81611
rect 662416 81599 662422 81611
rect 647786 81571 662422 81599
rect 647786 81559 647792 81571
rect 662416 81559 662422 81571
rect 662474 81559 662480 81611
rect 647920 80745 647926 80797
rect 647978 80785 647984 80797
rect 662512 80785 662518 80797
rect 647978 80757 662518 80785
rect 647978 80745 647984 80757
rect 662512 80745 662518 80757
rect 662570 80745 662576 80797
rect 149296 80597 149302 80649
rect 149354 80637 149360 80649
rect 184432 80637 184438 80649
rect 149354 80609 184438 80637
rect 149354 80597 149360 80609
rect 184432 80597 184438 80609
rect 184490 80597 184496 80649
rect 162448 80523 162454 80575
rect 162506 80563 162512 80575
rect 184528 80563 184534 80575
rect 162506 80535 184534 80563
rect 162506 80523 162512 80535
rect 184528 80523 184534 80535
rect 184586 80523 184592 80575
rect 165232 80449 165238 80501
rect 165290 80489 165296 80501
rect 184336 80489 184342 80501
rect 165290 80461 184342 80489
rect 165290 80449 165296 80461
rect 184336 80449 184342 80461
rect 184394 80449 184400 80501
rect 179920 80375 179926 80427
rect 179978 80415 179984 80427
rect 184624 80415 184630 80427
rect 179978 80387 184630 80415
rect 179978 80375 179984 80387
rect 184624 80375 184630 80387
rect 184682 80375 184688 80427
rect 149392 77711 149398 77763
rect 149450 77751 149456 77763
rect 184624 77751 184630 77763
rect 149450 77723 184630 77751
rect 149450 77711 149456 77723
rect 184624 77711 184630 77723
rect 184682 77711 184688 77763
rect 647056 77711 647062 77763
rect 647114 77751 647120 77763
rect 658288 77751 658294 77763
rect 647114 77723 658294 77751
rect 647114 77711 647120 77723
rect 658288 77711 658294 77723
rect 658346 77711 658352 77763
rect 149680 77637 149686 77689
rect 149738 77677 149744 77689
rect 184432 77677 184438 77689
rect 149738 77649 184438 77677
rect 149738 77637 149744 77649
rect 184432 77637 184438 77649
rect 184490 77637 184496 77689
rect 646480 77637 646486 77689
rect 646538 77677 646544 77689
rect 659536 77677 659542 77689
rect 646538 77649 659542 77677
rect 646538 77637 646544 77649
rect 659536 77637 659542 77649
rect 659594 77637 659600 77689
rect 156496 77563 156502 77615
rect 156554 77603 156560 77615
rect 184528 77603 184534 77615
rect 156554 77575 184534 77603
rect 156554 77563 156560 77575
rect 184528 77563 184534 77575
rect 184586 77563 184592 77615
rect 646576 77563 646582 77615
rect 646634 77603 646640 77615
rect 661744 77603 661750 77615
rect 646634 77575 661750 77603
rect 646634 77563 646640 77575
rect 661744 77563 661750 77575
rect 661802 77563 661808 77615
rect 159760 77489 159766 77541
rect 159818 77529 159824 77541
rect 184336 77529 184342 77541
rect 159818 77501 184342 77529
rect 159818 77489 159824 77501
rect 184336 77489 184342 77501
rect 184394 77489 184400 77541
rect 647920 77489 647926 77541
rect 647978 77529 647984 77541
rect 656944 77529 656950 77541
rect 647978 77501 656950 77529
rect 647978 77489 647984 77501
rect 656944 77489 656950 77501
rect 657002 77489 657008 77541
rect 646288 75639 646294 75691
rect 646346 75679 646352 75691
rect 657520 75679 657526 75691
rect 646346 75651 657526 75679
rect 646346 75639 646352 75651
rect 657520 75639 657526 75651
rect 657578 75639 657584 75691
rect 647152 74899 647158 74951
rect 647210 74939 647216 74951
rect 660112 74939 660118 74951
rect 647210 74911 660118 74939
rect 647210 74899 647216 74911
rect 660112 74899 660118 74911
rect 660170 74899 660176 74951
rect 148432 74825 148438 74877
rect 148490 74865 148496 74877
rect 184528 74865 184534 74877
rect 148490 74837 184534 74865
rect 148490 74825 148496 74837
rect 184528 74825 184534 74837
rect 184586 74825 184592 74877
rect 149200 74751 149206 74803
rect 149258 74791 149264 74803
rect 184624 74791 184630 74803
rect 149258 74763 184630 74791
rect 149258 74751 149264 74763
rect 184624 74751 184630 74763
rect 184682 74751 184688 74803
rect 151120 74677 151126 74729
rect 151178 74717 151184 74729
rect 184432 74717 184438 74729
rect 151178 74689 184438 74717
rect 151178 74677 151184 74689
rect 184432 74677 184438 74689
rect 184490 74677 184496 74729
rect 154096 74603 154102 74655
rect 154154 74643 154160 74655
rect 184336 74643 184342 74655
rect 154154 74615 184342 74643
rect 154154 74603 154160 74615
rect 184336 74603 184342 74615
rect 184394 74603 184400 74655
rect 149200 74011 149206 74063
rect 149258 74051 149264 74063
rect 149392 74051 149398 74063
rect 149258 74023 149398 74051
rect 149258 74011 149264 74023
rect 149392 74011 149398 74023
rect 149450 74011 149456 74063
rect 647920 72087 647926 72139
rect 647978 72127 647984 72139
rect 660688 72127 660694 72139
rect 647978 72099 660694 72127
rect 647978 72087 647984 72099
rect 660688 72087 660694 72099
rect 660746 72087 660752 72139
rect 148336 71939 148342 71991
rect 148394 71979 148400 71991
rect 184336 71979 184342 71991
rect 148394 71951 184342 71979
rect 148394 71939 148400 71951
rect 184336 71939 184342 71951
rect 184394 71939 184400 71991
rect 149392 71865 149398 71917
rect 149450 71905 149456 71917
rect 184432 71905 184438 71917
rect 149450 71877 184438 71905
rect 149450 71865 149456 71877
rect 184432 71865 184438 71877
rect 184490 71865 184496 71917
rect 149584 71791 149590 71843
rect 149642 71831 149648 71843
rect 184528 71831 184534 71843
rect 149642 71803 184534 71831
rect 149642 71791 149648 71803
rect 184528 71791 184534 71803
rect 184586 71791 184592 71843
rect 647920 69571 647926 69623
rect 647978 69611 647984 69623
rect 661168 69611 661174 69623
rect 647978 69583 661174 69611
rect 647978 69571 647984 69583
rect 661168 69571 661174 69583
rect 661226 69571 661232 69623
rect 149584 69053 149590 69105
rect 149642 69093 149648 69105
rect 184528 69093 184534 69105
rect 149642 69065 184534 69093
rect 149642 69053 149648 69065
rect 184528 69053 184534 69065
rect 184586 69053 184592 69105
rect 148816 68979 148822 69031
rect 148874 69019 148880 69031
rect 184336 69019 184342 69031
rect 148874 68991 184342 69019
rect 148874 68979 148880 68991
rect 184336 68979 184342 68991
rect 184394 68979 184400 69031
rect 149296 68905 149302 68957
rect 149354 68945 149360 68957
rect 184432 68945 184438 68957
rect 149354 68917 184438 68945
rect 149354 68905 149360 68917
rect 184432 68905 184438 68917
rect 184490 68905 184496 68957
rect 149200 68831 149206 68883
rect 149258 68871 149264 68883
rect 184336 68871 184342 68883
rect 149258 68843 184342 68871
rect 149258 68831 149264 68843
rect 184336 68831 184342 68843
rect 184394 68831 184400 68883
rect 149104 66167 149110 66219
rect 149162 66207 149168 66219
rect 184528 66207 184534 66219
rect 149162 66179 184534 66207
rect 149162 66167 149168 66179
rect 184528 66167 184534 66179
rect 184586 66167 184592 66219
rect 646000 66167 646006 66219
rect 646058 66207 646064 66219
rect 652336 66207 652342 66219
rect 646058 66179 652342 66207
rect 646058 66167 646064 66179
rect 652336 66167 652342 66179
rect 652394 66167 652400 66219
rect 149680 66093 149686 66145
rect 149738 66133 149744 66145
rect 184336 66133 184342 66145
rect 149738 66105 184342 66133
rect 149738 66093 149744 66105
rect 184336 66093 184342 66105
rect 184394 66093 184400 66145
rect 149488 66019 149494 66071
rect 149546 66059 149552 66071
rect 184432 66059 184438 66071
rect 149546 66031 184438 66059
rect 149546 66019 149552 66031
rect 184432 66019 184438 66031
rect 184490 66019 184496 66071
rect 149392 65945 149398 65997
rect 149450 65985 149456 65997
rect 184336 65985 184342 65997
rect 149450 65957 184342 65985
rect 149450 65945 149456 65957
rect 184336 65945 184342 65957
rect 184394 65945 184400 65997
rect 647920 63429 647926 63481
rect 647978 63469 647984 63481
rect 663184 63469 663190 63481
rect 647978 63441 663190 63469
rect 647978 63429 647984 63441
rect 663184 63429 663190 63441
rect 663242 63429 663248 63481
rect 149296 63281 149302 63333
rect 149354 63321 149360 63333
rect 184432 63321 184438 63333
rect 149354 63293 184438 63321
rect 149354 63281 149360 63293
rect 184432 63281 184438 63293
rect 184490 63281 184496 63333
rect 149392 63207 149398 63259
rect 149450 63247 149456 63259
rect 184624 63247 184630 63259
rect 149450 63219 184630 63247
rect 149450 63207 149456 63219
rect 184624 63207 184630 63219
rect 184682 63207 184688 63259
rect 149200 63133 149206 63185
rect 149258 63173 149264 63185
rect 184336 63173 184342 63185
rect 149258 63145 184342 63173
rect 149258 63133 149264 63145
rect 184336 63133 184342 63145
rect 184394 63133 184400 63185
rect 149488 63059 149494 63111
rect 149546 63099 149552 63111
rect 184528 63099 184534 63111
rect 149546 63071 184534 63099
rect 149546 63059 149552 63071
rect 184528 63059 184534 63071
rect 184586 63059 184592 63111
rect 647920 60987 647926 61039
rect 647978 61027 647984 61039
rect 663472 61027 663478 61039
rect 647978 60999 663478 61027
rect 647978 60987 647984 60999
rect 663472 60987 663478 60999
rect 663530 60987 663536 61039
rect 149392 60395 149398 60447
rect 149450 60435 149456 60447
rect 184432 60435 184438 60447
rect 149450 60407 184438 60435
rect 149450 60395 149456 60407
rect 184432 60395 184438 60407
rect 184490 60395 184496 60447
rect 149584 60321 149590 60373
rect 149642 60361 149648 60373
rect 184336 60361 184342 60373
rect 149642 60333 184342 60361
rect 149642 60321 149648 60333
rect 184336 60321 184342 60333
rect 184394 60321 184400 60373
rect 149296 60247 149302 60299
rect 149354 60287 149360 60299
rect 184528 60287 184534 60299
rect 149354 60259 184534 60287
rect 149354 60247 149360 60259
rect 184528 60247 184534 60259
rect 184586 60247 184592 60299
rect 646000 59063 646006 59115
rect 646058 59103 646064 59115
rect 652240 59103 652246 59115
rect 646058 59075 652246 59103
rect 646058 59063 646064 59075
rect 652240 59063 652246 59075
rect 652298 59063 652304 59115
rect 149392 58989 149398 59041
rect 149450 59029 149456 59041
rect 184336 59029 184342 59041
rect 149450 59001 184342 59029
rect 149450 58989 149456 59001
rect 184336 58989 184342 59001
rect 184394 58989 184400 59041
rect 149392 57509 149398 57561
rect 149450 57549 149456 57561
rect 184336 57549 184342 57561
rect 149450 57521 184342 57549
rect 149450 57509 149456 57521
rect 184336 57509 184342 57521
rect 184394 57509 184400 57561
rect 149488 56177 149494 56229
rect 149546 56217 149552 56229
rect 184336 56217 184342 56229
rect 149546 56189 184342 56217
rect 149546 56177 149552 56189
rect 184336 56177 184342 56189
rect 184394 56177 184400 56229
rect 149392 56103 149398 56155
rect 149450 56143 149456 56155
rect 184432 56143 184438 56155
rect 149450 56115 184438 56143
rect 149450 56103 149456 56115
rect 184432 56103 184438 56115
rect 184490 56103 184496 56155
rect 149680 54623 149686 54675
rect 149738 54663 149744 54675
rect 184336 54663 184342 54675
rect 149738 54635 184342 54663
rect 149738 54623 149744 54635
rect 184336 54623 184342 54635
rect 184394 54623 184400 54675
rect 149392 53217 149398 53269
rect 149450 53257 149456 53269
rect 184336 53257 184342 53269
rect 149450 53229 184342 53257
rect 149450 53217 149456 53229
rect 184336 53217 184342 53229
rect 184394 53217 184400 53269
rect 643600 51885 643606 51937
rect 643658 51925 643664 51937
rect 654064 51925 654070 51937
rect 643658 51897 654070 51925
rect 643658 51885 643664 51897
rect 654064 51885 654070 51897
rect 654122 51885 654128 51937
rect 311152 48037 311158 48089
rect 311210 48077 311216 48089
rect 354832 48077 354838 48089
rect 311210 48049 354838 48077
rect 311210 48037 311216 48049
rect 354832 48037 354838 48049
rect 354890 48037 354896 48089
rect 311056 47963 311062 48015
rect 311114 48003 311120 48015
rect 371920 48003 371926 48015
rect 311114 47975 371926 48003
rect 311114 47963 311120 47975
rect 371920 47963 371926 47975
rect 371978 47963 371984 48015
rect 405520 47963 405526 48015
rect 405578 48003 405584 48015
rect 441328 48003 441334 48015
rect 405578 47975 441334 48003
rect 405578 47963 405584 47975
rect 441328 47963 441334 47975
rect 441386 47963 441392 48015
rect 460336 47963 460342 48015
rect 460394 48003 460400 48015
rect 510352 48003 510358 48015
rect 460394 47975 510358 48003
rect 460394 47963 460400 47975
rect 510352 47963 510358 47975
rect 510410 47963 510416 48015
rect 320176 47889 320182 47941
rect 320234 47929 320240 47941
rect 529264 47929 529270 47941
rect 320234 47901 529270 47929
rect 320234 47889 320240 47901
rect 529264 47889 529270 47901
rect 529322 47889 529328 47941
rect 302896 47815 302902 47867
rect 302954 47855 302960 47867
rect 521104 47855 521110 47867
rect 302954 47827 521110 47855
rect 302954 47815 302960 47827
rect 521104 47815 521110 47827
rect 521162 47815 521168 47867
rect 285808 47741 285814 47793
rect 285866 47781 285872 47793
rect 515536 47781 515542 47793
rect 285866 47753 515542 47781
rect 285866 47741 285872 47753
rect 515536 47741 515542 47753
rect 515594 47741 515600 47793
rect 268528 47667 268534 47719
rect 268586 47707 268592 47719
rect 503920 47707 503926 47719
rect 268586 47679 503926 47707
rect 268586 47667 268592 47679
rect 503920 47667 503926 47679
rect 503978 47667 503984 47719
rect 233680 47593 233686 47645
rect 233738 47633 233744 47645
rect 233738 47605 468062 47633
rect 233738 47593 233744 47605
rect 250960 47519 250966 47571
rect 251018 47559 251024 47571
rect 468034 47559 468062 47605
rect 475216 47593 475222 47645
rect 475274 47633 475280 47645
rect 492976 47633 492982 47645
rect 475274 47605 492982 47633
rect 475274 47593 475280 47605
rect 492976 47593 492982 47605
rect 493034 47593 493040 47645
rect 475600 47559 475606 47571
rect 251018 47531 457934 47559
rect 468034 47531 475606 47559
rect 251018 47519 251024 47531
rect 457906 47411 457934 47531
rect 475600 47519 475606 47531
rect 475658 47519 475664 47571
rect 521200 47559 521206 47571
rect 478066 47531 521206 47559
rect 478066 47411 478094 47531
rect 521200 47519 521206 47531
rect 521258 47519 521264 47571
rect 457906 47383 478094 47411
rect 145360 47075 145366 47127
rect 145418 47115 145424 47127
rect 199120 47115 199126 47127
rect 145418 47087 199126 47115
rect 145418 47075 145424 47087
rect 199120 47075 199126 47087
rect 199178 47075 199184 47127
rect 334096 46927 334102 46979
rect 334154 46967 334160 46979
rect 337456 46967 337462 46979
rect 334154 46939 337462 46967
rect 334154 46927 334160 46939
rect 337456 46927 337462 46939
rect 337514 46927 337520 46979
rect 636496 46705 636502 46757
rect 636554 46745 636560 46757
rect 643600 46745 643606 46757
rect 636554 46717 643606 46745
rect 636554 46705 636560 46717
rect 643600 46705 643606 46717
rect 643658 46705 643664 46757
rect 403216 46335 403222 46387
rect 403274 46375 403280 46387
rect 406768 46375 406774 46387
rect 403274 46347 406774 46375
rect 403274 46335 403280 46347
rect 406768 46335 406774 46347
rect 406826 46335 406832 46387
rect 207376 46113 207382 46165
rect 207434 46153 207440 46165
rect 216400 46153 216406 46165
rect 207434 46125 216406 46153
rect 207434 46113 207440 46125
rect 216400 46113 216406 46125
rect 216458 46113 216464 46165
rect 522832 46113 522838 46165
rect 522890 46153 522896 46165
rect 527920 46153 527926 46165
rect 522890 46125 527926 46153
rect 522890 46113 522896 46125
rect 527920 46113 527926 46125
rect 527978 46113 527984 46165
rect 521104 44781 521110 44833
rect 521162 44821 521168 44833
rect 525904 44821 525910 44833
rect 521162 44793 525910 44821
rect 521162 44781 521168 44793
rect 525904 44781 525910 44793
rect 525962 44781 525968 44833
rect 515536 44633 515542 44685
rect 515594 44673 515600 44685
rect 524944 44673 524950 44685
rect 515594 44645 524950 44673
rect 515594 44633 515600 44645
rect 524944 44633 524950 44645
rect 525002 44633 525008 44685
rect 541456 43301 541462 43353
rect 541514 43341 541520 43353
rect 545200 43341 545206 43353
rect 541514 43313 545206 43341
rect 541514 43301 541520 43313
rect 545200 43301 545206 43313
rect 545258 43301 545264 43353
rect 503920 43227 503926 43279
rect 503978 43267 503984 43279
rect 503978 43239 520382 43267
rect 503978 43227 503984 43239
rect 520354 43205 520382 43239
rect 520336 43153 520342 43205
rect 520394 43153 520400 43205
rect 506800 41969 506806 42021
rect 506858 42009 506864 42021
rect 506858 41981 518414 42009
rect 506858 41969 506864 41981
rect 307216 41895 307222 41947
rect 307274 41935 307280 41947
rect 311056 41935 311062 41947
rect 307274 41907 311062 41935
rect 307274 41895 307280 41907
rect 311056 41895 311062 41907
rect 311114 41895 311120 41947
rect 394576 41895 394582 41947
rect 394634 41935 394640 41947
rect 424048 41935 424054 41947
rect 394634 41907 424054 41935
rect 394634 41895 394640 41907
rect 424048 41895 424054 41907
rect 424106 41895 424112 41947
rect 449296 41895 449302 41947
rect 449354 41935 449360 41947
rect 475216 41935 475222 41947
rect 449354 41907 475222 41935
rect 449354 41895 449360 41907
rect 475216 41895 475222 41907
rect 475274 41895 475280 41947
rect 514000 41895 514006 41947
rect 514058 41935 514064 41947
rect 514864 41935 514870 41947
rect 514058 41907 514870 41935
rect 514058 41895 514064 41907
rect 514864 41895 514870 41907
rect 514922 41895 514928 41947
rect 518386 41935 518414 41981
rect 562480 41935 562486 41947
rect 518386 41907 562486 41935
rect 562480 41895 562486 41907
rect 562538 41895 562544 41947
rect 145072 41821 145078 41873
rect 145130 41861 145136 41873
rect 636496 41861 636502 41873
rect 145130 41833 636502 41861
rect 145130 41821 145136 41833
rect 636496 41821 636502 41833
rect 636554 41821 636560 41873
rect 187600 41747 187606 41799
rect 187658 41747 187664 41799
rect 194320 41747 194326 41799
rect 194378 41787 194384 41799
rect 640720 41787 640726 41799
rect 194378 41759 640726 41787
rect 194378 41747 194384 41759
rect 640720 41747 640726 41759
rect 640778 41747 640784 41799
rect 187618 41491 187646 41747
rect 207376 41491 207382 41503
rect 187618 41463 207382 41491
rect 207376 41451 207382 41463
rect 207434 41451 207440 41503
rect 365872 37381 365878 37433
rect 365930 37421 365936 37433
rect 394576 37421 394582 37433
rect 365930 37393 394582 37421
rect 365930 37381 365936 37393
rect 394576 37381 394582 37393
rect 394634 37381 394640 37433
rect 420688 37381 420694 37433
rect 420746 37421 420752 37433
rect 449296 37421 449302 37433
rect 420746 37393 449302 37421
rect 420746 37381 420752 37393
rect 449296 37381 449302 37393
rect 449354 37381 449360 37433
rect 475600 37381 475606 37433
rect 475658 37421 475664 37433
rect 514000 37421 514006 37433
rect 475658 37393 514006 37421
rect 475658 37381 475664 37393
rect 514000 37381 514006 37393
rect 514058 37381 514064 37433
rect 475504 37307 475510 37359
rect 475562 37347 475568 37359
rect 506800 37347 506806 37359
rect 475562 37319 506806 37347
rect 475562 37307 475568 37319
rect 506800 37307 506806 37319
rect 506858 37307 506864 37359
<< via1 >>
rect 483670 1005153 483722 1005205
rect 529846 1005153 529898 1005205
rect 535030 1005153 535082 1005205
rect 561622 1005153 561674 1005205
rect 636886 1005153 636938 1005205
rect 649366 1005153 649418 1005205
rect 529846 999381 529898 999433
rect 561622 999381 561674 999433
rect 571894 999381 571946 999433
rect 532822 999307 532874 999359
rect 655414 892969 655466 893021
rect 676246 892969 676298 893021
rect 655222 892895 655274 892947
rect 676150 892895 676202 892947
rect 655126 892821 655178 892873
rect 676054 892821 676106 892873
rect 673846 892377 673898 892429
rect 676054 892377 676106 892429
rect 670966 891415 671018 891467
rect 676054 891415 676106 891467
rect 670870 890379 670922 890431
rect 676054 890379 676106 890431
rect 674038 887863 674090 887915
rect 676246 887863 676298 887915
rect 674230 887123 674282 887175
rect 676054 887123 676106 887175
rect 674422 887049 674474 887101
rect 676246 887049 676298 887101
rect 674134 885051 674186 885103
rect 676054 885051 676106 885103
rect 674326 884237 674378 884289
rect 676054 884237 676106 884289
rect 674902 884163 674954 884215
rect 676246 884163 676298 884215
rect 675286 883201 675338 883253
rect 679990 883201 680042 883253
rect 674518 883053 674570 883105
rect 680182 883053 680234 883105
rect 674998 882831 675050 882883
rect 679702 882831 679754 882883
rect 674710 881499 674762 881551
rect 675958 881499 676010 881551
rect 649462 881425 649514 881477
rect 679702 881425 679754 881477
rect 655318 881351 655370 881403
rect 675478 881351 675530 881403
rect 674806 881277 674858 881329
rect 676054 881277 676106 881329
rect 674614 881203 674666 881255
rect 680086 881203 680138 881255
rect 675190 880093 675242 880145
rect 679798 880093 679850 880145
rect 679894 878465 679946 878517
rect 675094 877947 675146 877999
rect 674998 877207 675050 877259
rect 675478 877207 675530 877259
rect 674614 876689 674666 876741
rect 675286 876689 675338 876741
rect 674518 876615 674570 876667
rect 675382 876615 675434 876667
rect 674230 876393 674282 876445
rect 674518 876393 674570 876445
rect 674038 876245 674090 876297
rect 674230 876245 674282 876297
rect 674806 872989 674858 873041
rect 675286 872989 675338 873041
rect 674710 872915 674762 872967
rect 675190 872915 675242 872967
rect 654166 872619 654218 872671
rect 675094 872619 675146 872671
rect 674614 870547 674666 870599
rect 675478 870547 675530 870599
rect 674326 869733 674378 869785
rect 675286 869733 675338 869785
rect 674518 869659 674570 869711
rect 674998 869659 675050 869711
rect 674134 867365 674186 867417
rect 675478 867365 675530 867417
rect 674230 865737 674282 865789
rect 675190 865737 675242 865789
rect 653782 863961 653834 864013
rect 675094 863961 675146 864013
rect 41782 817933 41834 817985
rect 47446 817933 47498 817985
rect 41782 817267 41834 817319
rect 44854 817267 44906 817319
rect 41590 816527 41642 816579
rect 44950 816527 45002 816579
rect 41782 815787 41834 815839
rect 43222 815787 43274 815839
rect 41782 814825 41834 814877
rect 44662 814825 44714 814877
rect 41590 813567 41642 813619
rect 44758 813567 44810 813619
rect 41590 812383 41642 812435
rect 42646 812383 42698 812435
rect 41782 809423 41834 809475
rect 43030 809423 43082 809475
rect 41590 807055 41642 807107
rect 42934 807055 42986 807107
rect 41974 806981 42026 807033
rect 43126 806981 43178 807033
rect 41590 806611 41642 806663
rect 42646 806611 42698 806663
rect 41782 806389 41834 806441
rect 42742 806389 42794 806441
rect 41590 805131 41642 805183
rect 44566 805131 44618 805183
rect 42358 800691 42410 800743
rect 57718 800691 57770 800743
rect 42454 800617 42506 800669
rect 57622 800617 57674 800669
rect 41974 800173 42026 800225
rect 41974 799951 42026 800003
rect 42358 796843 42410 796895
rect 42742 796843 42794 796895
rect 42550 795067 42602 795119
rect 42550 794845 42602 794897
rect 42454 794401 42506 794453
rect 42838 794401 42890 794453
rect 42070 794253 42122 794305
rect 42934 794253 42986 794305
rect 42454 793143 42506 793195
rect 43030 793143 43082 793195
rect 655126 792033 655178 792085
rect 675382 792033 675434 792085
rect 42166 790627 42218 790679
rect 43126 790627 43178 790679
rect 42166 790109 42218 790161
rect 42838 790109 42890 790161
rect 42166 789443 42218 789495
rect 42742 789443 42794 789495
rect 42454 789147 42506 789199
rect 58198 789147 58250 789199
rect 44950 789073 45002 789125
rect 58390 789073 58442 789125
rect 42166 788703 42218 788755
rect 42646 788703 42698 788755
rect 42166 787001 42218 787053
rect 42550 787001 42602 787053
rect 42166 786409 42218 786461
rect 42358 786409 42410 786461
rect 44854 785521 44906 785573
rect 59158 785521 59210 785573
rect 47446 785373 47498 785425
rect 59638 785373 59690 785425
rect 656566 783375 656618 783427
rect 675190 783375 675242 783427
rect 654358 780489 654410 780541
rect 675094 780489 675146 780541
rect 674902 778565 674954 778617
rect 675286 778565 675338 778617
rect 674806 777307 674858 777359
rect 675478 777307 675530 777359
rect 41782 774643 41834 774695
rect 47446 774643 47498 774695
rect 674326 774273 674378 774325
rect 675094 774273 675146 774325
rect 41590 773903 41642 773955
rect 44950 773903 45002 773955
rect 41782 773459 41834 773511
rect 45046 773459 45098 773511
rect 41590 773385 41642 773437
rect 43222 773385 43274 773437
rect 41782 772571 41834 772623
rect 43222 772571 43274 772623
rect 43126 772127 43178 772179
rect 62038 772127 62090 772179
rect 41590 771905 41642 771957
rect 61846 771905 61898 771957
rect 41782 767539 41834 767591
rect 42742 767539 42794 767591
rect 41590 767095 41642 767147
rect 42646 767095 42698 767147
rect 674422 767095 674474 767147
rect 675094 767095 675146 767147
rect 41782 766577 41834 766629
rect 42550 766577 42602 766629
rect 41590 765393 41642 765445
rect 42838 765393 42890 765445
rect 41782 764727 41834 764779
rect 42934 764727 42986 764779
rect 41590 763395 41642 763447
rect 43030 763395 43082 763447
rect 42070 763247 42122 763299
rect 43126 763247 43178 763299
rect 41590 761915 41642 761967
rect 44854 761915 44906 761967
rect 42454 757623 42506 757675
rect 43318 757623 43370 757675
rect 42454 757475 42506 757527
rect 58678 757475 58730 757527
rect 43126 757253 43178 757305
rect 43510 757253 43562 757305
rect 42646 757179 42698 757231
rect 43414 757179 43466 757231
rect 42550 757105 42602 757157
rect 43126 757105 43178 757157
rect 41878 757031 41930 757083
rect 42646 757031 42698 757083
rect 41782 756957 41834 757009
rect 42550 756957 42602 757009
rect 42262 756883 42314 756935
rect 42358 756661 42410 756713
rect 42358 753627 42410 753679
rect 42838 753627 42890 753679
rect 42838 753479 42890 753531
rect 43318 753479 43370 753531
rect 42358 751777 42410 751829
rect 43030 751777 43082 751829
rect 42454 751703 42506 751755
rect 43318 751703 43370 751755
rect 43030 751629 43082 751681
rect 43414 751629 43466 751681
rect 42454 751555 42506 751607
rect 42934 751555 42986 751607
rect 42262 750593 42314 750645
rect 43510 750593 43562 750645
rect 42070 749927 42122 749979
rect 42742 749927 42794 749979
rect 655702 748817 655754 748869
rect 675382 748817 675434 748869
rect 42070 746079 42122 746131
rect 43126 746079 43178 746131
rect 42646 745931 42698 745983
rect 54646 745931 54698 745983
rect 54742 745931 54794 745983
rect 57622 745931 57674 745983
rect 42166 745487 42218 745539
rect 43030 745487 43082 745539
rect 45046 745413 45098 745465
rect 58102 745413 58154 745465
rect 43318 744969 43370 745021
rect 58582 744969 58634 745021
rect 42166 743785 42218 743837
rect 42838 743785 42890 743837
rect 47446 742971 47498 743023
rect 59638 742971 59690 743023
rect 44950 742897 45002 742949
rect 59734 742897 59786 742949
rect 674710 742749 674762 742801
rect 675382 742749 675434 742801
rect 673654 737865 673706 737917
rect 675382 737865 675434 737917
rect 654070 737421 654122 737473
rect 674998 737421 675050 737473
rect 654166 737347 654218 737399
rect 675094 737347 675146 737399
rect 675190 735719 675242 735771
rect 675286 735497 675338 735549
rect 675094 733869 675146 733921
rect 675382 733869 675434 733921
rect 673462 733721 673514 733773
rect 675478 733721 675530 733773
rect 674230 732315 674282 732367
rect 675478 732315 675530 732367
rect 674998 732019 675050 732071
rect 675382 732019 675434 732071
rect 41782 731427 41834 731479
rect 47542 731427 47594 731479
rect 41590 730687 41642 730739
rect 44950 730687 45002 730739
rect 674710 730465 674762 730517
rect 675478 730465 675530 730517
rect 41782 730317 41834 730369
rect 45046 730317 45098 730369
rect 41590 730169 41642 730221
rect 43222 730169 43274 730221
rect 41782 729355 41834 729407
rect 43510 729355 43562 729407
rect 41782 728763 41834 728815
rect 43318 728763 43370 728815
rect 40438 728689 40490 728741
rect 62230 728689 62282 728741
rect 42262 728615 42314 728667
rect 62422 728615 62474 728667
rect 674614 728615 674666 728667
rect 675382 728615 675434 728667
rect 41782 727875 41834 727927
rect 43414 727875 43466 727927
rect 41782 726543 41834 726595
rect 42934 726543 42986 726595
rect 41782 726395 41834 726447
rect 42838 726395 42890 726447
rect 41782 722991 41834 723043
rect 43030 722991 43082 723043
rect 673846 722917 673898 722969
rect 679702 722917 679754 722969
rect 41590 720919 41642 720971
rect 42550 720919 42602 720971
rect 41782 720549 41834 720601
rect 43126 720549 43178 720601
rect 41590 720327 41642 720379
rect 42646 720327 42698 720379
rect 41782 720179 41834 720231
rect 42742 720179 42794 720231
rect 41590 718699 41642 718751
rect 47446 718699 47498 718751
rect 655606 714703 655658 714755
rect 676246 714703 676298 714755
rect 655414 714555 655466 714607
rect 676150 714555 676202 714607
rect 655222 714407 655274 714459
rect 676342 714407 676394 714459
rect 42358 714259 42410 714311
rect 59638 714259 59690 714311
rect 41974 713889 42026 713941
rect 43222 713889 43274 713941
rect 41782 713815 41834 713867
rect 41878 713815 41930 713867
rect 43606 713815 43658 713867
rect 669718 713075 669770 713127
rect 670966 713075 671018 713127
rect 676054 713075 676106 713127
rect 42262 712853 42314 712905
rect 42838 712853 42890 712905
rect 42838 712705 42890 712757
rect 670678 712631 670730 712683
rect 676054 712631 676106 712683
rect 669526 711891 669578 711943
rect 670870 711891 670922 711943
rect 676246 711891 676298 711943
rect 42166 711669 42218 711721
rect 42934 711669 42986 711721
rect 43222 711595 43274 711647
rect 42262 711447 42314 711499
rect 42358 711373 42410 711425
rect 43030 711373 43082 711425
rect 670582 711521 670634 711573
rect 676054 711521 676106 711573
rect 43318 711373 43370 711425
rect 43510 711373 43562 711425
rect 42166 711299 42218 711351
rect 42934 711299 42986 711351
rect 674326 711299 674378 711351
rect 676054 711299 676106 711351
rect 42838 711225 42890 711277
rect 42262 711077 42314 711129
rect 42166 710855 42218 710907
rect 42454 710855 42506 710907
rect 674422 710485 674474 710537
rect 676054 710485 676106 710537
rect 42166 709893 42218 709945
rect 42550 709893 42602 709945
rect 42070 708487 42122 708539
rect 43510 708487 43562 708539
rect 675286 708413 675338 708465
rect 676054 708413 676106 708465
rect 42070 708339 42122 708391
rect 42742 708339 42794 708391
rect 674902 708339 674954 708391
rect 676246 708339 676298 708391
rect 42262 708191 42314 708243
rect 42742 708191 42794 708243
rect 42454 708043 42506 708095
rect 43126 708043 43178 708095
rect 674806 708043 674858 708095
rect 676054 708043 676106 708095
rect 43126 707895 43178 707947
rect 43606 707895 43658 707947
rect 42454 707377 42506 707429
rect 42646 707377 42698 707429
rect 42454 706711 42506 706763
rect 43030 706711 43082 706763
rect 42166 704269 42218 704321
rect 43126 704269 43178 704321
rect 42070 703677 42122 703729
rect 42934 703677 42986 703729
rect 42262 702937 42314 702989
rect 42646 702937 42698 702989
rect 42070 702863 42122 702915
rect 42742 702863 42794 702915
rect 654742 702789 654794 702841
rect 675382 702789 675434 702841
rect 42454 702715 42506 702767
rect 58870 702715 58922 702767
rect 649462 702715 649514 702767
rect 679990 702715 680042 702767
rect 43510 702641 43562 702693
rect 58774 702641 58826 702693
rect 45046 702567 45098 702619
rect 58678 702567 58730 702619
rect 42070 700569 42122 700621
rect 42838 700569 42890 700621
rect 42166 699903 42218 699955
rect 42550 699903 42602 699955
rect 670774 699829 670826 699881
rect 679702 699829 679754 699881
rect 47542 699755 47594 699807
rect 59254 699755 59306 699807
rect 44950 699681 45002 699733
rect 58870 699681 58922 699733
rect 654166 694131 654218 694183
rect 675286 694131 675338 694183
rect 673750 692873 673802 692925
rect 675382 692873 675434 692925
rect 654070 691245 654122 691297
rect 675094 691245 675146 691297
rect 674902 690431 674954 690483
rect 675478 690431 675530 690483
rect 675190 689765 675242 689817
rect 675382 689765 675434 689817
rect 674806 689099 674858 689151
rect 675382 689099 675434 689151
rect 673558 688729 673610 688781
rect 675478 688729 675530 688781
rect 41782 688211 41834 688263
rect 50326 688211 50378 688263
rect 41590 687471 41642 687523
rect 47638 687471 47690 687523
rect 41782 687175 41834 687227
rect 47734 687175 47786 687227
rect 41590 686953 41642 687005
rect 43318 686953 43370 687005
rect 674326 686731 674378 686783
rect 675286 686731 675338 686783
rect 41590 685991 41642 686043
rect 43510 685991 43562 686043
rect 41782 685325 41834 685377
rect 43222 685325 43274 685377
rect 45046 685325 45098 685377
rect 41782 684141 41834 684193
rect 43414 684141 43466 684193
rect 44950 684141 45002 684193
rect 674422 683623 674474 683675
rect 675478 683623 675530 683675
rect 674518 682809 674570 682861
rect 675190 682809 675242 682861
rect 41782 681625 41834 681677
rect 42646 681625 42698 681677
rect 41782 679923 41834 679975
rect 42742 679923 42794 679975
rect 41782 679701 41834 679753
rect 42838 679701 42890 679753
rect 41782 677851 41834 677903
rect 43126 677851 43178 677903
rect 42454 677555 42506 677607
rect 42838 677555 42890 677607
rect 41782 677407 41834 677459
rect 43030 677407 43082 677459
rect 41590 677259 41642 677311
rect 42838 677259 42890 677311
rect 41782 677037 41834 677089
rect 42646 677037 42698 677089
rect 41782 675705 41834 675757
rect 47542 675705 47594 675757
rect 42454 671043 42506 671095
rect 59638 671043 59690 671095
rect 42742 670895 42794 670947
rect 42166 670747 42218 670799
rect 42742 670747 42794 670799
rect 42262 670451 42314 670503
rect 42262 670229 42314 670281
rect 42358 670229 42410 670281
rect 670774 669193 670826 669245
rect 676054 669193 676106 669245
rect 42166 668527 42218 668579
rect 42550 668527 42602 668579
rect 655510 668527 655562 668579
rect 676150 668527 676202 668579
rect 655318 668379 655370 668431
rect 676246 668379 676298 668431
rect 675094 668231 675146 668283
rect 676054 668231 676106 668283
rect 655126 668157 655178 668209
rect 676342 668157 676394 668209
rect 674710 668083 674762 668135
rect 676054 668083 676106 668135
rect 670678 668009 670730 668061
rect 675958 668009 676010 668061
rect 42166 667861 42218 667913
rect 42454 667861 42506 667913
rect 670870 667639 670922 667691
rect 675958 667639 676010 667691
rect 652246 666751 652298 666803
rect 670582 666751 670634 666803
rect 676246 666751 676298 666803
rect 42166 666677 42218 666729
rect 42838 666677 42890 666729
rect 649750 666677 649802 666729
rect 670678 666677 670730 666729
rect 670966 666307 671018 666359
rect 676246 666307 676298 666359
rect 42166 665271 42218 665323
rect 45142 665271 45194 665323
rect 674998 665197 675050 665249
rect 676246 665197 676298 665249
rect 42166 665123 42218 665175
rect 42646 665123 42698 665175
rect 674614 665123 674666 665175
rect 676054 665123 676106 665175
rect 42166 664827 42218 664879
rect 43126 664827 43178 664879
rect 42070 664161 42122 664213
rect 43030 664161 43082 664213
rect 42166 663347 42218 663399
rect 42358 663347 42410 663399
rect 674230 662311 674282 662363
rect 676054 662311 676106 662363
rect 42070 661053 42122 661105
rect 42550 661053 42602 661105
rect 673654 660609 673706 660661
rect 676054 660609 676106 660661
rect 42070 660387 42122 660439
rect 42454 660387 42506 660439
rect 42166 659869 42218 659921
rect 42934 659869 42986 659921
rect 673462 659869 673514 659921
rect 676246 659869 676298 659921
rect 42454 659499 42506 659551
rect 57718 659499 57770 659551
rect 47734 659425 47786 659477
rect 59158 659425 59210 659477
rect 45142 659351 45194 659403
rect 58774 659351 58826 659403
rect 42070 659055 42122 659107
rect 42646 659055 42698 659107
rect 654166 656761 654218 656813
rect 675382 656761 675434 656813
rect 42166 656687 42218 656739
rect 42550 656687 42602 656739
rect 649558 656687 649610 656739
rect 679798 656687 679850 656739
rect 50326 656613 50378 656665
rect 58198 656613 58250 656665
rect 47638 656539 47690 656591
rect 58390 656539 58442 656591
rect 655798 648177 655850 648229
rect 675190 648177 675242 648229
rect 673846 648029 673898 648081
rect 675286 648029 675338 648081
rect 655990 645143 656042 645195
rect 675094 645143 675146 645195
rect 41590 644847 41642 644899
rect 50326 644847 50378 644899
rect 673078 644551 673130 644603
rect 675286 644551 675338 644603
rect 41590 644255 41642 644307
rect 47734 644255 47786 644307
rect 41782 643959 41834 644011
rect 47830 643959 47882 644011
rect 673270 643885 673322 643937
rect 675286 643885 675338 643937
rect 41590 643737 41642 643789
rect 43510 643737 43562 643789
rect 673174 643367 673226 643419
rect 675286 643367 675338 643419
rect 41590 642775 41642 642827
rect 43414 642775 43466 642827
rect 41494 642479 41546 642531
rect 61942 642479 61994 642531
rect 673366 642257 673418 642309
rect 675190 642257 675242 642309
rect 41590 641295 41642 641347
rect 43318 641295 43370 641347
rect 41782 640555 41834 640607
rect 42838 640555 42890 640607
rect 674230 639075 674282 639127
rect 675094 639075 675146 639127
rect 41782 636707 41834 636759
rect 43030 636707 43082 636759
rect 41782 636041 41834 636093
rect 42550 636041 42602 636093
rect 41590 635375 41642 635427
rect 43126 635375 43178 635427
rect 674998 635005 675050 635057
rect 679702 635005 679754 635057
rect 41590 634487 41642 634539
rect 42838 634487 42890 634539
rect 41590 634191 41642 634243
rect 42742 634191 42794 634243
rect 41686 633895 41738 633947
rect 42934 633895 42986 633947
rect 41782 632489 41834 632541
rect 47638 632489 47690 632541
rect 43126 629307 43178 629359
rect 43510 629307 43562 629359
rect 42934 629159 42986 629211
rect 43318 629159 43370 629211
rect 674134 629085 674186 629137
rect 675094 629085 675146 629137
rect 42166 628789 42218 628841
rect 42838 628789 42890 628841
rect 42070 628715 42122 628767
rect 42742 628715 42794 628767
rect 42166 628123 42218 628175
rect 42646 628123 42698 628175
rect 42454 627975 42506 628027
rect 42646 627975 42698 628027
rect 42454 627827 42506 627879
rect 54646 627827 54698 627879
rect 42166 627383 42218 627435
rect 42262 626495 42314 626547
rect 42358 625385 42410 625437
rect 42166 625311 42218 625363
rect 42358 625237 42410 625289
rect 43318 625237 43370 625289
rect 655606 624941 655658 624993
rect 676246 624941 676298 624993
rect 54646 624793 54698 624845
rect 58966 624793 59018 624845
rect 42166 624645 42218 624697
rect 42454 624645 42506 624697
rect 42166 623461 42218 623513
rect 42550 623461 42602 623513
rect 672790 623387 672842 623439
rect 676054 623387 676106 623439
rect 669622 623091 669674 623143
rect 670870 623091 670922 623143
rect 676054 623091 676106 623143
rect 655414 622499 655466 622551
rect 676246 622499 676298 622551
rect 670774 622425 670826 622477
rect 676054 622425 676106 622477
rect 655222 622351 655274 622403
rect 676150 622351 676202 622403
rect 42166 622055 42218 622107
rect 47926 622055 47978 622107
rect 42070 621981 42122 622033
rect 42646 621981 42698 622033
rect 674518 621981 674570 622033
rect 676246 621981 676298 622033
rect 670966 621907 671018 621959
rect 676054 621907 676106 621959
rect 42262 621833 42314 621885
rect 42646 621833 42698 621885
rect 42454 621611 42506 621663
rect 42934 621611 42986 621663
rect 42358 621537 42410 621589
rect 43030 621537 43082 621589
rect 42934 621463 42986 621515
rect 43510 621463 43562 621515
rect 670870 621315 670922 621367
rect 676054 621315 676106 621367
rect 42454 620353 42506 620405
rect 43126 620353 43178 620405
rect 669814 619983 669866 620035
rect 670966 619983 671018 620035
rect 674902 619021 674954 619073
rect 676054 619021 676106 619073
rect 674422 618799 674474 618851
rect 676246 618799 676298 618851
rect 674326 618577 674378 618629
rect 676054 618577 676106 618629
rect 42262 617319 42314 617371
rect 42934 617319 42986 617371
rect 42166 616653 42218 616705
rect 42838 616653 42890 616705
rect 42262 616579 42314 616631
rect 42742 616579 42794 616631
rect 42934 616357 42986 616409
rect 58198 616357 58250 616409
rect 47830 616283 47882 616335
rect 58966 616283 59018 616335
rect 674806 616283 674858 616335
rect 676054 616283 676106 616335
rect 47926 616209 47978 616261
rect 59638 616209 59690 616261
rect 673750 615617 673802 615669
rect 676246 615617 676298 615669
rect 673558 614433 673610 614485
rect 676054 614433 676106 614485
rect 655798 613471 655850 613523
rect 675382 613471 675434 613523
rect 50326 613397 50378 613449
rect 59638 613397 59690 613449
rect 47734 613323 47786 613375
rect 59542 613323 59594 613375
rect 42070 612805 42122 612857
rect 42838 612805 42890 612857
rect 649654 610585 649706 610637
rect 679990 610585 680042 610637
rect 673750 603259 673802 603311
rect 675382 603259 675434 603311
rect 673654 602667 673706 602719
rect 675382 602667 675434 602719
rect 656566 602075 656618 602127
rect 674902 602075 674954 602127
rect 653974 602001 654026 602053
rect 674998 602001 675050 602053
rect 41590 601631 41642 601683
rect 50326 601631 50378 601683
rect 41782 601335 41834 601387
rect 47734 601335 47786 601387
rect 41782 600743 41834 600795
rect 47830 600743 47882 600795
rect 41782 600373 41834 600425
rect 43318 600373 43370 600425
rect 41782 599781 41834 599833
rect 43606 599781 43658 599833
rect 673462 599781 673514 599833
rect 675382 599781 675434 599833
rect 41782 599263 41834 599315
rect 43414 599263 43466 599315
rect 673558 599263 673610 599315
rect 675094 599263 675146 599315
rect 39862 599041 39914 599093
rect 41686 599041 41738 599093
rect 672886 598375 672938 598427
rect 675190 598375 675242 598427
rect 41782 598301 41834 598353
rect 43510 598301 43562 598353
rect 41782 597857 41834 597909
rect 43222 597857 43274 597909
rect 41590 596599 41642 596651
rect 42742 596599 42794 596651
rect 672982 596525 673034 596577
rect 675094 596525 675146 596577
rect 43222 596155 43274 596207
rect 45142 596155 45194 596207
rect 41590 595045 41642 595097
rect 43126 595045 43178 595097
rect 41782 594897 41834 594949
rect 42934 594897 42986 594949
rect 41590 593639 41642 593691
rect 42838 593639 42890 593691
rect 41686 592159 41738 592211
rect 42646 592159 42698 592211
rect 41974 590827 42026 590879
rect 43030 590827 43082 590879
rect 41590 590679 41642 590731
rect 42550 590679 42602 590731
rect 672790 590309 672842 590361
rect 679702 590309 679754 590361
rect 42166 587571 42218 587623
rect 43126 587571 43178 587623
rect 41590 587497 41642 587549
rect 56086 587497 56138 587549
rect 42454 587423 42506 587475
rect 42742 587423 42794 587475
rect 42838 587423 42890 587475
rect 43318 587423 43370 587475
rect 41878 587053 41930 587105
rect 43126 587053 43178 587105
rect 674614 586387 674666 586439
rect 675094 586387 675146 586439
rect 42742 585795 42794 585847
rect 43222 585795 43274 585847
rect 42262 585055 42314 585107
rect 42550 585055 42602 585107
rect 42358 584907 42410 584959
rect 43030 584907 43082 584959
rect 42454 584685 42506 584737
rect 58966 584685 59018 584737
rect 41782 584167 41834 584219
rect 42070 584167 42122 584219
rect 42646 584167 42698 584219
rect 41782 583945 41834 583997
rect 42262 582243 42314 582295
rect 42358 582021 42410 582073
rect 42358 581059 42410 581111
rect 42358 580689 42410 580741
rect 42358 579875 42410 579927
rect 42550 579801 42602 579853
rect 42454 578987 42506 579039
rect 47926 578987 47978 579039
rect 42358 578913 42410 578965
rect 42934 578913 42986 578965
rect 42934 578765 42986 578817
rect 43318 578765 43370 578817
rect 42262 578543 42314 578595
rect 42742 578543 42794 578595
rect 42262 577729 42314 577781
rect 42838 577729 42890 577781
rect 42454 576619 42506 576671
rect 43030 576619 43082 576671
rect 655510 576619 655562 576671
rect 676246 576619 676298 576671
rect 655318 576471 655370 576523
rect 676150 576471 676202 576523
rect 655126 576323 655178 576375
rect 676342 576323 676394 576375
rect 672790 576175 672842 576227
rect 676246 576175 676298 576227
rect 674230 575953 674282 576005
rect 676054 575953 676106 576005
rect 670774 575879 670826 575931
rect 675958 575879 676010 575931
rect 672598 575435 672650 575487
rect 675958 575435 676010 575487
rect 670870 574917 670922 574969
rect 675958 574917 676010 574969
rect 672694 574103 672746 574155
rect 676246 574103 676298 574155
rect 42070 573215 42122 573267
rect 42934 573215 42986 573267
rect 669910 573215 669962 573267
rect 670870 573215 670922 573267
rect 42454 573141 42506 573193
rect 58198 573141 58250 573193
rect 670102 573141 670154 573193
rect 670774 573141 670826 573193
rect 47830 573067 47882 573119
rect 58966 573067 59018 573119
rect 674134 573067 674186 573119
rect 676054 573067 676106 573119
rect 47926 572993 47978 573045
rect 59638 572993 59690 573045
rect 42166 572623 42218 572675
rect 42838 572623 42890 572675
rect 42070 570995 42122 571047
rect 43126 570995 43178 571047
rect 42358 570403 42410 570455
rect 42550 570403 42602 570455
rect 50326 570181 50378 570233
rect 59350 570181 59402 570233
rect 47734 570107 47786 570159
rect 59542 570107 59594 570159
rect 673366 569515 673418 569567
rect 676054 569515 676106 569567
rect 673270 569145 673322 569197
rect 676246 569145 676298 569197
rect 673846 568405 673898 568457
rect 676054 568405 676106 568457
rect 673078 567961 673130 568013
rect 676054 567961 676106 568013
rect 673174 567665 673226 567717
rect 676246 567665 676298 567717
rect 655702 567443 655754 567495
rect 675382 567443 675434 567495
rect 649846 564483 649898 564535
rect 679798 564483 679850 564535
rect 674038 559525 674090 559577
rect 675382 559525 675434 559577
rect 656566 558785 656618 558837
rect 675190 558785 675242 558837
rect 674806 558045 674858 558097
rect 675382 558045 675434 558097
rect 654166 555825 654218 555877
rect 675094 555825 675146 555877
rect 674326 555233 674378 555285
rect 675478 555233 675530 555285
rect 674998 553753 675050 553805
rect 675478 553753 675530 553805
rect 673846 553309 673898 553361
rect 675382 553309 675434 553361
rect 674230 551903 674282 551955
rect 675478 551903 675530 551955
rect 674518 548869 674570 548921
rect 675094 548869 675146 548921
rect 672790 547167 672842 547219
rect 679702 547167 679754 547219
rect 674422 543615 674474 543667
rect 675094 543615 675146 543667
rect 42358 541543 42410 541595
rect 57718 541543 57770 541595
rect 42454 541469 42506 541521
rect 57622 541469 57674 541521
rect 655606 533403 655658 533455
rect 676054 533403 676106 533455
rect 655414 533255 655466 533307
rect 676246 533255 676298 533307
rect 655222 533107 655274 533159
rect 676150 533107 676202 533159
rect 674710 532737 674762 532789
rect 676054 532737 676106 532789
rect 672598 532663 672650 532715
rect 675958 532663 676010 532715
rect 672406 531479 672458 531531
rect 672694 531479 672746 531531
rect 676246 531479 676298 531531
rect 42550 529925 42602 529977
rect 58198 529925 58250 529977
rect 674614 529851 674666 529903
rect 676054 529851 676106 529903
rect 673750 526669 673802 526721
rect 676054 526669 676106 526721
rect 672982 526299 673034 526351
rect 676054 526299 676106 526351
rect 673558 525929 673610 525981
rect 676246 525929 676298 525981
rect 42070 525707 42122 525759
rect 42550 525707 42602 525759
rect 673654 525189 673706 525241
rect 676054 525189 676106 525241
rect 673462 524819 673514 524871
rect 676054 524819 676106 524871
rect 672886 524449 672938 524501
rect 676246 524449 676298 524501
rect 50326 524301 50378 524353
rect 58582 524301 58634 524353
rect 47734 524227 47786 524279
rect 59350 524227 59402 524279
rect 42262 522229 42314 522281
rect 42454 522229 42506 522281
rect 649942 521267 649994 521319
rect 679798 521267 679850 521319
rect 676534 498253 676586 498305
rect 679702 498253 679754 498305
rect 655510 490039 655562 490091
rect 676246 490039 676298 490091
rect 655318 489891 655370 489943
rect 676246 489891 676298 489943
rect 655126 489743 655178 489795
rect 676150 489743 676202 489795
rect 676246 488707 676298 488759
rect 676726 488707 676778 488759
rect 670294 488115 670346 488167
rect 676054 488115 676106 488167
rect 676630 488115 676682 488167
rect 670486 487079 670538 487131
rect 676246 487079 676298 487131
rect 672502 486783 672554 486835
rect 676054 486783 676106 486835
rect 674518 486635 674570 486687
rect 676054 486635 676106 486687
rect 674038 486561 674090 486613
rect 676246 486561 676298 486613
rect 674326 485673 674378 485725
rect 676054 485673 676106 485725
rect 674806 483749 674858 483801
rect 676054 483749 676106 483801
rect 674422 483675 674474 483727
rect 675958 483675 676010 483727
rect 674998 483601 675050 483653
rect 676246 483601 676298 483653
rect 674230 482121 674282 482173
rect 676054 482121 676106 482173
rect 673846 480049 673898 480101
rect 676246 480049 676298 480101
rect 650038 478125 650090 478177
rect 679894 478125 679946 478177
rect 41863 476053 41915 476105
rect 50326 476053 50378 476105
rect 41850 475535 41902 475587
rect 47734 475535 47786 475587
rect 42041 474573 42093 474625
rect 43606 474573 43658 474625
rect 41782 472353 41834 472405
rect 58966 472353 59018 472405
rect 41782 463547 41834 463599
rect 47734 463547 47786 463599
rect 34486 463103 34538 463155
rect 41782 463103 41834 463155
rect 673846 440607 673898 440659
rect 675286 440607 675338 440659
rect 25846 437721 25898 437773
rect 39670 437795 39722 437847
rect 62518 437795 62570 437847
rect 670966 434909 671018 434961
rect 672502 434909 672554 434961
rect 41590 428443 41642 428495
rect 48022 428443 48074 428495
rect 41782 428073 41834 428125
rect 47926 428073 47978 428125
rect 39766 427629 39818 427681
rect 41590 427629 41642 427681
rect 41782 427555 41834 427607
rect 48118 427555 48170 427607
rect 41782 426519 41834 426571
rect 43222 426519 43274 426571
rect 41590 424965 41642 425017
rect 62614 423365 62666 423417
rect 40150 419119 40202 419171
rect 42454 419119 42506 419171
rect 39958 419045 40010 419097
rect 42934 419045 42986 419097
rect 39862 418971 39914 419023
rect 43030 418971 43082 419023
rect 41590 418083 41642 418135
rect 42742 418083 42794 418135
rect 34486 417713 34538 417765
rect 42358 417713 42410 417765
rect 41782 417195 41834 417247
rect 42838 417195 42890 417247
rect 41590 416455 41642 416507
rect 42646 416455 42698 416507
rect 41782 416085 41834 416137
rect 47830 416085 47882 416137
rect 42166 409453 42218 409505
rect 42454 409453 42506 409505
rect 42358 408121 42410 408173
rect 42838 408121 42890 408173
rect 42166 408047 42218 408099
rect 42550 408047 42602 408099
rect 42070 407973 42122 408025
rect 42454 407973 42506 408025
rect 42070 407455 42122 407507
rect 42742 407455 42794 407507
rect 42166 407011 42218 407063
rect 42646 407011 42698 407063
rect 42262 406049 42314 406101
rect 58486 406049 58538 406101
rect 42166 403163 42218 403215
rect 43030 403163 43082 403215
rect 42454 403015 42506 403067
rect 58774 403015 58826 403067
rect 673750 400573 673802 400625
rect 675958 400573 676010 400625
rect 655510 400499 655562 400551
rect 676054 400499 676106 400551
rect 655318 400425 655370 400477
rect 676246 400425 676298 400477
rect 655126 400351 655178 400403
rect 676150 400351 676202 400403
rect 48022 400277 48074 400329
rect 58198 400277 58250 400329
rect 672502 400277 672554 400329
rect 673846 400277 673898 400329
rect 676246 400277 676298 400329
rect 48118 400203 48170 400255
rect 58774 400203 58826 400255
rect 47926 400129 47978 400181
rect 59734 400129 59786 400181
rect 670966 399019 671018 399071
rect 676054 399019 676106 399071
rect 42070 394505 42122 394557
rect 57622 394505 57674 394557
rect 675190 392507 675242 392559
rect 676246 392507 676298 392559
rect 674998 391693 675050 391745
rect 676246 391693 676298 391745
rect 650134 388807 650186 388859
rect 679798 388807 679850 388859
rect 41590 385921 41642 385973
rect 48022 385921 48074 385973
rect 675094 385921 675146 385973
rect 675382 385921 675434 385973
rect 41590 385255 41642 385307
rect 48214 385255 48266 385307
rect 41878 384959 41930 385011
rect 48118 384959 48170 385011
rect 41590 384737 41642 384789
rect 43222 384737 43274 384789
rect 41590 383775 41642 383827
rect 43318 383775 43370 383827
rect 41590 382295 41642 382347
rect 43222 382295 43274 382347
rect 656566 381555 656618 381607
rect 675094 381555 675146 381607
rect 41782 379483 41834 379535
rect 42934 379483 42986 379535
rect 41590 377263 41642 377315
rect 42838 377263 42890 377315
rect 41494 374303 41546 374355
rect 42742 374303 42794 374355
rect 41782 374007 41834 374059
rect 43030 374007 43082 374059
rect 37366 373859 37418 373911
rect 41782 373859 41834 373911
rect 41590 373415 41642 373467
rect 42550 373415 42602 373467
rect 41590 373267 41642 373319
rect 47926 373267 47978 373319
rect 39958 372453 40010 372505
rect 42262 372453 42314 372505
rect 41686 371935 41738 371987
rect 42646 371935 42698 371987
rect 41782 370159 41834 370211
rect 41782 369937 41834 369989
rect 42166 366533 42218 366585
rect 42454 366533 42506 366585
rect 42262 364979 42314 365031
rect 42550 364979 42602 365031
rect 42262 364461 42314 364513
rect 42742 364461 42794 364513
rect 42166 363795 42218 363847
rect 42646 363795 42698 363847
rect 42262 363721 42314 363773
rect 43030 363721 43082 363773
rect 42070 362907 42122 362959
rect 42934 362907 42986 362959
rect 42454 362833 42506 362885
rect 58486 362833 58538 362885
rect 42358 359947 42410 359999
rect 59158 359947 59210 359999
rect 655318 357283 655370 357335
rect 676150 357283 676202 357335
rect 655222 357209 655274 357261
rect 676246 357209 676298 357261
rect 655126 357135 655178 357187
rect 676054 357135 676106 357187
rect 48022 357061 48074 357113
rect 58198 357061 58250 357113
rect 48118 356987 48170 357039
rect 59638 356987 59690 357039
rect 48214 356913 48266 356965
rect 58582 356913 58634 356965
rect 673750 356765 673802 356817
rect 676054 356765 676106 356817
rect 674518 352399 674570 352451
rect 676054 352399 676106 352451
rect 674806 351363 674858 351415
rect 676054 351363 676106 351415
rect 42166 351289 42218 351341
rect 57622 351289 57674 351341
rect 674134 348551 674186 348603
rect 676246 348551 676298 348603
rect 675190 348477 675242 348529
rect 676054 348477 676106 348529
rect 650230 345813 650282 345865
rect 679894 345813 679946 345865
rect 674902 345739 674954 345791
rect 675958 345739 676010 345791
rect 674998 345665 675050 345717
rect 676054 345665 676106 345717
rect 675094 345591 675146 345643
rect 676246 345591 676298 345643
rect 41782 342779 41834 342831
rect 48022 342779 48074 342831
rect 41782 342261 41834 342313
rect 48118 342261 48170 342313
rect 41782 341743 41834 341795
rect 48214 341743 48266 341795
rect 41782 341373 41834 341425
rect 43318 341373 43370 341425
rect 675766 341373 675818 341425
rect 675766 340707 675818 340759
rect 667798 340633 667850 340685
rect 675478 340633 675530 340685
rect 41590 340559 41642 340611
rect 43510 340559 43562 340611
rect 41782 340263 41834 340315
rect 43414 340263 43466 340315
rect 674806 339745 674858 339797
rect 675286 339745 675338 339797
rect 674518 339523 674570 339575
rect 675382 339523 675434 339575
rect 41590 339079 41642 339131
rect 43318 339079 43370 339131
rect 674134 336563 674186 336615
rect 675382 336563 675434 336615
rect 41590 334195 41642 334247
rect 42934 334195 42986 334247
rect 41878 334121 41930 334173
rect 43030 334121 43082 334173
rect 41494 331087 41546 331139
rect 42742 331087 42794 331139
rect 41398 331013 41450 331065
rect 42838 331013 42890 331065
rect 39766 330643 39818 330695
rect 42262 330643 42314 330695
rect 41878 330347 41930 330399
rect 45238 330347 45290 330399
rect 41590 328571 41642 328623
rect 42550 328571 42602 328623
rect 41686 328497 41738 328549
rect 42646 328497 42698 328549
rect 654166 328275 654218 328327
rect 667798 328275 667850 328327
rect 41782 327017 41834 327069
rect 41782 326721 41834 326773
rect 42070 323317 42122 323369
rect 42454 323317 42506 323369
rect 42262 321763 42314 321815
rect 42550 321763 42602 321815
rect 42262 321245 42314 321297
rect 42646 321245 42698 321297
rect 42166 321023 42218 321075
rect 42742 321023 42794 321075
rect 42262 319913 42314 319965
rect 42934 319913 42986 319965
rect 42454 319617 42506 319669
rect 58486 319617 58538 319669
rect 42454 319395 42506 319447
rect 42838 319395 42890 319447
rect 42454 316879 42506 316931
rect 43030 316879 43082 316931
rect 42550 316731 42602 316783
rect 59158 316731 59210 316783
rect 48214 313845 48266 313897
rect 59638 313845 59690 313897
rect 48022 313771 48074 313823
rect 58870 313771 58922 313823
rect 48118 313697 48170 313749
rect 59638 313697 59690 313749
rect 654262 311181 654314 311233
rect 676246 311181 676298 311233
rect 654166 311107 654218 311159
rect 676150 311107 676202 311159
rect 654070 311033 654122 311085
rect 676342 311033 676394 311085
rect 42166 308073 42218 308125
rect 59158 308073 59210 308125
rect 674134 305261 674186 305313
rect 676246 305261 676298 305313
rect 673942 302523 673994 302575
rect 675958 302523 676010 302575
rect 674038 302449 674090 302501
rect 676054 302449 676106 302501
rect 674230 302375 674282 302427
rect 676246 302375 676298 302427
rect 43414 300895 43466 300947
rect 63286 300895 63338 300947
rect 39766 299637 39818 299689
rect 43414 299637 43466 299689
rect 41782 299563 41834 299615
rect 43126 299563 43178 299615
rect 650326 299563 650378 299615
rect 679990 299563 680042 299615
rect 41782 299119 41834 299171
rect 51478 299119 51530 299171
rect 41782 298157 41834 298209
rect 43510 298157 43562 298209
rect 43222 298083 43274 298135
rect 61654 298083 61706 298135
rect 41782 297565 41834 297617
rect 43414 297565 43466 297617
rect 41782 297047 41834 297099
rect 43318 297047 43370 297099
rect 39958 296677 40010 296729
rect 43222 296677 43274 296729
rect 674134 295937 674186 295989
rect 675286 295937 675338 295989
rect 41590 295863 41642 295915
rect 43222 295863 43274 295915
rect 674230 295715 674282 295767
rect 675190 295715 675242 295767
rect 674038 294235 674090 294287
rect 675190 294235 675242 294287
rect 39670 293717 39722 293769
rect 58198 293717 58250 293769
rect 673942 291719 673994 291771
rect 675190 291719 675242 291771
rect 43126 291571 43178 291623
rect 59638 291571 59690 291623
rect 41590 291423 41642 291475
rect 43126 291423 43178 291475
rect 41590 290905 41642 290957
rect 42934 290905 42986 290957
rect 53302 290905 53354 290957
rect 59446 290905 59498 290957
rect 656566 290831 656618 290883
rect 675094 290831 675146 290883
rect 51478 288315 51530 288367
rect 58870 288315 58922 288367
rect 48022 288019 48074 288071
rect 59158 288019 59210 288071
rect 40246 287945 40298 287997
rect 42646 287945 42698 287997
rect 41494 287871 41546 287923
rect 42742 287871 42794 287923
rect 41878 287131 41930 287183
rect 45526 287131 45578 287183
rect 41590 285207 41642 285259
rect 42454 285207 42506 285259
rect 53206 285133 53258 285185
rect 59254 285133 59306 285185
rect 653782 284245 653834 284297
rect 658006 284245 658058 284297
rect 41782 283801 41834 283853
rect 41782 283505 41834 283557
rect 50326 282321 50378 282373
rect 58870 282321 58922 282373
rect 56182 282247 56234 282299
rect 57622 282247 57674 282299
rect 42166 281729 42218 281781
rect 42646 281729 42698 281781
rect 42070 280101 42122 280153
rect 42838 280101 42890 280153
rect 42166 279879 42218 279931
rect 42358 279879 42410 279931
rect 45334 279435 45386 279487
rect 59542 279435 59594 279487
rect 654166 279435 654218 279487
rect 663766 279435 663818 279487
rect 45430 279361 45482 279413
rect 59254 279361 59306 279413
rect 42166 278473 42218 278525
rect 43030 278473 43082 278525
rect 314902 278251 314954 278303
rect 408310 278251 408362 278303
rect 316630 278177 316682 278229
rect 411862 278177 411914 278229
rect 319510 278103 319562 278155
rect 418966 278103 419018 278155
rect 320950 278029 321002 278081
rect 422518 278029 422570 278081
rect 392278 277955 392330 278007
rect 599830 277955 599882 278007
rect 675094 277955 675146 278007
rect 679798 277955 679850 278007
rect 323830 277881 323882 277933
rect 429622 277881 429674 277933
rect 42166 277807 42218 277859
rect 42550 277807 42602 277859
rect 322102 277807 322154 277859
rect 426358 277807 426410 277859
rect 317878 277733 317930 277785
rect 415702 277733 415754 277785
rect 329302 277659 329354 277711
rect 444118 277659 444170 277711
rect 332374 277585 332426 277637
rect 451222 277585 451274 277637
rect 334966 277511 335018 277563
rect 458230 277511 458282 277563
rect 337846 277437 337898 277489
rect 465334 277437 465386 277489
rect 341014 277363 341066 277415
rect 472438 277363 472490 277415
rect 343894 277289 343946 277341
rect 479542 277289 479594 277341
rect 373846 277215 373898 277267
rect 554038 277215 554090 277267
rect 375094 277141 375146 277193
rect 557590 277141 557642 277193
rect 376822 277067 376874 277119
rect 561142 277067 561194 277119
rect 377974 276993 378026 277045
rect 564694 276993 564746 277045
rect 379414 276919 379466 276971
rect 568246 276919 568298 276971
rect 381046 276845 381098 276897
rect 571702 276845 571754 276897
rect 42358 276771 42410 276823
rect 43126 276771 43178 276823
rect 382294 276771 382346 276823
rect 575254 276771 575306 276823
rect 42550 276697 42602 276749
rect 42934 276697 42986 276749
rect 383638 276697 383690 276749
rect 578806 276697 578858 276749
rect 386518 276623 386570 276675
rect 585910 276623 585962 276675
rect 385366 276549 385418 276601
rect 582358 276549 582410 276601
rect 326422 276475 326474 276527
rect 437014 276475 437066 276527
rect 42838 276401 42890 276453
rect 59350 276401 59402 276453
rect 286102 276401 286154 276453
rect 336502 276401 336554 276453
rect 359158 276401 359210 276453
rect 517366 276401 517418 276453
rect 288694 276327 288746 276379
rect 343606 276327 343658 276379
rect 361750 276327 361802 276379
rect 524470 276327 524522 276379
rect 287350 276253 287402 276305
rect 340054 276253 340106 276305
rect 364630 276253 364682 276305
rect 531574 276253 531626 276305
rect 291862 276179 291914 276231
rect 350710 276179 350762 276231
rect 367702 276179 367754 276231
rect 538678 276179 538730 276231
rect 290326 276105 290378 276157
rect 347158 276105 347210 276157
rect 370294 276105 370346 276157
rect 545782 276105 545834 276157
rect 293014 276031 293066 276083
rect 354262 276031 354314 276083
rect 371062 276031 371114 276083
rect 546934 276031 546986 276083
rect 294646 275957 294698 276009
rect 357814 275957 357866 276009
rect 371926 275957 371978 276009
rect 549334 275957 549386 276009
rect 297334 275883 297386 275935
rect 364918 275883 364970 275935
rect 373462 275883 373514 275935
rect 552790 275883 552842 275935
rect 295894 275809 295946 275861
rect 361366 275809 361418 275861
rect 374614 275809 374666 275861
rect 556342 275809 556394 275861
rect 296470 275735 296522 275787
rect 362518 275735 362570 275787
rect 377494 275735 377546 275787
rect 563446 275735 563498 275787
rect 298966 275661 299018 275713
rect 368470 275661 368522 275713
rect 376246 275661 376298 275713
rect 559894 275661 559946 275713
rect 297814 275587 297866 275639
rect 366070 275587 366122 275639
rect 380566 275587 380618 275639
rect 570550 275587 570602 275639
rect 300214 275513 300266 275565
rect 372022 275513 372074 275565
rect 381814 275513 381866 275565
rect 574102 275513 574154 275565
rect 299158 275439 299210 275491
rect 369622 275439 369674 275491
rect 388918 275439 388970 275491
rect 591862 275439 591914 275491
rect 303286 275365 303338 275417
rect 379126 275365 379178 275417
rect 389590 275365 389642 275417
rect 593014 275365 593066 275417
rect 304438 275291 304490 275343
rect 382582 275291 382634 275343
rect 391990 275291 392042 275343
rect 598966 275291 599018 275343
rect 307318 275217 307370 275269
rect 389686 275217 389738 275269
rect 396310 275217 396362 275269
rect 609526 275217 609578 275269
rect 310390 275143 310442 275195
rect 396790 275143 396842 275195
rect 404950 275143 405002 275195
rect 314710 275069 314762 275121
rect 407446 275069 407498 275121
rect 311638 274995 311690 275047
rect 400342 274995 400394 275047
rect 407734 275143 407786 275195
rect 623734 275143 623786 275195
rect 408406 275069 408458 275121
rect 635542 275069 635594 275121
rect 630838 274995 630890 275047
rect 284470 274921 284522 274973
rect 332950 274921 333002 274973
rect 356182 274921 356234 274973
rect 510262 274921 510314 274973
rect 283030 274847 283082 274899
rect 329398 274847 329450 274899
rect 344566 274847 344618 274899
rect 481942 274847 481994 274899
rect 281782 274773 281834 274825
rect 325846 274773 325898 274825
rect 339094 274773 339146 274825
rect 467734 274773 467786 274825
rect 336022 274699 336074 274751
rect 460630 274699 460682 274751
rect 333142 274625 333194 274677
rect 453526 274625 453578 274677
rect 330454 274551 330506 274603
rect 446422 274551 446474 274603
rect 328822 274477 328874 274529
rect 442870 274477 442922 274529
rect 325942 274403 325994 274455
rect 435862 274403 435914 274455
rect 323350 274329 323402 274381
rect 428758 274329 428810 274381
rect 320182 274255 320234 274307
rect 421654 274255 421706 274307
rect 315958 274181 316010 274233
rect 410998 274181 411050 274233
rect 317302 274107 317354 274159
rect 414550 274107 414602 274159
rect 348502 274033 348554 274085
rect 401494 274033 401546 274085
rect 401782 274033 401834 274085
rect 407734 274033 407786 274085
rect 326806 273959 326858 274011
rect 373174 273959 373226 274011
rect 342166 273885 342218 273937
rect 387382 273885 387434 273937
rect 334294 273811 334346 273863
rect 380278 273811 380330 273863
rect 347062 273737 347114 273789
rect 394486 273737 394538 273789
rect 331222 273663 331274 273715
rect 376726 273663 376778 273715
rect 43030 273515 43082 273567
rect 59158 273515 59210 273567
rect 160438 273515 160490 273567
rect 207478 273515 207530 273567
rect 228982 273515 229034 273567
rect 242422 273515 242474 273567
rect 271030 273515 271082 273567
rect 299926 273515 299978 273567
rect 308374 273515 308426 273567
rect 344758 273515 344810 273567
rect 350038 273515 350090 273567
rect 494902 273515 494954 273567
rect 521302 273515 521354 273567
rect 631990 273515 632042 273567
rect 130870 273441 130922 273493
rect 190102 273441 190154 273493
rect 193558 273441 193610 273493
rect 221494 273441 221546 273493
rect 277078 273441 277130 273493
rect 314038 273441 314090 273493
rect 349462 273441 349514 273493
rect 493750 273441 493802 273493
rect 529846 273441 529898 273493
rect 624982 273441 625034 273493
rect 108406 273367 108458 273419
rect 109366 273367 109418 273419
rect 122614 273367 122666 273419
rect 123766 273367 123818 273419
rect 142678 273367 142730 273419
rect 209590 273367 209642 273419
rect 277750 273367 277802 273419
rect 316438 273367 316490 273419
rect 352438 273367 352490 273419
rect 500854 273367 500906 273419
rect 135574 273293 135626 273345
rect 209782 273293 209834 273345
rect 279670 273293 279722 273345
rect 321142 273293 321194 273345
rect 352630 273293 352682 273345
rect 502006 273293 502058 273345
rect 68278 273219 68330 273271
rect 142486 273219 142538 273271
rect 153334 273219 153386 273271
rect 207382 273219 207434 273271
rect 219574 273219 219626 273271
rect 238678 273219 238730 273271
rect 278230 273219 278282 273271
rect 317590 273219 317642 273271
rect 355510 273219 355562 273271
rect 509110 273219 509162 273271
rect 509206 273219 509258 273271
rect 548086 273219 548138 273271
rect 132022 273145 132074 273197
rect 209878 273145 209930 273197
rect 220726 273145 220778 273197
rect 239158 273145 239210 273197
rect 285622 273145 285674 273197
rect 335350 273145 335402 273197
rect 355030 273145 355082 273197
rect 507958 273145 508010 273197
rect 508246 273145 508298 273197
rect 639094 273145 639146 273197
rect 127318 273071 127370 273123
rect 209974 273071 210026 273123
rect 218326 273071 218378 273123
rect 238102 273071 238154 273123
rect 286774 273071 286826 273123
rect 338902 273071 338954 273123
rect 358582 273071 358634 273123
rect 125014 272997 125066 273049
rect 207286 272997 207338 273049
rect 217174 272997 217226 273049
rect 237622 272997 237674 273049
rect 284950 272997 285002 273049
rect 334198 272997 334250 273049
rect 360982 272997 361034 273049
rect 374806 272997 374858 273049
rect 374998 273071 375050 273123
rect 514966 273071 515018 273123
rect 516214 272997 516266 273049
rect 516310 272997 516362 273049
rect 580054 272997 580106 273049
rect 128470 272923 128522 272975
rect 210166 272923 210218 272975
rect 216022 272923 216074 272975
rect 236950 272923 237002 272975
rect 274198 272923 274250 272975
rect 306934 272923 306986 272975
rect 307030 272923 307082 272975
rect 358966 272923 359018 272975
rect 361270 272923 361322 272975
rect 523318 272923 523370 272975
rect 123670 272849 123722 272901
rect 209014 272849 209066 272901
rect 116662 272775 116714 272827
rect 207094 272775 207146 272827
rect 214774 272775 214826 272827
rect 236470 272849 236522 272901
rect 289942 272849 289994 272901
rect 346006 272849 346058 272901
rect 363574 272849 363626 272901
rect 120214 272701 120266 272753
rect 207862 272701 207914 272753
rect 212470 272701 212522 272753
rect 225910 272701 225962 272753
rect 113110 272627 113162 272679
rect 206038 272627 206090 272679
rect 213622 272627 213674 272679
rect 236278 272775 236330 272827
rect 292246 272775 292298 272827
rect 351862 272775 351914 272827
rect 364150 272775 364202 272827
rect 374806 272849 374858 272901
rect 522070 272849 522122 272901
rect 523030 272849 523082 272901
rect 583606 272849 583658 272901
rect 233686 272701 233738 272753
rect 244054 272701 244106 272753
rect 292726 272701 292778 272753
rect 353110 272701 353162 272753
rect 366550 272701 366602 272753
rect 374518 272701 374570 272753
rect 529174 272775 529226 272827
rect 530422 272701 530474 272753
rect 295414 272627 295466 272679
rect 360214 272627 360266 272679
rect 367126 272627 367178 272679
rect 537430 272627 537482 272679
rect 96598 272553 96650 272605
rect 106678 272553 106730 272605
rect 110806 272553 110858 272605
rect 205750 272553 205802 272605
rect 211222 272553 211274 272605
rect 235030 272553 235082 272605
rect 270262 272553 270314 272605
rect 297526 272553 297578 272605
rect 298294 272553 298346 272605
rect 367222 272553 367274 272605
rect 372694 272553 372746 272605
rect 106102 272479 106154 272531
rect 204022 272479 204074 272531
rect 210070 272479 210122 272531
rect 234550 272479 234602 272531
rect 270550 272479 270602 272531
rect 298678 272479 298730 272531
rect 301366 272479 301418 272531
rect 374326 272479 374378 272531
rect 374518 272553 374570 272605
rect 536278 272553 536330 272605
rect 551638 272479 551690 272531
rect 103702 272405 103754 272457
rect 203542 272405 203594 272457
rect 208918 272405 208970 272457
rect 234358 272405 234410 272457
rect 234934 272405 234986 272457
rect 244822 272405 244874 272457
rect 272758 272405 272810 272457
rect 303478 272405 303530 272457
rect 303958 272405 304010 272457
rect 381430 272405 381482 272457
rect 381526 272405 381578 272457
rect 572950 272405 573002 272457
rect 98998 272331 99050 272383
rect 199126 272331 199178 272383
rect 232534 272331 232586 272383
rect 243670 272331 243722 272383
rect 273430 272331 273482 272383
rect 305782 272331 305834 272383
rect 306838 272331 306890 272383
rect 388534 272331 388586 272383
rect 407446 272331 407498 272383
rect 587158 272331 587210 272383
rect 76534 272257 76586 272309
rect 84790 272183 84842 272235
rect 86326 272183 86378 272235
rect 104854 272183 104906 272235
rect 106486 272183 106538 272235
rect 106678 272257 106730 272309
rect 201622 272257 201674 272309
rect 207670 272257 207722 272309
rect 233878 272257 233930 272309
rect 236086 272257 236138 272309
rect 245302 272257 245354 272309
rect 275350 272257 275402 272309
rect 310486 272257 310538 272309
rect 195670 272183 195722 272235
rect 198262 272183 198314 272235
rect 224374 272183 224426 272235
rect 225910 272183 225962 272235
rect 235702 272183 235754 272235
rect 275158 272183 275210 272235
rect 309334 272183 309386 272235
rect 309910 272183 309962 272235
rect 395638 272257 395690 272309
rect 395926 272257 395978 272309
rect 608374 272257 608426 272309
rect 312790 272183 312842 272235
rect 402742 272183 402794 272235
rect 402934 272183 402986 272235
rect 622582 272183 622634 272235
rect 194710 272109 194762 272161
rect 224470 272109 224522 272161
rect 227830 272109 227882 272161
rect 242134 272109 242186 272161
rect 276310 272109 276362 272161
rect 312886 272109 312938 272161
rect 315478 272109 315530 272161
rect 409846 272109 409898 272161
rect 413686 272109 413738 272161
rect 643894 272109 643946 272161
rect 119062 272035 119114 272087
rect 120886 272035 120938 272087
rect 165142 272035 165194 272087
rect 166966 272035 167018 272087
rect 167542 272035 167594 272087
rect 210646 272035 210698 272087
rect 230134 272035 230186 272087
rect 242902 272035 242954 272087
rect 299446 272035 299498 272087
rect 174646 271961 174698 272013
rect 210550 271961 210602 272013
rect 231382 271961 231434 272013
rect 243094 271961 243146 272013
rect 159286 271887 159338 271939
rect 192982 271887 193034 271939
rect 195862 271887 195914 271939
rect 221686 271887 221738 271939
rect 272278 271887 272330 271939
rect 301942 271961 301994 272013
rect 306646 272035 306698 272087
rect 328246 272035 328298 272087
rect 346966 272035 347018 272087
rect 487798 272035 487850 272087
rect 327094 271961 327146 272013
rect 346486 271961 346538 272013
rect 486646 271961 486698 272013
rect 301078 271887 301130 271939
rect 324694 271887 324746 271939
rect 344086 271887 344138 271939
rect 480694 271887 480746 271939
rect 191158 271813 191210 271865
rect 227158 271813 227210 271865
rect 299350 271813 299402 271865
rect 306646 271813 306698 271865
rect 341494 271813 341546 271865
rect 473686 271813 473738 271865
rect 147382 271739 147434 271791
rect 149686 271739 149738 271791
rect 192310 271739 192362 271791
rect 224566 271739 224618 271791
rect 338614 271739 338666 271791
rect 466582 271739 466634 271791
rect 166294 271665 166346 271717
rect 198646 271665 198698 271717
rect 199414 271665 199466 271717
rect 221590 271665 221642 271717
rect 335446 271665 335498 271717
rect 459478 271665 459530 271717
rect 75286 271591 75338 271643
rect 77686 271591 77738 271643
rect 129718 271591 129770 271643
rect 132406 271591 132458 271643
rect 181750 271591 181802 271643
rect 210454 271591 210506 271643
rect 332566 271591 332618 271643
rect 452374 271591 452426 271643
rect 89494 271517 89546 271569
rect 92086 271517 92138 271569
rect 150934 271517 150986 271569
rect 152374 271517 152426 271569
rect 180502 271517 180554 271569
rect 205174 271517 205226 271569
rect 329974 271517 330026 271569
rect 445270 271517 445322 271569
rect 185206 271443 185258 271495
rect 210358 271443 210410 271495
rect 326902 271443 326954 271495
rect 438166 271443 438218 271495
rect 173398 271369 173450 271421
rect 200470 271369 200522 271421
rect 201814 271369 201866 271421
rect 223702 271369 223754 271421
rect 324022 271369 324074 271421
rect 431062 271369 431114 271421
rect 184054 271295 184106 271347
rect 205942 271295 205994 271347
rect 321430 271295 321482 271347
rect 423958 271295 424010 271347
rect 161590 271221 161642 271273
rect 163894 271221 163946 271273
rect 188758 271221 188810 271273
rect 210262 271221 210314 271273
rect 237238 271221 237290 271273
rect 245590 271221 245642 271273
rect 318358 271221 318410 271273
rect 416950 271221 417002 271273
rect 175798 271147 175850 271199
rect 178294 271147 178346 271199
rect 187606 271147 187658 271199
rect 205846 271147 205898 271199
rect 238486 271147 238538 271199
rect 246070 271147 246122 271199
rect 357910 271147 357962 271199
rect 374998 271147 375050 271199
rect 387286 271147 387338 271199
rect 407446 271147 407498 271199
rect 85942 271073 85994 271125
rect 198550 271073 198602 271125
rect 205366 271073 205418 271125
rect 232630 271073 232682 271125
rect 240790 271073 240842 271125
rect 247222 271073 247274 271125
rect 221878 270999 221930 271051
rect 239350 270999 239402 271051
rect 239542 270999 239594 271051
rect 241270 270999 241322 271051
rect 241942 270999 241994 271051
rect 247702 270999 247754 271051
rect 223030 270925 223082 270977
rect 240022 270925 240074 270977
rect 243190 270925 243242 270977
rect 247990 270925 248042 270977
rect 342742 270925 342794 270977
rect 348310 270925 348362 270977
rect 224278 270851 224330 270903
rect 240502 270851 240554 270903
rect 244342 270851 244394 270903
rect 248662 270851 248714 270903
rect 334102 270851 334154 270903
rect 337750 270851 337802 270903
rect 225430 270777 225482 270829
rect 241078 270777 241130 270829
rect 245494 270777 245546 270829
rect 249142 270777 249194 270829
rect 351382 270777 351434 270829
rect 355414 270777 355466 270829
rect 94198 270703 94250 270755
rect 94966 270703 95018 270755
rect 101302 270703 101354 270755
rect 103606 270703 103658 270755
rect 115510 270703 115562 270755
rect 118006 270703 118058 270755
rect 133270 270703 133322 270755
rect 135286 270703 135338 270755
rect 136822 270703 136874 270755
rect 138166 270703 138218 270755
rect 154486 270703 154538 270755
rect 155446 270703 155498 270755
rect 168694 270703 168746 270755
rect 169846 270703 169898 270755
rect 179350 270703 179402 270755
rect 181366 270703 181418 270755
rect 182902 270703 182954 270755
rect 184246 270703 184298 270755
rect 185494 270703 185546 270755
rect 186454 270703 186506 270755
rect 226582 270703 226634 270755
rect 239542 270703 239594 270755
rect 239638 270703 239690 270755
rect 246454 270703 246506 270755
rect 246742 270703 246794 270755
rect 249622 270703 249674 270755
rect 337942 270703 337994 270755
rect 341302 270703 341354 270755
rect 408982 270703 409034 270755
rect 413398 270703 413450 270755
rect 146230 270629 146282 270681
rect 214966 270629 215018 270681
rect 269686 270629 269738 270681
rect 296374 270629 296426 270681
rect 141526 270555 141578 270607
rect 213814 270555 213866 270607
rect 284374 270555 284426 270607
rect 284662 270555 284714 270607
rect 137974 270481 138026 270533
rect 212662 270481 212714 270533
rect 262966 270481 263018 270533
rect 279766 270481 279818 270533
rect 280150 270481 280202 270533
rect 293974 270555 294026 270607
rect 356662 270629 356714 270681
rect 371254 270629 371306 270681
rect 509206 270629 509258 270681
rect 296566 270555 296618 270607
rect 315286 270555 315338 270607
rect 345430 270555 345482 270607
rect 484246 270555 484298 270607
rect 322390 270481 322442 270533
rect 348406 270481 348458 270533
rect 491350 270481 491402 270533
rect 134422 270407 134474 270459
rect 211894 270407 211946 270459
rect 253942 270407 253994 270459
rect 257302 270407 257354 270459
rect 262486 270407 262538 270459
rect 278614 270407 278666 270459
rect 279286 270407 279338 270459
rect 284278 270407 284330 270459
rect 284758 270407 284810 270459
rect 318838 270407 318890 270459
rect 348118 270407 348170 270459
rect 490198 270407 490250 270459
rect 121462 270333 121514 270385
rect 208342 270333 208394 270385
rect 278902 270333 278954 270385
rect 284374 270333 284426 270385
rect 284854 270333 284906 270385
rect 323542 270333 323594 270385
rect 350710 270333 350762 270385
rect 497302 270333 497354 270385
rect 117910 270259 117962 270311
rect 207574 270259 207626 270311
rect 255286 270259 255338 270311
rect 260854 270259 260906 270311
rect 262006 270259 262058 270311
rect 277462 270259 277514 270311
rect 114358 270185 114410 270237
rect 206422 270185 206474 270237
rect 210550 270185 210602 270237
rect 222838 270185 222890 270237
rect 264886 270185 264938 270237
rect 284566 270259 284618 270311
rect 284662 270259 284714 270311
rect 319990 270259 320042 270311
rect 351286 270259 351338 270311
rect 498454 270259 498506 270311
rect 283702 270185 283754 270237
rect 330646 270185 330698 270237
rect 354070 270185 354122 270237
rect 505558 270185 505610 270237
rect 109558 270111 109610 270163
rect 205270 270111 205322 270163
rect 210358 270111 210410 270163
rect 225526 270111 225578 270163
rect 264694 270111 264746 270163
rect 283318 270111 283370 270163
rect 284182 270111 284234 270163
rect 331798 270111 331850 270163
rect 353686 270111 353738 270163
rect 504406 270111 504458 270163
rect 107254 270037 107306 270089
rect 204694 270037 204746 270089
rect 210262 270037 210314 270089
rect 226678 270037 226730 270089
rect 265366 270037 265418 270089
rect 285718 270037 285770 270089
rect 286294 270037 286346 270089
rect 334102 270037 334154 270089
rect 356758 270037 356810 270089
rect 511510 270037 511562 270089
rect 102550 269963 102602 270015
rect 203350 269963 203402 270015
rect 210454 269963 210506 270015
rect 224758 269963 224810 270015
rect 267094 269963 267146 270015
rect 289270 269963 289322 270015
rect 100150 269889 100202 269941
rect 202870 269889 202922 269941
rect 205174 269889 205226 269941
rect 224086 269889 224138 269941
rect 256246 269889 256298 269941
rect 263254 269889 263306 269941
rect 266518 269889 266570 269941
rect 95446 269815 95498 269867
rect 185590 269815 185642 269867
rect 93046 269741 93098 269793
rect 200950 269815 201002 269867
rect 205942 269815 205994 269867
rect 225238 269815 225290 269867
rect 261814 269815 261866 269867
rect 276214 269815 276266 269867
rect 280630 269889 280682 269941
rect 284854 269889 284906 269941
rect 288502 269889 288554 269941
rect 342454 269963 342506 270015
rect 356950 269963 357002 270015
rect 512662 269963 512714 270015
rect 288022 269815 288074 269867
rect 90646 269667 90698 269719
rect 199702 269741 199754 269793
rect 205846 269741 205898 269793
rect 226006 269741 226058 269793
rect 255766 269741 255818 269793
rect 262102 269741 262154 269793
rect 267286 269741 267338 269793
rect 290422 269741 290474 269793
rect 83638 269593 83690 269645
rect 198070 269667 198122 269719
rect 200470 269667 200522 269719
rect 222358 269667 222410 269719
rect 287926 269667 287978 269719
rect 337942 269889 337994 269941
rect 359830 269889 359882 269941
rect 519766 269889 519818 269941
rect 290614 269815 290666 269867
rect 342742 269815 342794 269867
rect 359350 269815 359402 269867
rect 518518 269815 518570 269867
rect 291094 269741 291146 269793
rect 349558 269741 349610 269793
rect 362806 269741 362858 269793
rect 526870 269741 526922 269793
rect 362230 269667 362282 269719
rect 525622 269667 525674 269719
rect 198646 269593 198698 269645
rect 220534 269593 220586 269645
rect 249046 269593 249098 269645
rect 250294 269593 250346 269645
rect 259894 269593 259946 269645
rect 271510 269593 271562 269645
rect 276502 269593 276554 269645
rect 291574 269593 291626 269645
rect 293494 269593 293546 269645
rect 351382 269593 351434 269645
rect 365302 269593 365354 269645
rect 532726 269593 532778 269645
rect 82390 269519 82442 269571
rect 197398 269519 197450 269571
rect 206518 269519 206570 269571
rect 233398 269519 233450 269571
rect 269206 269519 269258 269571
rect 295126 269519 295178 269571
rect 297046 269519 297098 269571
rect 363670 269519 363722 269571
rect 365686 269519 365738 269571
rect 533878 269519 533930 269571
rect 87190 269445 87242 269497
rect 199030 269445 199082 269497
rect 202966 269445 203018 269497
rect 231958 269445 232010 269497
rect 268630 269445 268682 269497
rect 293878 269445 293930 269497
rect 299638 269445 299690 269497
rect 370774 269445 370826 269497
rect 379894 269445 379946 269497
rect 569398 269445 569450 269497
rect 81238 269371 81290 269423
rect 196822 269371 196874 269423
rect 204118 269371 204170 269423
rect 232150 269371 232202 269423
rect 258646 269371 258698 269423
rect 269110 269371 269162 269423
rect 272950 269371 273002 269423
rect 304630 269371 304682 269423
rect 308278 269371 308330 269423
rect 392086 269371 392138 269423
rect 394390 269371 394442 269423
rect 604822 269371 604874 269423
rect 74134 269297 74186 269349
rect 194998 269297 195050 269349
rect 200662 269297 200714 269349
rect 230998 269297 231050 269349
rect 274678 269297 274730 269349
rect 308182 269297 308234 269349
rect 311158 269297 311210 269349
rect 399190 269297 399242 269349
rect 399958 269297 400010 269349
rect 619030 269297 619082 269349
rect 67030 269223 67082 269275
rect 192598 269223 192650 269275
rect 197110 269223 197162 269275
rect 229558 269223 229610 269275
rect 260566 269223 260618 269275
rect 273910 269223 273962 269275
rect 275830 269223 275882 269275
rect 311734 269223 311786 269275
rect 314230 269223 314282 269275
rect 406294 269223 406346 269275
rect 145078 269149 145130 269201
rect 214486 269149 214538 269201
rect 149782 269075 149834 269127
rect 216214 269075 216266 269127
rect 253366 269075 253418 269127
rect 256150 269075 256202 269127
rect 257014 269075 257066 269127
rect 264406 269075 264458 269127
rect 266038 269075 266090 269127
rect 286870 269149 286922 269201
rect 286966 269149 287018 269201
rect 292822 269149 292874 269201
rect 306358 269149 306410 269201
rect 342166 269149 342218 269201
rect 345238 269149 345290 269201
rect 483094 269149 483146 269201
rect 281302 269075 281354 269127
rect 301078 269075 301130 269127
rect 303766 269075 303818 269127
rect 334294 269075 334346 269127
rect 342646 269075 342698 269127
rect 477142 269075 477194 269127
rect 148630 269001 148682 269053
rect 215734 269001 215786 269053
rect 282070 269001 282122 269053
rect 299446 269001 299498 269053
rect 305686 269001 305738 269053
rect 384982 269001 385034 269053
rect 406582 269001 406634 269053
rect 408406 269001 408458 269053
rect 152182 268927 152234 268979
rect 216694 268927 216746 268979
rect 253174 268927 253226 268979
rect 254998 268927 255050 268979
rect 259414 268927 259466 268979
rect 270358 268927 270410 268979
rect 277558 268927 277610 268979
rect 296566 268927 296618 268979
rect 302038 268927 302090 268979
rect 331222 268927 331274 268979
rect 339766 268927 339818 268979
rect 470134 268927 470186 268979
rect 156886 268853 156938 268905
rect 218134 268853 218186 268905
rect 260086 268853 260138 268905
rect 272662 268853 272714 268905
rect 300694 268853 300746 268905
rect 326806 268853 326858 268905
rect 336886 268853 336938 268905
rect 463030 268853 463082 268905
rect 163990 268779 164042 268831
rect 219958 268779 220010 268831
rect 258166 268779 258218 268831
rect 267958 268779 268010 268831
rect 268438 268779 268490 268831
rect 286966 268779 287018 268831
rect 289174 268779 289226 268831
rect 308374 268779 308426 268831
rect 334294 268779 334346 268831
rect 455926 268779 455978 268831
rect 155734 268705 155786 268757
rect 217366 268705 217418 268757
rect 257686 268705 257738 268757
rect 266806 268705 266858 268757
rect 295222 268705 295274 268757
rect 307030 268705 307082 268757
rect 331222 268705 331274 268757
rect 448822 268705 448874 268757
rect 162838 268631 162890 268683
rect 219286 268631 219338 268683
rect 254614 268631 254666 268683
rect 258550 268631 258602 268683
rect 271510 268631 271562 268683
rect 300982 268631 301034 268683
rect 328342 268631 328394 268683
rect 441718 268631 441770 268683
rect 171094 268557 171146 268609
rect 221782 268557 221834 268609
rect 325750 268557 325802 268609
rect 434614 268557 434666 268609
rect 169750 268483 169802 268535
rect 221206 268483 221258 268535
rect 261238 268483 261290 268535
rect 275062 268483 275114 268535
rect 322582 268483 322634 268535
rect 427510 268483 427562 268535
rect 176950 268409 177002 268461
rect 223414 268409 223466 268461
rect 319702 268409 319754 268461
rect 420502 268409 420554 268461
rect 178198 268335 178250 268387
rect 223606 268335 223658 268387
rect 247894 268335 247946 268387
rect 249814 268335 249866 268387
rect 255094 268335 255146 268387
rect 259702 268335 259754 268387
rect 317110 268335 317162 268387
rect 408982 268335 409034 268387
rect 185590 268261 185642 268313
rect 201142 268261 201194 268313
rect 207478 268261 207530 268313
rect 212470 268261 212522 268313
rect 221494 268261 221546 268313
rect 227830 268261 227882 268313
rect 312310 268261 312362 268313
rect 348502 268261 348554 268313
rect 192982 268187 193034 268239
rect 218614 268187 218666 268239
rect 224374 268187 224426 268239
rect 230038 268187 230090 268239
rect 257494 268187 257546 268239
rect 265654 268187 265706 268239
rect 309238 268187 309290 268239
rect 347062 268187 347114 268239
rect 408502 268187 408554 268239
rect 640342 268187 640394 268239
rect 190102 268113 190154 268165
rect 210742 268113 210794 268165
rect 223702 268113 223754 268165
rect 231478 268113 231530 268165
rect 264118 268113 264170 268165
rect 282166 268113 282218 268165
rect 302614 268113 302666 268165
rect 377878 268113 377930 268165
rect 384118 268113 384170 268165
rect 516310 268113 516362 268165
rect 207382 268039 207434 268091
rect 216886 268039 216938 268091
rect 221590 268039 221642 268091
rect 230518 268039 230570 268091
rect 252694 268039 252746 268091
rect 253750 268039 253802 268091
rect 342166 268039 342218 268091
rect 359446 268039 359498 268091
rect 209878 267965 209930 268017
rect 211414 267965 211466 268017
rect 221686 267965 221738 268017
rect 229078 267965 229130 268017
rect 333622 267965 333674 268017
rect 351382 267965 351434 268017
rect 210646 267891 210698 267943
rect 221014 267891 221066 267943
rect 224470 267891 224522 267943
rect 228406 267891 228458 267943
rect 263638 267891 263690 267943
rect 281014 267891 281066 267943
rect 282550 267891 282602 267943
rect 299350 267891 299402 267943
rect 336694 267891 336746 267943
rect 354262 267891 354314 267943
rect 199126 267817 199178 267869
rect 202294 267817 202346 267869
rect 207286 267817 207338 267869
rect 209494 267817 209546 267869
rect 209782 267817 209834 267869
rect 212374 267817 212426 267869
rect 212470 267817 212522 267869
rect 218902 267817 218954 267869
rect 224566 267817 224618 267869
rect 227638 267817 227690 267869
rect 339286 267817 339338 267869
rect 360406 267817 360458 267869
rect 401302 267817 401354 267869
rect 402934 267817 402986 267869
rect 409942 267817 409994 267869
rect 413686 267817 413738 267869
rect 351958 267743 352010 267795
rect 499606 267743 499658 267795
rect 354838 267669 354890 267721
rect 506710 267669 506762 267721
rect 357430 267595 357482 267647
rect 513814 267595 513866 267647
rect 360310 267521 360362 267573
rect 520918 267521 520970 267573
rect 363382 267447 363434 267499
rect 528022 267447 528074 267499
rect 365974 267373 366026 267425
rect 535126 267373 535178 267425
rect 368950 267299 369002 267351
rect 542230 267299 542282 267351
rect 372502 267225 372554 267277
rect 550486 267225 550538 267277
rect 384886 267151 384938 267203
rect 581206 267151 581258 267203
rect 386038 267077 386090 267129
rect 584758 267077 584810 267129
rect 387766 267003 387818 267055
rect 588310 267003 588362 267055
rect 301846 266929 301898 266981
rect 375286 266929 375338 266981
rect 394678 266929 394730 266981
rect 606070 266929 606122 266981
rect 306166 266855 306218 266907
rect 386134 266855 386186 266907
rect 393238 266855 393290 266907
rect 602518 266855 602570 266907
rect 305014 266781 305066 266833
rect 383830 266781 383882 266833
rect 397558 266781 397610 266833
rect 613078 266781 613130 266833
rect 308758 266707 308810 266759
rect 392950 266707 393002 266759
rect 398230 266707 398282 266759
rect 614326 266707 614378 266759
rect 308086 266633 308138 266685
rect 390934 266633 390986 266685
rect 400630 266633 400682 266685
rect 620182 266633 620234 266685
rect 310678 266559 310730 266611
rect 398038 266559 398090 266611
rect 403222 266559 403274 266611
rect 627286 266559 627338 266611
rect 313558 266485 313610 266537
rect 405046 266485 405098 266537
rect 406102 266485 406154 266537
rect 634390 266485 634442 266537
rect 313078 266411 313130 266463
rect 403894 266411 403946 266463
rect 409174 266411 409226 266463
rect 641494 266411 641546 266463
rect 45046 266337 45098 266389
rect 673750 266337 673802 266389
rect 348886 266263 348938 266315
rect 492598 266263 492650 266315
rect 346006 266189 346058 266241
rect 485494 266189 485546 266241
rect 343318 266115 343370 266167
rect 478390 266115 478442 266167
rect 340246 266041 340298 266093
rect 471286 266041 471338 266093
rect 337366 265967 337418 266019
rect 464182 265967 464234 266019
rect 334774 265893 334826 265945
rect 457078 265893 457130 265945
rect 331894 265819 331946 265871
rect 449974 265819 450026 265871
rect 327574 265745 327626 265797
rect 439318 265745 439370 265797
rect 324502 265671 324554 265723
rect 432310 265671 432362 265723
rect 321622 265597 321674 265649
rect 425206 265597 425258 265649
rect 408022 265523 408074 265575
rect 508246 265523 508298 265575
rect 319030 265449 319082 265501
rect 418102 265449 418154 265501
rect 656566 265375 656618 265427
rect 676054 265375 676106 265427
rect 656278 265227 656330 265279
rect 676246 265227 676298 265279
rect 656086 265079 656138 265131
rect 676150 265079 676202 265131
rect 23062 265005 23114 265057
rect 43510 265005 43562 265057
rect 673750 265005 673802 265057
rect 676054 265005 676106 265057
rect 42166 264931 42218 264983
rect 53302 264931 53354 264983
rect 45718 264783 45770 264835
rect 669814 264931 669866 264983
rect 46006 264709 46058 264761
rect 669622 264857 669674 264909
rect 359446 264783 359498 264835
rect 475990 264783 476042 264835
rect 328054 264709 328106 264761
rect 440566 264709 440618 264761
rect 331126 264635 331178 264687
rect 447670 264635 447722 264687
rect 354262 264561 354314 264613
rect 461782 264561 461834 264613
rect 360406 264487 360458 264539
rect 468886 264487 468938 264539
rect 351382 264413 351434 264465
rect 454774 264413 454826 264465
rect 399382 264117 399434 264169
rect 410998 264117 411050 264169
rect 267718 264043 267770 264095
rect 276502 264043 276554 264095
rect 324982 264043 325034 264095
rect 433462 264043 433514 264095
rect 387958 263969 388010 264021
rect 589462 263969 589514 264021
rect 390838 263895 390890 263947
rect 596566 263895 596618 263947
rect 393910 263821 393962 263873
rect 603670 263821 603722 263873
rect 396790 263747 396842 263799
rect 610774 263747 610826 263799
rect 401110 263673 401162 263725
rect 23350 263599 23402 263651
rect 43318 263599 43370 263651
rect 46006 263599 46058 263651
rect 403990 263599 404042 263651
rect 410998 263673 411050 263725
rect 617878 263673 617930 263725
rect 23254 263525 23306 263577
rect 43222 263525 43274 263577
rect 45718 263525 45770 263577
rect 409654 263525 409706 263577
rect 621430 263599 621482 263651
rect 628438 263525 628490 263577
rect 642646 263451 642698 263503
rect 23158 262119 23210 262171
rect 43318 262119 43370 262171
rect 420406 262119 420458 262171
rect 606166 262119 606218 262171
rect 674806 262119 674858 262171
rect 676246 262119 676298 262171
rect 187222 260639 187274 260691
rect 189718 260639 189770 260691
rect 674614 259381 674666 259433
rect 676054 259381 676106 259433
rect 420406 259233 420458 259285
rect 606262 259233 606314 259285
rect 675190 259233 675242 259285
rect 676054 259233 676106 259285
rect 674518 256939 674570 256991
rect 676054 256939 676106 256991
rect 674710 256421 674762 256473
rect 676054 256421 676106 256473
rect 40246 256347 40298 256399
rect 59062 256347 59114 256399
rect 420406 256347 420458 256399
rect 606358 256347 606410 256399
rect 674998 256347 675050 256399
rect 676246 256347 676298 256399
rect 41782 255385 41834 255437
rect 53206 255385 53258 255437
rect 47926 255089 47978 255141
rect 186262 255089 186314 255141
rect 47734 255015 47786 255067
rect 186070 255015 186122 255067
rect 41782 254941 41834 254993
rect 43414 254941 43466 254993
rect 47830 254941 47882 254993
rect 186454 254941 186506 254993
rect 44854 254867 44906 254919
rect 185974 254867 186026 254919
rect 41782 254423 41834 254475
rect 43222 254423 43274 254475
rect 41590 253609 41642 253661
rect 56182 253609 56234 253661
rect 674902 253535 674954 253587
rect 676054 253535 676106 253587
rect 44950 253461 45002 253513
rect 58966 253461 59018 253513
rect 420406 253461 420458 253513
rect 603286 253461 603338 253513
rect 646678 253461 646730 253513
rect 679702 253461 679754 253513
rect 106486 252277 106538 252329
rect 156886 252277 156938 252329
rect 92086 252203 92138 252255
rect 145366 252203 145418 252255
rect 109366 252129 109418 252181
rect 171286 252129 171338 252181
rect 97846 252055 97898 252107
rect 182806 252055 182858 252107
rect 56086 251981 56138 252033
rect 186646 251981 186698 252033
rect 665878 250649 665930 250701
rect 675382 250649 675434 250701
rect 420406 250575 420458 250627
rect 603382 250575 603434 250627
rect 674806 250205 674858 250257
rect 675286 250205 675338 250257
rect 120886 249909 120938 249961
rect 145654 249909 145706 249961
rect 132406 249835 132458 249887
rect 159862 249835 159914 249887
rect 135286 249761 135338 249813
rect 168502 249761 168554 249813
rect 138166 249687 138218 249739
rect 171478 249687 171530 249739
rect 141046 249613 141098 249665
rect 180022 249613 180074 249665
rect 123766 249539 123818 249591
rect 165718 249539 165770 249591
rect 126646 249465 126698 249517
rect 177046 249465 177098 249517
rect 94966 249391 95018 249443
rect 154006 249391 154058 249443
rect 118006 249317 118058 249369
rect 182902 249317 182954 249369
rect 77686 249243 77738 249295
rect 145462 249243 145514 249295
rect 80566 249169 80618 249221
rect 162646 249169 162698 249221
rect 86326 249095 86378 249147
rect 174166 249095 174218 249147
rect 674614 249095 674666 249147
rect 675286 249095 675338 249147
rect 41878 247837 41930 247889
rect 42838 247837 42890 247889
rect 420310 247763 420362 247815
rect 603478 247763 603530 247815
rect 420406 247689 420458 247741
rect 629206 247689 629258 247741
rect 655894 247615 655946 247667
rect 665878 247615 665930 247667
rect 674518 247467 674570 247519
rect 675094 247467 675146 247519
rect 103606 246727 103658 246779
rect 165526 246727 165578 246779
rect 112246 246653 112298 246705
rect 185782 246653 185834 246705
rect 47542 246579 47594 246631
rect 186358 246579 186410 246631
rect 47446 246505 47498 246557
rect 186550 246505 186602 246557
rect 47638 246431 47690 246483
rect 186742 246431 186794 246483
rect 45526 246357 45578 246409
rect 186838 246357 186890 246409
rect 44566 246283 44618 246335
rect 186166 246283 186218 246335
rect 45238 246209 45290 246261
rect 187030 246209 187082 246261
rect 41590 245099 41642 245151
rect 145750 245099 145802 245151
rect 41590 244951 41642 245003
rect 145558 244951 145610 245003
rect 44758 244877 44810 244929
rect 186934 244877 186986 244929
rect 420406 244803 420458 244855
rect 629302 244803 629354 244855
rect 40246 244729 40298 244781
rect 42454 244729 42506 244781
rect 41494 244655 41546 244707
rect 42646 244655 42698 244707
rect 34486 243545 34538 243597
rect 42358 243545 42410 243597
rect 41686 243175 41738 243227
rect 42934 243175 42986 243227
rect 44662 242805 44714 242857
rect 185590 242805 185642 242857
rect 44854 242731 44906 242783
rect 185878 242731 185930 242783
rect 674710 242731 674762 242783
rect 675382 242731 675434 242783
rect 44566 242657 44618 242709
rect 185686 242657 185738 242709
rect 41590 242583 41642 242635
rect 142582 242583 142634 242635
rect 41878 241917 41930 241969
rect 43126 241917 43178 241969
rect 420406 241917 420458 241969
rect 600406 241917 600458 241969
rect 41782 240585 41834 240637
rect 41782 240363 41834 240415
rect 380854 239919 380906 239971
rect 412054 239919 412106 239971
rect 409558 239845 409610 239897
rect 412150 239845 412202 239897
rect 357142 239771 357194 239823
rect 434614 239771 434666 239823
rect 377302 239697 377354 239749
rect 446710 239697 446762 239749
rect 385366 239623 385418 239675
rect 470902 239623 470954 239675
rect 374422 239549 374474 239601
rect 488278 239549 488330 239601
rect 334294 239475 334346 239527
rect 458806 239475 458858 239527
rect 394678 239401 394730 239453
rect 532822 239401 532874 239453
rect 397942 239327 397994 239379
rect 541462 239327 541514 239379
rect 406006 239253 406058 239305
rect 550870 239253 550922 239305
rect 420406 239179 420458 239231
rect 599158 239179 599210 239231
rect 350422 239105 350474 239157
rect 508630 239105 508682 239157
rect 368566 239031 368618 239083
rect 544822 239031 544874 239083
rect 324406 238957 324458 239009
rect 455158 238957 455210 239009
rect 323926 238883 323978 238935
rect 455062 238883 455114 238935
rect 326710 238809 326762 238861
rect 462550 238809 462602 238861
rect 328918 238735 328970 238787
rect 464758 238735 464810 238787
rect 329878 238661 329930 238713
rect 468598 238661 468650 238713
rect 332662 238587 332714 238639
rect 474646 238587 474698 238639
rect 42166 238513 42218 238565
rect 42454 238513 42506 238565
rect 335734 238513 335786 238565
rect 480694 238513 480746 238565
rect 336694 238439 336746 238491
rect 478102 238439 478154 238491
rect 42550 238365 42602 238417
rect 338998 238365 339050 238417
rect 486742 238365 486794 238417
rect 341782 238291 341834 238343
rect 492790 238291 492842 238343
rect 345334 238217 345386 238269
rect 500278 238217 500330 238269
rect 346678 238143 346730 238195
rect 503350 238143 503402 238195
rect 42550 238069 42602 238121
rect 349942 238069 349994 238121
rect 509398 238069 509450 238121
rect 353494 237995 353546 238047
rect 514678 237995 514730 238047
rect 352726 237921 352778 237973
rect 512758 237921 512810 237973
rect 355702 237847 355754 237899
rect 522166 237847 522218 237899
rect 363094 237773 363146 237825
rect 535126 237773 535178 237825
rect 275350 237699 275402 237751
rect 357526 237699 357578 237751
rect 361750 237699 361802 237751
rect 533494 237699 533546 237751
rect 277078 237625 277130 237677
rect 363670 237625 363722 237677
rect 364438 237625 364490 237677
rect 535798 237625 535850 237677
rect 365878 237551 365930 237603
rect 541078 237551 541130 237603
rect 320854 237477 320906 237529
rect 450454 237477 450506 237529
rect 317590 237403 317642 237455
rect 444502 237403 444554 237455
rect 317110 237329 317162 237381
rect 440662 237329 440714 237381
rect 314806 237255 314858 237307
rect 438358 237255 438410 237307
rect 311542 237181 311594 237233
rect 432406 237181 432458 237233
rect 308566 237107 308618 237159
rect 426358 237107 426410 237159
rect 310774 237033 310826 237085
rect 428662 237033 428714 237085
rect 305782 236959 305834 237011
rect 420310 236959 420362 237011
rect 298966 236885 299018 236937
rect 404470 236885 404522 236937
rect 405910 236885 405962 236937
rect 414454 236885 414506 236937
rect 279862 236811 279914 236863
rect 370486 236811 370538 236863
rect 386998 236811 387050 236863
rect 387574 236811 387626 236863
rect 397846 236811 397898 236863
rect 413590 236811 413642 236863
rect 278422 236737 278474 236789
rect 366742 236737 366794 236789
rect 382390 236737 382442 236789
rect 398038 236737 398090 236789
rect 397078 236663 397130 236715
rect 397750 236663 397802 236715
rect 397462 236589 397514 236641
rect 413398 236589 413450 236641
rect 387190 236515 387242 236567
rect 387862 236515 387914 236567
rect 397462 236441 397514 236493
rect 397942 236441 397994 236493
rect 378166 236367 378218 236419
rect 397366 236367 397418 236419
rect 410710 236367 410762 236419
rect 442198 236367 442250 236419
rect 387094 236293 387146 236345
rect 387478 236293 387530 236345
rect 390742 236293 390794 236345
rect 492022 236293 492074 236345
rect 394582 236219 394634 236271
rect 505654 236219 505706 236271
rect 400342 236145 400394 236197
rect 523798 236145 523850 236197
rect 251062 236071 251114 236123
rect 273622 236071 273674 236123
rect 277558 236071 277610 236123
rect 313942 236071 313994 236123
rect 326134 236071 326186 236123
rect 334294 236071 334346 236123
rect 341206 236071 341258 236123
rect 374422 236071 374474 236123
rect 376342 236071 376394 236123
rect 208438 235997 208490 236049
rect 223222 235997 223274 236049
rect 247990 235997 248042 236049
rect 209686 235923 209738 235975
rect 226198 235923 226250 235975
rect 243286 235923 243338 235975
rect 271030 235923 271082 235975
rect 276118 235997 276170 236049
rect 310198 235997 310250 236049
rect 313846 235997 313898 236049
rect 357142 235997 357194 236049
rect 371830 235997 371882 236049
rect 406006 235997 406058 236049
rect 276214 235923 276266 235975
rect 280630 235923 280682 235975
rect 322006 235923 322058 235975
rect 386710 235923 386762 235975
rect 405622 235923 405674 235975
rect 410038 236071 410090 236123
rect 584566 236071 584618 236123
rect 406294 235997 406346 236049
rect 415414 235997 415466 236049
rect 413878 235923 413930 235975
rect 208918 235849 208970 235901
rect 226966 235849 227018 235901
rect 234262 235849 234314 235901
rect 264694 235849 264746 235901
rect 279286 235849 279338 235901
rect 318262 235849 318314 235901
rect 326230 235849 326282 235901
rect 460246 235849 460298 235901
rect 208822 235775 208874 235827
rect 224758 235775 224810 235827
rect 237526 235775 237578 235827
rect 268150 235775 268202 235827
rect 290326 235775 290378 235827
rect 334102 235775 334154 235827
rect 343510 235775 343562 235827
rect 495766 235775 495818 235827
rect 211222 235701 211274 235753
rect 229270 235701 229322 235753
rect 231190 235701 231242 235753
rect 259030 235701 259082 235753
rect 262870 235701 262922 235753
rect 305014 235701 305066 235753
rect 317206 235701 317258 235753
rect 410710 235701 410762 235753
rect 411862 235701 411914 235753
rect 413686 235701 413738 235753
rect 210646 235627 210698 235679
rect 230038 235627 230090 235679
rect 239350 235627 239402 235679
rect 210070 235553 210122 235605
rect 227830 235553 227882 235605
rect 236470 235553 236522 235605
rect 282934 235553 282986 235605
rect 287062 235627 287114 235679
rect 318454 235627 318506 235679
rect 358006 235627 358058 235679
rect 400342 235627 400394 235679
rect 287350 235553 287402 235605
rect 311158 235553 311210 235605
rect 408982 235627 409034 235679
rect 409174 235627 409226 235679
rect 588886 235627 588938 235679
rect 405622 235553 405674 235605
rect 411862 235553 411914 235605
rect 412150 235553 412202 235605
rect 590518 235553 590570 235605
rect 212950 235479 213002 235531
rect 232342 235479 232394 235531
rect 238006 235479 238058 235531
rect 285910 235479 285962 235531
rect 299830 235479 299882 235531
rect 354262 235479 354314 235531
rect 394966 235479 395018 235531
rect 587350 235479 587402 235531
rect 42166 235405 42218 235457
rect 42550 235405 42602 235457
rect 211990 235405 212042 235457
rect 233014 235405 233066 235457
rect 242134 235405 242186 235457
rect 293398 235405 293450 235457
rect 294838 235405 294890 235457
rect 338902 235405 338954 235457
rect 339478 235405 339530 235457
rect 395062 235405 395114 235457
rect 396790 235405 396842 235457
rect 588406 235405 588458 235457
rect 214198 235331 214250 235383
rect 220534 235331 220586 235383
rect 220630 235331 220682 235383
rect 241846 235331 241898 235383
rect 249718 235331 249770 235383
rect 302326 235331 302378 235383
rect 304822 235331 304874 235383
rect 362326 235331 362378 235383
rect 393430 235331 393482 235383
rect 587062 235331 587114 235383
rect 209302 235257 209354 235309
rect 228502 235257 228554 235309
rect 229750 235257 229802 235309
rect 253558 235257 253610 235309
rect 257494 235257 257546 235309
rect 308182 235257 308234 235309
rect 334966 235257 335018 235309
rect 391702 235257 391754 235309
rect 396310 235257 396362 235309
rect 587638 235257 587690 235309
rect 42262 235183 42314 235235
rect 42454 235183 42506 235235
rect 211606 235109 211658 235161
rect 230710 235183 230762 235235
rect 232918 235183 232970 235235
rect 223894 235109 223946 235161
rect 244726 235109 244778 235161
rect 288886 235183 288938 235235
rect 345718 235183 345770 235235
rect 392182 235183 392234 235235
rect 587254 235183 587306 235235
rect 262006 235109 262058 235161
rect 266134 235109 266186 235161
rect 324118 235109 324170 235161
rect 332182 235109 332234 235161
rect 385366 235109 385418 235161
rect 387670 235109 387722 235161
rect 583414 235109 583466 235161
rect 207478 235035 207530 235087
rect 223990 235035 224042 235087
rect 246646 235035 246698 235087
rect 299254 235035 299306 235087
rect 309334 235035 309386 235087
rect 370582 235035 370634 235087
rect 394870 235035 394922 235087
rect 596086 235035 596138 235087
rect 211030 234961 211082 235013
rect 231574 234961 231626 235013
rect 243862 234961 243914 235013
rect 296470 234961 296522 235013
rect 298006 234961 298058 235013
rect 362422 234961 362474 235013
rect 362518 234961 362570 235013
rect 394678 234961 394730 235013
rect 398998 234961 399050 235013
rect 605974 234961 606026 235013
rect 213430 234887 213482 234939
rect 204406 234813 204458 234865
rect 210166 234813 210218 234865
rect 204790 234739 204842 234791
rect 210454 234739 210506 234791
rect 220534 234887 220586 234939
rect 235318 234887 235370 234939
rect 235702 234887 235754 234939
rect 265078 234887 265130 234939
rect 268918 234887 268970 234939
rect 331414 234887 331466 234939
rect 333430 234887 333482 234939
rect 394774 234887 394826 234939
rect 398614 234887 398666 234939
rect 605302 234887 605354 234939
rect 225526 234813 225578 234865
rect 260182 234813 260234 234865
rect 260278 234813 260330 234865
rect 323158 234813 323210 234865
rect 327670 234813 327722 234865
rect 392470 234813 392522 234865
rect 403606 234813 403658 234865
rect 615862 234813 615914 234865
rect 236086 234739 236138 234791
rect 254230 234739 254282 234791
rect 306742 234739 306794 234791
rect 321622 234739 321674 234791
rect 387286 234739 387338 234791
rect 406678 234739 406730 234791
rect 621814 234739 621866 234791
rect 206518 234665 206570 234717
rect 222454 234665 222506 234717
rect 225142 234665 225194 234717
rect 247702 234665 247754 234717
rect 251158 234665 251210 234717
rect 304150 234665 304202 234717
rect 315286 234665 315338 234717
rect 394678 234665 394730 234717
rect 408118 234665 408170 234717
rect 624886 234665 624938 234717
rect 202870 234591 202922 234643
rect 214870 234591 214922 234643
rect 222262 234591 222314 234643
rect 202006 234517 202058 234569
rect 213430 234517 213482 234569
rect 240214 234591 240266 234643
rect 263830 234591 263882 234643
rect 267478 234591 267530 234643
rect 282358 234591 282410 234643
rect 286678 234591 286730 234643
rect 325750 234591 325802 234643
rect 329302 234591 329354 234643
rect 449302 234591 449354 234643
rect 243958 234517 244010 234569
rect 206134 234443 206186 234495
rect 211990 234443 212042 234495
rect 235606 234443 235658 234495
rect 250582 234517 250634 234569
rect 255286 234517 255338 234569
rect 278038 234517 278090 234569
rect 283894 234517 283946 234569
rect 322198 234517 322250 234569
rect 323542 234517 323594 234569
rect 434902 234517 434954 234569
rect 250486 234443 250538 234495
rect 267958 234443 268010 234495
rect 273046 234443 273098 234495
rect 305110 234443 305162 234495
rect 314422 234443 314474 234495
rect 426166 234443 426218 234495
rect 206998 234369 207050 234421
rect 221782 234369 221834 234421
rect 237046 234369 237098 234421
rect 258934 234369 258986 234421
rect 262486 234369 262538 234421
rect 290902 234369 290954 234421
rect 292918 234369 292970 234421
rect 311158 234369 311210 234421
rect 312694 234369 312746 234421
rect 407446 234369 407498 234421
rect 203254 234295 203306 234347
rect 206806 234295 206858 234347
rect 206902 234295 206954 234347
rect 220246 234295 220298 234347
rect 239830 234295 239882 234347
rect 260950 234295 261002 234347
rect 271606 234295 271658 234347
rect 302134 234295 302186 234347
rect 308470 234295 308522 234347
rect 414742 234295 414794 234347
rect 42262 234221 42314 234273
rect 42934 234221 42986 234273
rect 201526 234221 201578 234273
rect 211894 234221 211946 234273
rect 211990 234221 212042 234273
rect 221014 234221 221066 234273
rect 242902 234221 242954 234273
rect 261142 234221 261194 234273
rect 261238 234221 261290 234273
rect 288022 234221 288074 234273
rect 295222 234221 295274 234273
rect 348694 234221 348746 234273
rect 352150 234221 352202 234273
rect 398134 234221 398186 234273
rect 398230 234221 398282 234273
rect 406006 234221 406058 234273
rect 407254 234221 407306 234273
rect 503926 234221 503978 234273
rect 200278 234147 200330 234199
rect 210358 234147 210410 234199
rect 210454 234147 210506 234199
rect 219382 234147 219434 234199
rect 256534 234147 256586 234199
rect 279286 234147 279338 234199
rect 283990 234147 284042 234199
rect 311350 234147 311402 234199
rect 318358 234147 318410 234199
rect 371638 234147 371690 234199
rect 378550 234147 378602 234199
rect 399190 234147 399242 234199
rect 403510 234147 403562 234199
rect 495382 234147 495434 234199
rect 200182 234073 200234 234125
rect 208822 234073 208874 234125
rect 198742 233999 198794 234051
rect 207382 233999 207434 234051
rect 207862 233999 207914 234051
rect 225526 234073 225578 234125
rect 244342 234073 244394 234125
rect 264886 234073 264938 234125
rect 268534 234073 268586 234125
rect 293782 234073 293834 234125
rect 295702 234073 295754 234125
rect 341206 234073 341258 234125
rect 345910 234073 345962 234125
rect 400150 234073 400202 234125
rect 401782 234073 401834 234125
rect 484630 234073 484682 234125
rect 247414 233999 247466 234051
rect 266326 233999 266378 234051
rect 267094 233999 267146 234051
rect 290998 233999 291050 234051
rect 301654 233999 301706 234051
rect 344086 233999 344138 234051
rect 344374 233999 344426 234051
rect 394870 233999 394922 234051
rect 396694 233999 396746 234051
rect 475222 233999 475274 234051
rect 198358 233925 198410 233977
rect 205942 233925 205994 233977
rect 206806 233925 206858 233977
rect 216502 233925 216554 233977
rect 259798 233925 259850 233977
rect 281206 233925 281258 233977
rect 305206 233925 305258 233977
rect 351382 233925 351434 233977
rect 361270 233925 361322 233977
rect 432022 233925 432074 233977
rect 197494 233851 197546 233903
rect 204310 233851 204362 233903
rect 205174 233851 205226 233903
rect 217174 233851 217226 233903
rect 258358 233851 258410 233903
rect 279190 233851 279242 233903
rect 296086 233851 296138 233903
rect 339094 233851 339146 233903
rect 370294 233851 370346 233903
rect 427894 233851 427946 233903
rect 196918 233777 196970 233829
rect 202870 233777 202922 233829
rect 204214 233777 204266 233829
rect 215542 233777 215594 233829
rect 253462 233777 253514 233829
rect 270838 233777 270890 233829
rect 285142 233777 285194 233829
rect 325366 233777 325418 233829
rect 354934 233777 354986 233829
rect 407350 233777 407402 233829
rect 407446 233777 407498 233829
rect 423286 233777 423338 233829
rect 196534 233703 196586 233755
rect 200566 233703 200618 233755
rect 201046 233703 201098 233755
rect 209686 233703 209738 233755
rect 210166 233703 210218 233755
rect 217942 233703 217994 233755
rect 294454 233703 294506 233755
rect 331222 233703 331274 233755
rect 338038 233703 338090 233755
rect 386134 233703 386186 233755
rect 398134 233703 398186 233755
rect 403030 233703 403082 233755
rect 408982 233703 409034 233755
rect 410614 233703 410666 233755
rect 195670 233629 195722 233681
rect 201334 233629 201386 233681
rect 202486 233629 202538 233681
rect 212566 233629 212618 233681
rect 306262 233629 306314 233681
rect 344470 233629 344522 233681
rect 363478 233629 363530 233681
rect 363766 233629 363818 233681
rect 383638 233629 383690 233681
rect 408118 233629 408170 233681
rect 194230 233555 194282 233607
rect 198358 233555 198410 233607
rect 199126 233555 199178 233607
rect 205078 233555 205130 233607
rect 205558 233555 205610 233607
rect 192886 233481 192938 233533
rect 195286 233481 195338 233533
rect 195574 233481 195626 233533
rect 199798 233481 199850 233533
rect 200662 233481 200714 233533
rect 208150 233481 208202 233533
rect 228406 233555 228458 233607
rect 238102 233555 238154 233607
rect 259894 233555 259946 233607
rect 267766 233555 267818 233607
rect 302902 233555 302954 233607
rect 337366 233555 337418 233607
rect 348886 233555 348938 233607
rect 394582 233555 394634 233607
rect 218710 233481 218762 233533
rect 240598 233481 240650 233533
rect 290422 233481 290474 233533
rect 297238 233481 297290 233533
rect 328342 233481 328394 233533
rect 338614 233481 338666 233533
rect 466486 233481 466538 233533
rect 42454 233407 42506 233459
rect 43126 233407 43178 233459
rect 193846 233407 193898 233459
rect 196822 233407 196874 233459
rect 197974 233407 198026 233459
rect 203638 233407 203690 233459
rect 203926 233407 203978 233459
rect 214198 233407 214250 233459
rect 264406 233407 264458 233459
rect 271798 233407 271850 233459
rect 287446 233407 287498 233459
rect 311254 233407 311306 233459
rect 320278 233407 320330 233459
rect 448246 233407 448298 233459
rect 193270 233333 193322 233385
rect 194614 233333 194666 233385
rect 195190 233333 195242 233385
rect 197494 233333 197546 233385
rect 197878 233333 197930 233385
rect 202102 233333 202154 233385
rect 202390 233333 202442 233385
rect 211126 233333 211178 233385
rect 226678 233333 226730 233385
rect 238966 233333 239018 233385
rect 261622 233333 261674 233385
rect 269014 233333 269066 233385
rect 270454 233333 270506 233385
rect 275062 233333 275114 233385
rect 288406 233333 288458 233385
rect 311062 233333 311114 233385
rect 324790 233333 324842 233385
rect 327286 233333 327338 233385
rect 335350 233333 335402 233385
rect 463606 233333 463658 233385
rect 192406 233259 192458 233311
rect 193750 233259 193802 233311
rect 194710 233259 194762 233311
rect 196054 233259 196106 233311
rect 196150 233259 196202 233311
rect 199126 233259 199178 233311
rect 199702 233259 199754 233311
rect 206614 233259 206666 233311
rect 253846 233259 253898 233311
rect 256246 233259 256298 233311
rect 257974 233259 258026 233311
rect 269110 233259 269162 233311
rect 270262 233259 270314 233311
rect 273526 233259 273578 233311
rect 297142 233259 297194 233311
rect 317878 233259 317930 233311
rect 319894 233259 319946 233311
rect 377302 233259 377354 233311
rect 380470 233259 380522 233311
rect 382966 233259 383018 233311
rect 395926 233259 395978 233311
rect 400246 233259 400298 233311
rect 401206 233259 401258 233311
rect 408886 233259 408938 233311
rect 258742 233185 258794 233237
rect 326710 233185 326762 233237
rect 340822 233185 340874 233237
rect 491254 233185 491306 233237
rect 495382 233185 495434 233237
rect 614998 233185 615050 233237
rect 260662 233111 260714 233163
rect 331318 233111 331370 233163
rect 347062 233111 347114 233163
rect 501046 233111 501098 233163
rect 262102 233037 262154 233089
rect 334198 233037 334250 233089
rect 350326 233037 350378 233089
rect 507094 233037 507146 233089
rect 265750 232963 265802 233015
rect 338038 232963 338090 233015
rect 353110 232963 353162 233015
rect 513142 232963 513194 233015
rect 281302 232889 281354 232941
rect 288982 232889 289034 232941
rect 289942 232889 289994 232941
rect 382774 232889 382826 232941
rect 410038 232889 410090 232941
rect 572086 232889 572138 232941
rect 263926 232815 263978 232867
rect 337270 232815 337322 232867
rect 356278 232815 356330 232867
rect 519190 232815 519242 232867
rect 216598 232741 216650 232793
rect 242134 232741 242186 232793
rect 265174 232741 265226 232793
rect 340246 232741 340298 232793
rect 359062 232741 359114 232793
rect 525238 232741 525290 232793
rect 237622 232667 237674 232719
rect 284374 232667 284426 232719
rect 295318 232667 295370 232719
rect 397366 232667 397418 232719
rect 399190 232667 399242 232719
rect 566710 232667 566762 232719
rect 219766 232593 219818 232645
rect 248086 232593 248138 232645
rect 266614 232593 266666 232645
rect 343222 232593 343274 232645
rect 362134 232593 362186 232645
rect 531286 232593 531338 232645
rect 218038 232519 218090 232571
rect 245110 232519 245162 232571
rect 268438 232519 268490 232571
rect 346294 232519 346346 232571
rect 346774 232519 346826 232571
rect 356086 232519 356138 232571
rect 365398 232519 365450 232571
rect 537238 232519 537290 232571
rect 221110 232445 221162 232497
rect 251158 232445 251210 232497
rect 269686 232445 269738 232497
rect 349366 232445 349418 232497
rect 365014 232445 365066 232497
rect 539542 232445 539594 232497
rect 222550 232371 222602 232423
rect 254230 232371 254282 232423
rect 271222 232371 271274 232423
rect 222934 232297 222986 232349
rect 255670 232297 255722 232349
rect 274870 232297 274922 232349
rect 346774 232297 346826 232349
rect 346966 232371 347018 232423
rect 361366 232371 361418 232423
rect 368182 232371 368234 232423
rect 543382 232371 543434 232423
rect 352342 232297 352394 232349
rect 366262 232297 366314 232349
rect 542614 232297 542666 232349
rect 224278 232223 224330 232275
rect 257206 232223 257258 232275
rect 274198 232223 274250 232275
rect 358294 232223 358346 232275
rect 369526 232223 369578 232275
rect 548566 232223 548618 232275
rect 147862 232149 147914 232201
rect 154102 232149 154154 232201
rect 226294 232149 226346 232201
rect 261718 232149 261770 232201
rect 272950 232149 273002 232201
rect 355318 232149 355370 232201
rect 372694 232149 372746 232201
rect 552406 232149 552458 232201
rect 227062 232075 227114 232127
rect 263254 232075 263306 232127
rect 277462 232075 277514 232127
rect 364438 232075 364490 232127
rect 368086 232075 368138 232127
rect 545590 232075 545642 232127
rect 233878 232001 233930 232053
rect 274486 232001 274538 232053
rect 275734 232001 275786 232053
rect 346966 232001 347018 232053
rect 354262 232001 354314 232053
rect 367126 232001 367178 232053
rect 372310 232001 372362 232053
rect 554710 232001 554762 232053
rect 234838 231927 234890 231979
rect 278326 231927 278378 231979
rect 280246 231927 280298 231979
rect 370390 231927 370442 231979
rect 374518 231927 374570 231979
rect 557014 231927 557066 231979
rect 233206 231853 233258 231905
rect 275350 231853 275402 231905
rect 278998 231853 279050 231905
rect 367414 231853 367466 231905
rect 375766 231853 375818 231905
rect 558358 231853 558410 231905
rect 235990 231779 236042 231831
rect 281302 231779 281354 231831
rect 281974 231779 282026 231831
rect 373462 231779 373514 231831
rect 378934 231779 378986 231831
rect 564502 231779 564554 231831
rect 259126 231705 259178 231757
rect 328150 231705 328202 231757
rect 337558 231705 337610 231757
rect 485206 231705 485258 231757
rect 257590 231631 257642 231683
rect 325174 231631 325226 231683
rect 334870 231631 334922 231683
rect 479158 231631 479210 231683
rect 255766 231557 255818 231609
rect 320662 231557 320714 231609
rect 327094 231557 327146 231609
rect 464086 231557 464138 231609
rect 248374 231483 248426 231535
rect 305494 231483 305546 231535
rect 312214 231483 312266 231535
rect 433846 231483 433898 231535
rect 290806 231409 290858 231461
rect 374614 231409 374666 231461
rect 403126 231409 403178 231461
rect 520726 231409 520778 231461
rect 292534 231335 292586 231387
rect 379990 231335 380042 231387
rect 400150 231335 400202 231387
rect 499606 231335 499658 231387
rect 245206 231261 245258 231313
rect 299446 231261 299498 231313
rect 300214 231261 300266 231313
rect 385846 231261 385898 231313
rect 395062 231261 395114 231313
rect 485974 231261 486026 231313
rect 293494 231187 293546 231239
rect 365590 231187 365642 231239
rect 394774 231187 394826 231239
rect 473878 231187 473930 231239
rect 256150 231113 256202 231165
rect 322102 231113 322154 231165
rect 337366 231113 337418 231165
rect 252982 231039 253034 231091
rect 314518 231039 314570 231091
rect 344470 231039 344522 231091
rect 308182 230965 308234 231017
rect 323638 230965 323690 231017
rect 328342 230965 328394 231017
rect 401398 230965 401450 231017
rect 323158 230891 323210 230943
rect 329590 230891 329642 230943
rect 331222 230891 331274 230943
rect 395350 230891 395402 230943
rect 414742 231113 414794 231165
rect 424054 231113 424106 231165
rect 415702 230965 415754 231017
rect 419542 230891 419594 230943
rect 325750 230817 325802 230869
rect 380278 230817 380330 230869
rect 387286 230817 387338 230869
rect 449686 230817 449738 230869
rect 290710 230743 290762 230795
rect 297334 230743 297386 230795
rect 313942 230743 313994 230795
rect 362134 230743 362186 230795
rect 362326 230743 362378 230795
rect 416470 230743 416522 230795
rect 318262 230669 318314 230721
rect 365110 230669 365162 230721
rect 367126 230669 367178 230721
rect 409654 230669 409706 230721
rect 302326 230595 302378 230647
rect 308566 230595 308618 230647
rect 322198 230595 322250 230647
rect 374134 230595 374186 230647
rect 306742 230521 306794 230573
rect 317590 230521 317642 230573
rect 325366 230521 325418 230573
rect 377110 230521 377162 230573
rect 149398 230447 149450 230499
rect 156982 230447 157034 230499
rect 299254 230447 299306 230499
rect 302518 230447 302570 230499
rect 304150 230447 304202 230499
rect 311638 230447 311690 230499
rect 322006 230447 322058 230499
rect 368182 230447 368234 230499
rect 426166 230447 426218 230499
rect 436150 230447 436202 230499
rect 246166 230373 246218 230425
rect 298678 230373 298730 230425
rect 324022 230373 324074 230425
rect 346966 230373 347018 230425
rect 369910 230373 369962 230425
rect 387286 230373 387338 230425
rect 434902 230373 434954 230425
rect 454294 230373 454346 230425
rect 245782 230299 245834 230351
rect 300982 230299 301034 230351
rect 314902 230299 314954 230351
rect 439990 230299 440042 230351
rect 248950 230225 249002 230277
rect 304822 230225 304874 230277
rect 317974 230225 318026 230277
rect 445942 230225 445994 230277
rect 247030 230151 247082 230203
rect 303958 230151 304010 230203
rect 313462 230151 313514 230203
rect 436918 230151 436970 230203
rect 449302 230151 449354 230203
rect 466390 230151 466442 230203
rect 248758 230077 248810 230129
rect 307030 230077 307082 230129
rect 325846 230077 325898 230129
rect 461014 230077 461066 230129
rect 463606 230077 463658 230129
rect 478390 230077 478442 230129
rect 251926 230003 251978 230055
rect 310774 230003 310826 230055
rect 328534 230003 328586 230055
rect 251542 229929 251594 229981
rect 313078 229929 313130 229981
rect 331606 229929 331658 229981
rect 346966 230003 347018 230055
rect 458038 230003 458090 230055
rect 466486 230003 466538 230055
rect 484438 230003 484490 230055
rect 503926 230003 503978 230055
rect 622678 230003 622730 230055
rect 227446 229855 227498 229907
rect 264790 229855 264842 229907
rect 290902 229855 290954 229907
rect 331894 229855 331946 229907
rect 467062 229929 467114 229981
rect 475222 229929 475274 229981
rect 601462 229929 601514 229981
rect 473110 229855 473162 229907
rect 480886 229855 480938 229907
rect 609046 229855 609098 229907
rect 254806 229781 254858 229833
rect 319126 229781 319178 229833
rect 336310 229781 336362 229833
rect 482134 229781 482186 229833
rect 484630 229781 484682 229833
rect 612118 229781 612170 229833
rect 220150 229707 220202 229759
rect 249718 229707 249770 229759
rect 253078 229707 253130 229759
rect 316150 229707 316202 229759
rect 348502 229707 348554 229759
rect 504022 229707 504074 229759
rect 244246 229633 244298 229685
rect 298006 229633 298058 229685
rect 298582 229633 298634 229685
rect 406774 229633 406826 229685
rect 409846 229633 409898 229685
rect 565942 229633 565994 229685
rect 221590 229559 221642 229611
rect 252598 229559 252650 229611
rect 255190 229559 255242 229611
rect 316822 229559 316874 229611
rect 351766 229559 351818 229611
rect 510166 229559 510218 229611
rect 264310 229485 264362 229537
rect 334966 229485 335018 229537
rect 354838 229485 354890 229537
rect 516118 229485 516170 229537
rect 228886 229411 228938 229463
rect 267862 229411 267914 229463
rect 283510 229411 283562 229463
rect 368854 229411 368906 229463
rect 380086 229411 380138 229463
rect 538870 229411 538922 229463
rect 230326 229337 230378 229389
rect 269302 229337 269354 229389
rect 273526 229337 273578 229389
rect 347062 229337 347114 229389
rect 357622 229337 357674 229389
rect 522166 229337 522218 229389
rect 233494 229263 233546 229315
rect 276790 229263 276842 229315
rect 284758 229263 284810 229315
rect 146902 229189 146954 229241
rect 151318 229189 151370 229241
rect 231958 229189 232010 229241
rect 273814 229189 273866 229241
rect 286294 229189 286346 229241
rect 293974 229189 294026 229241
rect 294166 229263 294218 229315
rect 371254 229263 371306 229315
rect 374230 229263 374282 229315
rect 371542 229189 371594 229241
rect 387286 229263 387338 229315
rect 546358 229263 546410 229315
rect 555286 229189 555338 229241
rect 235222 229115 235274 229167
rect 279862 229115 279914 229167
rect 287926 229115 287978 229167
rect 374422 229115 374474 229167
rect 377206 229115 377258 229167
rect 561430 229115 561482 229167
rect 238390 229041 238442 229093
rect 283606 229041 283658 229093
rect 291190 229041 291242 229093
rect 215254 228967 215306 229019
rect 239062 228967 239114 229019
rect 241078 228967 241130 229019
rect 291958 228967 292010 229019
rect 293974 229041 294026 229093
rect 374518 229041 374570 229093
rect 376822 229041 376874 229093
rect 563638 229041 563690 229093
rect 382870 228967 382922 229019
rect 382966 228967 383018 229019
rect 567382 228967 567434 229019
rect 242518 228893 242570 228945
rect 294934 228893 294986 228945
rect 308950 228893 309002 228945
rect 427798 228893 427850 228945
rect 427894 228893 427946 228945
rect 547894 228893 547946 228945
rect 239734 228819 239786 228871
rect 288886 228819 288938 228871
rect 241654 228745 241706 228797
rect 231862 228671 231914 228723
rect 272278 228671 272330 228723
rect 230614 228597 230666 228649
rect 270742 228597 270794 228649
rect 282166 228671 282218 228723
rect 294166 228819 294218 228871
rect 310678 228819 310730 228871
rect 430870 228819 430922 228871
rect 432022 228819 432074 228871
rect 529750 228819 529802 228871
rect 304438 228745 304490 228797
rect 418774 228745 418826 228797
rect 289366 228671 289418 228723
rect 289750 228597 289802 228649
rect 293878 228597 293930 228649
rect 295798 228597 295850 228649
rect 306166 228671 306218 228723
rect 421846 228671 421898 228723
rect 380086 228597 380138 228649
rect 407350 228597 407402 228649
rect 517654 228597 517706 228649
rect 190198 228523 190250 228575
rect 192310 228523 192362 228575
rect 228790 228523 228842 228575
rect 266230 228523 266282 228575
rect 266326 228523 266378 228575
rect 301750 228523 301802 228575
rect 303478 228523 303530 228575
rect 413494 228523 413546 228575
rect 455062 228523 455114 228575
rect 456502 228523 456554 228575
rect 535798 228523 535850 228575
rect 538006 228523 538058 228575
rect 544342 228523 544394 228575
rect 547126 228523 547178 228575
rect 556150 228523 556202 228575
rect 558454 228523 558506 228575
rect 224374 228449 224426 228501
rect 258742 228449 258794 228501
rect 270838 228449 270890 228501
rect 313846 228449 313898 228501
rect 317878 228449 317930 228501
rect 403702 228449 403754 228501
rect 405334 228449 405386 228501
rect 502582 228449 502634 228501
rect 264886 228375 264938 228427
rect 295702 228375 295754 228427
rect 295798 228375 295850 228427
rect 382966 228375 383018 228427
rect 391702 228375 391754 228427
rect 476950 228375 477002 228427
rect 535798 228375 535850 228427
rect 537910 228375 537962 228427
rect 267958 228301 268010 228353
rect 307702 228301 307754 228353
rect 311158 228301 311210 228353
rect 392374 228301 392426 228353
rect 392470 228301 392522 228353
rect 461878 228301 461930 228353
rect 261142 228227 261194 228279
rect 292630 228227 292682 228279
rect 311062 228227 311114 228279
rect 383254 228227 383306 228279
rect 394678 228227 394730 228279
rect 437686 228227 437738 228279
rect 269110 228153 269162 228205
rect 322966 228153 323018 228205
rect 344086 228153 344138 228205
rect 412726 228153 412778 228205
rect 250582 228079 250634 228131
rect 277558 228079 277610 228131
rect 290998 228079 291050 228131
rect 341014 228079 341066 228131
rect 341206 228079 341258 228131
rect 398326 228079 398378 228131
rect 260950 228005 261002 228057
rect 286678 228005 286730 228057
rect 305110 228005 305162 228057
rect 310102 228005 310154 228057
rect 310198 228005 310250 228057
rect 258934 227931 258986 227983
rect 280630 227931 280682 227983
rect 293782 227931 293834 227983
rect 343990 227931 344042 227983
rect 357526 228005 357578 228057
rect 359926 228005 359978 228057
rect 368950 228005 369002 228057
rect 370486 228005 370538 228057
rect 370582 228005 370634 228057
rect 425590 228005 425642 228057
rect 359158 227931 359210 227983
rect 302134 227857 302186 227909
rect 350038 227857 350090 227909
rect 250198 227783 250250 227835
rect 310006 227783 310058 227835
rect 310102 227783 310154 227835
rect 353110 227783 353162 227835
rect 281206 227709 281258 227761
rect 325846 227709 325898 227761
rect 279286 227635 279338 227687
rect 319894 227635 319946 227687
rect 321238 227635 321290 227687
rect 451990 227635 452042 227687
rect 149398 227561 149450 227613
rect 174262 227561 174314 227613
rect 288022 227561 288074 227613
rect 328918 227561 328970 227613
rect 387766 227561 387818 227613
rect 396406 227561 396458 227613
rect 423286 227561 423338 227613
rect 433174 227561 433226 227613
rect 187126 227487 187178 227539
rect 190774 227487 190826 227539
rect 217462 227487 217514 227539
rect 241270 227487 241322 227539
rect 244726 227487 244778 227539
rect 254902 227487 254954 227539
rect 215734 227413 215786 227465
rect 238390 227413 238442 227465
rect 217078 227339 217130 227391
rect 243574 227339 243626 227391
rect 249334 227339 249386 227391
rect 306262 227487 306314 227539
rect 311350 227487 311402 227539
rect 375766 227487 375818 227539
rect 388918 227487 388970 227539
rect 586390 227487 586442 227539
rect 591478 227487 591530 227539
rect 594646 227487 594698 227539
rect 606262 227487 606314 227539
rect 256246 227413 256298 227465
rect 315382 227413 315434 227465
rect 318454 227413 318506 227465
rect 381814 227413 381866 227465
rect 388534 227413 388586 227465
rect 585622 227413 585674 227465
rect 587638 227413 587690 227465
rect 600790 227413 600842 227465
rect 629302 227487 629354 227539
rect 634006 227487 634058 227539
rect 639190 227413 639242 227465
rect 278038 227339 278090 227391
rect 279286 227339 279338 227391
rect 311254 227339 311306 227391
rect 384022 227339 384074 227391
rect 390454 227339 390506 227391
rect 589366 227339 589418 227391
rect 590422 227339 590474 227391
rect 627862 227339 627914 227391
rect 219478 227265 219530 227317
rect 245878 227265 245930 227317
rect 275062 227265 275114 227317
rect 348598 227265 348650 227317
rect 390070 227265 390122 227317
rect 217846 227191 217898 227243
rect 242902 227191 242954 227243
rect 271990 227191 272042 227243
rect 351574 227191 351626 227243
rect 365590 227191 365642 227243
rect 367126 227191 367178 227243
rect 390838 227191 390890 227243
rect 396406 227265 396458 227317
rect 407446 227265 407498 227317
rect 587446 227265 587498 227317
rect 630166 227265 630218 227317
rect 220342 227117 220394 227169
rect 247414 227117 247466 227169
rect 263830 227117 263882 227169
rect 288118 227117 288170 227169
rect 288982 227117 289034 227169
rect 369622 227117 369674 227169
rect 392662 227117 392714 227169
rect 588598 227191 588650 227243
rect 588886 227191 588938 227243
rect 626422 227191 626474 227243
rect 238774 227043 238826 227095
rect 252118 227043 252170 227095
rect 275254 227043 275306 227095
rect 213046 226969 213098 227021
rect 233782 226969 233834 227021
rect 238102 226969 238154 227021
rect 264022 226969 264074 227021
rect 276694 226969 276746 227021
rect 359830 227043 359882 227095
rect 393142 227043 393194 227095
rect 221686 226895 221738 226947
rect 250390 226895 250442 226947
rect 253558 226895 253610 226947
rect 266998 226895 267050 226947
rect 273430 226895 273482 226947
rect 357622 226969 357674 227021
rect 365686 226969 365738 227021
rect 393814 226969 393866 227021
rect 590134 227117 590186 227169
rect 590902 227117 590954 227169
rect 630934 227117 630986 227169
rect 397654 227043 397706 227095
rect 407350 227043 407402 227095
rect 407446 227043 407498 227095
rect 584086 227043 584138 227095
rect 590518 227043 590570 227095
rect 632374 227043 632426 227095
rect 593974 226969 594026 227021
rect 599158 226969 599210 227021
rect 606358 226969 606410 227021
rect 638518 226969 638570 227021
rect 224854 226821 224906 226873
rect 256438 226821 256490 226873
rect 324118 226821 324170 226873
rect 339478 226821 339530 226873
rect 360598 226895 360650 226947
rect 367030 226895 367082 226947
rect 408214 226895 408266 226947
rect 587350 226895 587402 226947
rect 598486 226895 598538 226947
rect 633142 226895 633194 226947
rect 354550 226821 354602 226873
rect 355894 226821 355946 226873
rect 366838 226821 366890 226873
rect 367126 226821 367178 226873
rect 396118 226821 396170 226873
rect 223318 226747 223370 226799
rect 253462 226747 253514 226799
rect 257110 226747 257162 226799
rect 273238 226747 273290 226799
rect 279766 226747 279818 226799
rect 366742 226747 366794 226799
rect 386614 226747 386666 226799
rect 388726 226747 388778 226799
rect 395542 226747 395594 226799
rect 599158 226821 599210 226873
rect 600406 226821 600458 226873
rect 634678 226821 634730 226873
rect 397462 226747 397514 226799
rect 400630 226747 400682 226799
rect 407350 226747 407402 226799
rect 149398 226673 149450 226725
rect 159766 226673 159818 226725
rect 227926 226673 227978 226725
rect 262486 226673 262538 226725
rect 282550 226673 282602 226725
rect 372694 226673 372746 226725
rect 374614 226673 374666 226725
rect 391510 226673 391562 226725
rect 397174 226673 397226 226725
rect 602998 226673 603050 226725
rect 226582 226599 226634 226651
rect 259414 226599 259466 226651
rect 285718 226599 285770 226651
rect 378742 226599 378794 226651
rect 382966 226599 383018 226651
rect 397654 226599 397706 226651
rect 400822 226599 400874 226651
rect 603382 226747 603434 226799
rect 636886 226747 636938 226799
rect 603286 226673 603338 226725
rect 637750 226673 637802 226725
rect 229558 226525 229610 226577
rect 265558 226525 265610 226577
rect 271030 226525 271082 226577
rect 294262 226525 294314 226577
rect 297334 226525 297386 226577
rect 390070 226525 390122 226577
rect 402358 226525 402410 226577
rect 603670 226599 603722 226651
rect 606166 226599 606218 226651
rect 639958 226599 640010 226651
rect 247702 226451 247754 226503
rect 257974 226451 258026 226503
rect 268150 226451 268202 226503
rect 282070 226451 282122 226503
rect 288502 226451 288554 226503
rect 384790 226451 384842 226503
rect 385750 226451 385802 226503
rect 394774 226451 394826 226503
rect 402646 226451 402698 226503
rect 609814 226525 609866 226577
rect 232534 226377 232586 226429
rect 271606 226377 271658 226429
rect 284662 226377 284714 226429
rect 378070 226377 378122 226429
rect 382678 226377 382730 226429
rect 386998 226377 387050 226429
rect 404950 226377 405002 226429
rect 612790 226451 612842 226503
rect 147190 226303 147242 226355
rect 151222 226303 151274 226355
rect 213814 226303 213866 226355
rect 237526 226303 237578 226355
rect 241750 226303 241802 226355
rect 216406 226229 216458 226281
rect 239830 226229 239882 226281
rect 245014 226229 245066 226281
rect 252118 226303 252170 226355
rect 285142 226303 285194 226355
rect 291574 226303 291626 226355
rect 390838 226303 390890 226355
rect 407734 226303 407786 226355
rect 613558 226377 613610 226429
rect 629206 226377 629258 226429
rect 635446 226377 635498 226429
rect 215638 226155 215690 226207
rect 240598 226155 240650 226207
rect 246550 226155 246602 226207
rect 291190 226229 291242 226281
rect 297622 226229 297674 226281
rect 402838 226229 402890 226281
rect 410422 226229 410474 226281
rect 618070 226303 618122 226355
rect 151126 226081 151178 226133
rect 187126 226081 187178 226133
rect 218326 226081 218378 226133
rect 246646 226081 246698 226133
rect 297238 226155 297290 226207
rect 301270 226155 301322 226207
rect 411286 226155 411338 226207
rect 624118 226229 624170 226281
rect 629398 226155 629450 226207
rect 300214 226081 300266 226133
rect 300694 226081 300746 226133
rect 408982 226081 409034 226133
rect 411670 226081 411722 226133
rect 631702 226081 631754 226133
rect 214582 226007 214634 226059
rect 236854 226007 236906 226059
rect 238966 226007 239018 226059
rect 261046 226007 261098 226059
rect 271798 226007 271850 226059
rect 336406 226007 336458 226059
rect 379990 226007 380042 226059
rect 394582 226007 394634 226059
rect 394678 226007 394730 226059
rect 582646 226007 582698 226059
rect 584566 226007 584618 226059
rect 212374 225933 212426 225985
rect 234550 225933 234602 225985
rect 267766 225933 267818 225985
rect 218806 225859 218858 225911
rect 244342 225859 244394 225911
rect 262006 225859 262058 225911
rect 273046 225859 273098 225911
rect 273238 225933 273290 225985
rect 321334 225933 321386 225985
rect 374326 225933 374378 225985
rect 387766 225933 387818 225985
rect 388150 225933 388202 225985
rect 584854 225933 584906 225985
rect 587062 226007 587114 226059
rect 595414 226007 595466 226059
rect 628630 226007 628682 226059
rect 603478 225933 603530 225985
rect 636214 225933 636266 225985
rect 327382 225859 327434 225911
rect 331414 225859 331466 225911
rect 345526 225859 345578 225911
rect 269014 225785 269066 225837
rect 330454 225785 330506 225837
rect 345718 225785 345770 225837
rect 382678 225859 382730 225911
rect 382870 225859 382922 225911
rect 386422 225859 386474 225911
rect 387382 225859 387434 225911
rect 394678 225859 394730 225911
rect 394774 225859 394826 225911
rect 579574 225859 579626 225911
rect 374422 225785 374474 225837
rect 385558 225785 385610 225837
rect 388822 225785 388874 225837
rect 581110 225785 581162 225837
rect 588406 225785 588458 225837
rect 602230 225785 602282 225837
rect 231094 225711 231146 225763
rect 268534 225711 268586 225763
rect 279190 225711 279242 225763
rect 324406 225711 324458 225763
rect 338902 225711 338954 225763
rect 396886 225711 396938 225763
rect 408886 225711 408938 225763
rect 610486 225711 610538 225763
rect 265078 225637 265130 225689
rect 279094 225637 279146 225689
rect 279286 225637 279338 225689
rect 318358 225637 318410 225689
rect 321718 225637 321770 225689
rect 451222 225637 451274 225689
rect 587254 225637 587306 225689
rect 592342 225637 592394 225689
rect 241846 225563 241898 225615
rect 248854 225563 248906 225615
rect 42166 225415 42218 225467
rect 48022 225415 48074 225467
rect 259030 225415 259082 225467
rect 269974 225415 270026 225467
rect 273622 225415 273674 225467
rect 309334 225563 309386 225615
rect 315766 225563 315818 225615
rect 439126 225563 439178 225615
rect 309910 225489 309962 225541
rect 427030 225489 427082 225541
rect 306646 225415 306698 225467
rect 420982 225415 421034 225467
rect 264694 225341 264746 225393
rect 276118 225341 276170 225393
rect 276214 225341 276266 225393
rect 303190 225341 303242 225393
rect 303862 225341 303914 225393
rect 415030 225341 415082 225393
rect 302230 225267 302282 225319
rect 411958 225267 412010 225319
rect 282358 225193 282410 225245
rect 342550 225193 342602 225245
rect 351382 225193 351434 225245
rect 418006 225193 418058 225245
rect 243958 225119 244010 225171
rect 251926 225119 251978 225171
rect 305014 225119 305066 225171
rect 333526 225119 333578 225171
rect 339094 225119 339146 225171
rect 399958 225119 400010 225171
rect 252694 225045 252746 225097
rect 312310 225045 312362 225097
rect 348694 225045 348746 225097
rect 399094 225045 399146 225097
rect 399382 225045 399434 225097
rect 606742 225119 606794 225171
rect 368854 224971 368906 225023
rect 376438 224971 376490 225023
rect 378646 224971 378698 225023
rect 405142 224971 405194 225023
rect 362806 224897 362858 224949
rect 402166 224897 402218 224949
rect 149398 224823 149450 224875
rect 162742 224823 162794 224875
rect 277942 224823 277994 224875
rect 363670 224823 363722 224875
rect 371542 224823 371594 224875
rect 379510 224823 379562 224875
rect 380086 224823 380138 224875
rect 388630 224823 388682 224875
rect 334102 224749 334154 224801
rect 374326 224749 374378 224801
rect 374518 224749 374570 224801
rect 382582 224749 382634 224801
rect 385846 224749 385898 224801
rect 407446 224823 407498 224875
rect 392278 224749 392330 224801
rect 593110 224749 593162 224801
rect 362422 224675 362474 224727
rect 378646 224675 378698 224727
rect 382774 224675 382826 224727
rect 386326 224675 386378 224727
rect 386422 224675 386474 224727
rect 389302 224675 389354 224727
rect 389494 224675 389546 224727
rect 587158 224675 587210 224727
rect 596086 224675 596138 224727
rect 597718 224675 597770 224727
rect 316342 224601 316394 224653
rect 441430 224601 441482 224653
rect 319414 224527 319466 224579
rect 447478 224527 447530 224579
rect 323254 224453 323306 224505
rect 452758 224453 452810 224505
rect 322294 224379 322346 224431
rect 453430 224379 453482 224431
rect 325270 224305 325322 224357
rect 459574 224305 459626 224357
rect 331510 224231 331562 224283
rect 471574 224231 471626 224283
rect 330742 224157 330794 224209
rect 467830 224157 467882 224209
rect 553270 224157 553322 224209
rect 555382 224157 555434 224209
rect 328246 224083 328298 224135
rect 465622 224083 465674 224135
rect 334486 224009 334538 224061
rect 477622 224009 477674 224061
rect 337174 223935 337226 223987
rect 483766 223935 483818 223987
rect 340438 223861 340490 223913
rect 489718 223861 489770 223913
rect 343606 223787 343658 223839
rect 497302 223787 497354 223839
rect 263542 223713 263594 223765
rect 335734 223713 335786 223765
rect 346582 223713 346634 223765
rect 501814 223713 501866 223765
rect 261910 223639 261962 223691
rect 332662 223639 332714 223691
rect 349558 223639 349610 223691
rect 507862 223639 507914 223691
rect 266422 223565 266474 223617
rect 341782 223565 341834 223617
rect 348118 223565 348170 223617
rect 506326 223565 506378 223617
rect 268054 223491 268106 223543
rect 344854 223491 344906 223543
rect 348022 223491 348074 223543
rect 504790 223491 504842 223543
rect 264598 223417 264650 223469
rect 338710 223417 338762 223469
rect 352534 223417 352586 223469
rect 513910 223417 513962 223469
rect 270934 223343 270986 223395
rect 350806 223343 350858 223395
rect 351094 223343 351146 223395
rect 510838 223343 510890 223395
rect 269398 223269 269450 223321
rect 347734 223269 347786 223321
rect 351190 223269 351242 223321
rect 512374 223269 512426 223321
rect 272566 223195 272618 223247
rect 353878 223195 353930 223247
rect 353974 223195 354026 223247
rect 516982 223195 517034 223247
rect 313366 223121 313418 223173
rect 435382 223121 435434 223173
rect 310294 223047 310346 223099
rect 429334 223047 429386 223099
rect 312598 222973 312650 223025
rect 431542 222973 431594 223025
rect 307222 222899 307274 222951
rect 423286 222899 423338 222951
rect 304246 222825 304298 222877
rect 417238 222825 417290 222877
rect 307990 222751 308042 222803
rect 422518 222751 422570 222803
rect 286198 222677 286250 222729
rect 381046 222677 381098 222729
rect 403030 222677 403082 222729
rect 511606 222677 511658 222729
rect 302806 222603 302858 222655
rect 414262 222603 414314 222655
rect 302038 222529 302090 222581
rect 410518 222529 410570 222581
rect 410614 222529 410666 222581
rect 430102 222529 430154 222581
rect 283030 222455 283082 222507
rect 374998 222455 375050 222507
rect 394870 222455 394922 222507
rect 496534 222455 496586 222507
rect 281590 222381 281642 222433
rect 371926 222381 371978 222433
rect 386134 222381 386186 222433
rect 482902 222381 482954 222433
rect 274102 222307 274154 222359
rect 356854 222307 356906 222359
rect 371638 222307 371690 222359
rect 443734 222307 443786 222359
rect 149398 221863 149450 221915
rect 168406 221863 168458 221915
rect 149494 221789 149546 221841
rect 171382 221789 171434 221841
rect 656182 221789 656234 221841
rect 676246 221789 676298 221841
rect 145750 221715 145802 221767
rect 184342 221715 184394 221767
rect 478102 221715 478154 221767
rect 479974 221715 480026 221767
rect 512758 221715 512810 221767
rect 515398 221715 515450 221767
rect 146902 221419 146954 221471
rect 151414 221419 151466 221471
rect 673846 219495 673898 219547
rect 676054 219495 676106 219547
rect 655990 219199 656042 219251
rect 676246 219199 676298 219251
rect 147670 219051 147722 219103
rect 179926 219051 179978 219103
rect 655798 219051 655850 219103
rect 676150 219051 676202 219103
rect 149398 218977 149450 219029
rect 165622 218977 165674 219029
rect 143062 218829 143114 218881
rect 184342 218829 184394 218881
rect 149494 216091 149546 216143
rect 174358 216091 174410 216143
rect 149398 216017 149450 216069
rect 177142 216017 177194 216069
rect 675094 216017 675146 216069
rect 676054 216017 676106 216069
rect 149398 214389 149450 214441
rect 159958 214389 160010 214441
rect 147094 214019 147146 214071
rect 151702 214019 151754 214071
rect 41782 213279 41834 213331
rect 45430 213279 45482 213331
rect 674710 213279 674762 213331
rect 676246 213279 676298 213331
rect 674806 213205 674858 213257
rect 675958 213205 676010 213257
rect 675286 213131 675338 213183
rect 676054 213131 676106 213183
rect 41590 212909 41642 212961
rect 45334 212909 45386 212961
rect 146902 212835 146954 212887
rect 152086 212835 152138 212887
rect 41782 212169 41834 212221
rect 44950 212169 45002 212221
rect 674518 212095 674570 212147
rect 676054 212095 676106 212147
rect 41782 211725 41834 211777
rect 43222 211725 43274 211777
rect 41590 211429 41642 211481
rect 44854 211429 44906 211481
rect 41782 210689 41834 210741
rect 50614 210689 50666 210741
rect 674614 210393 674666 210445
rect 675958 210393 676010 210445
rect 147478 210319 147530 210371
rect 151606 210319 151658 210371
rect 674902 210319 674954 210371
rect 676246 210319 676298 210371
rect 147382 210245 147434 210297
rect 151798 210245 151850 210297
rect 674998 210245 675050 210297
rect 676054 210245 676106 210297
rect 41782 210171 41834 210223
rect 43318 210171 43370 210223
rect 41590 209949 41642 210001
rect 50422 209949 50474 210001
rect 41590 209357 41642 209409
rect 43510 209357 43562 209409
rect 147190 207877 147242 207929
rect 151510 207877 151562 207929
rect 41782 207507 41834 207559
rect 42934 207507 42986 207559
rect 146902 207359 146954 207411
rect 151894 207359 151946 207411
rect 646774 207359 646826 207411
rect 679798 207359 679850 207411
rect 147286 206101 147338 206153
rect 151990 206101 152042 206153
rect 675766 206101 675818 206153
rect 675094 205657 675146 205709
rect 675478 205657 675530 205709
rect 675766 205583 675818 205635
rect 149398 204473 149450 204525
rect 182998 204473 183050 204525
rect 674806 202031 674858 202083
rect 675190 202031 675242 202083
rect 41590 201735 41642 201787
rect 42550 201735 42602 201787
rect 149398 201735 149450 201787
rect 174454 201735 174506 201787
rect 41974 201661 42026 201713
rect 44758 201661 44810 201713
rect 149494 201661 149546 201713
rect 177238 201661 177290 201713
rect 41878 201587 41930 201639
rect 42742 201587 42794 201639
rect 149302 201587 149354 201639
rect 180118 201587 180170 201639
rect 41590 201513 41642 201565
rect 44566 201513 44618 201565
rect 143062 201513 143114 201565
rect 185974 201513 186026 201565
rect 655606 201513 655658 201565
rect 675094 201513 675146 201565
rect 674710 201291 674762 201343
rect 675382 201291 675434 201343
rect 41590 200921 41642 200973
rect 44662 200921 44714 200973
rect 34486 200403 34538 200455
rect 42646 200403 42698 200455
rect 34102 200329 34154 200381
rect 42838 200329 42890 200381
rect 34198 200255 34250 200307
rect 43030 200255 43082 200307
rect 34294 200181 34346 200233
rect 42358 200181 42410 200233
rect 34390 200107 34442 200159
rect 43126 200107 43178 200159
rect 147478 198775 147530 198827
rect 154198 198775 154250 198827
rect 149398 198701 149450 198753
rect 162838 198701 162890 198753
rect 181366 198553 181418 198605
rect 185974 198553 186026 198605
rect 178294 198479 178346 198531
rect 186070 198479 186122 198531
rect 674518 197147 674570 197199
rect 675190 197147 675242 197199
rect 149398 195963 149450 196015
rect 168598 195963 168650 196015
rect 149494 195889 149546 195941
rect 171574 195889 171626 195941
rect 149398 195815 149450 195867
rect 183094 195815 183146 195867
rect 166966 195741 167018 195793
rect 184534 195741 184586 195793
rect 169846 195667 169898 195719
rect 184438 195667 184490 195719
rect 172726 195593 172778 195645
rect 184342 195593 184394 195645
rect 42262 194779 42314 194831
rect 42934 194779 42986 194831
rect 149398 193151 149450 193203
rect 160054 193151 160106 193203
rect 149494 193003 149546 193055
rect 165814 193003 165866 193055
rect 152374 192929 152426 192981
rect 184630 192929 184682 192981
rect 42358 192855 42410 192907
rect 43126 192855 43178 192907
rect 155446 192855 155498 192907
rect 184534 192855 184586 192907
rect 158134 192781 158186 192833
rect 184342 192781 184394 192833
rect 163894 192707 163946 192759
rect 184438 192707 184490 192759
rect 42646 191597 42698 191649
rect 42934 191597 42986 191649
rect 147382 190191 147434 190243
rect 154294 190191 154346 190243
rect 149398 190117 149450 190169
rect 157078 190117 157130 190169
rect 143926 190043 143978 190095
rect 184534 190043 184586 190095
rect 149686 189969 149738 190021
rect 184342 189969 184394 190021
rect 171478 189895 171530 189947
rect 184438 189895 184490 189947
rect 180022 189821 180074 189873
rect 184342 189821 184394 189873
rect 159862 187157 159914 187209
rect 184438 187157 184490 187209
rect 165718 187083 165770 187135
rect 184534 187083 184586 187135
rect 168502 187009 168554 187061
rect 184342 187009 184394 187061
rect 177046 186935 177098 186987
rect 184630 186935 184682 186987
rect 149398 185751 149450 185803
rect 186070 185751 186122 185803
rect 145654 184271 145706 184323
rect 184342 184271 184394 184323
rect 171286 184197 171338 184249
rect 184438 184197 184490 184249
rect 182902 184123 182954 184175
rect 186742 184123 186794 184175
rect 645142 183087 645194 183139
rect 649366 183087 649418 183139
rect 149494 182939 149546 182991
rect 185974 182939 186026 182991
rect 149302 182865 149354 182917
rect 186166 182865 186218 182917
rect 149398 181459 149450 181511
rect 171478 181459 171530 181511
rect 182806 181385 182858 181437
rect 184630 181385 184682 181437
rect 156886 181311 156938 181363
rect 184342 181311 184394 181363
rect 165526 181237 165578 181289
rect 184438 181237 184490 181289
rect 154006 181163 154058 181215
rect 184534 181163 184586 181215
rect 149590 180053 149642 180105
rect 185302 180053 185354 180105
rect 149206 179979 149258 180031
rect 186454 179979 186506 180031
rect 645142 179387 645194 179439
rect 649462 179387 649514 179439
rect 149398 178721 149450 178773
rect 162934 178721 162986 178773
rect 149494 178647 149546 178699
rect 165718 178647 165770 178699
rect 149302 178573 149354 178625
rect 168502 178573 168554 178625
rect 42166 178499 42218 178551
rect 50326 178499 50378 178551
rect 145366 178499 145418 178551
rect 184438 178499 184490 178551
rect 162646 178425 162698 178477
rect 184534 178425 184586 178477
rect 174166 178351 174218 178403
rect 184342 178351 184394 178403
rect 149398 177241 149450 177293
rect 156886 177241 156938 177293
rect 655702 176131 655754 176183
rect 676150 176131 676202 176183
rect 147766 175983 147818 176035
rect 154006 175983 154058 176035
rect 655510 175983 655562 176035
rect 676246 175983 676298 176035
rect 655414 175835 655466 175887
rect 676342 175835 676394 175887
rect 145558 175613 145610 175665
rect 184438 175613 184490 175665
rect 145462 175539 145514 175591
rect 184342 175539 184394 175591
rect 645142 174873 645194 174925
rect 649558 174873 649610 174925
rect 148822 174281 148874 174333
rect 149686 174281 149738 174333
rect 149206 174207 149258 174259
rect 186262 174207 186314 174259
rect 149398 172801 149450 172853
rect 182806 172801 182858 172853
rect 148342 172727 148394 172779
rect 184630 172727 184682 172779
rect 148726 172653 148778 172705
rect 184438 172653 184490 172705
rect 148534 172579 148586 172631
rect 184342 172579 184394 172631
rect 149014 172505 149066 172557
rect 184534 172505 184586 172557
rect 645142 171025 645194 171077
rect 649654 171025 649706 171077
rect 675286 169915 675338 169967
rect 676054 169915 676106 169967
rect 148246 169841 148298 169893
rect 184438 169841 184490 169893
rect 148822 169767 148874 169819
rect 184630 169767 184682 169819
rect 148630 169693 148682 169745
rect 184342 169693 184394 169745
rect 149110 169619 149162 169671
rect 184534 169619 184586 169671
rect 645142 168213 645194 168265
rect 649846 168213 649898 168265
rect 674998 167103 675050 167155
rect 676246 167103 676298 167155
rect 675190 167029 675242 167081
rect 676054 167029 676106 167081
rect 148438 166955 148490 167007
rect 184342 166955 184394 167007
rect 149686 166881 149738 166933
rect 184438 166881 184490 166933
rect 154102 166807 154154 166859
rect 184534 166807 184586 166859
rect 647062 164291 647114 164343
rect 676246 164291 676298 164343
rect 646966 164217 647018 164269
rect 676150 164217 676202 164269
rect 646870 164143 646922 164195
rect 676054 164143 676106 164195
rect 151318 164069 151370 164121
rect 184534 164069 184586 164121
rect 156982 163995 157034 164047
rect 184342 163995 184394 164047
rect 159766 163921 159818 163973
rect 184438 163921 184490 163973
rect 174262 163847 174314 163899
rect 184342 163847 184394 163899
rect 645142 163329 645194 163381
rect 649942 163329 649994 163381
rect 151222 161183 151274 161235
rect 184438 161183 184490 161235
rect 162742 161109 162794 161161
rect 184534 161109 184586 161161
rect 675670 161109 675722 161161
rect 168406 161035 168458 161087
rect 184630 161035 184682 161087
rect 171382 160961 171434 161013
rect 184342 160961 184394 161013
rect 675670 160591 675722 160643
rect 670390 160443 670442 160495
rect 675382 160443 675434 160495
rect 645142 159703 645194 159755
rect 650038 159703 650090 159755
rect 147094 158445 147146 158497
rect 151318 158445 151370 158497
rect 151414 158371 151466 158423
rect 184342 158371 184394 158423
rect 165622 158297 165674 158349
rect 184438 158297 184490 158349
rect 179926 158223 179978 158275
rect 184534 158223 184586 158275
rect 177142 158149 177194 158201
rect 184630 158149 184682 158201
rect 146902 156151 146954 156203
rect 151222 156151 151274 156203
rect 645142 156003 645194 156055
rect 650134 156003 650186 156055
rect 149686 155633 149738 155685
rect 177046 155633 177098 155685
rect 148822 155559 148874 155611
rect 180022 155559 180074 155611
rect 151702 155485 151754 155537
rect 184534 155485 184586 155537
rect 658006 155485 658058 155537
rect 670390 155485 670442 155537
rect 152086 155411 152138 155463
rect 184630 155411 184682 155463
rect 159958 155337 160010 155389
rect 184438 155337 184490 155389
rect 174358 155263 174410 155315
rect 184342 155263 184394 155315
rect 148822 153191 148874 153243
rect 149494 153191 149546 153243
rect 149494 152747 149546 152799
rect 174166 152747 174218 152799
rect 149302 152673 149354 152725
rect 182902 152673 182954 152725
rect 151894 152599 151946 152651
rect 184534 152599 184586 152651
rect 151798 152525 151850 152577
rect 184342 152525 184394 152577
rect 645142 152525 645194 152577
rect 650230 152525 650282 152577
rect 151606 152451 151658 152503
rect 184438 152451 184490 152503
rect 149302 149935 149354 149987
rect 171382 149935 171434 149987
rect 149494 149861 149546 149913
rect 174262 149861 174314 149913
rect 149686 149787 149738 149839
rect 180214 149787 180266 149839
rect 182998 149713 183050 149765
rect 186742 149713 186794 149765
rect 151990 149639 152042 149691
rect 184438 149639 184490 149691
rect 180118 149565 180170 149617
rect 184534 149565 184586 149617
rect 151510 149491 151562 149543
rect 184342 149491 184394 149543
rect 645142 148159 645194 148211
rect 650326 148159 650378 148211
rect 149494 146975 149546 147027
rect 168406 146975 168458 147027
rect 149302 146901 149354 146953
rect 177142 146901 177194 146953
rect 154198 146827 154250 146879
rect 184534 146827 184586 146879
rect 162838 146753 162890 146805
rect 184438 146753 184490 146805
rect 174454 146679 174506 146731
rect 184342 146679 184394 146731
rect 177238 146605 177290 146657
rect 184630 146605 184682 146657
rect 147670 145717 147722 145769
rect 165526 145717 165578 145769
rect 147670 144015 147722 144067
rect 162742 144015 162794 144067
rect 183094 143941 183146 143993
rect 184630 143941 184682 143993
rect 168598 143867 168650 143919
rect 184438 143867 184490 143919
rect 171574 143793 171626 143845
rect 184342 143793 184394 143845
rect 165814 143719 165866 143771
rect 184534 143719 184586 143771
rect 147286 142461 147338 142513
rect 159862 142461 159914 142513
rect 147478 142165 147530 142217
rect 156982 142165 157034 142217
rect 149686 141203 149738 141255
rect 154102 141203 154154 141255
rect 154294 141055 154346 141107
rect 184534 141055 184586 141107
rect 157078 140981 157130 141033
rect 184438 140981 184490 141033
rect 160054 140907 160106 140959
rect 184342 140907 184394 140959
rect 147478 140315 147530 140367
rect 151126 140315 151178 140367
rect 147670 138243 147722 138295
rect 159766 138243 159818 138295
rect 148630 136911 148682 136963
rect 148342 136689 148394 136741
rect 149014 136837 149066 136889
rect 149206 136837 149258 136889
rect 148822 136763 148874 136815
rect 149206 136689 149258 136741
rect 149686 135431 149738 135483
rect 171286 135431 171338 135483
rect 149590 135357 149642 135409
rect 179926 135357 179978 135409
rect 168502 135283 168554 135335
rect 184438 135283 184490 135335
rect 171478 135209 171530 135261
rect 184342 135209 184394 135261
rect 177142 134321 177194 134373
rect 184726 134321 184778 134373
rect 149686 132471 149738 132523
rect 182998 132471 183050 132523
rect 154006 132397 154058 132449
rect 184630 132397 184682 132449
rect 156886 132323 156938 132375
rect 184534 132323 184586 132375
rect 162934 132249 162986 132301
rect 184438 132249 184490 132301
rect 165718 132175 165770 132227
rect 184342 132175 184394 132227
rect 655318 130103 655370 130155
rect 676150 130103 676202 130155
rect 655222 129955 655274 130007
rect 676246 129955 676298 130007
rect 655126 129807 655178 129859
rect 676342 129807 676394 129859
rect 147478 129659 147530 129711
rect 165622 129659 165674 129711
rect 149686 129585 149738 129637
rect 168502 129585 168554 129637
rect 180214 129585 180266 129637
rect 185686 129585 185738 129637
rect 645718 129585 645770 129637
rect 676246 129585 676298 129637
rect 182806 129511 182858 129563
rect 186742 129511 186794 129563
rect 149398 129437 149450 129489
rect 184438 129437 184490 129489
rect 149494 129363 149546 129415
rect 184534 129363 184586 129415
rect 149110 129289 149162 129341
rect 184342 129289 184394 129341
rect 147670 127291 147722 127343
rect 162646 127291 162698 127343
rect 646486 126847 646538 126899
rect 676246 126847 676298 126899
rect 646582 126773 646634 126825
rect 676150 126773 676202 126825
rect 674134 126699 674186 126751
rect 676054 126699 676106 126751
rect 149014 126625 149066 126677
rect 184438 126625 184490 126677
rect 148726 126551 148778 126603
rect 184534 126551 184586 126603
rect 149206 126477 149258 126529
rect 184342 126477 184394 126529
rect 674326 124627 674378 124679
rect 676054 124627 676106 124679
rect 149398 124035 149450 124087
rect 156886 124035 156938 124087
rect 674038 124035 674090 124087
rect 675958 124035 676010 124087
rect 674422 123961 674474 124013
rect 676054 123961 676106 124013
rect 675094 123887 675146 123939
rect 676246 123887 676298 123939
rect 148438 123813 148490 123865
rect 184534 123813 184586 123865
rect 148534 123739 148586 123791
rect 184342 123739 184394 123791
rect 148246 123665 148298 123717
rect 184438 123665 184490 123717
rect 148630 123591 148682 123643
rect 184342 123591 184394 123643
rect 174262 122407 174314 122459
rect 186166 122407 186218 122459
rect 674614 122111 674666 122163
rect 676054 122111 676106 122163
rect 674518 121149 674570 121201
rect 676054 121149 676106 121201
rect 674230 121075 674282 121127
rect 676246 121075 676298 121127
rect 674806 121001 674858 121053
rect 676054 121001 676106 121053
rect 148150 120927 148202 120979
rect 184342 120927 184394 120979
rect 148342 120853 148394 120905
rect 184438 120853 184490 120905
rect 171382 120779 171434 120831
rect 184534 120779 184586 120831
rect 147478 119891 147530 119943
rect 153142 119891 153194 119943
rect 647830 118337 647882 118389
rect 676246 118337 676298 118389
rect 149398 118189 149450 118241
rect 168598 118189 168650 118241
rect 647926 118189 647978 118241
rect 676150 118189 676202 118241
rect 149494 118115 149546 118167
rect 174262 118115 174314 118167
rect 645238 118115 645290 118167
rect 676054 118115 676106 118167
rect 159862 118041 159914 118093
rect 184630 118041 184682 118093
rect 162742 117967 162794 118019
rect 184534 117967 184586 118019
rect 165526 117893 165578 117945
rect 184438 117893 184490 117945
rect 168406 117819 168458 117871
rect 184342 117819 184394 117871
rect 675094 115377 675146 115429
rect 675286 115377 675338 115429
rect 149398 115303 149450 115355
rect 162838 115303 162890 115355
rect 149494 115229 149546 115281
rect 165718 115229 165770 115281
rect 647926 115229 647978 115281
rect 665302 115229 665354 115281
rect 151318 115155 151370 115207
rect 184534 115155 184586 115207
rect 663766 115155 663818 115207
rect 665206 115155 665258 115207
rect 154102 115081 154154 115133
rect 184438 115081 184490 115133
rect 156982 115007 157034 115059
rect 184342 115007 184394 115059
rect 674422 114933 674474 114985
rect 675190 114933 675242 114985
rect 674614 114563 674666 114615
rect 180022 114341 180074 114393
rect 184630 114341 184682 114393
rect 675286 114341 675338 114393
rect 674134 114119 674186 114171
rect 675382 114119 675434 114171
rect 149494 113009 149546 113061
rect 159862 113009 159914 113061
rect 674326 112491 674378 112543
rect 675382 112491 675434 112543
rect 149398 112343 149450 112395
rect 177142 112343 177194 112395
rect 151222 112269 151274 112321
rect 184342 112269 184394 112321
rect 665206 112269 665258 112321
rect 675094 112269 675146 112321
rect 182902 112195 182954 112247
rect 184534 112195 184586 112247
rect 177046 112121 177098 112173
rect 184438 112121 184490 112173
rect 674518 112121 674570 112173
rect 675094 112121 675146 112173
rect 674038 111677 674090 111729
rect 675382 111677 675434 111729
rect 149398 110789 149450 110841
rect 156982 110789 157034 110841
rect 674230 110049 674282 110101
rect 675094 110049 675146 110101
rect 148630 109531 148682 109583
rect 154006 109531 154058 109583
rect 159766 109383 159818 109435
rect 184438 109383 184490 109435
rect 174166 109309 174218 109361
rect 184342 109309 184394 109361
rect 147190 108347 147242 108399
rect 151126 108347 151178 108399
rect 182998 106497 183050 106549
rect 184534 106497 184586 106549
rect 171286 106423 171338 106475
rect 184342 106423 184394 106475
rect 179926 106349 179978 106401
rect 185302 106349 185354 106401
rect 149014 106275 149066 106327
rect 184438 106275 184490 106327
rect 153142 105091 153194 105143
rect 184726 105091 184778 105143
rect 654070 104499 654122 104551
rect 665206 104499 665258 104551
rect 647926 103907 647978 103959
rect 661174 103907 661226 103959
rect 646102 103833 646154 103885
rect 657526 103833 657578 103885
rect 643606 103685 643658 103737
rect 665590 103685 665642 103737
rect 148822 103611 148874 103663
rect 184438 103611 184490 103663
rect 149590 103537 149642 103589
rect 184630 103537 184682 103589
rect 165622 103463 165674 103515
rect 184534 103463 184586 103515
rect 168502 103389 168554 103441
rect 184342 103389 184394 103441
rect 645142 102057 645194 102109
rect 652438 102057 652490 102109
rect 149398 100799 149450 100851
rect 171286 100799 171338 100851
rect 149302 100725 149354 100777
rect 184438 100725 184490 100777
rect 149686 100651 149738 100703
rect 184534 100651 184586 100703
rect 156886 100577 156938 100629
rect 184630 100577 184682 100629
rect 162646 100503 162698 100555
rect 184342 100503 184394 100555
rect 149398 97987 149450 98039
rect 184246 97987 184298 98039
rect 149494 97913 149546 97965
rect 186166 97913 186218 97965
rect 647926 97913 647978 97965
rect 662518 97913 662570 97965
rect 148918 97839 148970 97891
rect 184438 97839 184490 97891
rect 149206 97765 149258 97817
rect 184342 97765 184394 97817
rect 645430 95915 645482 95967
rect 653686 95915 653738 95967
rect 149494 95101 149546 95153
rect 168214 95101 168266 95153
rect 149398 95027 149450 95079
rect 179926 95027 179978 95079
rect 162838 94953 162890 95005
rect 184630 94953 184682 95005
rect 165718 94879 165770 94931
rect 184534 94879 184586 94931
rect 168598 94805 168650 94857
rect 184438 94805 184490 94857
rect 174262 94731 174314 94783
rect 184342 94731 184394 94783
rect 646774 92659 646826 92711
rect 663094 92659 663146 92711
rect 646390 92363 646442 92415
rect 660694 92363 660746 92415
rect 646678 92289 646730 92341
rect 661750 92289 661802 92341
rect 149398 92215 149450 92267
rect 162454 92215 162506 92267
rect 646870 92215 646922 92267
rect 659830 92215 659882 92267
rect 149494 92141 149546 92193
rect 165238 92141 165290 92193
rect 646966 92141 647018 92193
rect 658870 92141 658922 92193
rect 148438 92067 148490 92119
rect 184438 92067 184490 92119
rect 156982 91993 157034 92045
rect 184534 91993 184586 92045
rect 159862 91919 159914 91971
rect 184342 91919 184394 91971
rect 177142 91845 177194 91897
rect 184630 91845 184682 91897
rect 149398 90069 149450 90121
rect 159766 90069 159818 90121
rect 148342 89181 148394 89233
rect 184534 89181 184586 89233
rect 148630 89107 148682 89159
rect 184630 89107 184682 89159
rect 151126 89033 151178 89085
rect 184438 89033 184490 89085
rect 154006 88959 154058 89011
rect 184342 88959 184394 89011
rect 645910 87479 645962 87531
rect 650902 87479 650954 87531
rect 647926 87257 647978 87309
rect 658006 87257 658058 87309
rect 647158 87035 647210 87087
rect 663286 87035 663338 87087
rect 149494 86739 149546 86791
rect 156502 86739 156554 86791
rect 148630 86443 148682 86495
rect 154102 86443 154154 86495
rect 148246 86369 148298 86421
rect 184438 86369 184490 86421
rect 148534 86295 148586 86347
rect 184534 86295 184586 86347
rect 148726 86221 148778 86273
rect 184342 86221 184394 86273
rect 640726 84963 640778 85015
rect 643606 84963 643658 85015
rect 645718 84149 645770 84201
rect 657046 84149 657098 84201
rect 146998 83557 147050 83609
rect 151126 83557 151178 83609
rect 646774 83557 646826 83609
rect 653686 83557 653738 83609
rect 168214 83483 168266 83535
rect 184438 83483 184490 83535
rect 171286 83409 171338 83461
rect 184342 83409 184394 83461
rect 647926 81855 647978 81907
rect 663286 81855 663338 81907
rect 647830 81781 647882 81833
rect 663382 81781 663434 81833
rect 657046 81633 657098 81685
rect 658582 81633 658634 81685
rect 647734 81559 647786 81611
rect 662422 81559 662474 81611
rect 647926 80745 647978 80797
rect 662518 80745 662570 80797
rect 149302 80597 149354 80649
rect 184438 80597 184490 80649
rect 162454 80523 162506 80575
rect 184534 80523 184586 80575
rect 165238 80449 165290 80501
rect 184342 80449 184394 80501
rect 179926 80375 179978 80427
rect 184630 80375 184682 80427
rect 149398 77711 149450 77763
rect 184630 77711 184682 77763
rect 647062 77711 647114 77763
rect 658294 77711 658346 77763
rect 149686 77637 149738 77689
rect 184438 77637 184490 77689
rect 646486 77637 646538 77689
rect 659542 77637 659594 77689
rect 156502 77563 156554 77615
rect 184534 77563 184586 77615
rect 646582 77563 646634 77615
rect 661750 77563 661802 77615
rect 159766 77489 159818 77541
rect 184342 77489 184394 77541
rect 647926 77489 647978 77541
rect 656950 77489 657002 77541
rect 646294 75639 646346 75691
rect 657526 75639 657578 75691
rect 647158 74899 647210 74951
rect 660118 74899 660170 74951
rect 148438 74825 148490 74877
rect 184534 74825 184586 74877
rect 149206 74751 149258 74803
rect 184630 74751 184682 74803
rect 151126 74677 151178 74729
rect 184438 74677 184490 74729
rect 154102 74603 154154 74655
rect 184342 74603 184394 74655
rect 149206 74011 149258 74063
rect 149398 74011 149450 74063
rect 647926 72087 647978 72139
rect 660694 72087 660746 72139
rect 148342 71939 148394 71991
rect 184342 71939 184394 71991
rect 149398 71865 149450 71917
rect 184438 71865 184490 71917
rect 149590 71791 149642 71843
rect 184534 71791 184586 71843
rect 647926 69571 647978 69623
rect 661174 69571 661226 69623
rect 149590 69053 149642 69105
rect 184534 69053 184586 69105
rect 148822 68979 148874 69031
rect 184342 68979 184394 69031
rect 149302 68905 149354 68957
rect 184438 68905 184490 68957
rect 149206 68831 149258 68883
rect 184342 68831 184394 68883
rect 149110 66167 149162 66219
rect 184534 66167 184586 66219
rect 646006 66167 646058 66219
rect 652342 66167 652394 66219
rect 149686 66093 149738 66145
rect 184342 66093 184394 66145
rect 149494 66019 149546 66071
rect 184438 66019 184490 66071
rect 149398 65945 149450 65997
rect 184342 65945 184394 65997
rect 647926 63429 647978 63481
rect 663190 63429 663242 63481
rect 149302 63281 149354 63333
rect 184438 63281 184490 63333
rect 149398 63207 149450 63259
rect 184630 63207 184682 63259
rect 149206 63133 149258 63185
rect 184342 63133 184394 63185
rect 149494 63059 149546 63111
rect 184534 63059 184586 63111
rect 647926 60987 647978 61039
rect 663478 60987 663530 61039
rect 149398 60395 149450 60447
rect 184438 60395 184490 60447
rect 149590 60321 149642 60373
rect 184342 60321 184394 60373
rect 149302 60247 149354 60299
rect 184534 60247 184586 60299
rect 646006 59063 646058 59115
rect 652246 59063 652298 59115
rect 149398 58989 149450 59041
rect 184342 58989 184394 59041
rect 149398 57509 149450 57561
rect 184342 57509 184394 57561
rect 149494 56177 149546 56229
rect 184342 56177 184394 56229
rect 149398 56103 149450 56155
rect 184438 56103 184490 56155
rect 149686 54623 149738 54675
rect 184342 54623 184394 54675
rect 149398 53217 149450 53269
rect 184342 53217 184394 53269
rect 643606 51885 643658 51937
rect 654070 51885 654122 51937
rect 311158 48037 311210 48089
rect 354838 48037 354890 48089
rect 311062 47963 311114 48015
rect 371926 47963 371978 48015
rect 405526 47963 405578 48015
rect 441334 47963 441386 48015
rect 460342 47963 460394 48015
rect 510358 47963 510410 48015
rect 320182 47889 320234 47941
rect 529270 47889 529322 47941
rect 302902 47815 302954 47867
rect 521110 47815 521162 47867
rect 285814 47741 285866 47793
rect 515542 47741 515594 47793
rect 268534 47667 268586 47719
rect 503926 47667 503978 47719
rect 233686 47593 233738 47645
rect 250966 47519 251018 47571
rect 475222 47593 475274 47645
rect 492982 47593 493034 47645
rect 475606 47519 475658 47571
rect 521206 47519 521258 47571
rect 145366 47075 145418 47127
rect 199126 47075 199178 47127
rect 334102 46927 334154 46979
rect 337462 46927 337514 46979
rect 636502 46705 636554 46757
rect 643606 46705 643658 46757
rect 403222 46335 403274 46387
rect 406774 46335 406826 46387
rect 207382 46113 207434 46165
rect 216406 46113 216458 46165
rect 522838 46113 522890 46165
rect 527926 46113 527978 46165
rect 521110 44781 521162 44833
rect 525910 44781 525962 44833
rect 515542 44633 515594 44685
rect 524950 44633 525002 44685
rect 541462 43301 541514 43353
rect 545206 43301 545258 43353
rect 503926 43227 503978 43279
rect 520342 43153 520394 43205
rect 506806 41969 506858 42021
rect 307222 41895 307274 41947
rect 311062 41895 311114 41947
rect 394582 41895 394634 41947
rect 424054 41895 424106 41947
rect 449302 41895 449354 41947
rect 475222 41895 475274 41947
rect 514006 41895 514058 41947
rect 514870 41895 514922 41947
rect 562486 41895 562538 41947
rect 145078 41821 145130 41873
rect 636502 41821 636554 41873
rect 187606 41747 187658 41799
rect 194326 41747 194378 41799
rect 640726 41747 640778 41799
rect 207382 41451 207434 41503
rect 365878 37381 365930 37433
rect 394582 37381 394634 37433
rect 420694 37381 420746 37433
rect 449302 37381 449354 37433
rect 475606 37381 475658 37433
rect 514006 37381 514058 37433
rect 475510 37307 475562 37359
rect 506806 37307 506858 37359
<< metal2 >>
rect 483670 1005205 483722 1005211
rect 483668 1005170 483670 1005179
rect 529846 1005205 529898 1005211
rect 483722 1005170 483724 1005179
rect 535030 1005205 535082 1005211
rect 529846 1005147 529898 1005153
rect 535028 1005170 535030 1005179
rect 561622 1005205 561674 1005211
rect 535082 1005170 535084 1005179
rect 483668 1005105 483724 1005114
rect 529858 999439 529886 1005147
rect 636886 1005205 636938 1005211
rect 561622 1005147 561674 1005153
rect 636884 1005170 636886 1005179
rect 649366 1005205 649418 1005211
rect 636938 1005170 636940 1005179
rect 535028 1005105 535084 1005114
rect 561634 999439 561662 1005147
rect 649366 1005147 649418 1005153
rect 636884 1005105 636940 1005114
rect 529846 999433 529898 999439
rect 529846 999375 529898 999381
rect 561622 999433 561674 999439
rect 561622 999375 561674 999381
rect 571894 999433 571946 999439
rect 571894 999375 571946 999381
rect 532822 999359 532874 999365
rect 532822 999301 532874 999307
rect 532834 997925 532862 999301
rect 571906 998463 571934 999375
rect 649378 998964 649406 1005147
rect 233218 997740 233246 997742
rect 240514 997740 240542 997742
rect 649378 961644 649406 977732
rect 671074 976210 671102 977732
rect 679714 964183 679742 967171
rect 679700 964174 679756 964183
rect 679700 964109 679756 964118
rect 649460 961658 649516 961667
rect 649378 961616 649460 961644
rect 649460 961593 649516 961602
rect 676148 894170 676204 894179
rect 676148 894105 676204 894114
rect 676052 893430 676108 893439
rect 676052 893365 676108 893374
rect 655414 893021 655466 893027
rect 655414 892963 655466 892969
rect 655222 892947 655274 892953
rect 655222 892889 655274 892895
rect 655126 892873 655178 892879
rect 655126 892815 655178 892821
rect 649462 881477 649514 881483
rect 649462 881419 649514 881425
rect 649474 861134 649502 881419
rect 654166 872671 654218 872677
rect 654166 872613 654218 872619
rect 653782 864013 653834 864019
rect 654178 863987 654206 872613
rect 655138 866503 655166 892815
rect 655234 867687 655262 892889
rect 655318 881403 655370 881409
rect 655318 881345 655370 881351
rect 655220 867678 655276 867687
rect 655220 867613 655276 867622
rect 655124 866494 655180 866503
rect 655124 866429 655180 866438
rect 655330 865319 655358 881345
rect 655426 868871 655454 892963
rect 676066 892879 676094 893365
rect 676162 892953 676190 894105
rect 676244 893578 676300 893587
rect 676244 893513 676300 893522
rect 676258 893027 676286 893513
rect 676246 893021 676298 893027
rect 676246 892963 676298 892969
rect 676150 892947 676202 892953
rect 676150 892889 676202 892895
rect 676054 892873 676106 892879
rect 676054 892815 676106 892821
rect 676052 892468 676108 892477
rect 673846 892429 673898 892435
rect 676052 892403 676054 892412
rect 673846 892371 673898 892377
rect 676106 892403 676108 892412
rect 676054 892371 676106 892377
rect 670966 891467 671018 891473
rect 670966 891409 671018 891415
rect 670870 890431 670922 890437
rect 670870 890373 670922 890379
rect 655412 868862 655468 868871
rect 655412 868797 655468 868806
rect 655316 865310 655372 865319
rect 655316 865245 655372 865254
rect 653782 863955 653834 863961
rect 654164 863978 654220 863987
rect 653794 862951 653822 863955
rect 654164 863913 654220 863922
rect 653780 862942 653836 862951
rect 653780 862877 653836 862886
rect 649378 861106 649502 861134
rect 41782 817985 41834 817991
rect 41780 817950 41782 817959
rect 47446 817985 47498 817991
rect 41834 817950 41836 817959
rect 47446 817927 47498 817933
rect 41780 817885 41836 817894
rect 41780 817358 41836 817367
rect 41780 817293 41782 817302
rect 41834 817293 41836 817302
rect 44854 817319 44906 817325
rect 41782 817261 41834 817267
rect 44854 817261 44906 817267
rect 41588 816618 41644 816627
rect 41588 816553 41590 816562
rect 41642 816553 41644 816562
rect 41590 816521 41642 816527
rect 41780 815878 41836 815887
rect 41780 815813 41782 815822
rect 41834 815813 41836 815822
rect 43222 815839 43274 815845
rect 41782 815781 41834 815787
rect 43222 815781 43274 815787
rect 41780 814916 41836 814925
rect 41780 814851 41782 814860
rect 41834 814851 41836 814860
rect 41782 814819 41834 814825
rect 41588 813658 41644 813667
rect 41588 813593 41590 813602
rect 41642 813593 41644 813602
rect 41590 813561 41642 813567
rect 41588 813214 41644 813223
rect 41588 813149 41644 813158
rect 40244 812474 40300 812483
rect 41602 812441 41630 813149
rect 42260 812918 42316 812927
rect 42260 812853 42316 812862
rect 40244 812409 40300 812418
rect 41590 812435 41642 812441
rect 28820 805666 28876 805675
rect 28820 805601 28876 805610
rect 28834 805231 28862 805601
rect 28820 805222 28876 805231
rect 28820 805157 28876 805166
rect 40258 802323 40286 812409
rect 41590 812377 41642 812383
rect 41492 811734 41548 811743
rect 41492 811669 41548 811678
rect 40244 802314 40300 802323
rect 40244 802249 40300 802258
rect 41506 800495 41534 811669
rect 41780 811364 41836 811373
rect 41780 811299 41836 811308
rect 41794 809481 41822 811299
rect 41876 810846 41932 810855
rect 41876 810781 41932 810790
rect 41782 809475 41834 809481
rect 41782 809417 41834 809423
rect 41780 808922 41836 808931
rect 41780 808857 41836 808866
rect 41588 808182 41644 808191
rect 41588 808117 41644 808126
rect 41602 807113 41630 808117
rect 41590 807107 41642 807113
rect 41590 807049 41642 807055
rect 41588 806702 41644 806711
rect 41588 806637 41590 806646
rect 41642 806637 41644 806646
rect 41590 806605 41642 806611
rect 41794 806447 41822 808857
rect 41890 806836 41918 810781
rect 42164 809810 42220 809819
rect 42164 809745 42220 809754
rect 42068 809366 42124 809375
rect 42068 809301 42124 809310
rect 41972 807886 42028 807895
rect 41972 807821 42028 807830
rect 41986 807039 42014 807821
rect 41974 807033 42026 807039
rect 41974 806975 42026 806981
rect 41890 806808 42014 806836
rect 41782 806441 41834 806447
rect 41782 806383 41834 806389
rect 41588 806110 41644 806119
rect 41588 806045 41644 806054
rect 41602 805231 41630 806045
rect 41588 805222 41644 805231
rect 41588 805157 41590 805166
rect 41642 805157 41644 805166
rect 41590 805125 41642 805131
rect 41492 800486 41548 800495
rect 41492 800421 41548 800430
rect 41986 800231 42014 806808
rect 42082 800347 42110 809301
rect 42178 800495 42206 809745
rect 42164 800486 42220 800495
rect 42164 800421 42220 800430
rect 42068 800338 42124 800347
rect 42068 800273 42124 800282
rect 41974 800225 42026 800231
rect 41974 800167 42026 800173
rect 41974 800003 42026 800009
rect 41974 799945 42026 799951
rect 41986 799422 42014 799945
rect 42274 797619 42302 812853
rect 42646 812435 42698 812441
rect 42646 812377 42698 812383
rect 42658 812174 42686 812377
rect 42562 812146 42686 812174
rect 42358 800743 42410 800749
rect 42358 800685 42410 800691
rect 42192 797591 42302 797619
rect 42370 796994 42398 800685
rect 42454 800669 42506 800675
rect 42454 800611 42506 800617
rect 42178 796920 42206 796980
rect 42274 796966 42398 796994
rect 42274 796920 42302 796966
rect 42178 796892 42302 796920
rect 42358 796895 42410 796901
rect 42358 796837 42410 796843
rect 42370 795779 42398 796837
rect 42192 795751 42398 795779
rect 42466 795144 42494 800611
rect 42192 795116 42494 795144
rect 42562 795125 42590 812146
rect 43030 809475 43082 809481
rect 43030 809417 43082 809423
rect 42836 807442 42892 807451
rect 42836 807377 42892 807386
rect 42646 806663 42698 806669
rect 42646 806605 42698 806611
rect 42550 795119 42602 795125
rect 42550 795061 42602 795067
rect 42658 794996 42686 806605
rect 42742 806441 42794 806447
rect 42742 806383 42794 806389
rect 42754 796901 42782 806383
rect 42742 796895 42794 796901
rect 42742 796837 42794 796843
rect 42740 796786 42796 796795
rect 42740 796721 42796 796730
rect 42466 794968 42686 794996
rect 42466 794583 42494 794968
rect 42550 794897 42602 794903
rect 42550 794839 42602 794845
rect 42192 794555 42494 794583
rect 42454 794453 42506 794459
rect 42454 794395 42506 794401
rect 42070 794305 42122 794311
rect 42070 794247 42122 794253
rect 42082 793946 42110 794247
rect 42466 793294 42494 794395
rect 42192 793266 42494 793294
rect 42454 793195 42506 793201
rect 42454 793137 42506 793143
rect 42466 792743 42494 793137
rect 42192 792715 42494 792743
rect 42260 791902 42316 791911
rect 42260 791837 42316 791846
rect 42166 790679 42218 790685
rect 42166 790621 42218 790627
rect 42178 790246 42206 790621
rect 42166 790161 42218 790167
rect 42166 790103 42218 790109
rect 42178 789580 42206 790103
rect 42166 789495 42218 789501
rect 42166 789437 42218 789443
rect 42178 788957 42206 789437
rect 42166 788755 42218 788761
rect 42166 788697 42218 788703
rect 42178 788396 42206 788697
rect 42166 787053 42218 787059
rect 42166 786995 42218 787001
rect 42178 786546 42206 786995
rect 42166 786461 42218 786467
rect 42166 786403 42218 786409
rect 42178 785921 42206 786403
rect 42274 786264 42302 791837
rect 42356 791754 42412 791763
rect 42356 791689 42412 791698
rect 42370 786467 42398 791689
rect 42454 789199 42506 789205
rect 42454 789141 42506 789147
rect 42358 786461 42410 786467
rect 42358 786403 42410 786409
rect 42274 786236 42398 786264
rect 42370 785302 42398 786236
rect 42192 785274 42398 785302
rect 42466 784739 42494 789141
rect 42562 787059 42590 794839
rect 42644 794418 42700 794427
rect 42644 794353 42700 794362
rect 42658 793072 42686 794353
rect 42754 793220 42782 796721
rect 42850 794459 42878 807377
rect 42934 807107 42986 807113
rect 42934 807049 42986 807055
rect 42838 794453 42890 794459
rect 42838 794395 42890 794401
rect 42946 794311 42974 807049
rect 42934 794305 42986 794311
rect 42934 794247 42986 794253
rect 42754 793192 42878 793220
rect 43042 793201 43070 809417
rect 43126 807033 43178 807039
rect 43126 806975 43178 806981
rect 42658 793044 42782 793072
rect 42644 792938 42700 792947
rect 42644 792873 42700 792882
rect 42658 788761 42686 792873
rect 42754 789501 42782 793044
rect 42850 790167 42878 793192
rect 43030 793195 43082 793201
rect 43030 793137 43082 793143
rect 43138 790685 43166 806975
rect 43126 790679 43178 790685
rect 43126 790621 43178 790627
rect 42838 790161 42890 790167
rect 42838 790103 42890 790109
rect 42742 789495 42794 789501
rect 42742 789437 42794 789443
rect 42646 788755 42698 788761
rect 42646 788697 42698 788703
rect 42550 787053 42602 787059
rect 42550 786995 42602 787001
rect 42192 784711 42494 784739
rect 41780 774734 41836 774743
rect 41780 774669 41782 774678
rect 41834 774669 41836 774678
rect 41782 774637 41834 774643
rect 41588 773994 41644 774003
rect 41588 773929 41590 773938
rect 41642 773929 41644 773938
rect 41590 773897 41642 773903
rect 41780 773550 41836 773559
rect 41780 773485 41782 773494
rect 41834 773485 41836 773494
rect 41782 773453 41834 773459
rect 43234 773443 43262 815781
rect 44662 814877 44714 814883
rect 44662 814819 44714 814825
rect 44566 805183 44618 805189
rect 44566 805125 44618 805131
rect 41590 773437 41642 773443
rect 41588 773402 41590 773411
rect 43222 773437 43274 773443
rect 41642 773402 41644 773411
rect 43222 773379 43274 773385
rect 41588 773337 41644 773346
rect 41780 772662 41836 772671
rect 41780 772597 41782 772606
rect 41834 772597 41836 772606
rect 43222 772623 43274 772629
rect 41782 772565 41834 772571
rect 43222 772565 43274 772571
rect 41588 772366 41644 772375
rect 41588 772301 41644 772310
rect 41602 771963 41630 772301
rect 43126 772179 43178 772185
rect 43126 772121 43178 772127
rect 41590 771957 41642 771963
rect 43138 771931 43166 772121
rect 41590 771899 41642 771905
rect 43124 771922 43180 771931
rect 41602 770895 41630 771899
rect 43124 771857 43180 771866
rect 41588 770886 41644 770895
rect 41588 770821 41644 770830
rect 42452 770146 42508 770155
rect 42452 770081 42508 770090
rect 41972 769702 42028 769711
rect 41972 769637 42028 769646
rect 38804 768962 38860 768971
rect 38804 768897 38860 768906
rect 33044 767038 33100 767047
rect 33044 766973 33100 766982
rect 28820 762450 28876 762459
rect 28820 762385 28876 762394
rect 28834 762015 28862 762385
rect 28820 762006 28876 762015
rect 28820 761941 28876 761950
rect 33058 758907 33086 766973
rect 33044 758898 33100 758907
rect 33044 758833 33100 758842
rect 38818 757575 38846 768897
rect 41588 768518 41644 768527
rect 41588 768453 41644 768462
rect 41602 767153 41630 768453
rect 41780 768222 41836 768231
rect 41780 768157 41836 768166
rect 41794 767597 41822 768157
rect 41782 767591 41834 767597
rect 41782 767533 41834 767539
rect 41590 767147 41642 767153
rect 41590 767089 41642 767095
rect 41780 766668 41836 766677
rect 41780 766603 41782 766612
rect 41834 766603 41836 766612
rect 41782 766571 41834 766577
rect 41876 766150 41932 766159
rect 41876 766085 41932 766094
rect 41588 765558 41644 765567
rect 41588 765493 41644 765502
rect 41602 765451 41630 765493
rect 41590 765445 41642 765451
rect 41590 765387 41642 765393
rect 41780 765188 41836 765197
rect 41780 765123 41836 765132
rect 41794 764785 41822 765123
rect 41782 764779 41834 764785
rect 41782 764721 41834 764727
rect 41780 764670 41836 764679
rect 41780 764605 41836 764614
rect 41588 763486 41644 763495
rect 41588 763421 41590 763430
rect 41642 763421 41644 763430
rect 41590 763389 41642 763395
rect 41588 762894 41644 762903
rect 41588 762829 41644 762838
rect 41602 762015 41630 762829
rect 41588 762006 41644 762015
rect 41588 761941 41590 761950
rect 41642 761941 41644 761950
rect 41590 761909 41642 761915
rect 38804 757566 38860 757575
rect 38804 757501 38860 757510
rect 41794 757015 41822 764605
rect 41890 757089 41918 766085
rect 41986 760334 42014 769637
rect 42356 767630 42412 767639
rect 42356 767565 42412 767574
rect 42068 764226 42124 764235
rect 42068 764161 42124 764170
rect 42082 763305 42110 764161
rect 42070 763299 42122 763305
rect 42070 763241 42122 763247
rect 41986 760306 42302 760334
rect 41878 757083 41930 757089
rect 41878 757025 41930 757031
rect 41782 757009 41834 757015
rect 41782 756951 41834 756957
rect 42274 756941 42302 760306
rect 42262 756935 42314 756941
rect 42262 756877 42314 756883
rect 42370 756812 42398 767565
rect 42466 757681 42494 770081
rect 42742 767591 42794 767597
rect 42742 767533 42794 767539
rect 42646 767147 42698 767153
rect 42646 767089 42698 767095
rect 42550 766629 42602 766635
rect 42550 766571 42602 766577
rect 42454 757675 42506 757681
rect 42454 757617 42506 757623
rect 42454 757527 42506 757533
rect 42454 757469 42506 757475
rect 42178 756784 42398 756812
rect 42178 756245 42206 756784
rect 42358 756713 42410 756719
rect 42358 756655 42410 756661
rect 42370 754444 42398 756655
rect 42178 754296 42206 754430
rect 42274 754416 42398 754444
rect 42274 754296 42302 754416
rect 42178 754268 42302 754296
rect 42466 753778 42494 757469
rect 42562 757163 42590 766571
rect 42658 757237 42686 767089
rect 42646 757231 42698 757237
rect 42646 757173 42698 757179
rect 42550 757157 42602 757163
rect 42550 757099 42602 757105
rect 42646 757083 42698 757089
rect 42646 757025 42698 757031
rect 42550 757009 42602 757015
rect 42550 756951 42602 756957
rect 42192 753750 42494 753778
rect 42358 753679 42410 753685
rect 42358 753621 42410 753627
rect 42370 752594 42398 753621
rect 42178 752520 42206 752580
rect 42274 752566 42398 752594
rect 42274 752520 42302 752566
rect 42178 752492 42302 752520
rect 42192 751900 42494 751928
rect 42358 751829 42410 751835
rect 42358 751771 42410 751777
rect 42370 751410 42398 751771
rect 42466 751761 42494 751900
rect 42454 751755 42506 751761
rect 42454 751697 42506 751703
rect 42454 751607 42506 751613
rect 42454 751549 42506 751555
rect 42178 751336 42206 751396
rect 42274 751382 42398 751410
rect 42274 751336 42302 751382
rect 42178 751308 42302 751336
rect 42466 750744 42494 751549
rect 42192 750716 42494 750744
rect 42262 750645 42314 750651
rect 42262 750587 42314 750593
rect 42274 750448 42302 750587
rect 42178 750420 42302 750448
rect 42178 750064 42206 750420
rect 42070 749979 42122 749985
rect 42070 749921 42122 749927
rect 42082 749546 42110 749921
rect 42562 747488 42590 756951
rect 42178 747460 42590 747488
rect 42178 747030 42206 747460
rect 42658 746415 42686 757025
rect 42754 749985 42782 767533
rect 42838 765445 42890 765451
rect 42838 765387 42890 765393
rect 42850 753685 42878 765387
rect 42934 764779 42986 764785
rect 42934 764721 42986 764727
rect 42838 753679 42890 753685
rect 42838 753621 42890 753627
rect 42838 753531 42890 753537
rect 42838 753473 42890 753479
rect 42742 749979 42794 749985
rect 42742 749921 42794 749927
rect 42192 746387 42686 746415
rect 42356 746318 42412 746327
rect 42356 746253 42412 746262
rect 42070 746131 42122 746137
rect 42070 746073 42122 746079
rect 42082 745772 42110 746073
rect 42166 745539 42218 745545
rect 42166 745481 42218 745487
rect 42178 745180 42206 745481
rect 42166 743837 42218 743843
rect 42166 743779 42218 743785
rect 42178 743365 42206 743779
rect 42370 742752 42398 746253
rect 42548 746022 42604 746031
rect 42548 745957 42604 745966
rect 42646 745983 42698 745989
rect 42178 742604 42206 742738
rect 42274 742724 42398 742752
rect 42274 742604 42302 742724
rect 42178 742576 42302 742604
rect 42562 742086 42590 745957
rect 42646 745925 42698 745931
rect 42192 742058 42590 742086
rect 42658 741568 42686 745925
rect 42850 743843 42878 753473
rect 42946 751613 42974 764721
rect 43030 763447 43082 763453
rect 43030 763389 43082 763395
rect 43042 751835 43070 763389
rect 43126 763299 43178 763305
rect 43126 763241 43178 763247
rect 43138 757311 43166 763241
rect 43126 757305 43178 757311
rect 43126 757247 43178 757253
rect 43126 757157 43178 757163
rect 43126 757099 43178 757105
rect 43030 751829 43082 751835
rect 43030 751771 43082 751777
rect 43030 751681 43082 751687
rect 43030 751623 43082 751629
rect 42934 751607 42986 751613
rect 42934 751549 42986 751555
rect 43042 745545 43070 751623
rect 43138 746137 43166 757099
rect 43126 746131 43178 746137
rect 43126 746073 43178 746079
rect 43030 745539 43082 745545
rect 43030 745481 43082 745487
rect 42838 743837 42890 743843
rect 42838 743779 42890 743785
rect 42562 741540 42686 741568
rect 42562 741539 42590 741540
rect 42192 741511 42590 741539
rect 41780 731518 41836 731527
rect 41780 731453 41782 731462
rect 41834 731453 41836 731462
rect 41782 731421 41834 731427
rect 41588 730778 41644 730787
rect 41588 730713 41590 730722
rect 41642 730713 41644 730722
rect 41590 730681 41642 730687
rect 41780 730408 41836 730417
rect 41780 730343 41782 730352
rect 41834 730343 41836 730352
rect 41782 730311 41834 730317
rect 43234 730227 43262 772565
rect 43318 757675 43370 757681
rect 43318 757617 43370 757623
rect 43330 753537 43358 757617
rect 43510 757305 43562 757311
rect 43510 757247 43562 757253
rect 43414 757231 43466 757237
rect 43414 757173 43466 757179
rect 43318 753531 43370 753537
rect 43318 753473 43370 753479
rect 43318 751755 43370 751761
rect 43318 751697 43370 751703
rect 43330 745027 43358 751697
rect 43426 751687 43454 757173
rect 43414 751681 43466 751687
rect 43414 751623 43466 751629
rect 43522 750651 43550 757247
rect 43510 750645 43562 750651
rect 43510 750587 43562 750593
rect 43318 745021 43370 745027
rect 43318 744963 43370 744969
rect 41590 730221 41642 730227
rect 41588 730186 41590 730195
rect 43222 730221 43274 730227
rect 41642 730186 41644 730195
rect 43222 730163 43274 730169
rect 41588 730121 41644 730130
rect 41780 729446 41836 729455
rect 41780 729381 41782 729390
rect 41834 729381 41836 729390
rect 43510 729407 43562 729413
rect 41782 729349 41834 729355
rect 43510 729349 43562 729355
rect 42260 729298 42316 729307
rect 42260 729233 42316 729242
rect 41780 728854 41836 728863
rect 41780 728789 41782 728798
rect 41834 728789 41836 728798
rect 41782 728757 41834 728763
rect 40438 728741 40490 728747
rect 40436 728706 40438 728715
rect 40490 728706 40492 728715
rect 42274 728673 42302 729233
rect 43318 728815 43370 728821
rect 43318 728757 43370 728763
rect 40436 728641 40492 728650
rect 42262 728667 42314 728673
rect 42262 728609 42314 728615
rect 41780 727966 41836 727975
rect 41780 727901 41782 727910
rect 41834 727901 41836 727910
rect 41782 727869 41834 727875
rect 41780 727004 41836 727013
rect 41780 726939 41836 726948
rect 41794 726601 41822 726939
rect 41782 726595 41834 726601
rect 41782 726537 41834 726543
rect 42934 726595 42986 726601
rect 42934 726537 42986 726543
rect 41780 726486 41836 726495
rect 41780 726421 41782 726430
rect 41834 726421 41836 726430
rect 42838 726447 42890 726453
rect 41782 726389 41834 726395
rect 42838 726389 42890 726395
rect 40244 725746 40300 725755
rect 40244 725681 40300 725690
rect 34484 723822 34540 723831
rect 34484 723757 34540 723766
rect 28820 719234 28876 719243
rect 28820 719169 28876 719178
rect 28834 718799 28862 719169
rect 28820 718790 28876 718799
rect 28820 718725 28876 718734
rect 34498 715839 34526 723757
rect 40258 717373 40286 725681
rect 41684 725302 41740 725311
rect 41684 725237 41740 725246
rect 41588 722342 41644 722351
rect 41588 722277 41644 722286
rect 41602 720977 41630 722277
rect 41590 720971 41642 720977
rect 41590 720913 41642 720919
rect 41588 720862 41644 720871
rect 41588 720797 41644 720806
rect 41602 720385 41630 720797
rect 41590 720379 41642 720385
rect 41590 720321 41642 720327
rect 41698 720108 41726 725237
rect 41972 725006 42028 725015
rect 41972 724941 42028 724950
rect 41780 723526 41836 723535
rect 41780 723461 41836 723470
rect 41794 723049 41822 723461
rect 41782 723043 41834 723049
rect 41782 722985 41834 722991
rect 41780 721972 41836 721981
rect 41780 721907 41836 721916
rect 41794 720607 41822 721907
rect 41876 721454 41932 721463
rect 41876 721389 41932 721398
rect 41782 720601 41834 720607
rect 41782 720543 41834 720549
rect 41780 720492 41836 720501
rect 41780 720427 41836 720436
rect 41794 720237 41822 720427
rect 41782 720231 41834 720237
rect 41782 720173 41834 720179
rect 41698 720080 41822 720108
rect 41588 718790 41644 718799
rect 41588 718725 41590 718734
rect 41642 718725 41644 718734
rect 41590 718693 41642 718699
rect 40244 717364 40300 717373
rect 40244 717299 40300 717308
rect 34484 715830 34540 715839
rect 34484 715765 34540 715774
rect 41794 713873 41822 720080
rect 41890 713873 41918 721389
rect 41986 713947 42014 724941
rect 42260 724414 42316 724423
rect 42260 724349 42316 724358
rect 41974 713941 42026 713947
rect 41974 713883 42026 713889
rect 41782 713867 41834 713873
rect 41782 713809 41834 713815
rect 41878 713867 41930 713873
rect 41878 713809 41930 713815
rect 42178 713004 42206 713064
rect 42274 713004 42302 724349
rect 42452 722934 42508 722943
rect 42452 722869 42508 722878
rect 42358 714311 42410 714317
rect 42358 714253 42410 714259
rect 42178 712976 42302 713004
rect 42262 712905 42314 712911
rect 42262 712847 42314 712853
rect 42166 711721 42218 711727
rect 42166 711663 42218 711669
rect 42178 711357 42206 711663
rect 42274 711505 42302 712847
rect 42370 711524 42398 714253
rect 42466 711695 42494 722869
rect 42550 720971 42602 720977
rect 42550 720913 42602 720919
rect 42452 711686 42508 711695
rect 42452 711621 42508 711630
rect 42262 711499 42314 711505
rect 42370 711496 42494 711524
rect 42262 711441 42314 711447
rect 42358 711425 42410 711431
rect 42358 711367 42410 711373
rect 42166 711351 42218 711357
rect 42166 711293 42218 711299
rect 42370 711228 42398 711367
rect 42192 711200 42398 711228
rect 42262 711129 42314 711135
rect 42262 711071 42314 711077
rect 42356 711094 42412 711103
rect 42166 710907 42218 710913
rect 42166 710849 42218 710855
rect 42178 710548 42206 710849
rect 42166 709945 42218 709951
rect 42166 709887 42218 709893
rect 42178 709364 42206 709887
rect 42082 708545 42110 708698
rect 42070 708539 42122 708545
rect 42070 708481 42122 708487
rect 42070 708391 42122 708397
rect 42070 708333 42122 708339
rect 42082 708180 42110 708333
rect 42274 708249 42302 711071
rect 42356 711029 42412 711038
rect 42370 710636 42398 711029
rect 42466 710913 42494 711496
rect 42454 710907 42506 710913
rect 42454 710849 42506 710855
rect 42370 710608 42494 710636
rect 42466 708268 42494 710608
rect 42562 709951 42590 720913
rect 42646 720379 42698 720385
rect 42646 720321 42698 720327
rect 42550 709945 42602 709951
rect 42550 709887 42602 709893
rect 42262 708243 42314 708249
rect 42466 708240 42590 708268
rect 42262 708185 42314 708191
rect 42454 708095 42506 708101
rect 42454 708037 42506 708043
rect 42466 707528 42494 708037
rect 42192 707500 42494 707528
rect 42454 707429 42506 707435
rect 42454 707371 42506 707377
rect 42466 706895 42494 707371
rect 42562 707084 42590 708240
rect 42658 707435 42686 720321
rect 42742 720231 42794 720237
rect 42742 720173 42794 720179
rect 42754 708397 42782 720173
rect 42850 712911 42878 726389
rect 42838 712905 42890 712911
rect 42838 712847 42890 712853
rect 42838 712757 42890 712763
rect 42838 712699 42890 712705
rect 42850 711397 42878 712699
rect 42946 711727 42974 726537
rect 43030 723043 43082 723049
rect 43030 722985 43082 722991
rect 42934 711721 42986 711727
rect 42934 711663 42986 711669
rect 43042 711524 43070 722985
rect 43126 720601 43178 720607
rect 43126 720543 43178 720549
rect 42946 711496 43070 711524
rect 42836 711388 42892 711397
rect 42946 711357 42974 711496
rect 43030 711425 43082 711431
rect 43030 711367 43082 711373
rect 42836 711323 42892 711332
rect 42934 711351 42986 711357
rect 42934 711293 42986 711299
rect 42838 711277 42890 711283
rect 42838 711219 42890 711225
rect 42932 711242 42988 711251
rect 42742 708391 42794 708397
rect 42742 708333 42794 708339
rect 42742 708243 42794 708249
rect 42742 708185 42794 708191
rect 42646 707429 42698 707435
rect 42646 707371 42698 707377
rect 42562 707056 42686 707084
rect 42192 706867 42494 706895
rect 42454 706763 42506 706769
rect 42454 706705 42506 706711
rect 42466 706344 42494 706705
rect 42192 706316 42494 706344
rect 42166 704321 42218 704327
rect 42166 704263 42218 704269
rect 42178 703845 42206 704263
rect 42070 703729 42122 703735
rect 42070 703671 42122 703677
rect 42082 703222 42110 703671
rect 42658 702995 42686 707056
rect 42262 702989 42314 702995
rect 42646 702989 42698 702995
rect 42262 702931 42314 702937
rect 42356 702954 42412 702963
rect 42070 702915 42122 702921
rect 42070 702857 42122 702863
rect 42082 702556 42110 702857
rect 42274 702019 42302 702931
rect 42646 702931 42698 702937
rect 42754 702921 42782 708185
rect 42356 702889 42412 702898
rect 42742 702915 42794 702921
rect 42192 701991 42302 702019
rect 42070 700621 42122 700627
rect 42070 700563 42122 700569
rect 42082 700188 42110 700563
rect 42166 699955 42218 699961
rect 42166 699897 42218 699903
rect 42178 699522 42206 699897
rect 42178 698916 42302 698944
rect 42178 698856 42206 698916
rect 42274 698870 42302 698916
rect 42370 698870 42398 702889
rect 42742 702857 42794 702863
rect 42548 702806 42604 702815
rect 42454 702767 42506 702773
rect 42548 702741 42604 702750
rect 42454 702709 42506 702715
rect 42274 698842 42398 698870
rect 42466 698352 42494 702709
rect 42562 699961 42590 702741
rect 42850 700627 42878 711219
rect 42932 711177 42988 711186
rect 42946 703735 42974 711177
rect 43042 706769 43070 711367
rect 43138 708101 43166 720543
rect 43222 713941 43274 713947
rect 43222 713883 43274 713889
rect 43234 711653 43262 713883
rect 43222 711647 43274 711653
rect 43222 711589 43274 711595
rect 43330 711524 43358 728757
rect 43414 727927 43466 727933
rect 43414 727869 43466 727875
rect 43234 711496 43358 711524
rect 43126 708095 43178 708101
rect 43126 708037 43178 708043
rect 43126 707947 43178 707953
rect 43126 707889 43178 707895
rect 43030 706763 43082 706769
rect 43030 706705 43082 706711
rect 43138 704327 43166 707889
rect 43126 704321 43178 704327
rect 43126 704263 43178 704269
rect 42934 703729 42986 703735
rect 42934 703671 42986 703677
rect 42838 700621 42890 700627
rect 42838 700563 42890 700569
rect 42550 699955 42602 699961
rect 42550 699897 42602 699903
rect 42192 698324 42494 698352
rect 41780 688302 41836 688311
rect 41780 688237 41782 688246
rect 41834 688237 41836 688246
rect 41782 688205 41834 688211
rect 41588 687562 41644 687571
rect 41588 687497 41590 687506
rect 41642 687497 41644 687506
rect 41590 687465 41642 687471
rect 41780 687266 41836 687275
rect 41780 687201 41782 687210
rect 41834 687201 41836 687210
rect 41782 687169 41834 687175
rect 41590 687005 41642 687011
rect 41588 686970 41590 686979
rect 41642 686970 41644 686979
rect 41588 686905 41644 686914
rect 41588 686082 41644 686091
rect 41588 686017 41590 686026
rect 41642 686017 41644 686026
rect 41590 685985 41642 685991
rect 43234 685383 43262 711496
rect 43318 711425 43370 711431
rect 43318 711367 43370 711373
rect 43330 687011 43358 711367
rect 43318 687005 43370 687011
rect 43318 686947 43370 686953
rect 41782 685377 41834 685383
rect 41780 685342 41782 685351
rect 43222 685377 43274 685383
rect 41834 685342 41836 685351
rect 43222 685319 43274 685325
rect 41780 685277 41836 685286
rect 43426 684199 43454 727869
rect 43522 711431 43550 729349
rect 43606 713867 43658 713873
rect 43606 713809 43658 713815
rect 43510 711425 43562 711431
rect 43510 711367 43562 711373
rect 43510 708539 43562 708545
rect 43510 708481 43562 708487
rect 43522 702699 43550 708481
rect 43618 707953 43646 713809
rect 43606 707947 43658 707953
rect 43606 707889 43658 707895
rect 43510 702693 43562 702699
rect 43510 702635 43562 702641
rect 43510 686043 43562 686049
rect 43510 685985 43562 685991
rect 41782 684193 41834 684199
rect 41780 684158 41782 684167
rect 43414 684193 43466 684199
rect 41834 684158 41836 684167
rect 43414 684135 43466 684141
rect 41780 684093 41836 684102
rect 42068 683862 42124 683871
rect 42068 683797 42124 683806
rect 39860 682530 39916 682539
rect 39860 682465 39916 682474
rect 34484 680606 34540 680615
rect 34484 680541 34540 680550
rect 28820 676018 28876 676027
rect 28820 675953 28876 675962
rect 28834 675583 28862 675953
rect 28820 675574 28876 675583
rect 28820 675509 28876 675518
rect 34498 672925 34526 680541
rect 34484 672916 34540 672925
rect 34484 672851 34540 672860
rect 39874 671143 39902 682465
rect 41780 681790 41836 681799
rect 41780 681725 41836 681734
rect 41794 681683 41822 681725
rect 41782 681677 41834 681683
rect 41782 681619 41834 681625
rect 41780 680310 41836 680319
rect 41780 680245 41836 680254
rect 41794 679981 41822 680245
rect 41782 679975 41834 679981
rect 41782 679917 41834 679923
rect 41782 679753 41834 679759
rect 41780 679718 41782 679727
rect 41834 679718 41836 679727
rect 41780 679653 41836 679662
rect 41588 679126 41644 679135
rect 41588 679061 41644 679070
rect 41602 677317 41630 679061
rect 41780 678830 41836 678839
rect 41780 678765 41836 678774
rect 41794 677909 41822 678765
rect 41972 678238 42028 678247
rect 41972 678173 42028 678182
rect 41782 677903 41834 677909
rect 41782 677845 41834 677851
rect 41780 677794 41836 677803
rect 41780 677729 41836 677738
rect 41794 677465 41822 677729
rect 41782 677459 41834 677465
rect 41782 677401 41834 677407
rect 41590 677311 41642 677317
rect 41590 677253 41642 677259
rect 41780 677276 41836 677285
rect 41780 677211 41836 677220
rect 41794 677095 41822 677211
rect 41782 677089 41834 677095
rect 41782 677031 41834 677037
rect 41780 676758 41836 676767
rect 41780 676693 41836 676702
rect 41794 675805 41822 676693
rect 41780 675796 41836 675805
rect 41780 675731 41782 675740
rect 41834 675731 41836 675740
rect 41782 675699 41834 675705
rect 39860 671134 39916 671143
rect 39860 671069 39916 671078
rect 41986 670699 42014 678173
rect 41972 670690 42028 670699
rect 42082 670676 42110 683797
rect 42548 683270 42604 683279
rect 42548 683205 42604 683214
rect 42164 682234 42220 682243
rect 42164 682169 42220 682178
rect 42178 670805 42206 682169
rect 42356 681198 42412 681207
rect 42356 681133 42412 681142
rect 42166 670799 42218 670805
rect 42166 670741 42218 670747
rect 42082 670648 42302 670676
rect 41972 670625 42028 670634
rect 42274 670509 42302 670648
rect 42262 670503 42314 670509
rect 42262 670445 42314 670451
rect 42370 670380 42398 681133
rect 42454 677607 42506 677613
rect 42454 677549 42506 677555
rect 42466 671291 42494 677549
rect 42452 671282 42508 671291
rect 42452 671217 42508 671226
rect 42454 671095 42506 671101
rect 42454 671037 42506 671043
rect 42178 670352 42398 670380
rect 42178 669848 42206 670352
rect 42262 670281 42314 670287
rect 42262 670223 42314 670229
rect 42358 670281 42410 670287
rect 42358 670223 42410 670229
rect 42166 668579 42218 668585
rect 42166 668521 42218 668527
rect 42178 667998 42206 668521
rect 42166 667913 42218 667919
rect 42166 667855 42218 667861
rect 42178 667361 42206 667855
rect 42166 666729 42218 666735
rect 42166 666671 42218 666677
rect 42178 666148 42206 666671
rect 42178 665329 42206 665521
rect 42166 665323 42218 665329
rect 42166 665265 42218 665271
rect 42166 665175 42218 665181
rect 42166 665117 42218 665123
rect 42178 664964 42206 665117
rect 42166 664879 42218 664885
rect 42166 664821 42218 664827
rect 42178 664298 42206 664821
rect 42070 664213 42122 664219
rect 42070 664155 42122 664161
rect 42082 663706 42110 664155
rect 42166 663399 42218 663405
rect 42166 663341 42218 663347
rect 42178 663114 42206 663341
rect 42070 661105 42122 661111
rect 42070 661047 42122 661053
rect 42082 660672 42110 661047
rect 42070 660439 42122 660445
rect 42070 660381 42122 660387
rect 42082 660006 42110 660381
rect 42166 659921 42218 659927
rect 42166 659863 42218 659869
rect 42178 659340 42206 659863
rect 42070 659107 42122 659113
rect 42070 659049 42122 659055
rect 42082 658822 42110 659049
rect 42274 656986 42302 670223
rect 42370 663405 42398 670223
rect 42466 667919 42494 671037
rect 42562 668585 42590 683205
rect 42646 681677 42698 681683
rect 42646 681619 42698 681625
rect 42658 677188 42686 681619
rect 42742 679975 42794 679981
rect 42742 679917 42794 679923
rect 42754 677484 42782 679917
rect 42838 679753 42890 679759
rect 42838 679695 42890 679701
rect 42850 677613 42878 679695
rect 43126 677903 43178 677909
rect 43126 677845 43178 677851
rect 42838 677607 42890 677613
rect 42838 677549 42890 677555
rect 42754 677456 42974 677484
rect 42838 677311 42890 677317
rect 42838 677253 42890 677259
rect 42658 677160 42782 677188
rect 42646 677089 42698 677095
rect 42646 677031 42698 677037
rect 42550 668579 42602 668585
rect 42550 668521 42602 668527
rect 42548 668470 42604 668479
rect 42548 668405 42604 668414
rect 42454 667913 42506 667919
rect 42454 667855 42506 667861
rect 42452 667730 42508 667739
rect 42452 667665 42508 667674
rect 42358 663399 42410 663405
rect 42358 663341 42410 663347
rect 42466 660445 42494 667665
rect 42562 661111 42590 668405
rect 42658 665181 42686 677031
rect 42754 670953 42782 677160
rect 42742 670947 42794 670953
rect 42742 670889 42794 670895
rect 42742 670799 42794 670805
rect 42742 670741 42794 670747
rect 42646 665175 42698 665181
rect 42646 665117 42698 665123
rect 42550 661105 42602 661111
rect 42550 661047 42602 661053
rect 42548 660922 42604 660931
rect 42548 660857 42604 660866
rect 42454 660439 42506 660445
rect 42454 660381 42506 660387
rect 42454 659551 42506 659557
rect 42454 659493 42506 659499
rect 42356 659442 42412 659451
rect 42356 659377 42412 659386
rect 42192 656958 42302 656986
rect 42166 656739 42218 656745
rect 42166 656681 42218 656687
rect 42178 656306 42206 656681
rect 42370 655691 42398 659377
rect 42192 655663 42398 655691
rect 42466 655136 42494 659493
rect 42562 656745 42590 660857
rect 42754 659534 42782 670741
rect 42850 666735 42878 677253
rect 42838 666729 42890 666735
rect 42838 666671 42890 666677
rect 42946 659927 42974 677456
rect 43030 677459 43082 677465
rect 43030 677401 43082 677407
rect 43042 664219 43070 677401
rect 43138 664885 43166 677845
rect 43126 664879 43178 664885
rect 43126 664821 43178 664827
rect 43030 664213 43082 664219
rect 43030 664155 43082 664161
rect 42934 659921 42986 659927
rect 42934 659863 42986 659869
rect 42658 659506 42782 659534
rect 42658 659113 42686 659506
rect 42646 659107 42698 659113
rect 42646 659049 42698 659055
rect 42550 656739 42602 656745
rect 42550 656681 42602 656687
rect 42192 655108 42494 655136
rect 41588 644938 41644 644947
rect 41588 644873 41590 644882
rect 41642 644873 41644 644882
rect 41590 644841 41642 644847
rect 41492 644790 41548 644799
rect 41492 644725 41548 644734
rect 41506 642537 41534 644725
rect 41588 644346 41644 644355
rect 41588 644281 41590 644290
rect 41642 644281 41644 644290
rect 41590 644249 41642 644255
rect 41780 644050 41836 644059
rect 41780 643985 41782 643994
rect 41834 643985 41836 643994
rect 41782 643953 41834 643959
rect 43522 643795 43550 685985
rect 41590 643789 41642 643795
rect 41588 643754 41590 643763
rect 43510 643789 43562 643795
rect 41642 643754 41644 643763
rect 43510 643731 43562 643737
rect 41588 643689 41644 643698
rect 41588 642866 41644 642875
rect 41588 642801 41590 642810
rect 41642 642801 41644 642810
rect 43414 642827 43466 642833
rect 41590 642769 41642 642775
rect 43414 642769 43466 642775
rect 41494 642531 41546 642537
rect 41494 642473 41546 642479
rect 41506 641247 41534 642473
rect 41588 641386 41644 641395
rect 41588 641321 41590 641330
rect 41642 641321 41644 641330
rect 43318 641347 43370 641353
rect 41590 641289 41642 641295
rect 43318 641289 43370 641295
rect 41492 641238 41548 641247
rect 41492 641173 41548 641182
rect 41780 640646 41836 640655
rect 41780 640581 41782 640590
rect 41834 640581 41836 640590
rect 42838 640607 42890 640613
rect 41782 640549 41834 640555
rect 42838 640549 42890 640555
rect 42164 640054 42220 640063
rect 42164 639989 42220 639998
rect 42178 639374 42206 639989
rect 42850 639374 42878 640549
rect 43330 639374 43358 641289
rect 42178 639346 42302 639374
rect 39860 639314 39916 639323
rect 39860 639249 39916 639258
rect 34484 637390 34540 637399
rect 34484 637325 34540 637334
rect 28820 632802 28876 632811
rect 28820 632737 28876 632746
rect 28834 632367 28862 632737
rect 28820 632358 28876 632367
rect 28820 632293 28876 632302
rect 34498 627927 34526 637325
rect 39874 628075 39902 639249
rect 42068 639166 42124 639175
rect 42068 639101 42124 639110
rect 41780 638574 41836 638583
rect 41780 638509 41836 638518
rect 41794 636765 41822 638509
rect 41876 637982 41932 637991
rect 41876 637917 41932 637926
rect 41782 636759 41834 636765
rect 41782 636701 41834 636707
rect 41588 636354 41644 636363
rect 41588 636289 41644 636298
rect 41602 635433 41630 636289
rect 41780 636132 41836 636141
rect 41780 636067 41782 636076
rect 41834 636067 41836 636076
rect 41782 636035 41834 636041
rect 41590 635427 41642 635433
rect 41590 635369 41642 635375
rect 41588 635318 41644 635327
rect 41588 635253 41644 635262
rect 41602 634545 41630 635253
rect 41684 634874 41740 634883
rect 41684 634809 41740 634818
rect 41590 634539 41642 634545
rect 41590 634481 41642 634487
rect 41588 634430 41644 634439
rect 41588 634365 41644 634374
rect 41602 634249 41630 634365
rect 41590 634243 41642 634249
rect 41590 634185 41642 634191
rect 41698 633953 41726 634809
rect 41686 633947 41738 633953
rect 41686 633889 41738 633895
rect 41780 633542 41836 633551
rect 41780 633477 41836 633486
rect 41794 632589 41822 633477
rect 41780 632580 41836 632589
rect 41780 632515 41782 632524
rect 41834 632515 41836 632524
rect 41782 632483 41834 632489
rect 41890 628644 41918 637917
rect 42082 628773 42110 639101
rect 42164 637094 42220 637103
rect 42164 637029 42220 637038
rect 42178 628847 42206 637029
rect 42166 628841 42218 628847
rect 42166 628783 42218 628789
rect 42274 628792 42302 639346
rect 42658 639346 42878 639374
rect 43234 639346 43358 639374
rect 42550 636093 42602 636099
rect 42550 636035 42602 636041
rect 42356 634134 42412 634143
rect 42356 634069 42412 634078
rect 42370 630734 42398 634069
rect 42370 630706 42494 630734
rect 42070 628767 42122 628773
rect 42274 628764 42398 628792
rect 42070 628709 42122 628715
rect 41890 628616 42302 628644
rect 42166 628175 42218 628181
rect 42166 628117 42218 628123
rect 39860 628066 39916 628075
rect 39860 628001 39916 628010
rect 34484 627918 34540 627927
rect 34484 627853 34540 627862
rect 42178 627441 42206 628117
rect 42166 627435 42218 627441
rect 42166 627377 42218 627383
rect 42274 626646 42302 628616
rect 42192 626618 42302 626646
rect 42262 626547 42314 626553
rect 42262 626489 42314 626495
rect 42166 625363 42218 625369
rect 42166 625305 42218 625311
rect 42178 624782 42206 625305
rect 42166 624697 42218 624703
rect 42166 624639 42218 624645
rect 42178 624161 42206 624639
rect 42166 623513 42218 623519
rect 42166 623455 42218 623461
rect 42178 622965 42206 623455
rect 42178 622113 42206 622340
rect 42166 622107 42218 622113
rect 42166 622049 42218 622055
rect 42070 622033 42122 622039
rect 42070 621975 42122 621981
rect 42082 621748 42110 621975
rect 42274 621891 42302 626489
rect 42370 625443 42398 628764
rect 42466 628033 42494 630706
rect 42454 628027 42506 628033
rect 42454 627969 42506 627975
rect 42454 627879 42506 627885
rect 42454 627821 42506 627827
rect 42358 625437 42410 625443
rect 42358 625379 42410 625385
rect 42358 625289 42410 625295
rect 42358 625231 42410 625237
rect 42370 624204 42398 625231
rect 42466 624703 42494 627821
rect 42454 624697 42506 624703
rect 42454 624639 42506 624645
rect 42370 624176 42494 624204
rect 42262 621885 42314 621891
rect 42262 621827 42314 621833
rect 42466 621762 42494 624176
rect 42562 623519 42590 636035
rect 42658 628181 42686 639346
rect 43030 636759 43082 636765
rect 43030 636701 43082 636707
rect 42838 634539 42890 634545
rect 42838 634481 42890 634487
rect 42742 634243 42794 634249
rect 42742 634185 42794 634191
rect 42754 628940 42782 634185
rect 42850 629088 42878 634481
rect 42934 633947 42986 633953
rect 42934 633889 42986 633895
rect 42946 629217 42974 633889
rect 43042 629236 43070 636701
rect 43126 635427 43178 635433
rect 43126 635369 43178 635375
rect 43138 629365 43166 635369
rect 43126 629359 43178 629365
rect 43126 629301 43178 629307
rect 42934 629211 42986 629217
rect 43042 629208 43166 629236
rect 42934 629153 42986 629159
rect 42850 629060 43070 629088
rect 42754 628912 42974 628940
rect 42838 628841 42890 628847
rect 42838 628783 42890 628789
rect 42742 628767 42794 628773
rect 42742 628709 42794 628715
rect 42646 628175 42698 628181
rect 42646 628117 42698 628123
rect 42646 628027 42698 628033
rect 42646 627969 42698 627975
rect 42550 623513 42602 623519
rect 42550 623455 42602 623461
rect 42658 622039 42686 627969
rect 42646 622033 42698 622039
rect 42646 621975 42698 621981
rect 42646 621885 42698 621891
rect 42646 621827 42698 621833
rect 42466 621734 42590 621762
rect 42454 621663 42506 621669
rect 42454 621605 42506 621611
rect 42358 621589 42410 621595
rect 42358 621531 42410 621537
rect 42370 621139 42398 621531
rect 42192 621111 42398 621139
rect 42466 620504 42494 621605
rect 42192 620476 42494 620504
rect 42454 620405 42506 620411
rect 42454 620347 42506 620353
rect 42466 619943 42494 620347
rect 42192 619915 42494 619943
rect 42562 619320 42590 621734
rect 42274 619292 42590 619320
rect 42274 617470 42302 619292
rect 42192 617442 42302 617470
rect 42262 617371 42314 617377
rect 42262 617313 42314 617319
rect 42274 616804 42302 617313
rect 42192 616776 42302 616804
rect 42166 616705 42218 616711
rect 42166 616647 42218 616653
rect 42178 616157 42206 616647
rect 42262 616631 42314 616637
rect 42262 616573 42314 616579
rect 42274 615620 42302 616573
rect 42658 615768 42686 621827
rect 42754 616637 42782 628709
rect 42850 616711 42878 628783
rect 42946 621669 42974 628912
rect 42934 621663 42986 621669
rect 42934 621605 42986 621611
rect 43042 621595 43070 629060
rect 43030 621589 43082 621595
rect 43030 621531 43082 621537
rect 42934 621515 42986 621521
rect 42934 621457 42986 621463
rect 42946 617377 42974 621457
rect 43138 620411 43166 629208
rect 43126 620405 43178 620411
rect 43126 620347 43178 620353
rect 42934 617371 42986 617377
rect 42934 617313 42986 617319
rect 42838 616705 42890 616711
rect 42838 616647 42890 616653
rect 42742 616631 42794 616637
rect 42742 616573 42794 616579
rect 42836 616522 42892 616531
rect 42836 616457 42892 616466
rect 42740 616374 42796 616383
rect 42740 616309 42796 616318
rect 42192 615592 42302 615620
rect 42562 615740 42686 615768
rect 42562 613844 42590 615740
rect 42274 613816 42590 613844
rect 42274 613770 42302 613816
rect 42192 613742 42302 613770
rect 42754 613135 42782 616309
rect 42192 613107 42782 613135
rect 42850 612863 42878 616457
rect 42934 616409 42986 616415
rect 42934 616351 42986 616357
rect 42070 612857 42122 612863
rect 42070 612799 42122 612805
rect 42838 612857 42890 612863
rect 42838 612799 42890 612805
rect 42082 612498 42110 612799
rect 42946 612216 42974 616351
rect 42178 612188 42974 612216
rect 42178 611906 42206 612188
rect 41684 602166 41740 602175
rect 41684 602101 41740 602110
rect 41588 601722 41644 601731
rect 41588 601657 41590 601666
rect 41642 601657 41644 601666
rect 41590 601625 41642 601631
rect 41698 599099 41726 602101
rect 41780 601426 41836 601435
rect 41780 601361 41782 601370
rect 41834 601361 41836 601370
rect 41782 601329 41834 601335
rect 41780 600834 41836 600843
rect 41780 600769 41782 600778
rect 41834 600769 41836 600778
rect 41782 600737 41834 600743
rect 41782 600425 41834 600431
rect 41780 600390 41782 600399
rect 41834 600390 41836 600399
rect 41780 600325 41836 600334
rect 41780 599872 41836 599881
rect 41780 599807 41782 599816
rect 41834 599807 41836 599816
rect 41782 599775 41834 599781
rect 41780 599354 41836 599363
rect 41780 599289 41782 599298
rect 41834 599289 41836 599298
rect 41782 599257 41834 599263
rect 39862 599093 39914 599099
rect 39862 599035 39914 599041
rect 41686 599093 41738 599099
rect 41686 599035 41738 599041
rect 39874 598771 39902 599035
rect 39860 598762 39916 598771
rect 39860 598697 39916 598706
rect 41780 598392 41836 598401
rect 41780 598327 41782 598336
rect 41834 598327 41836 598336
rect 41782 598295 41834 598301
rect 43234 597915 43262 639346
rect 43318 629211 43370 629217
rect 43318 629153 43370 629159
rect 43330 625295 43358 629153
rect 43318 625289 43370 625295
rect 43318 625231 43370 625237
rect 43426 610574 43454 642769
rect 43510 629359 43562 629365
rect 43510 629301 43562 629307
rect 43522 621521 43550 629301
rect 43510 621515 43562 621521
rect 43510 621457 43562 621463
rect 43330 610546 43454 610574
rect 43330 600431 43358 610546
rect 43318 600425 43370 600431
rect 43318 600367 43370 600373
rect 43606 599833 43658 599839
rect 43606 599775 43658 599781
rect 43414 599315 43466 599321
rect 43414 599257 43466 599263
rect 41782 597909 41834 597915
rect 41780 597874 41782 597883
rect 43222 597909 43274 597915
rect 41834 597874 41836 597883
rect 43222 597851 43274 597857
rect 41780 597809 41836 597818
rect 41876 597430 41932 597439
rect 41876 597365 41932 597374
rect 41588 596690 41644 596699
rect 41588 596625 41590 596634
rect 41642 596625 41644 596634
rect 41590 596593 41642 596599
rect 34388 596098 34444 596107
rect 34388 596033 34444 596042
rect 28820 589586 28876 589595
rect 28820 589521 28876 589530
rect 28834 589151 28862 589521
rect 28820 589142 28876 589151
rect 28820 589077 28876 589086
rect 34402 585985 34430 596033
rect 41780 595950 41836 595959
rect 41780 595885 41836 595894
rect 41588 595210 41644 595219
rect 41588 595145 41644 595154
rect 41602 595103 41630 595145
rect 41590 595097 41642 595103
rect 41590 595039 41642 595045
rect 41794 594955 41822 595885
rect 41782 594949 41834 594955
rect 41782 594891 41834 594897
rect 41780 594840 41836 594849
rect 41780 594775 41836 594784
rect 34484 594174 34540 594183
rect 34484 594109 34540 594118
rect 34498 586281 34526 594109
rect 41588 593730 41644 593739
rect 41588 593665 41590 593674
rect 41642 593665 41644 593674
rect 41590 593633 41642 593639
rect 41684 592250 41740 592259
rect 41684 592185 41686 592194
rect 41738 592185 41740 592194
rect 41686 592153 41738 592159
rect 41588 591214 41644 591223
rect 41588 591149 41644 591158
rect 41602 590737 41630 591149
rect 41590 590731 41642 590737
rect 41590 590673 41642 590679
rect 41588 589142 41644 589151
rect 41588 589077 41644 589086
rect 41602 587555 41630 589077
rect 41590 587549 41642 587555
rect 41590 587491 41642 587497
rect 34484 586272 34540 586281
rect 34484 586207 34540 586216
rect 34388 585976 34444 585985
rect 34388 585911 34444 585920
rect 41794 584225 41822 594775
rect 41890 587111 41918 597365
rect 42742 596651 42794 596657
rect 42742 596593 42794 596599
rect 42068 593360 42124 593369
rect 42068 593295 42124 593304
rect 41972 590918 42028 590927
rect 41972 590853 41974 590862
rect 42026 590853 42028 590862
rect 41974 590821 42026 590827
rect 41878 587105 41930 587111
rect 41878 587047 41930 587053
rect 42082 584225 42110 593295
rect 42260 592990 42316 592999
rect 42260 592925 42316 592934
rect 42166 587623 42218 587629
rect 42166 587565 42218 587571
rect 42178 584244 42206 587565
rect 42274 585113 42302 592925
rect 42646 592211 42698 592217
rect 42646 592153 42698 592159
rect 42356 591806 42412 591815
rect 42356 591741 42412 591750
rect 42262 585107 42314 585113
rect 42262 585049 42314 585055
rect 42370 584965 42398 591741
rect 42550 590731 42602 590737
rect 42550 590673 42602 590679
rect 42454 587475 42506 587481
rect 42454 587417 42506 587423
rect 42358 584959 42410 584965
rect 42358 584901 42410 584907
rect 42466 584836 42494 587417
rect 42562 587204 42590 590673
rect 42658 587352 42686 592153
rect 42754 587481 42782 596593
rect 43234 596213 43262 597851
rect 43222 596207 43274 596213
rect 43222 596149 43274 596155
rect 43126 595097 43178 595103
rect 43126 595039 43178 595045
rect 42934 594949 42986 594955
rect 42934 594891 42986 594897
rect 42838 593691 42890 593697
rect 42838 593633 42890 593639
rect 42850 587481 42878 593633
rect 42946 587523 42974 594891
rect 43030 590879 43082 590885
rect 43030 590821 43082 590827
rect 42932 587514 42988 587523
rect 42742 587475 42794 587481
rect 42742 587417 42794 587423
rect 42838 587475 42890 587481
rect 42932 587449 42988 587458
rect 42838 587417 42890 587423
rect 43042 587352 43070 590821
rect 43138 587629 43166 595039
rect 43126 587623 43178 587629
rect 43126 587565 43178 587571
rect 43318 587475 43370 587481
rect 43318 587417 43370 587423
rect 42658 587324 42974 587352
rect 43042 587324 43166 587352
rect 42562 587176 42878 587204
rect 42742 585847 42794 585853
rect 42742 585789 42794 585795
rect 42550 585107 42602 585113
rect 42550 585049 42602 585055
rect 42370 584808 42494 584836
rect 41782 584219 41834 584225
rect 41782 584161 41834 584167
rect 42070 584219 42122 584225
rect 42178 584216 42302 584244
rect 42070 584161 42122 584167
rect 41782 583997 41834 584003
rect 41782 583939 41834 583945
rect 41794 583445 41822 583939
rect 42274 582301 42302 584216
rect 42262 582295 42314 582301
rect 42262 582237 42314 582243
rect 42370 582172 42398 584808
rect 42454 584737 42506 584743
rect 42454 584679 42506 584685
rect 42178 582144 42398 582172
rect 42178 581605 42206 582144
rect 42358 582073 42410 582079
rect 42358 582015 42410 582021
rect 42370 581117 42398 582015
rect 42358 581111 42410 581117
rect 42358 581053 42410 581059
rect 42466 580988 42494 584679
rect 42192 580960 42494 580988
rect 42358 580741 42410 580747
rect 42358 580683 42410 580689
rect 42370 579933 42398 580683
rect 42562 579952 42590 585049
rect 42646 584219 42698 584225
rect 42646 584161 42698 584167
rect 42358 579927 42410 579933
rect 42358 579869 42410 579875
rect 42466 579924 42590 579952
rect 42466 579804 42494 579924
rect 42178 579656 42206 579790
rect 42274 579776 42494 579804
rect 42550 579853 42602 579859
rect 42550 579795 42602 579801
rect 42274 579656 42302 579776
rect 42178 579628 42302 579656
rect 42192 579110 42494 579138
rect 42466 579045 42494 579110
rect 42454 579039 42506 579045
rect 42454 578981 42506 578987
rect 42358 578965 42410 578971
rect 42358 578907 42410 578913
rect 42262 578595 42314 578601
rect 42192 578555 42262 578583
rect 42262 578537 42314 578543
rect 42370 577954 42398 578907
rect 42178 577880 42206 577940
rect 42274 577926 42398 577954
rect 42274 577880 42302 577926
rect 42178 577852 42302 577880
rect 42262 577781 42314 577787
rect 42262 577723 42314 577729
rect 42274 577288 42302 577723
rect 42192 577260 42302 577288
rect 42562 576770 42590 579795
rect 42658 578472 42686 584161
rect 42754 578601 42782 585789
rect 42742 578595 42794 578601
rect 42742 578537 42794 578543
rect 42658 578444 42782 578472
rect 42178 576696 42206 576756
rect 42274 576742 42590 576770
rect 42274 576696 42302 576742
rect 42178 576668 42302 576696
rect 42454 576671 42506 576677
rect 42454 576613 42506 576619
rect 42466 574254 42494 576613
rect 42192 574226 42494 574254
rect 42754 574180 42782 578444
rect 42850 577787 42878 587176
rect 42946 578971 42974 587324
rect 43138 587204 43166 587324
rect 43138 587176 43262 587204
rect 43126 587105 43178 587111
rect 43126 587047 43178 587053
rect 43030 584959 43082 584965
rect 43030 584901 43082 584907
rect 42934 578965 42986 578971
rect 42934 578907 42986 578913
rect 42934 578817 42986 578823
rect 42934 578759 42986 578765
rect 42838 577781 42890 577787
rect 42838 577723 42890 577729
rect 42836 577302 42892 577311
rect 42836 577237 42892 577246
rect 42178 574152 42782 574180
rect 42178 573574 42206 574152
rect 42260 574046 42316 574055
rect 42260 573981 42316 573990
rect 42070 573267 42122 573273
rect 42070 573209 42122 573215
rect 42082 572982 42110 573209
rect 42166 572675 42218 572681
rect 42166 572617 42218 572623
rect 42178 572390 42206 572617
rect 42070 571047 42122 571053
rect 42070 570989 42122 570995
rect 42082 570540 42110 570989
rect 42274 570254 42302 573981
rect 42548 573898 42604 573907
rect 42548 573833 42604 573842
rect 42454 573193 42506 573199
rect 42454 573135 42506 573141
rect 42358 570455 42410 570461
rect 42358 570397 42410 570403
rect 42082 570226 42302 570254
rect 42082 569948 42110 570226
rect 42370 569296 42398 570397
rect 42192 569268 42398 569296
rect 42466 568739 42494 573135
rect 42562 570461 42590 573833
rect 42850 572681 42878 577237
rect 42946 573273 42974 578759
rect 43042 576677 43070 584901
rect 43030 576671 43082 576677
rect 43030 576613 43082 576619
rect 42934 573267 42986 573273
rect 42934 573209 42986 573215
rect 42838 572675 42890 572681
rect 42838 572617 42890 572623
rect 43138 571053 43166 587047
rect 43234 585853 43262 587176
rect 43222 585847 43274 585853
rect 43222 585789 43274 585795
rect 43330 578823 43358 587417
rect 43318 578817 43370 578823
rect 43318 578759 43370 578765
rect 43126 571047 43178 571053
rect 43126 570989 43178 570995
rect 42550 570455 42602 570461
rect 42550 570397 42602 570403
rect 42192 568711 42494 568739
rect 42358 541595 42410 541601
rect 42358 541537 42410 541543
rect 41794 539867 41822 540245
rect 41780 539858 41836 539867
rect 41780 539793 41836 539802
rect 41794 538091 41822 538424
rect 41780 538082 41836 538091
rect 41780 538017 41836 538026
rect 42370 537772 42398 541537
rect 42454 541521 42506 541527
rect 42454 541463 42506 541469
rect 42192 537744 42398 537772
rect 41794 536315 41822 536574
rect 41780 536306 41836 536315
rect 41780 536241 41836 536250
rect 42466 535922 42494 541463
rect 42192 535894 42494 535922
rect 41794 535131 41822 535390
rect 41780 535122 41836 535131
rect 41780 535057 41836 535066
rect 41794 534243 41822 534724
rect 41780 534234 41836 534243
rect 41780 534169 41836 534178
rect 41794 533947 41822 534058
rect 41780 533938 41836 533947
rect 41780 533873 41836 533882
rect 41890 533059 41918 533540
rect 41876 533050 41932 533059
rect 41876 532985 41932 532994
rect 41794 530839 41822 531024
rect 41780 530830 41836 530839
rect 41780 530765 41836 530774
rect 41794 530099 41822 530401
rect 41780 530090 41836 530099
rect 41780 530025 41836 530034
rect 42550 529977 42602 529983
rect 42550 529919 42602 529925
rect 42178 529359 42206 529766
rect 42164 529350 42220 529359
rect 42164 529285 42220 529294
rect 42192 529191 42302 529219
rect 42178 527287 42206 527365
rect 42164 527278 42220 527287
rect 42164 527213 42220 527222
rect 42274 527139 42302 529191
rect 42260 527130 42316 527139
rect 42260 527065 42316 527074
rect 42192 526718 42494 526746
rect 42192 526052 42302 526080
rect 42070 525759 42122 525765
rect 42070 525701 42122 525707
rect 42082 525548 42110 525701
rect 42274 522287 42302 526052
rect 42466 525932 42494 526718
rect 42370 525904 42494 525932
rect 42262 522281 42314 522287
rect 42262 522223 42314 522229
rect 41479 476049 41488 476109
rect 41548 476093 41557 476109
rect 41857 476093 41863 476105
rect 41548 476065 41863 476093
rect 41548 476049 41557 476065
rect 41857 476053 41863 476065
rect 41915 476053 41921 476105
rect 41502 475531 41511 475591
rect 41571 475575 41580 475591
rect 41850 475587 41902 475593
rect 41571 475547 41850 475575
rect 41571 475531 41580 475547
rect 41850 475529 41902 475535
rect 41098 475009 41158 475018
rect 41098 474940 41158 474949
rect 41114 474285 41142 474940
rect 41460 474569 41469 474629
rect 41529 474613 41538 474629
rect 42041 474625 42093 474631
rect 41529 474585 42041 474613
rect 41529 474569 41538 474585
rect 42041 474567 42093 474573
rect 41114 474257 41822 474285
rect 40340 473850 40396 473859
rect 40340 473785 40396 473794
rect 39764 473258 39820 473267
rect 39764 473193 39820 473202
rect 39668 472370 39724 472379
rect 39668 472305 39724 472314
rect 34484 464378 34540 464387
rect 34484 464313 34540 464322
rect 23060 463786 23116 463795
rect 23060 463721 23116 463730
rect 23074 463351 23102 463721
rect 23060 463342 23116 463351
rect 23060 463277 23116 463286
rect 34498 463161 34526 464313
rect 34486 463155 34538 463161
rect 34486 463097 34538 463103
rect 39682 437853 39710 472305
rect 39670 437847 39722 437853
rect 39670 437789 39722 437795
rect 25846 437773 25898 437779
rect 25846 437715 25898 437721
rect 25858 424991 25886 437715
rect 39778 427687 39806 473193
rect 39766 427681 39818 427687
rect 39766 427623 39818 427629
rect 40354 426915 40382 473785
rect 41794 472411 41822 474257
rect 41782 472405 41834 472411
rect 41782 472347 41834 472353
rect 42260 472222 42316 472231
rect 42260 472157 42316 472166
rect 42274 470011 42302 472157
rect 42260 470002 42316 470011
rect 42260 469937 42316 469946
rect 42370 468679 42398 525904
rect 42562 525765 42590 529919
rect 42550 525759 42602 525765
rect 42550 525701 42602 525707
rect 42454 522281 42506 522287
rect 42454 522223 42506 522229
rect 42466 470603 42494 522223
rect 43426 498254 43454 599257
rect 43510 598353 43562 598359
rect 43510 598295 43562 598301
rect 43234 498226 43454 498254
rect 43234 478151 43262 498226
rect 43522 489614 43550 598295
rect 43330 489586 43550 489614
rect 43212 478142 43268 478151
rect 43212 478077 43268 478086
rect 43124 472222 43180 472231
rect 43330 472208 43358 489586
rect 43618 474631 43646 599775
rect 43606 474625 43658 474631
rect 43606 474567 43658 474573
rect 43180 472180 43358 472208
rect 43124 472157 43180 472166
rect 42452 470594 42508 470603
rect 42452 470529 42508 470538
rect 42356 468670 42412 468679
rect 42356 468605 42412 468614
rect 41780 463638 41836 463647
rect 41780 463573 41782 463582
rect 41834 463573 41836 463582
rect 41782 463541 41834 463547
rect 41794 463161 41822 463541
rect 41782 463155 41834 463161
rect 41782 463097 41834 463103
rect 41588 428534 41644 428543
rect 41588 428469 41590 428478
rect 41642 428469 41644 428478
rect 41590 428437 41642 428443
rect 41780 428164 41836 428173
rect 41780 428099 41782 428108
rect 41834 428099 41836 428108
rect 41782 428067 41834 428073
rect 41590 427681 41642 427687
rect 41590 427623 41642 427629
rect 41780 427646 41836 427655
rect 40340 426906 40396 426915
rect 40340 426841 40396 426850
rect 34292 425870 34348 425879
rect 34292 425805 34348 425814
rect 25844 424982 25900 424991
rect 25844 424917 25900 424926
rect 34306 420847 34334 425805
rect 41602 425435 41630 427623
rect 41780 427581 41782 427590
rect 41834 427581 41836 427590
rect 41782 427549 41834 427555
rect 41780 426610 41836 426619
rect 41780 426545 41782 426554
rect 41834 426545 41836 426554
rect 43222 426571 43274 426577
rect 41782 426513 41834 426519
rect 43222 426513 43274 426519
rect 41588 425426 41644 425435
rect 41588 425361 41644 425370
rect 41602 425023 41630 425361
rect 41590 425017 41642 425023
rect 41590 424959 41642 424965
rect 34484 424834 34540 424843
rect 34484 424769 34540 424778
rect 34388 423502 34444 423511
rect 34388 423437 34444 423446
rect 34292 420838 34348 420847
rect 34292 420773 34348 420782
rect 34402 419214 34430 423437
rect 34498 423363 34526 424769
rect 34484 423354 34540 423363
rect 34484 423289 34540 423298
rect 42260 421578 42316 421587
rect 42260 421513 42316 421522
rect 39956 420394 40012 420403
rect 39956 420329 40012 420338
rect 39860 419950 39916 419959
rect 39860 419885 39916 419894
rect 34402 419186 34526 419214
rect 34498 417771 34526 419186
rect 39874 419029 39902 419885
rect 39970 419103 39998 420329
rect 40148 419506 40204 419515
rect 40148 419441 40204 419450
rect 40162 419177 40190 419441
rect 40150 419171 40202 419177
rect 40150 419113 40202 419119
rect 39958 419097 40010 419103
rect 39958 419039 40010 419045
rect 39862 419023 39914 419029
rect 39862 418965 39914 418971
rect 41588 418914 41644 418923
rect 41588 418849 41644 418858
rect 41602 418141 41630 418849
rect 41780 418618 41836 418627
rect 41780 418553 41836 418562
rect 41590 418135 41642 418141
rect 41590 418077 41642 418083
rect 41588 418026 41644 418035
rect 41588 417961 41644 417970
rect 34486 417765 34538 417771
rect 34486 417707 34538 417713
rect 41602 416513 41630 417961
rect 41794 417253 41822 418553
rect 41782 417247 41834 417253
rect 41782 417189 41834 417195
rect 41780 417138 41836 417147
rect 41780 417073 41836 417082
rect 41590 416507 41642 416513
rect 41590 416449 41642 416455
rect 23060 416398 23116 416407
rect 23060 416333 23116 416342
rect 23074 415963 23102 416333
rect 41794 416185 41822 417073
rect 41780 416176 41836 416185
rect 41780 416111 41782 416120
rect 41834 416111 41836 416120
rect 41782 416079 41834 416085
rect 23060 415954 23116 415963
rect 23060 415889 23116 415898
rect 42274 413156 42302 421513
rect 42454 419171 42506 419177
rect 42454 419113 42506 419119
rect 42358 417765 42410 417771
rect 42358 417707 42410 417713
rect 42178 413128 42302 413156
rect 42178 412624 42206 413128
rect 42370 410819 42398 417707
rect 42192 410791 42398 410819
rect 42178 409752 42206 410182
rect 42178 409724 42398 409752
rect 42166 409505 42218 409511
rect 42166 409447 42218 409453
rect 42178 408965 42206 409447
rect 42082 408031 42110 408332
rect 42370 408272 42398 409724
rect 42466 409511 42494 419113
rect 42934 419097 42986 419103
rect 42934 419039 42986 419045
rect 42742 418135 42794 418141
rect 42742 418077 42794 418083
rect 42548 417730 42604 417739
rect 42548 417665 42604 417674
rect 42454 409505 42506 409511
rect 42454 409447 42506 409453
rect 42274 408244 42398 408272
rect 42166 408099 42218 408105
rect 42166 408041 42218 408047
rect 42070 408025 42122 408031
rect 42070 407967 42122 407973
rect 42178 407769 42206 408041
rect 42070 407507 42122 407513
rect 42070 407449 42122 407455
rect 42082 407148 42110 407449
rect 42166 407063 42218 407069
rect 42166 407005 42218 407011
rect 42178 406482 42206 407005
rect 42274 406107 42302 408244
rect 42358 408173 42410 408179
rect 42358 408115 42410 408121
rect 42262 406101 42314 406107
rect 42068 406066 42124 406075
rect 42262 406043 42314 406049
rect 42068 406001 42124 406010
rect 42082 405929 42110 406001
rect 42370 403462 42398 408115
rect 42562 408105 42590 417665
rect 42646 416507 42698 416513
rect 42646 416449 42698 416455
rect 42550 408099 42602 408105
rect 42550 408041 42602 408047
rect 42454 408025 42506 408031
rect 42454 407967 42506 407973
rect 42192 403434 42398 403462
rect 42166 403215 42218 403221
rect 42166 403157 42218 403163
rect 42178 402782 42206 403157
rect 42466 403073 42494 407967
rect 42658 407069 42686 416449
rect 42754 407513 42782 418077
rect 42838 417247 42890 417253
rect 42838 417189 42890 417195
rect 42850 408179 42878 417189
rect 42838 408173 42890 408179
rect 42838 408115 42890 408121
rect 42742 407507 42794 407513
rect 42742 407449 42794 407455
rect 42646 407063 42698 407069
rect 42646 407005 42698 407011
rect 42454 403067 42506 403073
rect 42454 403009 42506 403015
rect 42946 402171 42974 419039
rect 43030 419023 43082 419029
rect 43030 418965 43082 418971
rect 43042 403221 43070 418965
rect 43030 403215 43082 403221
rect 43030 403157 43082 403163
rect 42192 402143 42974 402171
rect 41780 402070 41836 402079
rect 41780 402005 41836 402014
rect 41794 401598 41822 402005
rect 41780 400146 41836 400155
rect 41780 400081 41836 400090
rect 41794 399748 41822 400081
rect 41780 399554 41836 399563
rect 41780 399489 41836 399498
rect 41794 399121 41822 399489
rect 41780 398814 41836 398823
rect 41780 398749 41836 398758
rect 41794 398490 41822 398749
rect 42082 394563 42110 397898
rect 42070 394557 42122 394563
rect 42070 394499 42122 394505
rect 41780 388140 41836 388149
rect 41780 388075 41836 388084
rect 41794 386095 41822 388075
rect 41780 386086 41836 386095
rect 41780 386021 41836 386030
rect 41590 385973 41642 385979
rect 41588 385938 41590 385947
rect 41642 385938 41644 385947
rect 41588 385873 41644 385882
rect 41588 385346 41644 385355
rect 41588 385281 41590 385290
rect 41642 385281 41644 385290
rect 41590 385249 41642 385255
rect 41590 384789 41642 384795
rect 41588 384754 41590 384763
rect 41642 384754 41644 384763
rect 41588 384689 41644 384698
rect 41588 383866 41644 383875
rect 41588 383801 41590 383810
rect 41642 383801 41644 383810
rect 41590 383769 41642 383775
rect 34484 383274 34540 383283
rect 34484 383209 34540 383218
rect 34498 378843 34526 383209
rect 41794 383135 41822 386021
rect 41876 385050 41932 385059
rect 41876 384985 41878 384994
rect 41930 384985 41932 384994
rect 41878 384953 41930 384959
rect 43234 384795 43262 426513
rect 43222 384789 43274 384795
rect 43222 384731 43274 384737
rect 43318 383827 43370 383833
rect 43318 383769 43370 383775
rect 41876 383274 41932 383283
rect 41876 383209 41932 383218
rect 41780 383126 41836 383135
rect 41780 383061 41836 383070
rect 41588 382386 41644 382395
rect 41588 382321 41590 382330
rect 41642 382321 41644 382330
rect 41590 382289 41642 382295
rect 41890 382025 41918 383209
rect 43222 382347 43274 382353
rect 43222 382289 43274 382295
rect 41876 382016 41932 382025
rect 41876 381951 41932 381960
rect 39956 380906 40012 380915
rect 39956 380841 40012 380850
rect 37364 379278 37420 379287
rect 37364 379213 37420 379222
rect 34484 378834 34540 378843
rect 34484 378769 34540 378778
rect 37378 373917 37406 379213
rect 37366 373911 37418 373917
rect 37366 373853 37418 373859
rect 28820 373802 28876 373811
rect 28820 373737 28876 373746
rect 28834 373367 28862 373737
rect 28820 373358 28876 373367
rect 28820 373293 28876 373302
rect 39970 372511 39998 380841
rect 41780 379574 41836 379583
rect 41780 379509 41782 379518
rect 41834 379509 41836 379518
rect 42934 379535 42986 379541
rect 41782 379477 41834 379483
rect 42934 379477 42986 379483
rect 41588 377354 41644 377363
rect 41588 377289 41590 377298
rect 41642 377289 41644 377298
rect 42838 377315 42890 377321
rect 41590 377257 41642 377263
rect 42838 377257 42890 377263
rect 42452 377058 42508 377067
rect 42452 376993 42508 377002
rect 41492 376318 41548 376327
rect 41492 376253 41548 376262
rect 41506 374361 41534 376253
rect 41780 376022 41836 376031
rect 41780 375957 41836 375966
rect 41684 375430 41740 375439
rect 41684 375365 41740 375374
rect 41588 374838 41644 374847
rect 41588 374773 41644 374782
rect 41494 374355 41546 374361
rect 41494 374297 41546 374303
rect 41602 373473 41630 374773
rect 41590 373467 41642 373473
rect 41590 373409 41642 373415
rect 41588 373358 41644 373367
rect 41588 373293 41590 373302
rect 41642 373293 41644 373302
rect 41590 373261 41642 373267
rect 39958 372505 40010 372511
rect 39958 372447 40010 372453
rect 41698 371993 41726 375365
rect 41794 374065 41822 375957
rect 41782 374059 41834 374065
rect 41782 374001 41834 374007
rect 41782 373911 41834 373917
rect 41782 373853 41834 373859
rect 41686 371987 41738 371993
rect 41686 371929 41738 371935
rect 41794 370217 41822 373853
rect 42262 372505 42314 372511
rect 42262 372447 42314 372453
rect 41782 370211 41834 370217
rect 41782 370153 41834 370159
rect 41782 369989 41834 369995
rect 41782 369931 41834 369937
rect 41794 369445 41822 369931
rect 42178 367572 42206 367632
rect 42274 367572 42302 372447
rect 42178 367544 42302 367572
rect 42178 366591 42206 366966
rect 42466 366832 42494 376993
rect 42742 374355 42794 374361
rect 42742 374297 42794 374303
rect 42550 373467 42602 373473
rect 42550 373409 42602 373415
rect 42370 366804 42494 366832
rect 42166 366585 42218 366591
rect 42166 366527 42218 366533
rect 42370 365796 42398 366804
rect 42454 366585 42506 366591
rect 42454 366527 42506 366533
rect 42178 365648 42206 365782
rect 42274 365768 42398 365796
rect 42274 365648 42302 365768
rect 42178 365620 42302 365648
rect 42192 365102 42398 365130
rect 42262 365031 42314 365037
rect 42262 364973 42314 364979
rect 42274 364583 42302 364973
rect 42192 364555 42302 364583
rect 42262 364513 42314 364519
rect 42262 364455 42314 364461
rect 42274 363946 42302 364455
rect 42192 363918 42302 363946
rect 42166 363847 42218 363853
rect 42166 363789 42218 363795
rect 42178 363266 42206 363789
rect 42262 363773 42314 363779
rect 42262 363715 42314 363721
rect 42070 362959 42122 362965
rect 42070 362901 42122 362907
rect 42082 362748 42110 362901
rect 42274 360246 42302 363715
rect 42192 360218 42302 360246
rect 42370 360005 42398 365102
rect 42466 362891 42494 366527
rect 42562 365037 42590 373409
rect 42646 371987 42698 371993
rect 42646 371929 42698 371935
rect 42550 365031 42602 365037
rect 42550 364973 42602 364979
rect 42658 363853 42686 371929
rect 42754 364519 42782 374297
rect 42742 364513 42794 364519
rect 42742 364455 42794 364461
rect 42646 363847 42698 363853
rect 42646 363789 42698 363795
rect 42454 362885 42506 362891
rect 42454 362827 42506 362833
rect 42358 359999 42410 360005
rect 42358 359941 42410 359947
rect 42850 359615 42878 377257
rect 42946 362965 42974 379477
rect 43030 374059 43082 374065
rect 43030 374001 43082 374007
rect 43042 363779 43070 374001
rect 43030 363773 43082 363779
rect 43030 363715 43082 363721
rect 42934 362959 42986 362965
rect 42934 362901 42986 362907
rect 42192 359587 42878 359615
rect 41780 359298 41836 359307
rect 41780 359233 41836 359242
rect 41794 358974 41822 359233
rect 41780 358854 41836 358863
rect 41780 358789 41836 358798
rect 41794 358382 41822 358789
rect 41780 356930 41836 356939
rect 41780 356865 41836 356874
rect 41794 356565 41822 356865
rect 41780 356486 41836 356495
rect 41780 356421 41836 356430
rect 41794 355940 41822 356421
rect 41780 355598 41836 355607
rect 41780 355533 41836 355542
rect 41794 355274 41822 355533
rect 42178 351347 42206 354725
rect 42166 351341 42218 351347
rect 42166 351283 42218 351289
rect 41684 343166 41740 343175
rect 41684 343101 41740 343110
rect 41588 340650 41644 340659
rect 41588 340585 41590 340594
rect 41642 340585 41644 340594
rect 41590 340553 41642 340559
rect 41698 340067 41726 343101
rect 41780 342870 41836 342879
rect 41780 342805 41782 342814
rect 41834 342805 41836 342814
rect 41782 342773 41834 342779
rect 41780 342352 41836 342361
rect 41780 342287 41782 342296
rect 41834 342287 41836 342296
rect 41782 342255 41834 342261
rect 41780 341834 41836 341843
rect 41780 341769 41782 341778
rect 41834 341769 41836 341778
rect 41782 341737 41834 341743
rect 41782 341425 41834 341431
rect 41780 341390 41782 341399
rect 41834 341390 41836 341399
rect 41780 341325 41836 341334
rect 41780 340354 41836 340363
rect 41780 340289 41782 340298
rect 41834 340289 41836 340298
rect 41782 340257 41834 340263
rect 41684 340058 41740 340067
rect 41684 339993 41740 340002
rect 41588 339170 41644 339179
rect 41588 339105 41590 339114
rect 41642 339105 41644 339114
rect 41590 339073 41642 339079
rect 43124 338874 43180 338883
rect 43234 338860 43262 382289
rect 43330 341431 43358 383769
rect 43318 341425 43370 341431
rect 43318 341367 43370 341373
rect 43510 340611 43562 340617
rect 43510 340553 43562 340559
rect 43414 340315 43466 340321
rect 43414 340257 43466 340263
rect 43318 339131 43370 339137
rect 43318 339073 43370 339079
rect 43180 338832 43262 338860
rect 43124 338809 43180 338818
rect 39764 337690 39820 337699
rect 39764 337625 39820 337634
rect 39778 330701 39806 337625
rect 41588 336210 41644 336219
rect 41588 336145 41644 336154
rect 41602 334253 41630 336145
rect 41780 335766 41836 335775
rect 41780 335701 41836 335710
rect 41590 334247 41642 334253
rect 41590 334189 41642 334195
rect 41492 333102 41548 333111
rect 41492 333037 41548 333046
rect 41396 332658 41452 332667
rect 41396 332593 41452 332602
rect 41410 331071 41438 332593
rect 41506 331145 41534 333037
rect 41684 332214 41740 332223
rect 41684 332149 41740 332158
rect 41588 331622 41644 331631
rect 41588 331557 41644 331566
rect 41494 331139 41546 331145
rect 41494 331081 41546 331087
rect 41398 331065 41450 331071
rect 41398 331007 41450 331013
rect 39766 330695 39818 330701
rect 39766 330637 39818 330643
rect 28820 330586 28876 330595
rect 28820 330521 28876 330530
rect 28834 330151 28862 330521
rect 28820 330142 28876 330151
rect 28820 330077 28876 330086
rect 41602 328629 41630 331557
rect 41590 328623 41642 328629
rect 41590 328565 41642 328571
rect 41698 328555 41726 332149
rect 41686 328549 41738 328555
rect 41686 328491 41738 328497
rect 41794 327075 41822 335701
rect 41876 334286 41932 334295
rect 41876 334221 41932 334230
rect 42934 334247 42986 334253
rect 41890 334179 41918 334221
rect 42934 334189 42986 334195
rect 41878 334173 41930 334179
rect 41878 334115 41930 334121
rect 42452 333842 42508 333851
rect 42452 333777 42508 333786
rect 42262 330695 42314 330701
rect 42262 330637 42314 330643
rect 41876 330438 41932 330447
rect 41876 330373 41878 330382
rect 41930 330373 41932 330382
rect 41878 330341 41930 330347
rect 41782 327069 41834 327075
rect 41782 327011 41834 327017
rect 41782 326773 41834 326779
rect 41782 326715 41834 326721
rect 41794 326266 41822 326715
rect 42274 324430 42302 330637
rect 42192 324402 42302 324430
rect 42082 323375 42110 323750
rect 42466 323616 42494 333777
rect 42742 331139 42794 331145
rect 42742 331081 42794 331087
rect 42550 328623 42602 328629
rect 42550 328565 42602 328571
rect 42370 323588 42494 323616
rect 42070 323369 42122 323375
rect 42070 323311 42122 323317
rect 42370 322580 42398 323588
rect 42454 323369 42506 323375
rect 42454 323311 42506 323317
rect 42192 322552 42398 322580
rect 42178 321960 42302 321988
rect 42178 321900 42206 321960
rect 42274 321914 42302 321960
rect 42274 321886 42398 321914
rect 42262 321815 42314 321821
rect 42262 321757 42314 321763
rect 42274 321396 42302 321757
rect 42192 321368 42302 321396
rect 42262 321297 42314 321303
rect 42262 321239 42314 321245
rect 42166 321075 42218 321081
rect 42166 321017 42218 321023
rect 42178 320716 42206 321017
rect 42274 320095 42302 321239
rect 42192 320067 42302 320095
rect 42262 319965 42314 319971
rect 42262 319907 42314 319913
rect 42274 319546 42302 319907
rect 42192 319518 42302 319546
rect 42370 319546 42398 321886
rect 42466 319675 42494 323311
rect 42562 321821 42590 328565
rect 42646 328549 42698 328555
rect 42646 328491 42698 328497
rect 42550 321815 42602 321821
rect 42550 321757 42602 321763
rect 42658 321303 42686 328491
rect 42646 321297 42698 321303
rect 42646 321239 42698 321245
rect 42754 321081 42782 331081
rect 42838 331065 42890 331071
rect 42838 331007 42890 331013
rect 42742 321075 42794 321081
rect 42742 321017 42794 321023
rect 42454 319669 42506 319675
rect 42454 319611 42506 319617
rect 42370 319518 42590 319546
rect 42454 319447 42506 319453
rect 42454 319389 42506 319395
rect 42466 317059 42494 319389
rect 42192 317031 42494 317059
rect 42454 316931 42506 316937
rect 42454 316873 42506 316879
rect 42466 316438 42494 316873
rect 42562 316789 42590 319518
rect 42850 319453 42878 331007
rect 42946 319971 42974 334189
rect 43030 334173 43082 334179
rect 43030 334115 43082 334121
rect 42934 319965 42986 319971
rect 42934 319907 42986 319913
rect 42838 319447 42890 319453
rect 42838 319389 42890 319395
rect 43042 316937 43070 334115
rect 43030 316931 43082 316937
rect 43030 316873 43082 316879
rect 43330 316814 43358 339073
rect 42550 316783 42602 316789
rect 42550 316725 42602 316731
rect 43234 316786 43358 316814
rect 42178 316364 42206 316424
rect 42274 316410 42494 316438
rect 42274 316364 42302 316410
rect 42178 316336 42302 316364
rect 41780 316230 41836 316239
rect 41780 316165 41836 316174
rect 41794 315758 41822 316165
rect 41780 315490 41836 315499
rect 41780 315425 41836 315434
rect 41794 315205 41822 315425
rect 41780 313714 41836 313723
rect 41780 313649 41836 313658
rect 41794 313390 41822 313649
rect 41780 313270 41836 313279
rect 41780 313205 41836 313214
rect 41794 312724 41822 313205
rect 41780 312382 41836 312391
rect 41780 312317 41836 312326
rect 41794 312058 41822 312317
rect 42178 308131 42206 311540
rect 42166 308125 42218 308131
rect 42166 308067 42218 308073
rect 39766 299689 39818 299695
rect 39766 299631 39818 299637
rect 41780 299654 41836 299663
rect 39668 298766 39724 298775
rect 39668 298701 39724 298710
rect 39682 293775 39710 298701
rect 39778 296555 39806 299631
rect 41780 299589 41782 299598
rect 41834 299589 41836 299598
rect 43126 299615 43178 299621
rect 41782 299557 41834 299563
rect 43126 299557 43178 299563
rect 41780 299210 41836 299219
rect 41780 299145 41782 299154
rect 41834 299145 41836 299154
rect 41782 299113 41834 299119
rect 41782 298209 41834 298215
rect 41780 298174 41782 298183
rect 41834 298174 41836 298183
rect 41780 298109 41836 298118
rect 41780 297656 41836 297665
rect 41780 297591 41782 297600
rect 41834 297591 41836 297600
rect 41782 297559 41834 297565
rect 41780 297138 41836 297147
rect 41780 297073 41782 297082
rect 41834 297073 41836 297082
rect 41782 297041 41834 297047
rect 39958 296729 40010 296735
rect 39958 296671 40010 296677
rect 39764 296546 39820 296555
rect 39764 296481 39820 296490
rect 39970 295963 39998 296671
rect 39956 295954 40012 295963
rect 39956 295889 40012 295898
rect 41588 295954 41644 295963
rect 41588 295889 41590 295898
rect 41642 295889 41644 295898
rect 41590 295857 41642 295863
rect 40244 294474 40300 294483
rect 40244 294409 40300 294418
rect 39670 293769 39722 293775
rect 39670 293711 39722 293717
rect 40258 288003 40286 294409
rect 41588 292994 41644 293003
rect 41588 292929 41644 292938
rect 41602 291481 41630 292929
rect 41780 292624 41836 292633
rect 41780 292559 41836 292568
rect 41590 291475 41642 291481
rect 41590 291417 41642 291423
rect 41590 290957 41642 290963
rect 41588 290922 41590 290931
rect 41642 290922 41644 290931
rect 41588 290857 41644 290866
rect 41492 289442 41548 289451
rect 41492 289377 41548 289386
rect 40246 287997 40298 288003
rect 40246 287939 40298 287945
rect 41506 287929 41534 289377
rect 41588 288998 41644 289007
rect 41588 288933 41644 288942
rect 41494 287923 41546 287929
rect 41494 287865 41546 287871
rect 28820 287370 28876 287379
rect 28820 287305 28876 287314
rect 28834 286935 28862 287305
rect 28820 286926 28876 286935
rect 28820 286861 28876 286870
rect 41602 285265 41630 288933
rect 41590 285259 41642 285265
rect 41590 285201 41642 285207
rect 41794 283859 41822 292559
rect 43138 291629 43166 299557
rect 43234 298141 43262 316786
rect 43426 300953 43454 340257
rect 43414 300947 43466 300953
rect 43414 300889 43466 300895
rect 43426 299695 43454 300889
rect 43414 299689 43466 299695
rect 43414 299631 43466 299637
rect 43522 298215 43550 340553
rect 43510 298209 43562 298215
rect 43510 298151 43562 298157
rect 43222 298135 43274 298141
rect 43222 298077 43274 298083
rect 43234 296735 43262 298077
rect 43414 297617 43466 297623
rect 43414 297559 43466 297565
rect 43318 297099 43370 297105
rect 43318 297041 43370 297047
rect 43222 296729 43274 296735
rect 43222 296671 43274 296677
rect 43222 295915 43274 295921
rect 43222 295857 43274 295863
rect 43126 291623 43178 291629
rect 43126 291565 43178 291571
rect 43126 291475 43178 291481
rect 43126 291417 43178 291423
rect 42934 290957 42986 290963
rect 42934 290899 42986 290905
rect 42356 290774 42412 290783
rect 42356 290709 42412 290718
rect 42260 288702 42316 288711
rect 42260 288637 42316 288646
rect 41876 287222 41932 287231
rect 41876 287157 41878 287166
rect 41930 287157 41932 287166
rect 41878 287125 41930 287131
rect 41782 283853 41834 283859
rect 41782 283795 41834 283801
rect 41782 283557 41834 283563
rect 41782 283499 41834 283505
rect 41794 283050 41822 283499
rect 42166 281781 42218 281787
rect 42166 281723 42218 281729
rect 42178 281200 42206 281723
rect 42082 280159 42110 280534
rect 42070 280153 42122 280159
rect 42070 280095 42122 280101
rect 42166 279931 42218 279937
rect 42166 279873 42218 279879
rect 42178 279350 42206 279873
rect 42178 278531 42206 278721
rect 42166 278525 42218 278531
rect 42166 278467 42218 278473
rect 42274 278180 42302 288637
rect 42370 279937 42398 290709
rect 42548 290182 42604 290191
rect 42548 290117 42604 290126
rect 42454 285259 42506 285265
rect 42454 285201 42506 285207
rect 42358 279931 42410 279937
rect 42358 279873 42410 279879
rect 42192 278152 42302 278180
rect 42166 277859 42218 277865
rect 42166 277801 42218 277807
rect 42178 277500 42206 277801
rect 42466 276922 42494 285201
rect 42562 277865 42590 290117
rect 42646 287997 42698 288003
rect 42646 287939 42698 287945
rect 42658 281787 42686 287939
rect 42742 287923 42794 287929
rect 42742 287865 42794 287871
rect 42646 281781 42698 281787
rect 42646 281723 42698 281729
rect 42550 277859 42602 277865
rect 42550 277801 42602 277807
rect 42178 276848 42206 276908
rect 42274 276894 42494 276922
rect 42274 276848 42302 276894
rect 42754 276848 42782 287865
rect 42838 280153 42890 280159
rect 42838 280095 42890 280101
rect 42178 276820 42302 276848
rect 42358 276823 42410 276829
rect 42358 276765 42410 276771
rect 42466 276820 42782 276848
rect 42370 276330 42398 276765
rect 42192 276302 42398 276330
rect 42466 273859 42494 276820
rect 42550 276749 42602 276755
rect 42550 276691 42602 276697
rect 42192 273831 42494 273859
rect 42562 273222 42590 276691
rect 42850 276459 42878 280095
rect 42946 276755 42974 290899
rect 43030 278525 43082 278531
rect 43030 278467 43082 278473
rect 42934 276749 42986 276755
rect 42934 276691 42986 276697
rect 42838 276453 42890 276459
rect 42838 276395 42890 276401
rect 43042 273573 43070 278467
rect 43138 276829 43166 291417
rect 43126 276823 43178 276829
rect 43126 276765 43178 276771
rect 43030 273567 43082 273573
rect 43030 273509 43082 273515
rect 42192 273194 42590 273222
rect 41780 273014 41836 273023
rect 41780 272949 41836 272958
rect 41794 272542 41822 272949
rect 41780 272422 41836 272431
rect 41780 272357 41836 272366
rect 41794 272024 41822 272357
rect 41780 270646 41836 270655
rect 41780 270581 41836 270590
rect 41794 270174 41822 270581
rect 41780 270054 41836 270063
rect 41780 269989 41836 269998
rect 41794 269508 41822 269989
rect 41780 269166 41836 269175
rect 41780 269101 41836 269110
rect 41794 268877 41822 269101
rect 23062 265057 23114 265063
rect 23062 264999 23114 265005
rect 23074 253339 23102 264999
rect 42178 264989 42206 268324
rect 42166 264983 42218 264989
rect 42166 264925 42218 264931
rect 23350 263651 23402 263657
rect 23350 263593 23402 263599
rect 23254 263577 23306 263583
rect 23254 263519 23306 263525
rect 23158 262171 23210 262177
rect 23158 262113 23210 262119
rect 23170 254227 23198 262113
rect 23156 254218 23212 254227
rect 23156 254153 23212 254162
rect 23060 253330 23116 253339
rect 23060 253265 23116 253274
rect 23266 252747 23294 263519
rect 23362 253339 23390 263593
rect 43234 263583 43262 295857
rect 43330 263657 43358 297041
rect 43318 263651 43370 263657
rect 43318 263593 43370 263599
rect 43222 263577 43274 263583
rect 43222 263519 43274 263525
rect 43318 262171 43370 262177
rect 43318 262113 43370 262119
rect 43330 261951 43358 262113
rect 43316 261942 43372 261951
rect 43316 261877 43372 261886
rect 40246 256399 40298 256405
rect 40246 256341 40298 256347
rect 40258 256299 40286 256341
rect 40244 256290 40300 256299
rect 40244 256225 40300 256234
rect 41588 255698 41644 255707
rect 41588 255633 41644 255642
rect 41602 253667 41630 255633
rect 41782 255437 41834 255443
rect 41780 255402 41782 255411
rect 41834 255402 41836 255411
rect 41780 255337 41836 255346
rect 41782 254993 41834 254999
rect 41780 254958 41782 254967
rect 41834 254958 41836 254967
rect 41780 254893 41836 254902
rect 41780 254514 41836 254523
rect 41780 254449 41782 254458
rect 41834 254449 41836 254458
rect 43222 254475 43274 254481
rect 41782 254417 41834 254423
rect 43222 254417 43274 254423
rect 41590 253661 41642 253667
rect 41590 253603 41642 253609
rect 23348 253330 23404 253339
rect 23348 253265 23404 253274
rect 23252 252738 23308 252747
rect 23252 252673 23308 252682
rect 40244 251258 40300 251267
rect 40244 251193 40300 251202
rect 34484 249778 34540 249787
rect 34484 249713 34540 249722
rect 34498 243603 34526 249713
rect 40258 244787 40286 251193
rect 41780 249482 41836 249491
rect 41780 249417 41836 249426
rect 41492 246670 41548 246679
rect 41492 246605 41548 246614
rect 40246 244781 40298 244787
rect 40246 244723 40298 244729
rect 41506 244713 41534 246605
rect 41684 245782 41740 245791
rect 41684 245717 41740 245726
rect 41588 245190 41644 245199
rect 41588 245125 41590 245134
rect 41642 245125 41644 245134
rect 41590 245093 41642 245099
rect 41590 245003 41642 245009
rect 41590 244945 41642 244951
rect 41602 244755 41630 244945
rect 41588 244746 41644 244755
rect 41494 244707 41546 244713
rect 41588 244681 41644 244690
rect 41494 244649 41546 244655
rect 41588 243710 41644 243719
rect 41588 243645 41644 243654
rect 34486 243597 34538 243603
rect 34486 243539 34538 243545
rect 41602 242641 41630 243645
rect 41698 243233 41726 245717
rect 41686 243227 41738 243233
rect 41686 243169 41738 243175
rect 41590 242635 41642 242641
rect 41590 242577 41642 242583
rect 41794 240643 41822 249417
rect 41876 247928 41932 247937
rect 41876 247863 41878 247872
rect 41930 247863 41932 247872
rect 42838 247889 42890 247895
rect 41878 247831 41930 247837
rect 42838 247831 42890 247837
rect 42260 247558 42316 247567
rect 42260 247493 42316 247502
rect 41876 246374 41932 246383
rect 41876 246309 41932 246318
rect 41890 241975 41918 246309
rect 41878 241969 41930 241975
rect 41878 241911 41930 241917
rect 41782 240637 41834 240643
rect 41782 240579 41834 240585
rect 41782 240415 41834 240421
rect 41782 240357 41834 240363
rect 41794 239834 41822 240357
rect 42166 238565 42218 238571
rect 42166 238507 42218 238513
rect 42178 237984 42206 238507
rect 42274 236179 42302 247493
rect 42548 245486 42604 245495
rect 42548 245421 42604 245430
rect 42454 244781 42506 244787
rect 42454 244723 42506 244729
rect 42358 243597 42410 243603
rect 42358 243539 42410 243545
rect 42192 236151 42302 236179
rect 42166 235457 42218 235463
rect 42166 235399 42218 235405
rect 42178 234950 42206 235399
rect 42262 235235 42314 235241
rect 42262 235177 42314 235183
rect 42274 234339 42302 235177
rect 42370 234520 42398 243539
rect 42466 238571 42494 244723
rect 42454 238565 42506 238571
rect 42454 238507 42506 238513
rect 42562 238423 42590 245421
rect 42646 244707 42698 244713
rect 42646 244649 42698 244655
rect 42550 238417 42602 238423
rect 42550 238359 42602 238365
rect 42658 238220 42686 244649
rect 42466 238192 42686 238220
rect 42466 235241 42494 238192
rect 42550 238121 42602 238127
rect 42550 238063 42602 238069
rect 42562 235463 42590 238063
rect 42850 237924 42878 247831
rect 42934 243227 42986 243233
rect 42934 243169 42986 243175
rect 42658 237896 42878 237924
rect 42550 235457 42602 235463
rect 42550 235399 42602 235405
rect 42454 235235 42506 235241
rect 42454 235177 42506 235183
rect 42370 234492 42494 234520
rect 42192 234311 42302 234339
rect 42262 234273 42314 234279
rect 42262 234215 42314 234221
rect 42274 233706 42302 234215
rect 42192 233678 42302 233706
rect 42466 233632 42494 234492
rect 42370 233604 42494 233632
rect 42370 233143 42398 233604
rect 42454 233459 42506 233465
rect 42454 233401 42506 233407
rect 42192 233115 42398 233143
rect 42466 230672 42494 233401
rect 42192 230644 42494 230672
rect 42658 230006 42686 237896
rect 42946 234279 42974 243169
rect 43126 241969 43178 241975
rect 43126 241911 43178 241917
rect 42934 234273 42986 234279
rect 42934 234215 42986 234221
rect 43138 233465 43166 241911
rect 43126 233459 43178 233465
rect 43126 233401 43178 233407
rect 42192 229978 42686 230006
rect 41780 229798 41836 229807
rect 41780 229733 41836 229742
rect 41794 229357 41822 229733
rect 41780 229206 41836 229215
rect 41780 229141 41836 229150
rect 41794 228808 41822 229141
rect 41780 227430 41836 227439
rect 41780 227365 41836 227374
rect 41794 226958 41822 227365
rect 41780 226838 41836 226847
rect 41780 226773 41836 226782
rect 41794 226321 41822 226773
rect 41780 225950 41836 225959
rect 41780 225885 41836 225894
rect 41794 225700 41822 225885
rect 42166 225467 42218 225473
rect 42166 225409 42218 225415
rect 42178 225108 42206 225409
rect 41782 213331 41834 213337
rect 41780 213296 41782 213305
rect 41834 213296 41836 213305
rect 41780 213231 41836 213240
rect 41590 212961 41642 212967
rect 41588 212926 41590 212935
rect 41642 212926 41644 212935
rect 41588 212861 41644 212870
rect 41782 212221 41834 212227
rect 41780 212186 41782 212195
rect 41834 212186 41836 212195
rect 41780 212121 41836 212130
rect 43234 211783 43262 254417
rect 41782 211777 41834 211783
rect 41780 211742 41782 211751
rect 43222 211777 43274 211783
rect 41834 211742 41836 211751
rect 43222 211719 43274 211725
rect 41780 211677 41836 211686
rect 41590 211481 41642 211487
rect 41588 211446 41590 211455
rect 41642 211446 41644 211455
rect 41588 211381 41644 211390
rect 41782 210741 41834 210747
rect 41780 210706 41782 210715
rect 41834 210706 41836 210715
rect 41780 210641 41836 210650
rect 41780 210262 41836 210271
rect 43330 210229 43358 261877
rect 43426 254999 43454 297559
rect 43508 266946 43564 266955
rect 43508 266881 43564 266890
rect 43522 265063 43550 266881
rect 43510 265057 43562 265063
rect 43510 264999 43562 265005
rect 43414 254993 43466 254999
rect 43414 254935 43466 254941
rect 41780 210197 41782 210206
rect 41834 210197 41836 210206
rect 43318 210223 43370 210229
rect 41782 210165 41834 210171
rect 43318 210165 43370 210171
rect 41590 210001 41642 210007
rect 41588 209966 41590 209975
rect 41642 209966 41644 209975
rect 41588 209901 41644 209910
rect 43522 209415 43550 264999
rect 44578 246341 44606 805125
rect 44674 267103 44702 814819
rect 44758 813619 44810 813625
rect 44758 813561 44810 813567
rect 44770 275391 44798 813561
rect 44866 785579 44894 817261
rect 44950 816579 45002 816585
rect 44950 816521 45002 816527
rect 44962 789131 44990 816521
rect 44950 789125 45002 789131
rect 44950 789067 45002 789073
rect 44854 785573 44906 785579
rect 44854 785515 44906 785521
rect 47458 785431 47486 817927
rect 57718 800743 57770 800749
rect 57718 800685 57770 800691
rect 57622 800669 57674 800675
rect 57622 800611 57674 800617
rect 57634 789691 57662 800611
rect 57730 790875 57758 800685
rect 57716 790866 57772 790875
rect 57716 790801 57772 790810
rect 57620 789682 57676 789691
rect 57620 789617 57676 789626
rect 58198 789199 58250 789205
rect 58198 789141 58250 789147
rect 58210 788507 58238 789141
rect 58390 789125 58442 789131
rect 58390 789067 58442 789073
rect 58196 788498 58252 788507
rect 58196 788433 58252 788442
rect 58402 787323 58430 789067
rect 58388 787314 58444 787323
rect 58388 787249 58444 787258
rect 59158 785573 59210 785579
rect 59158 785515 59210 785521
rect 59636 785538 59692 785547
rect 47446 785425 47498 785431
rect 47446 785367 47498 785373
rect 59170 784955 59198 785515
rect 59636 785473 59692 785482
rect 59650 785431 59678 785473
rect 59638 785425 59690 785431
rect 59638 785367 59690 785373
rect 59156 784946 59212 784955
rect 59156 784881 59212 784890
rect 47446 774695 47498 774701
rect 47446 774637 47498 774643
rect 44950 773955 45002 773961
rect 44950 773897 45002 773903
rect 44854 761967 44906 761973
rect 44854 761909 44906 761915
rect 44756 275382 44812 275391
rect 44756 275317 44812 275326
rect 44660 267094 44716 267103
rect 44660 267029 44716 267038
rect 44866 254925 44894 761909
rect 44962 742955 44990 773897
rect 45046 773511 45098 773517
rect 45046 773453 45098 773459
rect 45058 745471 45086 773453
rect 45046 745465 45098 745471
rect 45046 745407 45098 745413
rect 47458 743029 47486 774637
rect 62038 772179 62090 772185
rect 62038 772121 62090 772127
rect 61846 771957 61898 771963
rect 61846 771899 61898 771905
rect 58678 757527 58730 757533
rect 58678 757469 58730 757475
rect 58690 747659 58718 757469
rect 58676 747650 58732 747659
rect 58676 747585 58732 747594
rect 54740 746022 54796 746031
rect 54646 745983 54698 745989
rect 54740 745957 54742 745966
rect 54646 745925 54698 745931
rect 54794 745957 54796 745966
rect 57622 745983 57674 745989
rect 54742 745925 54794 745931
rect 57622 745925 57674 745931
rect 54658 745883 54686 745925
rect 54644 745874 54700 745883
rect 54644 745809 54700 745818
rect 57634 745291 57662 745925
rect 58102 745465 58154 745471
rect 58102 745407 58154 745413
rect 58580 745430 58636 745439
rect 57620 745282 57676 745291
rect 57620 745217 57676 745226
rect 58114 744107 58142 745407
rect 58580 745365 58636 745374
rect 58594 745027 58622 745365
rect 58582 745021 58634 745027
rect 58582 744963 58634 744969
rect 58100 744098 58156 744107
rect 58100 744033 58156 744042
rect 47446 743023 47498 743029
rect 47446 742965 47498 742971
rect 59638 743023 59690 743029
rect 59638 742965 59690 742971
rect 44950 742949 45002 742955
rect 59650 742923 59678 742965
rect 59734 742949 59786 742955
rect 44950 742891 45002 742897
rect 59636 742914 59692 742923
rect 59734 742891 59786 742897
rect 59636 742849 59692 742858
rect 59746 741739 59774 742891
rect 59732 741730 59788 741739
rect 59732 741665 59788 741674
rect 47542 731479 47594 731485
rect 47542 731421 47594 731427
rect 44950 730739 45002 730745
rect 44950 730681 45002 730687
rect 44962 699739 44990 730681
rect 45046 730369 45098 730375
rect 45046 730311 45098 730317
rect 45058 702625 45086 730311
rect 47446 718751 47498 718757
rect 47446 718693 47498 718699
rect 45046 702619 45098 702625
rect 45046 702561 45098 702567
rect 44950 699733 45002 699739
rect 44950 699675 45002 699681
rect 45046 685377 45098 685383
rect 45046 685319 45098 685325
rect 44950 684193 45002 684199
rect 44950 684135 45002 684141
rect 44962 261707 44990 684135
rect 45058 266395 45086 685319
rect 45142 665323 45194 665329
rect 45142 665265 45194 665271
rect 45154 659409 45182 665265
rect 45142 659403 45194 659409
rect 45142 659345 45194 659351
rect 45142 596207 45194 596213
rect 45142 596149 45194 596155
rect 45154 276279 45182 596149
rect 45238 330399 45290 330405
rect 45238 330341 45290 330347
rect 45140 276270 45196 276279
rect 45140 276205 45196 276214
rect 45046 266389 45098 266395
rect 45046 266331 45098 266337
rect 44948 261698 45004 261707
rect 44948 261633 45004 261642
rect 44854 254919 44906 254925
rect 44854 254861 44906 254867
rect 44950 253513 45002 253519
rect 44950 253455 45002 253461
rect 44566 246335 44618 246341
rect 44566 246277 44618 246283
rect 44758 244929 44810 244935
rect 44758 244871 44810 244877
rect 44662 242857 44714 242863
rect 44662 242799 44714 242805
rect 44566 242709 44618 242715
rect 44566 242651 44618 242657
rect 41590 209409 41642 209415
rect 41588 209374 41590 209383
rect 43510 209409 43562 209415
rect 41642 209374 41644 209383
rect 43510 209351 43562 209357
rect 41588 209309 41644 209318
rect 41780 208264 41836 208273
rect 41780 208199 41836 208208
rect 41794 207565 41822 208199
rect 41782 207559 41834 207565
rect 41782 207501 41834 207507
rect 42934 207559 42986 207565
rect 42934 207501 42986 207507
rect 34100 206562 34156 206571
rect 34100 206497 34156 206506
rect 34114 200387 34142 206497
rect 42260 206266 42316 206275
rect 42260 206201 42316 206210
rect 34196 204490 34252 204499
rect 34196 204425 34252 204434
rect 34102 200381 34154 200387
rect 34102 200323 34154 200329
rect 34210 200313 34238 204425
rect 34292 204046 34348 204055
rect 34292 203981 34348 203990
rect 34198 200307 34250 200313
rect 34198 200249 34250 200255
rect 34306 200239 34334 203981
rect 41588 203602 41644 203611
rect 41588 203537 41644 203546
rect 34484 203010 34540 203019
rect 34484 202945 34540 202954
rect 34388 201974 34444 201983
rect 34388 201909 34444 201918
rect 34294 200233 34346 200239
rect 34294 200175 34346 200181
rect 34402 200165 34430 201909
rect 34498 200461 34526 202945
rect 41602 201793 41630 203537
rect 41876 202862 41932 202871
rect 41876 202797 41932 202806
rect 41590 201787 41642 201793
rect 41590 201729 41642 201735
rect 41890 201645 41918 202797
rect 41974 201713 42026 201719
rect 41972 201678 41974 201687
rect 42026 201678 42028 201687
rect 41878 201639 41930 201645
rect 41972 201613 42028 201622
rect 41878 201581 41930 201587
rect 41590 201565 41642 201571
rect 41588 201530 41590 201539
rect 41642 201530 41644 201539
rect 41588 201465 41644 201474
rect 41590 200973 41642 200979
rect 41588 200938 41590 200947
rect 41642 200938 41644 200947
rect 41588 200873 41644 200882
rect 34486 200455 34538 200461
rect 34486 200397 34538 200403
rect 34390 200159 34442 200165
rect 34390 200101 34442 200107
rect 42274 197224 42302 206201
rect 42550 201787 42602 201793
rect 42550 201729 42602 201735
rect 42358 200233 42410 200239
rect 42358 200175 42410 200181
rect 42178 197196 42302 197224
rect 42178 196618 42206 197196
rect 42262 194831 42314 194837
rect 42192 194791 42262 194819
rect 42262 194773 42314 194779
rect 42370 193006 42398 200175
rect 42562 195854 42590 201729
rect 42742 201639 42794 201645
rect 42742 201581 42794 201587
rect 42646 200455 42698 200461
rect 42646 200397 42698 200403
rect 42178 192932 42206 192992
rect 42274 192978 42398 193006
rect 42466 195826 42590 195854
rect 42274 192932 42302 192978
rect 42178 192904 42302 192932
rect 42358 192907 42410 192913
rect 42358 192849 42410 192855
rect 42370 191783 42398 192849
rect 42192 191755 42398 191783
rect 42466 191156 42494 195826
rect 42658 191655 42686 200397
rect 42646 191649 42698 191655
rect 42646 191591 42698 191597
rect 42178 191008 42206 191142
rect 42274 191128 42494 191156
rect 42274 191008 42302 191128
rect 42178 190980 42302 191008
rect 42754 190564 42782 201581
rect 42838 200381 42890 200387
rect 42838 200323 42890 200329
rect 42562 190536 42782 190564
rect 42562 190490 42590 190536
rect 42192 190462 42590 190490
rect 42850 190120 42878 200323
rect 42946 194837 42974 207501
rect 44578 201571 44606 242651
rect 44566 201565 44618 201571
rect 44566 201507 44618 201513
rect 44674 200979 44702 242799
rect 44770 201719 44798 244871
rect 44854 242783 44906 242789
rect 44854 242725 44906 242731
rect 44866 211487 44894 242725
rect 44962 212227 44990 253455
rect 45250 246267 45278 330341
rect 45526 287183 45578 287189
rect 45526 287125 45578 287131
rect 45334 279487 45386 279493
rect 45334 279429 45386 279435
rect 45238 246261 45290 246267
rect 45238 246203 45290 246209
rect 45346 212967 45374 279429
rect 45430 279413 45482 279419
rect 45430 279355 45482 279361
rect 45442 213337 45470 279355
rect 45538 246415 45566 287125
rect 45718 264835 45770 264841
rect 45718 264777 45770 264783
rect 45730 263583 45758 264777
rect 46006 264761 46058 264767
rect 46006 264703 46058 264709
rect 46018 263657 46046 264703
rect 46006 263651 46058 263657
rect 46006 263593 46058 263599
rect 45718 263577 45770 263583
rect 45718 263519 45770 263525
rect 47458 246563 47486 718693
rect 47554 699813 47582 731421
rect 59638 714311 59690 714317
rect 59638 714253 59690 714259
rect 59650 704443 59678 714253
rect 59636 704434 59692 704443
rect 59636 704369 59692 704378
rect 58870 702767 58922 702773
rect 58870 702709 58922 702715
rect 58774 702693 58826 702699
rect 58772 702658 58774 702667
rect 58826 702658 58828 702667
rect 58678 702619 58730 702625
rect 58772 702593 58828 702602
rect 58678 702561 58730 702567
rect 58690 700891 58718 702561
rect 58882 702075 58910 702709
rect 58868 702066 58924 702075
rect 58868 702001 58924 702010
rect 58676 700882 58732 700891
rect 58676 700817 58732 700826
rect 47542 699807 47594 699813
rect 47542 699749 47594 699755
rect 59254 699807 59306 699813
rect 59254 699749 59306 699755
rect 58870 699733 58922 699739
rect 59266 699707 59294 699749
rect 58870 699675 58922 699681
rect 59252 699698 59308 699707
rect 58882 698523 58910 699675
rect 59252 699633 59308 699642
rect 58868 698514 58924 698523
rect 58868 698449 58924 698458
rect 50326 688263 50378 688269
rect 50326 688205 50378 688211
rect 47638 687523 47690 687529
rect 47638 687465 47690 687471
rect 47542 675757 47594 675763
rect 47542 675699 47594 675705
rect 47554 246637 47582 675699
rect 47650 656597 47678 687465
rect 47734 687227 47786 687233
rect 47734 687169 47786 687175
rect 47746 659483 47774 687169
rect 47734 659477 47786 659483
rect 47734 659419 47786 659425
rect 50338 656671 50366 688205
rect 59638 671095 59690 671101
rect 59638 671037 59690 671043
rect 59650 661227 59678 671037
rect 59636 661218 59692 661227
rect 59636 661153 59692 661162
rect 57718 659551 57770 659557
rect 57718 659493 57770 659499
rect 57730 658859 57758 659493
rect 59158 659477 59210 659483
rect 58772 659442 58828 659451
rect 59158 659419 59210 659425
rect 58772 659377 58774 659386
rect 58826 659377 58828 659386
rect 58774 659345 58826 659351
rect 57716 658850 57772 658859
rect 57716 658785 57772 658794
rect 59170 657675 59198 659419
rect 59156 657666 59212 657675
rect 59156 657601 59212 657610
rect 50326 656665 50378 656671
rect 50326 656607 50378 656613
rect 58198 656665 58250 656671
rect 58198 656607 58250 656613
rect 47638 656591 47690 656597
rect 47638 656533 47690 656539
rect 58210 656491 58238 656607
rect 58390 656591 58442 656597
rect 58390 656533 58442 656539
rect 58196 656482 58252 656491
rect 58196 656417 58252 656426
rect 58402 655307 58430 656533
rect 58388 655298 58444 655307
rect 58388 655233 58444 655242
rect 50326 644899 50378 644905
rect 50326 644841 50378 644847
rect 47734 644307 47786 644313
rect 47734 644249 47786 644255
rect 47638 632541 47690 632547
rect 47638 632483 47690 632489
rect 47542 246631 47594 246637
rect 47542 246573 47594 246579
rect 47446 246557 47498 246563
rect 47446 246499 47498 246505
rect 47650 246489 47678 632483
rect 47746 613381 47774 644249
rect 47830 644011 47882 644017
rect 47830 643953 47882 643959
rect 47842 616341 47870 643953
rect 47926 622107 47978 622113
rect 47926 622049 47978 622055
rect 47830 616335 47882 616341
rect 47830 616277 47882 616283
rect 47938 616267 47966 622049
rect 47926 616261 47978 616267
rect 47926 616203 47978 616209
rect 50338 613455 50366 644841
rect 54646 627879 54698 627885
rect 54646 627821 54698 627827
rect 54658 624851 54686 627821
rect 54646 624845 54698 624851
rect 54646 624787 54698 624793
rect 58966 624845 59018 624851
rect 58966 624787 59018 624793
rect 58978 618011 59006 624787
rect 58964 618002 59020 618011
rect 58964 617937 59020 617946
rect 58198 616409 58250 616415
rect 58198 616351 58250 616357
rect 58210 615643 58238 616351
rect 58966 616335 59018 616341
rect 58966 616277 59018 616283
rect 58196 615634 58252 615643
rect 58196 615569 58252 615578
rect 58978 614459 59006 616277
rect 59638 616261 59690 616267
rect 59636 616226 59638 616235
rect 59690 616226 59692 616235
rect 59636 616161 59692 616170
rect 58964 614450 59020 614459
rect 58964 614385 59020 614394
rect 50326 613449 50378 613455
rect 50326 613391 50378 613397
rect 59638 613449 59690 613455
rect 59638 613391 59690 613397
rect 47734 613375 47786 613381
rect 47734 613317 47786 613323
rect 59542 613375 59594 613381
rect 59542 613317 59594 613323
rect 59554 612091 59582 613317
rect 59650 613275 59678 613391
rect 59636 613266 59692 613275
rect 59636 613201 59692 613210
rect 59540 612082 59596 612091
rect 59540 612017 59596 612026
rect 50326 601683 50378 601689
rect 50326 601625 50378 601631
rect 47734 601387 47786 601393
rect 47734 601329 47786 601335
rect 47746 570165 47774 601329
rect 47830 600795 47882 600801
rect 47830 600737 47882 600743
rect 47842 573125 47870 600737
rect 47926 579039 47978 579045
rect 47926 578981 47978 578987
rect 47830 573119 47882 573125
rect 47830 573061 47882 573067
rect 47938 573051 47966 578981
rect 47926 573045 47978 573051
rect 47926 572987 47978 572993
rect 50338 570239 50366 601625
rect 56086 587549 56138 587555
rect 56086 587491 56138 587497
rect 50326 570233 50378 570239
rect 50326 570175 50378 570181
rect 47734 570159 47786 570165
rect 47734 570101 47786 570107
rect 50326 524353 50378 524359
rect 50326 524295 50378 524301
rect 47734 524279 47786 524285
rect 47734 524221 47786 524227
rect 47746 475593 47774 524221
rect 50338 476111 50366 524295
rect 50326 476105 50378 476111
rect 50326 476047 50378 476053
rect 47734 475587 47786 475593
rect 47734 475529 47786 475535
rect 47734 463599 47786 463605
rect 47734 463541 47786 463547
rect 47746 255073 47774 463541
rect 48022 428495 48074 428501
rect 48022 428437 48074 428443
rect 47926 428125 47978 428131
rect 47926 428067 47978 428073
rect 47830 416137 47882 416143
rect 47830 416079 47882 416085
rect 47734 255067 47786 255073
rect 47734 255009 47786 255015
rect 47842 254999 47870 416079
rect 47938 400187 47966 428067
rect 48034 400335 48062 428437
rect 48118 427607 48170 427613
rect 48118 427549 48170 427555
rect 48022 400329 48074 400335
rect 48022 400271 48074 400277
rect 48130 400261 48158 427549
rect 48118 400255 48170 400261
rect 48118 400197 48170 400203
rect 47926 400181 47978 400187
rect 47926 400123 47978 400129
rect 48022 385973 48074 385979
rect 48022 385915 48074 385921
rect 47926 373319 47978 373325
rect 47926 373261 47978 373267
rect 47938 255147 47966 373261
rect 48034 357119 48062 385915
rect 48214 385307 48266 385313
rect 48214 385249 48266 385255
rect 48118 385011 48170 385017
rect 48118 384953 48170 384959
rect 48022 357113 48074 357119
rect 48022 357055 48074 357061
rect 48130 357045 48158 384953
rect 48118 357039 48170 357045
rect 48118 356981 48170 356987
rect 48226 356971 48254 385249
rect 48214 356965 48266 356971
rect 48214 356907 48266 356913
rect 48022 342831 48074 342837
rect 48022 342773 48074 342779
rect 48034 313829 48062 342773
rect 48118 342313 48170 342319
rect 48118 342255 48170 342261
rect 48022 313823 48074 313829
rect 48022 313765 48074 313771
rect 48130 313755 48158 342255
rect 48214 341795 48266 341801
rect 48214 341737 48266 341743
rect 48226 313903 48254 341737
rect 48214 313897 48266 313903
rect 48214 313839 48266 313845
rect 48118 313749 48170 313755
rect 48118 313691 48170 313697
rect 51478 299171 51530 299177
rect 51478 299113 51530 299119
rect 51490 288373 51518 299113
rect 53302 290957 53354 290963
rect 53302 290899 53354 290905
rect 51478 288367 51530 288373
rect 51478 288309 51530 288315
rect 48022 288071 48074 288077
rect 48022 288013 48074 288019
rect 47926 255141 47978 255147
rect 47926 255083 47978 255089
rect 47830 254993 47882 254999
rect 47830 254935 47882 254941
rect 47638 246483 47690 246489
rect 47638 246425 47690 246431
rect 45526 246409 45578 246415
rect 45526 246351 45578 246357
rect 48034 225473 48062 288013
rect 53206 285185 53258 285191
rect 53206 285127 53258 285133
rect 50326 282373 50378 282379
rect 50326 282315 50378 282321
rect 48022 225467 48074 225473
rect 48022 225409 48074 225415
rect 45430 213331 45482 213337
rect 45430 213273 45482 213279
rect 45334 212961 45386 212967
rect 45334 212903 45386 212909
rect 44950 212221 45002 212227
rect 44950 212163 45002 212169
rect 44854 211481 44906 211487
rect 44854 211423 44906 211429
rect 44758 201713 44810 201719
rect 44758 201655 44810 201661
rect 44662 200973 44714 200979
rect 44662 200915 44714 200921
rect 43030 200307 43082 200313
rect 43030 200249 43082 200255
rect 42934 194831 42986 194837
rect 42934 194773 42986 194779
rect 42934 191649 42986 191655
rect 42934 191591 42986 191597
rect 42562 190092 42878 190120
rect 42562 189943 42590 190092
rect 42192 189915 42590 189943
rect 42946 187604 42974 191591
rect 42562 187576 42974 187604
rect 42562 187456 42590 187576
rect 42192 187428 42590 187456
rect 43042 186864 43070 200249
rect 43126 200159 43178 200165
rect 43126 200101 43178 200107
rect 43138 192913 43166 200101
rect 43126 192907 43178 192913
rect 43126 192849 43178 192855
rect 42178 186836 42302 186864
rect 42178 186776 42206 186836
rect 42274 186790 42302 186836
rect 42466 186836 43070 186864
rect 42466 186790 42494 186836
rect 42274 186762 42494 186790
rect 41780 186730 41836 186739
rect 41780 186665 41836 186674
rect 41794 186184 41822 186665
rect 41780 185842 41836 185851
rect 41780 185777 41836 185786
rect 41794 185592 41822 185777
rect 41780 184214 41836 184223
rect 41780 184149 41836 184158
rect 41794 183742 41822 184149
rect 41780 183622 41836 183631
rect 41780 183557 41836 183566
rect 41794 183121 41822 183557
rect 41780 182882 41836 182891
rect 41780 182817 41836 182826
rect 41794 182484 41822 182817
rect 42178 178557 42206 181925
rect 50338 178557 50366 282315
rect 50612 275234 50668 275243
rect 50612 275169 50668 275178
rect 50420 275086 50476 275095
rect 50420 275021 50476 275030
rect 50434 210007 50462 275021
rect 50626 210747 50654 275169
rect 53218 255443 53246 285127
rect 53314 264989 53342 290899
rect 53302 264983 53354 264989
rect 53302 264925 53354 264931
rect 53206 255437 53258 255443
rect 53206 255379 53258 255385
rect 56098 252039 56126 587491
rect 58966 584737 59018 584743
rect 58966 584679 59018 584685
rect 58978 574795 59006 584679
rect 58964 574786 59020 574795
rect 58964 574721 59020 574730
rect 58198 573193 58250 573199
rect 58198 573135 58250 573141
rect 58210 572427 58238 573135
rect 58966 573119 59018 573125
rect 58966 573061 59018 573067
rect 58196 572418 58252 572427
rect 58196 572353 58252 572362
rect 58978 571243 59006 573061
rect 59638 573045 59690 573051
rect 59636 573010 59638 573019
rect 59690 573010 59692 573019
rect 59636 572945 59692 572954
rect 58964 571234 59020 571243
rect 58964 571169 59020 571178
rect 59350 570233 59402 570239
rect 59350 570175 59402 570181
rect 59362 570059 59390 570175
rect 59542 570159 59594 570165
rect 59542 570101 59594 570107
rect 59348 570050 59404 570059
rect 59348 569985 59404 569994
rect 59554 568875 59582 570101
rect 59540 568866 59596 568875
rect 59540 568801 59596 568810
rect 57718 541595 57770 541601
rect 57718 541537 57770 541543
rect 57622 541521 57674 541527
rect 57622 541463 57674 541469
rect 57634 530543 57662 541463
rect 57730 531727 57758 541537
rect 57716 531718 57772 531727
rect 57716 531653 57772 531662
rect 57620 530534 57676 530543
rect 57620 530469 57676 530478
rect 58198 529977 58250 529983
rect 58198 529919 58250 529925
rect 58210 529359 58238 529919
rect 58196 529350 58252 529359
rect 58196 529285 58252 529294
rect 58964 527130 59020 527139
rect 58964 527065 59020 527074
rect 58580 525946 58636 525955
rect 58580 525881 58636 525890
rect 58594 524359 58622 525881
rect 58582 524353 58634 524359
rect 58582 524295 58634 524301
rect 58978 472411 59006 527065
rect 59348 524762 59404 524771
rect 59348 524697 59404 524706
rect 59362 524285 59390 524697
rect 59350 524279 59402 524285
rect 59350 524221 59402 524227
rect 58966 472405 59018 472411
rect 58966 472347 59018 472353
rect 58486 406101 58538 406107
rect 58486 406043 58538 406049
rect 58498 404151 58526 406043
rect 58484 404142 58540 404151
rect 58484 404077 58540 404086
rect 58774 403067 58826 403073
rect 58774 403009 58826 403015
rect 58786 402967 58814 403009
rect 58772 402958 58828 402967
rect 58772 402893 58828 402902
rect 57620 400590 57676 400599
rect 57620 400525 57676 400534
rect 57634 394563 57662 400525
rect 58198 400329 58250 400335
rect 58198 400271 58250 400277
rect 58210 399415 58238 400271
rect 58774 400255 58826 400261
rect 58774 400197 58826 400203
rect 58786 400007 58814 400197
rect 59734 400181 59786 400187
rect 59734 400123 59786 400129
rect 58772 399998 58828 400007
rect 58772 399933 58828 399942
rect 58196 399406 58252 399415
rect 58196 399341 58252 399350
rect 59746 398231 59774 400123
rect 59732 398222 59788 398231
rect 59732 398157 59788 398166
rect 57622 394557 57674 394563
rect 57622 394499 57674 394505
rect 58486 362885 58538 362891
rect 58486 362827 58538 362833
rect 58498 360935 58526 362827
rect 58484 360926 58540 360935
rect 58484 360861 58540 360870
rect 59158 359999 59210 360005
rect 59158 359941 59210 359947
rect 59170 359751 59198 359941
rect 59156 359742 59212 359751
rect 59156 359677 59212 359686
rect 57620 357522 57676 357531
rect 57620 357457 57676 357466
rect 57634 351347 57662 357457
rect 58198 357113 58250 357119
rect 58198 357055 58250 357061
rect 58210 356199 58238 357055
rect 59638 357039 59690 357045
rect 59638 356981 59690 356987
rect 58582 356965 58634 356971
rect 58582 356907 58634 356913
rect 58196 356190 58252 356199
rect 58196 356125 58252 356134
rect 58594 355015 58622 356907
rect 59650 356791 59678 356981
rect 59636 356782 59692 356791
rect 59636 356717 59692 356726
rect 58580 355006 58636 355015
rect 58580 354941 58636 354950
rect 57622 351341 57674 351347
rect 57622 351283 57674 351289
rect 58486 319669 58538 319675
rect 58486 319611 58538 319617
rect 58498 317719 58526 319611
rect 58484 317710 58540 317719
rect 58484 317645 58540 317654
rect 59158 316783 59210 316789
rect 59158 316725 59210 316731
rect 59170 316535 59198 316725
rect 59156 316526 59212 316535
rect 59156 316461 59212 316470
rect 59156 314158 59212 314167
rect 59156 314093 59212 314102
rect 58870 313823 58922 313829
rect 58870 313765 58922 313771
rect 58882 312983 58910 313765
rect 58868 312974 58924 312983
rect 58868 312909 58924 312918
rect 59170 308131 59198 314093
rect 59638 313897 59690 313903
rect 59636 313862 59638 313871
rect 59690 313862 59692 313871
rect 59636 313797 59692 313806
rect 59638 313749 59690 313755
rect 59638 313691 59690 313697
rect 59650 311799 59678 313691
rect 59636 311790 59692 311799
rect 59636 311725 59692 311734
rect 59158 308125 59210 308131
rect 59158 308067 59210 308073
rect 61654 298135 61706 298141
rect 61654 298077 61706 298083
rect 59348 295214 59404 295223
rect 59348 295149 59404 295158
rect 59252 294030 59308 294039
rect 59252 293965 59308 293974
rect 58198 293769 58250 293775
rect 58198 293711 58250 293717
rect 58210 292707 58238 293711
rect 58196 292698 58252 292707
rect 58196 292633 58252 292642
rect 58868 289294 58924 289303
rect 58868 289229 58924 289238
rect 58882 288373 58910 289229
rect 58870 288367 58922 288373
rect 58870 288309 58922 288315
rect 59156 288110 59212 288119
rect 59156 288045 59158 288054
rect 59210 288045 59212 288054
rect 59158 288013 59210 288019
rect 59266 287060 59294 293965
rect 59170 287032 59294 287060
rect 59060 285742 59116 285751
rect 59060 285677 59116 285686
rect 57620 284558 57676 284567
rect 57620 284493 57676 284502
rect 57634 282305 57662 284493
rect 58868 283374 58924 283383
rect 58868 283309 58924 283318
rect 58882 282379 58910 283309
rect 58870 282373 58922 282379
rect 58870 282315 58922 282321
rect 58964 282338 59020 282347
rect 56182 282299 56234 282305
rect 56182 282241 56234 282247
rect 57622 282299 57674 282305
rect 58964 282273 59020 282282
rect 57622 282241 57674 282247
rect 56194 253667 56222 282241
rect 56182 253661 56234 253667
rect 56182 253603 56234 253609
rect 58978 253519 59006 282273
rect 59074 256405 59102 285677
rect 59170 273573 59198 287032
rect 59252 286926 59308 286935
rect 59252 286861 59308 286870
rect 59266 285191 59294 286861
rect 59254 285185 59306 285191
rect 59254 285127 59306 285133
rect 59252 281006 59308 281015
rect 59252 280941 59308 280950
rect 59266 279419 59294 280941
rect 59254 279413 59306 279419
rect 59254 279355 59306 279361
rect 59362 276459 59390 295149
rect 59444 292846 59500 292855
rect 59444 292781 59500 292790
rect 59458 290963 59486 292781
rect 59638 291623 59690 291629
rect 59638 291565 59690 291571
rect 59650 291523 59678 291565
rect 59636 291514 59692 291523
rect 59636 291449 59692 291458
rect 59446 290957 59498 290963
rect 59446 290899 59498 290905
rect 59540 279822 59596 279831
rect 59540 279757 59596 279766
rect 59554 279493 59582 279757
rect 59542 279487 59594 279493
rect 59542 279429 59594 279435
rect 61666 277907 61694 298077
rect 61652 277898 61708 277907
rect 61652 277833 61708 277842
rect 59350 276453 59402 276459
rect 59350 276395 59402 276401
rect 59158 273567 59210 273573
rect 59158 273509 59210 273515
rect 61858 266659 61886 771899
rect 61942 642531 61994 642537
rect 61942 642473 61994 642479
rect 61954 278351 61982 642473
rect 61940 278342 61996 278351
rect 61940 278277 61996 278286
rect 62050 266807 62078 772121
rect 62230 728741 62282 728747
rect 62230 728683 62282 728689
rect 62132 602166 62188 602175
rect 62132 602101 62188 602110
rect 62146 278499 62174 602101
rect 62132 278490 62188 278499
rect 62132 278425 62188 278434
rect 62036 266798 62092 266807
rect 62036 266733 62092 266742
rect 61844 266650 61900 266659
rect 61844 266585 61900 266594
rect 62242 266363 62270 728683
rect 62422 728667 62474 728673
rect 62422 728609 62474 728615
rect 62324 537046 62380 537055
rect 62324 536981 62380 536990
rect 62338 270655 62366 536981
rect 62324 270646 62380 270655
rect 62324 270581 62380 270590
rect 62434 266511 62462 728609
rect 62518 437847 62570 437853
rect 62518 437789 62570 437795
rect 62530 278055 62558 437789
rect 62614 423417 62666 423423
rect 62614 423359 62666 423365
rect 62516 278046 62572 278055
rect 62516 277981 62572 277990
rect 62626 273467 62654 423359
rect 62708 386086 62764 386095
rect 62708 386021 62764 386030
rect 62722 277611 62750 386021
rect 62900 383274 62956 383283
rect 62900 383209 62956 383218
rect 62914 277759 62942 383209
rect 63092 343166 63148 343175
rect 63092 343101 63148 343110
rect 63106 278203 63134 343101
rect 63286 300947 63338 300953
rect 63286 300889 63338 300895
rect 63092 278194 63148 278203
rect 63092 278129 63148 278138
rect 62900 277750 62956 277759
rect 62900 277685 62956 277694
rect 62708 277602 62764 277611
rect 62708 277537 62764 277546
rect 63298 277463 63326 300889
rect 408322 278309 408624 278328
rect 314902 278303 314954 278309
rect 314902 278245 314954 278251
rect 408310 278303 408624 278309
rect 408362 278300 408624 278303
rect 408310 278245 408362 278251
rect 63284 277454 63340 277463
rect 63284 277389 63340 277398
rect 62612 273458 62668 273467
rect 62612 273393 62668 273402
rect 65890 269323 65918 278018
rect 65876 269314 65932 269323
rect 67042 269281 67070 278018
rect 68290 273277 68318 278018
rect 68278 273271 68330 273277
rect 68278 273213 68330 273219
rect 69442 269619 69470 278018
rect 70594 272135 70622 278018
rect 70580 272126 70636 272135
rect 70580 272061 70636 272070
rect 69428 269610 69484 269619
rect 69428 269545 69484 269554
rect 71746 269471 71774 278018
rect 72994 272283 73022 278018
rect 72980 272274 73036 272283
rect 72980 272209 73036 272218
rect 71732 269462 71788 269471
rect 71732 269397 71788 269406
rect 74146 269355 74174 278018
rect 75298 271649 75326 278018
rect 76546 272315 76574 278018
rect 77698 276494 77726 278018
rect 77602 276466 77726 276494
rect 76534 272309 76586 272315
rect 76534 272251 76586 272257
rect 75286 271643 75338 271649
rect 75286 271585 75338 271591
rect 77602 269767 77630 276466
rect 78850 272431 78878 278018
rect 80112 278004 80606 278032
rect 78836 272422 78892 272431
rect 78836 272357 78892 272366
rect 77686 271643 77738 271649
rect 77686 271585 77738 271591
rect 77588 269758 77644 269767
rect 77588 269693 77644 269702
rect 74134 269349 74186 269355
rect 74134 269291 74186 269297
rect 65876 269249 65932 269258
rect 67030 269275 67082 269281
rect 67030 269217 67082 269223
rect 62420 266502 62476 266511
rect 62420 266437 62476 266446
rect 62228 266354 62284 266363
rect 62228 266289 62284 266298
rect 59062 256399 59114 256405
rect 59062 256341 59114 256347
rect 58966 253513 59018 253519
rect 58966 253455 59018 253461
rect 56086 252033 56138 252039
rect 56086 251975 56138 251981
rect 77698 249301 77726 271585
rect 77686 249295 77738 249301
rect 77686 249237 77738 249243
rect 80578 249227 80606 278004
rect 81250 269429 81278 278018
rect 82402 269577 82430 278018
rect 83650 269651 83678 278018
rect 84802 272241 84830 278018
rect 84790 272235 84842 272241
rect 84790 272177 84842 272183
rect 85954 271131 85982 278018
rect 86326 272235 86378 272241
rect 86326 272177 86378 272183
rect 85942 271125 85994 271131
rect 85942 271067 85994 271073
rect 83638 269645 83690 269651
rect 83638 269587 83690 269593
rect 82390 269571 82442 269577
rect 82390 269513 82442 269519
rect 81238 269423 81290 269429
rect 81238 269365 81290 269371
rect 80566 249221 80618 249227
rect 80566 249163 80618 249169
rect 86338 249153 86366 272177
rect 87202 269503 87230 278018
rect 88354 272579 88382 278018
rect 88340 272570 88396 272579
rect 88340 272505 88396 272514
rect 89506 271575 89534 278018
rect 89494 271569 89546 271575
rect 89494 271511 89546 271517
rect 90658 269725 90686 278018
rect 91906 272727 91934 278018
rect 91892 272718 91948 272727
rect 91892 272653 91948 272662
rect 92086 271569 92138 271575
rect 92086 271511 92138 271517
rect 90646 269719 90698 269725
rect 90646 269661 90698 269667
rect 87190 269497 87242 269503
rect 87190 269439 87242 269445
rect 92098 252261 92126 271511
rect 93058 269799 93086 278018
rect 94210 270761 94238 278018
rect 94198 270755 94250 270761
rect 94198 270697 94250 270703
rect 94966 270755 95018 270761
rect 94966 270697 95018 270703
rect 93046 269793 93098 269799
rect 93046 269735 93098 269741
rect 92086 252255 92138 252261
rect 92086 252197 92138 252203
rect 94978 249449 95006 270697
rect 95458 269873 95486 278018
rect 96610 272611 96638 278018
rect 97776 278004 97886 278032
rect 96598 272605 96650 272611
rect 96598 272547 96650 272553
rect 95446 269867 95498 269873
rect 95446 269809 95498 269815
rect 97858 252113 97886 278004
rect 99010 272389 99038 278018
rect 98998 272383 99050 272389
rect 98998 272325 99050 272331
rect 100162 269947 100190 278018
rect 101314 270761 101342 278018
rect 101302 270755 101354 270761
rect 101302 270697 101354 270703
rect 102562 270021 102590 278018
rect 103714 272463 103742 278018
rect 103702 272457 103754 272463
rect 103702 272399 103754 272405
rect 104866 272241 104894 278018
rect 106114 272537 106142 278018
rect 106678 272605 106730 272611
rect 106678 272547 106730 272553
rect 106102 272531 106154 272537
rect 106102 272473 106154 272479
rect 106690 272315 106718 272547
rect 106678 272309 106730 272315
rect 106678 272251 106730 272257
rect 104854 272235 104906 272241
rect 104854 272177 104906 272183
rect 106486 272235 106538 272241
rect 106486 272177 106538 272183
rect 103606 270755 103658 270761
rect 103606 270697 103658 270703
rect 102550 270015 102602 270021
rect 102550 269957 102602 269963
rect 100150 269941 100202 269947
rect 100150 269883 100202 269889
rect 97846 252107 97898 252113
rect 97846 252049 97898 252055
rect 94966 249443 95018 249449
rect 94966 249385 95018 249391
rect 86326 249147 86378 249153
rect 86326 249089 86378 249095
rect 103618 246785 103646 270697
rect 106498 252335 106526 272177
rect 107266 270095 107294 278018
rect 108418 273425 108446 278018
rect 108406 273419 108458 273425
rect 108406 273361 108458 273367
rect 109366 273419 109418 273425
rect 109366 273361 109418 273367
rect 107254 270089 107306 270095
rect 107254 270031 107306 270037
rect 106486 252329 106538 252335
rect 106486 252271 106538 252277
rect 109378 252187 109406 273361
rect 109570 270169 109598 278018
rect 110818 272611 110846 278018
rect 111984 278004 112286 278032
rect 110806 272605 110858 272611
rect 110806 272547 110858 272553
rect 109558 270163 109610 270169
rect 109558 270105 109610 270111
rect 109366 252181 109418 252187
rect 109366 252123 109418 252129
rect 103606 246779 103658 246785
rect 103606 246721 103658 246727
rect 112258 246711 112286 278004
rect 113122 272685 113150 278018
rect 113110 272679 113162 272685
rect 113110 272621 113162 272627
rect 114370 270243 114398 278018
rect 115522 270761 115550 278018
rect 116674 272833 116702 278018
rect 116662 272827 116714 272833
rect 116662 272769 116714 272775
rect 115510 270755 115562 270761
rect 115510 270697 115562 270703
rect 117922 270317 117950 278018
rect 119074 272093 119102 278018
rect 120226 272759 120254 278018
rect 120214 272753 120266 272759
rect 120214 272695 120266 272701
rect 119062 272087 119114 272093
rect 119062 272029 119114 272035
rect 120886 272087 120938 272093
rect 120886 272029 120938 272035
rect 118006 270755 118058 270761
rect 118006 270697 118058 270703
rect 117910 270311 117962 270317
rect 117910 270253 117962 270259
rect 114358 270237 114410 270243
rect 114358 270179 114410 270185
rect 118018 249375 118046 270697
rect 120898 249967 120926 272029
rect 121474 270391 121502 278018
rect 122626 273425 122654 278018
rect 123778 276494 123806 278018
rect 123682 276466 123806 276494
rect 122614 273419 122666 273425
rect 122614 273361 122666 273367
rect 123682 272907 123710 276466
rect 123766 273419 123818 273425
rect 123766 273361 123818 273367
rect 123670 272901 123722 272907
rect 123670 272843 123722 272849
rect 121462 270385 121514 270391
rect 121462 270327 121514 270333
rect 120886 249961 120938 249967
rect 120886 249903 120938 249909
rect 123778 249597 123806 273361
rect 125026 273055 125054 278018
rect 126192 278004 126686 278032
rect 125014 273049 125066 273055
rect 125014 272991 125066 272997
rect 123766 249591 123818 249597
rect 123766 249533 123818 249539
rect 126658 249523 126686 278004
rect 127330 273129 127358 278018
rect 127318 273123 127370 273129
rect 127318 273065 127370 273071
rect 128482 272981 128510 278018
rect 128470 272975 128522 272981
rect 128470 272917 128522 272923
rect 129730 271649 129758 278018
rect 130882 273499 130910 278018
rect 130870 273493 130922 273499
rect 130870 273435 130922 273441
rect 132034 273203 132062 278018
rect 132022 273197 132074 273203
rect 132022 273139 132074 273145
rect 129718 271643 129770 271649
rect 129718 271585 129770 271591
rect 132406 271643 132458 271649
rect 132406 271585 132458 271591
rect 132418 249893 132446 271585
rect 133282 270761 133310 278018
rect 133270 270755 133322 270761
rect 133270 270697 133322 270703
rect 134434 270465 134462 278018
rect 135586 273351 135614 278018
rect 135574 273345 135626 273351
rect 135574 273287 135626 273293
rect 136834 270761 136862 278018
rect 135286 270755 135338 270761
rect 135286 270697 135338 270703
rect 136822 270755 136874 270761
rect 136822 270697 136874 270703
rect 134422 270459 134474 270465
rect 134422 270401 134474 270407
rect 132406 249887 132458 249893
rect 132406 249829 132458 249835
rect 135298 249819 135326 270697
rect 137986 270539 138014 278018
rect 138166 270755 138218 270761
rect 138166 270697 138218 270703
rect 137974 270533 138026 270539
rect 137974 270475 138026 270481
rect 135286 249813 135338 249819
rect 135286 249755 135338 249761
rect 138178 249745 138206 270697
rect 139138 269915 139166 278018
rect 140400 278004 141086 278032
rect 139124 269906 139180 269915
rect 139124 269841 139180 269850
rect 138166 249739 138218 249745
rect 138166 249681 138218 249687
rect 141058 249671 141086 278004
rect 141538 270613 141566 278018
rect 142690 273425 142718 278018
rect 142678 273419 142730 273425
rect 142678 273361 142730 273367
rect 142486 273271 142538 273277
rect 142486 273213 142538 273219
rect 141526 270607 141578 270613
rect 141526 270549 141578 270555
rect 141046 249665 141098 249671
rect 141046 249607 141098 249613
rect 126646 249517 126698 249523
rect 126646 249459 126698 249465
rect 118006 249369 118058 249375
rect 118006 249311 118058 249317
rect 112246 246705 112298 246711
rect 112246 246647 112298 246653
rect 142498 216014 142526 273213
rect 142582 242635 142634 242641
rect 142582 242577 142634 242583
rect 142594 236174 142622 242577
rect 142594 236146 143102 236174
rect 143074 218887 143102 236146
rect 143062 218881 143114 218887
rect 143062 218823 143114 218829
rect 142498 215986 143102 216014
rect 50614 210741 50666 210747
rect 50614 210683 50666 210689
rect 50422 210001 50474 210007
rect 50422 209943 50474 209949
rect 143074 201571 143102 215986
rect 143062 201565 143114 201571
rect 143062 201507 143114 201513
rect 143938 190101 143966 278018
rect 145090 269207 145118 278018
rect 146242 270687 146270 278018
rect 147394 271797 147422 278018
rect 147382 271791 147434 271797
rect 147382 271733 147434 271739
rect 146230 270681 146282 270687
rect 146230 270623 146282 270629
rect 145078 269201 145130 269207
rect 145078 269143 145130 269149
rect 148642 269059 148670 278018
rect 149686 271791 149738 271797
rect 149686 271733 149738 271739
rect 148630 269053 148682 269059
rect 148630 268995 148682 269001
rect 145366 252255 145418 252261
rect 145366 252197 145418 252203
rect 143926 190095 143978 190101
rect 143926 190037 143978 190043
rect 145378 178557 145406 252197
rect 145654 249961 145706 249967
rect 145654 249903 145706 249909
rect 145462 249295 145514 249301
rect 145462 249237 145514 249243
rect 42166 178551 42218 178557
rect 42166 178493 42218 178499
rect 50326 178551 50378 178557
rect 50326 178493 50378 178499
rect 145366 178551 145418 178557
rect 145366 178493 145418 178499
rect 145474 175597 145502 249237
rect 145558 245003 145610 245009
rect 145558 244945 145610 244951
rect 145570 175671 145598 244945
rect 145666 184329 145694 249903
rect 145750 245151 145802 245157
rect 145750 245093 145802 245099
rect 145762 221773 145790 245093
rect 148532 244598 148588 244607
rect 148532 244533 148588 244542
rect 148340 242082 148396 242091
rect 148340 242017 148396 242026
rect 148244 239714 148300 239723
rect 148244 239649 148300 239658
rect 147860 232314 147916 232323
rect 147860 232249 147916 232258
rect 147874 232207 147902 232249
rect 147862 232201 147914 232207
rect 147862 232143 147914 232149
rect 146900 229946 146956 229955
rect 146900 229881 146956 229890
rect 146914 229247 146942 229881
rect 146902 229241 146954 229247
rect 146902 229183 146954 229189
rect 147188 226394 147244 226403
rect 147188 226329 147190 226338
rect 147242 226329 147244 226338
rect 147190 226297 147242 226303
rect 145750 221767 145802 221773
rect 145750 221709 145802 221715
rect 146900 221510 146956 221519
rect 146900 221445 146902 221454
rect 146954 221445 146956 221454
rect 146902 221413 146954 221419
rect 147670 219103 147722 219109
rect 147670 219045 147722 219051
rect 147682 219003 147710 219045
rect 147668 218994 147724 219003
rect 147668 218929 147724 218938
rect 147092 214110 147148 214119
rect 147092 214045 147094 214054
rect 147146 214045 147148 214054
rect 147094 214013 147146 214019
rect 146900 212926 146956 212935
rect 146900 212861 146902 212870
rect 146954 212861 146956 212870
rect 146902 212829 146954 212835
rect 147380 211742 147436 211751
rect 147380 211677 147436 211686
rect 147394 210303 147422 211677
rect 147476 210410 147532 210419
rect 147476 210345 147478 210354
rect 147530 210345 147532 210354
rect 147478 210313 147530 210319
rect 147382 210297 147434 210303
rect 147382 210239 147434 210245
rect 146900 209226 146956 209235
rect 146900 209161 146956 209170
rect 146914 207417 146942 209161
rect 147188 208042 147244 208051
rect 147188 207977 147244 207986
rect 147202 207935 147230 207977
rect 147190 207929 147242 207935
rect 147190 207871 147242 207877
rect 146902 207411 146954 207417
rect 146902 207353 146954 207359
rect 147284 206414 147340 206423
rect 147284 206349 147340 206358
rect 147298 206159 147326 206349
rect 147286 206153 147338 206159
rect 147286 206095 147338 206101
rect 147476 199606 147532 199615
rect 147476 199541 147532 199550
rect 147490 198833 147518 199541
rect 147478 198827 147530 198833
rect 147478 198769 147530 198775
rect 147380 191022 147436 191031
rect 147380 190957 147436 190966
rect 147394 190249 147422 190957
rect 147382 190243 147434 190249
rect 147382 190185 147434 190191
rect 145654 184323 145706 184329
rect 145654 184265 145706 184271
rect 147764 176518 147820 176527
rect 147764 176453 147820 176462
rect 147778 176041 147806 176453
rect 147766 176035 147818 176041
rect 147766 175977 147818 175983
rect 145558 175665 145610 175671
rect 145558 175607 145610 175613
rect 145462 175591 145514 175597
rect 145462 175533 145514 175539
rect 148258 169899 148286 239649
rect 148354 172785 148382 242017
rect 148436 234830 148492 234839
rect 148436 234765 148492 234774
rect 148342 172779 148394 172785
rect 148342 172721 148394 172727
rect 148246 169893 148298 169899
rect 148246 169835 148298 169841
rect 148450 167013 148478 234765
rect 148546 172637 148574 244533
rect 148724 243414 148780 243423
rect 148724 243349 148780 243358
rect 148628 238530 148684 238539
rect 148628 238465 148684 238474
rect 148534 172631 148586 172637
rect 148534 172573 148586 172579
rect 148642 169751 148670 238465
rect 148738 172711 148766 243349
rect 149012 240898 149068 240907
rect 149012 240833 149068 240842
rect 148916 236754 148972 236763
rect 148916 236689 148972 236698
rect 148820 233646 148876 233655
rect 148820 233581 148876 233590
rect 148834 174339 148862 233581
rect 148822 174333 148874 174339
rect 148822 174275 148874 174281
rect 148930 174136 148958 236689
rect 148834 174108 148958 174136
rect 148726 172705 148778 172711
rect 148726 172647 148778 172653
rect 148834 169825 148862 174108
rect 148916 174002 148972 174011
rect 148916 173937 148972 173946
rect 148930 172360 148958 173937
rect 149026 172563 149054 240833
rect 149108 236014 149164 236023
rect 149108 235949 149164 235958
rect 149014 172557 149066 172563
rect 149014 172499 149066 172505
rect 148930 172332 149054 172360
rect 148822 169819 148874 169825
rect 148822 169761 148874 169767
rect 148630 169745 148682 169751
rect 148630 169687 148682 169693
rect 148916 168082 148972 168091
rect 148916 168017 148972 168026
rect 148438 167007 148490 167013
rect 148438 166949 148490 166955
rect 148532 166306 148588 166315
rect 148532 166241 148588 166250
rect 148340 165566 148396 165575
rect 148340 165501 148396 165510
rect 148244 161866 148300 161875
rect 148244 161801 148300 161810
rect 147092 159498 147148 159507
rect 147092 159433 147148 159442
rect 147106 158503 147134 159433
rect 147094 158497 147146 158503
rect 147094 158439 147146 158445
rect 146900 156982 146956 156991
rect 146900 156917 146956 156926
rect 146914 156209 146942 156917
rect 146902 156203 146954 156209
rect 146902 156145 146954 156151
rect 148258 146894 148286 161801
rect 148162 146866 148286 146894
rect 147668 146178 147724 146187
rect 147668 146113 147724 146122
rect 147682 145775 147710 146113
rect 147670 145769 147722 145775
rect 147670 145711 147722 145717
rect 147668 144550 147724 144559
rect 147668 144485 147724 144494
rect 147682 144073 147710 144485
rect 147670 144067 147722 144073
rect 147670 144009 147722 144015
rect 147284 143662 147340 143671
rect 147284 143597 147340 143606
rect 147298 142519 147326 143597
rect 147286 142513 147338 142519
rect 147286 142455 147338 142461
rect 147476 142478 147532 142487
rect 147476 142413 147532 142422
rect 147490 142223 147518 142413
rect 147478 142217 147530 142223
rect 147478 142159 147530 142165
rect 147478 140367 147530 140373
rect 147478 140309 147530 140315
rect 147490 139971 147518 140309
rect 147476 139962 147532 139971
rect 147476 139897 147532 139906
rect 147668 138778 147724 138787
rect 147668 138713 147724 138722
rect 147682 138301 147710 138713
rect 147670 138295 147722 138301
rect 147670 138237 147722 138243
rect 147476 130342 147532 130351
rect 147476 130277 147532 130286
rect 147490 129717 147518 130277
rect 147478 129711 147530 129717
rect 147478 129653 147530 129659
rect 147668 127974 147724 127983
rect 147668 127909 147724 127918
rect 147682 127349 147710 127909
rect 147670 127343 147722 127349
rect 147670 127285 147722 127291
rect 148162 120985 148190 146866
rect 148354 136840 148382 165501
rect 148436 163198 148492 163207
rect 148436 163133 148492 163142
rect 148258 136812 148382 136840
rect 148258 123723 148286 136812
rect 148342 136741 148394 136747
rect 148342 136683 148394 136689
rect 148246 123717 148298 123723
rect 148246 123659 148298 123665
rect 148150 120979 148202 120985
rect 148150 120921 148202 120927
rect 148354 120911 148382 136683
rect 148450 123871 148478 163133
rect 148438 123865 148490 123871
rect 148438 123807 148490 123813
rect 148546 123797 148574 166241
rect 148724 164382 148780 164391
rect 148724 164317 148780 164326
rect 148628 160682 148684 160691
rect 148628 160617 148684 160626
rect 148642 136969 148670 160617
rect 148630 136963 148682 136969
rect 148630 136905 148682 136911
rect 148738 136840 148766 164317
rect 148820 157722 148876 157731
rect 148820 157657 148876 157666
rect 148834 155617 148862 157657
rect 148822 155611 148874 155617
rect 148822 155553 148874 155559
rect 148822 153243 148874 153249
rect 148822 153185 148874 153191
rect 148642 136812 148766 136840
rect 148834 136821 148862 153185
rect 148822 136815 148874 136821
rect 148534 123791 148586 123797
rect 148534 123733 148586 123739
rect 148642 123649 148670 136812
rect 148822 136757 148874 136763
rect 148930 136692 148958 168017
rect 149026 166810 149054 172332
rect 149122 169677 149150 235949
rect 149396 231130 149452 231139
rect 149396 231065 149452 231074
rect 149410 230505 149438 231065
rect 149398 230499 149450 230505
rect 149398 230441 149450 230447
rect 149396 228170 149452 228179
rect 149396 228105 149452 228114
rect 149410 227619 149438 228105
rect 149398 227613 149450 227619
rect 149398 227555 149450 227561
rect 149396 227430 149452 227439
rect 149396 227365 149452 227374
rect 149410 226731 149438 227365
rect 149398 226725 149450 226731
rect 149398 226667 149450 226673
rect 149396 225210 149452 225219
rect 149396 225145 149452 225154
rect 149410 224881 149438 225145
rect 149398 224875 149450 224881
rect 149398 224817 149450 224823
rect 149492 223878 149548 223887
rect 149492 223813 149548 223822
rect 149396 222694 149452 222703
rect 149396 222629 149452 222638
rect 149410 221921 149438 222629
rect 149398 221915 149450 221921
rect 149398 221857 149450 221863
rect 149506 221847 149534 223813
rect 149494 221841 149546 221847
rect 149494 221783 149546 221789
rect 149396 219734 149452 219743
rect 149396 219669 149452 219678
rect 149410 219035 149438 219669
rect 149398 219029 149450 219035
rect 149398 218971 149450 218977
rect 149396 217810 149452 217819
rect 149396 217745 149452 217754
rect 149410 216075 149438 217745
rect 149492 216626 149548 216635
rect 149492 216561 149548 216570
rect 149506 216149 149534 216561
rect 149494 216143 149546 216149
rect 149494 216085 149546 216091
rect 149398 216069 149450 216075
rect 149398 216011 149450 216017
rect 149396 214850 149452 214859
rect 149396 214785 149452 214794
rect 149410 214447 149438 214785
rect 149398 214441 149450 214447
rect 149398 214383 149450 214389
rect 149396 205674 149452 205683
rect 149396 205609 149452 205618
rect 149410 204531 149438 205609
rect 149398 204525 149450 204531
rect 149300 204490 149356 204499
rect 149398 204467 149450 204473
rect 149300 204425 149356 204434
rect 149314 201645 149342 204425
rect 149492 203306 149548 203315
rect 149492 203241 149548 203250
rect 149396 201974 149452 201983
rect 149396 201909 149452 201918
rect 149410 201793 149438 201909
rect 149398 201787 149450 201793
rect 149398 201729 149450 201735
rect 149506 201719 149534 203241
rect 149494 201713 149546 201719
rect 149494 201655 149546 201661
rect 149302 201639 149354 201645
rect 149302 201581 149354 201587
rect 149396 200790 149452 200799
rect 149396 200725 149452 200734
rect 149410 198759 149438 200725
rect 149398 198753 149450 198759
rect 149398 198695 149450 198701
rect 149492 198422 149548 198431
rect 149492 198357 149548 198366
rect 149396 197090 149452 197099
rect 149396 197025 149452 197034
rect 149410 196021 149438 197025
rect 149398 196015 149450 196021
rect 149398 195957 149450 195963
rect 149506 195947 149534 198357
rect 149494 195941 149546 195947
rect 149396 195906 149452 195915
rect 149494 195883 149546 195889
rect 149396 195841 149398 195850
rect 149450 195841 149452 195850
rect 149398 195809 149450 195815
rect 149492 194722 149548 194731
rect 149492 194657 149548 194666
rect 149396 193390 149452 193399
rect 149396 193325 149452 193334
rect 149410 193209 149438 193325
rect 149398 193203 149450 193209
rect 149398 193145 149450 193151
rect 149506 193061 149534 194657
rect 149494 193055 149546 193061
rect 149494 192997 149546 193003
rect 149396 192206 149452 192215
rect 149396 192141 149452 192150
rect 149410 190175 149438 192141
rect 149398 190169 149450 190175
rect 149398 190111 149450 190117
rect 149698 190027 149726 271733
rect 149794 269133 149822 278018
rect 150946 271575 150974 278018
rect 150934 271569 150986 271575
rect 150934 271511 150986 271517
rect 149782 269127 149834 269133
rect 149782 269069 149834 269075
rect 152194 268985 152222 278018
rect 153346 273277 153374 278018
rect 153334 273271 153386 273277
rect 153334 273213 153386 273219
rect 152374 271569 152426 271575
rect 152374 271511 152426 271517
rect 152182 268979 152234 268985
rect 152182 268921 152234 268927
rect 151318 229241 151370 229247
rect 151318 229183 151370 229189
rect 151222 226355 151274 226361
rect 151222 226297 151274 226303
rect 151126 226133 151178 226139
rect 151126 226075 151178 226081
rect 149686 190021 149738 190027
rect 149686 189963 149738 189969
rect 149396 189838 149452 189847
rect 149396 189773 149452 189782
rect 149300 187470 149356 187479
rect 149300 187405 149356 187414
rect 149204 186286 149260 186295
rect 149204 186221 149260 186230
rect 149218 180037 149246 186221
rect 149314 182923 149342 187405
rect 149410 185809 149438 189773
rect 149492 188062 149548 188071
rect 149492 187997 149548 188006
rect 149398 185803 149450 185809
rect 149398 185745 149450 185751
rect 149396 183770 149452 183779
rect 149396 183705 149452 183714
rect 149302 182917 149354 182923
rect 149302 182859 149354 182865
rect 149410 181517 149438 183705
rect 149506 182997 149534 187997
rect 149588 184510 149644 184519
rect 149588 184445 149644 184454
rect 149494 182991 149546 182997
rect 149494 182933 149546 182939
rect 149492 182586 149548 182595
rect 149492 182521 149548 182530
rect 149398 181511 149450 181517
rect 149398 181453 149450 181459
rect 149300 181402 149356 181411
rect 149300 181337 149356 181346
rect 149206 180031 149258 180037
rect 149206 179973 149258 179979
rect 149314 178631 149342 181337
rect 149506 179908 149534 182521
rect 149602 180111 149630 184445
rect 149590 180105 149642 180111
rect 149590 180047 149642 180053
rect 149506 179880 149630 179908
rect 149492 179626 149548 179635
rect 149492 179561 149548 179570
rect 149396 178886 149452 178895
rect 149396 178821 149452 178830
rect 149410 178779 149438 178821
rect 149398 178773 149450 178779
rect 149398 178715 149450 178721
rect 149506 178705 149534 179561
rect 149494 178699 149546 178705
rect 149494 178641 149546 178647
rect 149302 178625 149354 178631
rect 149302 178567 149354 178573
rect 149396 177702 149452 177711
rect 149396 177637 149452 177646
rect 149410 177299 149438 177637
rect 149398 177293 149450 177299
rect 149398 177235 149450 177241
rect 149602 175694 149630 179880
rect 149218 175666 149630 175694
rect 149218 174265 149246 175666
rect 149396 175186 149452 175195
rect 149396 175121 149452 175130
rect 149206 174259 149258 174265
rect 149206 174201 149258 174207
rect 149410 172859 149438 175121
rect 149686 174333 149738 174339
rect 149686 174275 149738 174281
rect 149398 172853 149450 172859
rect 149300 172818 149356 172827
rect 149398 172795 149450 172801
rect 149300 172753 149356 172762
rect 149204 170302 149260 170311
rect 149204 170237 149260 170246
rect 149110 169671 149162 169677
rect 149110 169613 149162 169619
rect 149026 166782 149150 166810
rect 149014 136889 149066 136895
rect 149014 136831 149066 136837
rect 148738 136664 148958 136692
rect 148738 126609 148766 136664
rect 148916 133894 148972 133903
rect 148916 133829 148972 133838
rect 148820 132710 148876 132719
rect 148820 132645 148876 132654
rect 148726 126603 148778 126609
rect 148726 126545 148778 126551
rect 148630 123643 148682 123649
rect 148630 123585 148682 123591
rect 148342 120905 148394 120911
rect 148342 120847 148394 120853
rect 147476 120574 147532 120583
rect 147476 120509 147532 120518
rect 147490 119949 147518 120509
rect 147478 119943 147530 119949
rect 147478 119885 147530 119891
rect 148436 111990 148492 111999
rect 148436 111925 148492 111934
rect 147188 108438 147244 108447
rect 147188 108373 147190 108382
rect 147242 108373 147244 108382
rect 147190 108341 147242 108347
rect 148340 107254 148396 107263
rect 148340 107189 148396 107198
rect 148244 104738 148300 104747
rect 148244 104673 148300 104682
rect 148258 86427 148286 104673
rect 148354 89239 148382 107189
rect 148450 92125 148478 111925
rect 148628 109622 148684 109631
rect 148628 109557 148630 109566
rect 148682 109557 148684 109566
rect 148630 109525 148682 109531
rect 148628 106070 148684 106079
rect 148628 106005 148684 106014
rect 148532 102370 148588 102379
rect 148532 102305 148588 102314
rect 148438 92119 148490 92125
rect 148438 92061 148490 92067
rect 148342 89233 148394 89239
rect 148342 89175 148394 89181
rect 148246 86421 148298 86427
rect 148246 86363 148298 86369
rect 148546 86353 148574 102305
rect 148642 89165 148670 106005
rect 148834 103669 148862 132645
rect 148930 126480 148958 133829
rect 149026 126683 149054 136831
rect 149122 129347 149150 166782
rect 149218 136895 149246 170237
rect 149314 155636 149342 172753
rect 149588 171042 149644 171051
rect 149588 170977 149644 170986
rect 149492 169118 149548 169127
rect 149492 169053 149548 169062
rect 149314 155608 149438 155636
rect 149300 154614 149356 154623
rect 149300 154549 149356 154558
rect 149314 152731 149342 154549
rect 149302 152725 149354 152731
rect 149302 152667 149354 152673
rect 149302 149987 149354 149993
rect 149302 149929 149354 149935
rect 149314 149887 149342 149929
rect 149300 149878 149356 149887
rect 149300 149813 149356 149822
rect 149300 148546 149356 148555
rect 149300 148481 149356 148490
rect 149314 146959 149342 148481
rect 149302 146953 149354 146959
rect 149302 146895 149354 146901
rect 149206 136889 149258 136895
rect 149206 136831 149258 136837
rect 149206 136741 149258 136747
rect 149206 136683 149258 136689
rect 149110 129341 149162 129347
rect 149110 129283 149162 129289
rect 149108 129158 149164 129167
rect 149108 129093 149164 129102
rect 149014 126677 149066 126683
rect 149014 126619 149066 126625
rect 148930 126452 149054 126480
rect 148916 121758 148972 121767
rect 148916 121693 148972 121702
rect 148822 103663 148874 103669
rect 148822 103605 148874 103611
rect 148724 103554 148780 103563
rect 148724 103489 148780 103498
rect 148630 89159 148682 89165
rect 148630 89101 148682 89107
rect 148628 86534 148684 86543
rect 148628 86469 148630 86478
rect 148682 86469 148684 86478
rect 148630 86437 148682 86443
rect 148534 86347 148586 86353
rect 148534 86289 148586 86295
rect 148738 86279 148766 103489
rect 148930 97897 148958 121693
rect 149026 106333 149054 126452
rect 149122 115255 149150 129093
rect 149218 126535 149246 136683
rect 149410 129495 149438 155608
rect 149506 153249 149534 169053
rect 149494 153243 149546 153249
rect 149494 153185 149546 153191
rect 149492 153134 149548 153143
rect 149492 153069 149548 153078
rect 149506 152805 149534 153069
rect 149494 152799 149546 152805
rect 149494 152741 149546 152747
rect 149492 150914 149548 150923
rect 149492 150849 149548 150858
rect 149506 149919 149534 150849
rect 149494 149913 149546 149919
rect 149494 149855 149546 149861
rect 149492 147362 149548 147371
rect 149492 147297 149548 147306
rect 149506 147033 149534 147297
rect 149494 147027 149546 147033
rect 149494 146969 149546 146975
rect 149602 146894 149630 170977
rect 149698 166939 149726 174275
rect 149686 166933 149738 166939
rect 149686 166875 149738 166881
rect 149684 155798 149740 155807
rect 149684 155733 149740 155742
rect 149698 155691 149726 155733
rect 149686 155685 149738 155691
rect 149686 155627 149738 155633
rect 149684 152098 149740 152107
rect 149684 152033 149740 152042
rect 149698 149845 149726 152033
rect 149686 149839 149738 149845
rect 149686 149781 149738 149787
rect 149506 146866 149630 146894
rect 149398 129489 149450 129495
rect 149398 129431 149450 129437
rect 149506 129421 149534 146866
rect 149684 141294 149740 141303
rect 149684 141229 149686 141238
rect 149738 141229 149740 141238
rect 149686 141197 149738 141203
rect 151138 140373 151166 226075
rect 151234 161241 151262 226297
rect 151330 164127 151358 229183
rect 151414 221471 151466 221477
rect 151414 221413 151466 221419
rect 151318 164121 151370 164127
rect 151318 164063 151370 164069
rect 151222 161235 151274 161241
rect 151222 161177 151274 161183
rect 151318 158497 151370 158503
rect 151318 158439 151370 158445
rect 151222 156203 151274 156209
rect 151222 156145 151274 156151
rect 151126 140367 151178 140373
rect 151126 140309 151178 140315
rect 149588 137594 149644 137603
rect 149588 137529 149644 137538
rect 149602 135415 149630 137529
rect 149684 135966 149740 135975
rect 149684 135901 149740 135910
rect 149698 135489 149726 135901
rect 149686 135483 149738 135489
rect 149686 135425 149738 135431
rect 149590 135409 149642 135415
rect 149590 135351 149642 135357
rect 149684 135078 149740 135087
rect 149684 135013 149740 135022
rect 149698 132529 149726 135013
rect 149686 132523 149738 132529
rect 149686 132465 149738 132471
rect 149684 130934 149740 130943
rect 149684 130869 149740 130878
rect 149698 129643 149726 130869
rect 149686 129637 149738 129643
rect 149686 129579 149738 129585
rect 149494 129415 149546 129421
rect 149494 129357 149546 129363
rect 149300 126642 149356 126651
rect 149300 126577 149356 126586
rect 149206 126529 149258 126535
rect 149206 126471 149258 126477
rect 149204 122498 149260 122507
rect 149204 122433 149260 122442
rect 149108 115246 149164 115255
rect 149108 115181 149164 115190
rect 149014 106327 149066 106333
rect 149014 106269 149066 106275
rect 148918 97891 148970 97897
rect 148918 97833 148970 97839
rect 149218 97823 149246 122433
rect 149314 100783 149342 126577
rect 149588 125458 149644 125467
rect 149588 125393 149644 125402
rect 149396 124274 149452 124283
rect 149396 124209 149452 124218
rect 149410 124093 149438 124209
rect 149398 124087 149450 124093
rect 149398 124029 149450 124035
rect 149492 119390 149548 119399
rect 149492 119325 149548 119334
rect 149398 118241 149450 118247
rect 149396 118206 149398 118215
rect 149450 118206 149452 118215
rect 149506 118173 149534 119325
rect 149396 118141 149452 118150
rect 149494 118167 149546 118173
rect 149494 118109 149546 118115
rect 149492 116874 149548 116883
rect 149492 116809 149548 116818
rect 149396 115690 149452 115699
rect 149396 115625 149452 115634
rect 149410 115361 149438 115625
rect 149398 115355 149450 115361
rect 149398 115297 149450 115303
rect 149506 115287 149534 116809
rect 149494 115281 149546 115287
rect 149396 115246 149452 115255
rect 149494 115223 149546 115229
rect 149396 115181 149452 115190
rect 149602 115214 149630 125393
rect 149602 115186 149726 115214
rect 149410 114640 149438 115181
rect 149410 114612 149630 114640
rect 149492 114506 149548 114515
rect 149492 114441 149548 114450
rect 149396 113174 149452 113183
rect 149396 113109 149452 113118
rect 149410 112401 149438 113109
rect 149506 113067 149534 114441
rect 149494 113061 149546 113067
rect 149494 113003 149546 113009
rect 149398 112395 149450 112401
rect 149398 112337 149450 112343
rect 149396 110954 149452 110963
rect 149396 110889 149452 110898
rect 149410 110847 149438 110889
rect 149398 110841 149450 110847
rect 149398 110783 149450 110789
rect 149602 103595 149630 114612
rect 149590 103589 149642 103595
rect 149590 103531 149642 103537
rect 149396 100890 149452 100899
rect 149396 100825 149398 100834
rect 149450 100825 149452 100834
rect 149398 100793 149450 100799
rect 149302 100777 149354 100783
rect 149302 100719 149354 100725
rect 149698 100709 149726 115186
rect 151234 112327 151262 156145
rect 151330 115213 151358 158439
rect 151426 158429 151454 221413
rect 151702 214071 151754 214077
rect 151702 214013 151754 214019
rect 151606 210371 151658 210377
rect 151606 210313 151658 210319
rect 151510 207929 151562 207935
rect 151510 207871 151562 207877
rect 151414 158423 151466 158429
rect 151414 158365 151466 158371
rect 151522 149549 151550 207871
rect 151618 152509 151646 210313
rect 151714 155543 151742 214013
rect 152086 212887 152138 212893
rect 152086 212829 152138 212835
rect 151798 210297 151850 210303
rect 151798 210239 151850 210245
rect 151702 155537 151754 155543
rect 151702 155479 151754 155485
rect 151810 152583 151838 210239
rect 151894 207411 151946 207417
rect 151894 207353 151946 207359
rect 151906 152657 151934 207353
rect 151990 206153 152042 206159
rect 151990 206095 152042 206101
rect 151894 152651 151946 152657
rect 151894 152593 151946 152599
rect 151798 152577 151850 152583
rect 151798 152519 151850 152525
rect 151606 152503 151658 152509
rect 151606 152445 151658 152451
rect 152002 149697 152030 206095
rect 152098 155469 152126 212829
rect 152386 192987 152414 271511
rect 154498 270761 154526 278018
rect 154486 270755 154538 270761
rect 154486 270697 154538 270703
rect 155446 270755 155498 270761
rect 155446 270697 155498 270703
rect 154006 249443 154058 249449
rect 154006 249385 154058 249391
rect 152374 192981 152426 192987
rect 152374 192923 152426 192929
rect 154018 181221 154046 249385
rect 154102 232201 154154 232207
rect 154102 232143 154154 232149
rect 154006 181215 154058 181221
rect 154006 181157 154058 181163
rect 154006 176035 154058 176041
rect 154006 175977 154058 175983
rect 152086 155463 152138 155469
rect 152086 155405 152138 155411
rect 151990 149691 152042 149697
rect 151990 149633 152042 149639
rect 151510 149543 151562 149549
rect 151510 149485 151562 149491
rect 154018 132455 154046 175977
rect 154114 166865 154142 232143
rect 154198 198827 154250 198833
rect 154198 198769 154250 198775
rect 154102 166859 154154 166865
rect 154102 166801 154154 166807
rect 154210 146885 154238 198769
rect 155458 192913 155486 270697
rect 155746 268763 155774 278018
rect 156898 268911 156926 278018
rect 158050 276494 158078 278018
rect 158050 276466 158174 276494
rect 156886 268905 156938 268911
rect 156886 268847 156938 268853
rect 155734 268757 155786 268763
rect 155734 268699 155786 268705
rect 156886 252329 156938 252335
rect 156886 252271 156938 252277
rect 155446 192907 155498 192913
rect 155446 192849 155498 192855
rect 154294 190243 154346 190249
rect 154294 190185 154346 190191
rect 154198 146879 154250 146885
rect 154198 146821 154250 146827
rect 154102 141255 154154 141261
rect 154102 141197 154154 141203
rect 154006 132449 154058 132455
rect 154006 132391 154058 132397
rect 153142 119943 153194 119949
rect 153142 119885 153194 119891
rect 151318 115207 151370 115213
rect 151318 115149 151370 115155
rect 151222 112321 151274 112327
rect 151222 112263 151274 112269
rect 151126 108399 151178 108405
rect 151126 108341 151178 108347
rect 149686 100703 149738 100709
rect 149686 100645 149738 100651
rect 149492 99854 149548 99863
rect 149492 99789 149548 99798
rect 149396 98670 149452 98679
rect 149396 98605 149452 98614
rect 149410 98045 149438 98605
rect 149398 98039 149450 98045
rect 149398 97981 149450 97987
rect 149506 97971 149534 99789
rect 149494 97965 149546 97971
rect 149494 97907 149546 97913
rect 149206 97817 149258 97823
rect 149206 97759 149258 97765
rect 149492 97486 149548 97495
rect 149492 97421 149548 97430
rect 149396 95710 149452 95719
rect 149396 95645 149452 95654
rect 149410 95085 149438 95645
rect 149506 95159 149534 97421
rect 149494 95153 149546 95159
rect 149494 95095 149546 95101
rect 149398 95079 149450 95085
rect 149398 95021 149450 95027
rect 149300 94970 149356 94979
rect 149300 94905 149356 94914
rect 148726 86273 148778 86279
rect 148726 86215 148778 86221
rect 148436 85350 148492 85359
rect 148436 85285 148492 85294
rect 146996 84166 147052 84175
rect 146996 84101 147052 84110
rect 147010 83615 147038 84101
rect 146998 83609 147050 83615
rect 146998 83551 147050 83557
rect 148340 81650 148396 81659
rect 148340 81585 148396 81594
rect 148354 71997 148382 81585
rect 148450 74883 148478 85285
rect 149204 82390 149260 82399
rect 149204 82325 149260 82334
rect 148820 77950 148876 77959
rect 148820 77885 148876 77894
rect 148438 74877 148490 74883
rect 148438 74819 148490 74825
rect 148342 71991 148394 71997
rect 148342 71933 148394 71939
rect 148834 69037 148862 77885
rect 149218 74809 149246 82325
rect 149314 80655 149342 94905
rect 149492 93786 149548 93795
rect 149492 93721 149548 93730
rect 149396 92602 149452 92611
rect 149396 92537 149452 92546
rect 149410 92273 149438 92537
rect 149398 92267 149450 92273
rect 149398 92209 149450 92215
rect 149506 92199 149534 93721
rect 149494 92193 149546 92199
rect 149494 92135 149546 92141
rect 149684 91418 149740 91427
rect 149684 91353 149740 91362
rect 149396 90234 149452 90243
rect 149396 90169 149452 90178
rect 149410 90127 149438 90169
rect 149398 90121 149450 90127
rect 149398 90063 149450 90069
rect 149396 89050 149452 89059
rect 149396 88985 149452 88994
rect 149302 80649 149354 80655
rect 149302 80591 149354 80597
rect 149300 80466 149356 80475
rect 149300 80401 149356 80410
rect 149206 74803 149258 74809
rect 149206 74745 149258 74751
rect 149206 74063 149258 74069
rect 149206 74005 149258 74011
rect 149108 72030 149164 72039
rect 149108 71965 149164 71974
rect 148822 69031 148874 69037
rect 148822 68973 148874 68979
rect 149122 66225 149150 71965
rect 149218 68889 149246 74005
rect 149314 73940 149342 80401
rect 149410 77769 149438 88985
rect 149492 87274 149548 87283
rect 149492 87209 149548 87218
rect 149506 86797 149534 87209
rect 149494 86791 149546 86797
rect 149494 86733 149546 86739
rect 149588 79282 149644 79291
rect 149588 79217 149644 79226
rect 149398 77763 149450 77769
rect 149398 77705 149450 77711
rect 149396 76766 149452 76775
rect 149396 76701 149452 76710
rect 149410 74069 149438 76701
rect 149492 75582 149548 75591
rect 149492 75517 149548 75526
rect 149398 74063 149450 74069
rect 149398 74005 149450 74011
rect 149314 73912 149438 73940
rect 149300 73806 149356 73815
rect 149300 73741 149356 73750
rect 149314 68963 149342 73741
rect 149410 71923 149438 73912
rect 149398 71917 149450 71923
rect 149398 71859 149450 71865
rect 149506 70980 149534 75517
rect 149602 71849 149630 79217
rect 149698 77695 149726 91353
rect 151138 89091 151166 108341
rect 153154 105149 153182 119885
rect 154114 115139 154142 141197
rect 154306 141113 154334 190185
rect 156898 181369 156926 252271
rect 156982 230499 157034 230505
rect 156982 230441 157034 230447
rect 156886 181363 156938 181369
rect 156886 181305 156938 181311
rect 156886 177293 156938 177299
rect 156886 177235 156938 177241
rect 154294 141107 154346 141113
rect 154294 141049 154346 141055
rect 156898 132381 156926 177235
rect 156994 164053 157022 230441
rect 158146 192839 158174 276466
rect 159298 271945 159326 278018
rect 160450 273573 160478 278018
rect 160438 273567 160490 273573
rect 160438 273509 160490 273515
rect 159286 271939 159338 271945
rect 159286 271881 159338 271887
rect 161602 271279 161630 278018
rect 161590 271273 161642 271279
rect 161590 271215 161642 271221
rect 162850 268689 162878 278018
rect 163894 271273 163946 271279
rect 163894 271215 163946 271221
rect 162838 268683 162890 268689
rect 162838 268625 162890 268631
rect 159862 249887 159914 249893
rect 159862 249829 159914 249835
rect 159766 226725 159818 226731
rect 159766 226667 159818 226673
rect 158134 192833 158186 192839
rect 158134 192775 158186 192781
rect 157078 190169 157130 190175
rect 157078 190111 157130 190117
rect 156982 164047 157034 164053
rect 156982 163989 157034 163995
rect 156982 142217 157034 142223
rect 156982 142159 157034 142165
rect 156886 132375 156938 132381
rect 156886 132317 156938 132323
rect 156886 124087 156938 124093
rect 156886 124029 156938 124035
rect 154102 115133 154154 115139
rect 154102 115075 154154 115081
rect 154006 109583 154058 109589
rect 154006 109525 154058 109531
rect 153142 105143 153194 105149
rect 153142 105085 153194 105091
rect 151126 89085 151178 89091
rect 151126 89027 151178 89033
rect 154018 89017 154046 109525
rect 156898 100635 156926 124029
rect 156994 115065 157022 142159
rect 157090 141039 157118 190111
rect 159778 163979 159806 226667
rect 159874 187215 159902 249829
rect 162646 249221 162698 249227
rect 162646 249163 162698 249169
rect 159958 214441 160010 214447
rect 159958 214383 160010 214389
rect 159862 187209 159914 187215
rect 159862 187151 159914 187157
rect 159766 163973 159818 163979
rect 159766 163915 159818 163921
rect 159970 155395 159998 214383
rect 160054 193203 160106 193209
rect 160054 193145 160106 193151
rect 159958 155389 160010 155395
rect 159958 155331 160010 155337
rect 159862 142513 159914 142519
rect 159862 142455 159914 142461
rect 157078 141033 157130 141039
rect 157078 140975 157130 140981
rect 159766 138295 159818 138301
rect 159766 138237 159818 138243
rect 156982 115059 157034 115065
rect 156982 115001 157034 115007
rect 156982 110841 157034 110847
rect 156982 110783 157034 110789
rect 156886 100629 156938 100635
rect 156886 100571 156938 100577
rect 156994 92051 157022 110783
rect 159778 109441 159806 138237
rect 159874 118099 159902 142455
rect 160066 140965 160094 193145
rect 162658 178483 162686 249163
rect 162742 224875 162794 224881
rect 162742 224817 162794 224823
rect 162646 178477 162698 178483
rect 162646 178419 162698 178425
rect 162754 161167 162782 224817
rect 162838 198753 162890 198759
rect 162838 198695 162890 198701
rect 162742 161161 162794 161167
rect 162742 161103 162794 161109
rect 162850 146811 162878 198695
rect 163906 192765 163934 271215
rect 164002 268837 164030 278018
rect 165154 272093 165182 278018
rect 165142 272087 165194 272093
rect 165142 272029 165194 272035
rect 166306 271723 166334 278018
rect 167554 272093 167582 278018
rect 166966 272087 167018 272093
rect 166966 272029 167018 272035
rect 167542 272087 167594 272093
rect 167542 272029 167594 272035
rect 166294 271717 166346 271723
rect 166294 271659 166346 271665
rect 163990 268831 164042 268837
rect 163990 268773 164042 268779
rect 165718 249591 165770 249597
rect 165718 249533 165770 249539
rect 165526 246779 165578 246785
rect 165526 246721 165578 246727
rect 163894 192759 163946 192765
rect 163894 192701 163946 192707
rect 165538 181295 165566 246721
rect 165622 219029 165674 219035
rect 165622 218971 165674 218977
rect 165526 181289 165578 181295
rect 165526 181231 165578 181237
rect 162934 178773 162986 178779
rect 162934 178715 162986 178721
rect 162838 146805 162890 146811
rect 162838 146747 162890 146753
rect 162742 144067 162794 144073
rect 162742 144009 162794 144015
rect 160054 140959 160106 140965
rect 160054 140901 160106 140907
rect 162646 127343 162698 127349
rect 162646 127285 162698 127291
rect 159862 118093 159914 118099
rect 159862 118035 159914 118041
rect 159862 113061 159914 113067
rect 159862 113003 159914 113009
rect 159766 109435 159818 109441
rect 159766 109377 159818 109383
rect 156982 92045 157034 92051
rect 156982 91987 157034 91993
rect 159874 91977 159902 113003
rect 162658 100561 162686 127285
rect 162754 118025 162782 144009
rect 162946 132307 162974 178715
rect 165634 158355 165662 218971
rect 165730 187141 165758 249533
rect 166978 195799 167006 272029
rect 168706 270761 168734 278018
rect 169762 278004 169872 278032
rect 168694 270755 168746 270761
rect 168694 270697 168746 270703
rect 169762 268541 169790 278004
rect 169846 270755 169898 270761
rect 169846 270697 169898 270703
rect 169750 268535 169802 268541
rect 169750 268477 169802 268483
rect 168502 249813 168554 249819
rect 168502 249755 168554 249761
rect 168406 221915 168458 221921
rect 168406 221857 168458 221863
rect 166966 195793 167018 195799
rect 166966 195735 167018 195741
rect 165814 193055 165866 193061
rect 165814 192997 165866 193003
rect 165718 187135 165770 187141
rect 165718 187077 165770 187083
rect 165718 178699 165770 178705
rect 165718 178641 165770 178647
rect 165622 158349 165674 158355
rect 165622 158291 165674 158297
rect 165526 145769 165578 145775
rect 165526 145711 165578 145717
rect 162934 132301 162986 132307
rect 162934 132243 162986 132249
rect 162742 118019 162794 118025
rect 162742 117961 162794 117967
rect 165538 117951 165566 145711
rect 165730 132233 165758 178641
rect 165826 143777 165854 192997
rect 168418 161093 168446 221857
rect 168514 187067 168542 249755
rect 168598 196015 168650 196021
rect 168598 195957 168650 195963
rect 168502 187061 168554 187067
rect 168502 187003 168554 187009
rect 168502 178625 168554 178631
rect 168502 178567 168554 178573
rect 168406 161087 168458 161093
rect 168406 161029 168458 161035
rect 168406 147027 168458 147033
rect 168406 146969 168458 146975
rect 165814 143771 165866 143777
rect 165814 143713 165866 143719
rect 165718 132227 165770 132233
rect 165718 132169 165770 132175
rect 165622 129711 165674 129717
rect 165622 129653 165674 129659
rect 165526 117945 165578 117951
rect 165526 117887 165578 117893
rect 162838 115355 162890 115361
rect 162838 115297 162890 115303
rect 162646 100555 162698 100561
rect 162646 100497 162698 100503
rect 162850 95011 162878 115297
rect 165634 103521 165662 129653
rect 168418 117877 168446 146969
rect 168514 135341 168542 178567
rect 168610 143925 168638 195957
rect 169858 195725 169886 270697
rect 171106 268615 171134 278018
rect 172272 278004 172766 278032
rect 171094 268609 171146 268615
rect 171094 268551 171146 268557
rect 171286 252181 171338 252187
rect 171286 252123 171338 252129
rect 169846 195719 169898 195725
rect 169846 195661 169898 195667
rect 171298 184255 171326 252123
rect 171478 249739 171530 249745
rect 171478 249681 171530 249687
rect 171382 221841 171434 221847
rect 171382 221783 171434 221789
rect 171286 184249 171338 184255
rect 171286 184191 171338 184197
rect 171394 161019 171422 221783
rect 171490 189953 171518 249681
rect 171574 195941 171626 195947
rect 171574 195883 171626 195889
rect 171478 189947 171530 189953
rect 171478 189889 171530 189895
rect 171478 181511 171530 181517
rect 171478 181453 171530 181459
rect 171382 161013 171434 161019
rect 171382 160955 171434 160961
rect 171382 149987 171434 149993
rect 171382 149929 171434 149935
rect 168598 143919 168650 143925
rect 168598 143861 168650 143867
rect 171286 135483 171338 135489
rect 171286 135425 171338 135431
rect 168502 135335 168554 135341
rect 168502 135277 168554 135283
rect 168502 129637 168554 129643
rect 168502 129579 168554 129585
rect 168406 117871 168458 117877
rect 168406 117813 168458 117819
rect 165718 115281 165770 115287
rect 165718 115223 165770 115229
rect 165622 103515 165674 103521
rect 165622 103457 165674 103463
rect 162838 95005 162890 95011
rect 162838 94947 162890 94953
rect 165730 94937 165758 115223
rect 168514 103447 168542 129579
rect 168598 118241 168650 118247
rect 168598 118183 168650 118189
rect 168502 103441 168554 103447
rect 168502 103383 168554 103389
rect 168214 95153 168266 95159
rect 168214 95095 168266 95101
rect 165718 94931 165770 94937
rect 165718 94873 165770 94879
rect 162454 92267 162506 92273
rect 162454 92209 162506 92215
rect 159862 91971 159914 91977
rect 159862 91913 159914 91919
rect 159766 90121 159818 90127
rect 159766 90063 159818 90069
rect 154006 89011 154058 89017
rect 154006 88953 154058 88959
rect 156502 86791 156554 86797
rect 156502 86733 156554 86739
rect 154102 86495 154154 86501
rect 154102 86437 154154 86443
rect 151126 83609 151178 83615
rect 151126 83551 151178 83557
rect 149686 77689 149738 77695
rect 149686 77631 149738 77637
rect 151138 74735 151166 83551
rect 151126 74729 151178 74735
rect 151126 74671 151178 74677
rect 154114 74661 154142 86437
rect 156514 77621 156542 86733
rect 156502 77615 156554 77621
rect 156502 77557 156554 77563
rect 159778 77547 159806 90063
rect 162466 80581 162494 92209
rect 165238 92193 165290 92199
rect 165238 92135 165290 92141
rect 162454 80575 162506 80581
rect 162454 80517 162506 80523
rect 165250 80507 165278 92135
rect 168226 83541 168254 95095
rect 168610 94863 168638 118183
rect 171298 106481 171326 135425
rect 171394 120837 171422 149929
rect 171490 135267 171518 181453
rect 171586 143851 171614 195883
rect 172738 195651 172766 278004
rect 173410 271427 173438 278018
rect 174658 272019 174686 278018
rect 174646 272013 174698 272019
rect 174646 271955 174698 271961
rect 173398 271421 173450 271427
rect 173398 271363 173450 271369
rect 175810 271205 175838 278018
rect 175798 271199 175850 271205
rect 175798 271141 175850 271147
rect 176962 268467 176990 278018
rect 176950 268461 177002 268467
rect 176950 268403 177002 268409
rect 178210 268393 178238 278018
rect 178294 271199 178346 271205
rect 178294 271141 178346 271147
rect 178198 268387 178250 268393
rect 178198 268329 178250 268335
rect 177046 249517 177098 249523
rect 177046 249459 177098 249465
rect 174166 249147 174218 249153
rect 174166 249089 174218 249095
rect 172726 195645 172778 195651
rect 172726 195587 172778 195593
rect 174178 178409 174206 249089
rect 174262 227613 174314 227619
rect 174262 227555 174314 227561
rect 174166 178403 174218 178409
rect 174166 178345 174218 178351
rect 174274 163905 174302 227555
rect 174358 216143 174410 216149
rect 174358 216085 174410 216091
rect 174262 163899 174314 163905
rect 174262 163841 174314 163847
rect 174370 155321 174398 216085
rect 174454 201787 174506 201793
rect 174454 201729 174506 201735
rect 174358 155315 174410 155321
rect 174358 155257 174410 155263
rect 174166 152799 174218 152805
rect 174166 152741 174218 152747
rect 171574 143845 171626 143851
rect 171574 143787 171626 143793
rect 171478 135261 171530 135267
rect 171478 135203 171530 135209
rect 171382 120831 171434 120837
rect 171382 120773 171434 120779
rect 174178 109367 174206 152741
rect 174262 149913 174314 149919
rect 174262 149855 174314 149861
rect 174274 122465 174302 149855
rect 174466 146737 174494 201729
rect 177058 186993 177086 249459
rect 177142 216069 177194 216075
rect 177142 216011 177194 216017
rect 177046 186987 177098 186993
rect 177046 186929 177098 186935
rect 177154 158207 177182 216011
rect 177238 201713 177290 201719
rect 177238 201655 177290 201661
rect 177142 158201 177194 158207
rect 177142 158143 177194 158149
rect 177046 155685 177098 155691
rect 177046 155627 177098 155633
rect 174454 146731 174506 146737
rect 174454 146673 174506 146679
rect 174262 122459 174314 122465
rect 174262 122401 174314 122407
rect 174262 118167 174314 118173
rect 174262 118109 174314 118115
rect 174166 109361 174218 109367
rect 174166 109303 174218 109309
rect 171286 106475 171338 106481
rect 171286 106417 171338 106423
rect 171286 100851 171338 100857
rect 171286 100793 171338 100799
rect 168598 94857 168650 94863
rect 168598 94799 168650 94805
rect 168214 83535 168266 83541
rect 168214 83477 168266 83483
rect 171298 83467 171326 100793
rect 174274 94789 174302 118109
rect 177058 112179 177086 155627
rect 177142 146953 177194 146959
rect 177142 146895 177194 146901
rect 177154 134379 177182 146895
rect 177250 146663 177278 201655
rect 178306 198537 178334 271141
rect 179362 270761 179390 278018
rect 180514 271575 180542 278018
rect 181762 271649 181790 278018
rect 181750 271643 181802 271649
rect 181750 271585 181802 271591
rect 180502 271569 180554 271575
rect 180502 271511 180554 271517
rect 182914 270761 182942 278018
rect 184066 271353 184094 278018
rect 185218 271501 185246 278018
rect 185206 271495 185258 271501
rect 185206 271437 185258 271443
rect 184054 271347 184106 271353
rect 184054 271289 184106 271295
rect 186466 270761 186494 278018
rect 187618 271205 187646 278018
rect 188770 271279 188798 278018
rect 189730 278004 190032 278032
rect 188758 271273 188810 271279
rect 188758 271215 188810 271221
rect 187606 271199 187658 271205
rect 187606 271141 187658 271147
rect 179350 270755 179402 270761
rect 179350 270697 179402 270703
rect 181366 270755 181418 270761
rect 181366 270697 181418 270703
rect 182902 270755 182954 270761
rect 182902 270697 182954 270703
rect 184246 270755 184298 270761
rect 184246 270697 184298 270703
rect 185494 270755 185546 270761
rect 185494 270697 185546 270703
rect 186454 270755 186506 270761
rect 186454 270697 186506 270703
rect 180022 249665 180074 249671
rect 180022 249607 180074 249613
rect 179926 219103 179978 219109
rect 179926 219045 179978 219051
rect 178294 198531 178346 198537
rect 178294 198473 178346 198479
rect 179938 158281 179966 219045
rect 180034 189879 180062 249607
rect 180130 201645 180158 201697
rect 180118 201639 180170 201645
rect 180118 201581 180170 201587
rect 180022 189873 180074 189879
rect 180022 189815 180074 189821
rect 179926 158275 179978 158281
rect 179926 158217 179978 158223
rect 180022 155611 180074 155617
rect 180022 155553 180074 155559
rect 177238 146657 177290 146663
rect 177238 146599 177290 146605
rect 179926 135409 179978 135415
rect 179926 135351 179978 135357
rect 177142 134373 177194 134379
rect 177142 134315 177194 134321
rect 177142 112395 177194 112401
rect 177142 112337 177194 112343
rect 177046 112173 177098 112179
rect 177046 112115 177098 112121
rect 174262 94783 174314 94789
rect 174262 94725 174314 94731
rect 177154 91903 177182 112337
rect 179938 106407 179966 135351
rect 180034 114399 180062 155553
rect 180130 149623 180158 201581
rect 181378 198611 181406 270697
rect 182806 252107 182858 252113
rect 182806 252049 182858 252055
rect 181366 198605 181418 198611
rect 181366 198547 181418 198553
rect 182818 181443 182846 252049
rect 182902 249369 182954 249375
rect 182902 249311 182954 249317
rect 182914 184181 182942 249311
rect 182998 204525 183050 204531
rect 182998 204467 183050 204473
rect 182902 184175 182954 184181
rect 182902 184117 182954 184123
rect 182806 181437 182858 181443
rect 182806 181379 182858 181385
rect 182806 172853 182858 172859
rect 182806 172795 182858 172801
rect 180214 149839 180266 149845
rect 180214 149781 180266 149787
rect 180118 149617 180170 149623
rect 180118 149559 180170 149565
rect 180226 129643 180254 149781
rect 180214 129637 180266 129643
rect 180214 129579 180266 129585
rect 182818 129569 182846 172795
rect 182902 152725 182954 152731
rect 182902 152667 182954 152673
rect 182806 129563 182858 129569
rect 182806 129505 182858 129511
rect 180022 114393 180074 114399
rect 180022 114335 180074 114341
rect 182914 112253 182942 152667
rect 183010 149771 183038 204467
rect 184258 197691 184286 270697
rect 184342 221767 184394 221773
rect 184342 221709 184394 221715
rect 184354 219595 184382 221709
rect 184340 219586 184396 219595
rect 184340 219521 184396 219530
rect 184342 218881 184394 218887
rect 184340 218846 184342 218855
rect 184394 218846 184396 218855
rect 184340 218781 184396 218790
rect 185506 198283 185534 270697
rect 185590 269867 185642 269873
rect 185590 269809 185642 269815
rect 185602 268319 185630 269809
rect 185590 268313 185642 268319
rect 185590 268255 185642 268261
rect 189730 260697 189758 278004
rect 190102 273493 190154 273499
rect 190102 273435 190154 273441
rect 190114 268171 190142 273435
rect 191170 271871 191198 278018
rect 191158 271865 191210 271871
rect 191158 271807 191210 271813
rect 192322 271797 192350 278018
rect 193570 273499 193598 278018
rect 193558 273493 193610 273499
rect 193558 273435 193610 273441
rect 194420 272274 194476 272283
rect 194420 272209 194476 272218
rect 193748 272126 193804 272135
rect 193748 272061 193804 272070
rect 192982 271939 193034 271945
rect 192982 271881 193034 271887
rect 192310 271791 192362 271797
rect 192310 271733 192362 271739
rect 192404 269314 192460 269323
rect 192404 269249 192460 269258
rect 192598 269275 192650 269281
rect 190102 268165 190154 268171
rect 190102 268107 190154 268113
rect 192418 263810 192446 269249
rect 192598 269217 192650 269223
rect 192610 263824 192638 269217
rect 192994 268245 193022 271881
rect 193076 269610 193132 269619
rect 193076 269545 193132 269554
rect 192982 268239 193034 268245
rect 192982 268181 193034 268187
rect 193090 263824 193118 269545
rect 192610 263796 192864 263824
rect 193090 263796 193344 263824
rect 193762 263810 193790 272061
rect 194228 269462 194284 269471
rect 194228 269397 194284 269406
rect 194242 263810 194270 269397
rect 194434 263824 194462 272209
rect 194722 272167 194750 278018
rect 195670 272235 195722 272241
rect 195670 272177 195722 272183
rect 194710 272161 194762 272167
rect 194710 272103 194762 272109
rect 194998 269349 195050 269355
rect 194998 269291 195050 269297
rect 195010 263824 195038 269291
rect 194434 263796 194736 263824
rect 195010 263796 195264 263824
rect 195682 263810 195710 272177
rect 195874 271945 195902 278018
rect 196628 272422 196684 272431
rect 196628 272357 196684 272366
rect 195862 271939 195914 271945
rect 195862 271881 195914 271887
rect 196148 269758 196204 269767
rect 196148 269693 196204 269702
rect 196162 263810 196190 269693
rect 196642 263810 196670 272357
rect 196822 269423 196874 269429
rect 196822 269365 196874 269371
rect 196834 263824 196862 269365
rect 197122 269281 197150 278018
rect 198274 272241 198302 278018
rect 199220 272570 199276 272579
rect 199220 272505 199276 272514
rect 199126 272383 199178 272389
rect 199126 272325 199178 272331
rect 198262 272235 198314 272241
rect 198262 272177 198314 272183
rect 198646 271717 198698 271723
rect 198646 271659 198698 271665
rect 198550 271125 198602 271131
rect 198550 271067 198602 271073
rect 198070 269719 198122 269725
rect 198070 269661 198122 269667
rect 197398 269571 197450 269577
rect 197398 269513 197450 269519
rect 197110 269275 197162 269281
rect 197110 269217 197162 269223
rect 197410 263824 197438 269513
rect 196834 263796 197088 263824
rect 197410 263796 197664 263824
rect 198082 263810 198110 269661
rect 198562 263810 198590 271067
rect 198658 269651 198686 271659
rect 198646 269645 198698 269651
rect 198646 269587 198698 269593
rect 199030 269497 199082 269503
rect 199030 269439 199082 269445
rect 199042 263810 199070 269439
rect 199138 267875 199166 272325
rect 199126 267869 199178 267875
rect 199126 267811 199178 267817
rect 199234 263824 199262 272505
rect 199426 271723 199454 278018
rect 200180 272718 200236 272727
rect 200180 272653 200236 272662
rect 199414 271717 199466 271723
rect 199414 271659 199466 271665
rect 199702 269793 199754 269799
rect 199702 269735 199754 269741
rect 199714 263824 199742 269735
rect 200194 263824 200222 272653
rect 200470 271421 200522 271427
rect 200470 271363 200522 271369
rect 200482 269725 200510 271363
rect 200470 269719 200522 269725
rect 200470 269661 200522 269667
rect 200674 269355 200702 278018
rect 201622 272309 201674 272315
rect 201622 272251 201674 272257
rect 200950 269867 201002 269873
rect 200950 269809 201002 269815
rect 200662 269349 200714 269355
rect 200662 269291 200714 269297
rect 199234 263796 199488 263824
rect 199714 263796 199968 263824
rect 200194 263796 200496 263824
rect 200962 263810 200990 269809
rect 201142 268313 201194 268319
rect 201142 268255 201194 268261
rect 201154 263824 201182 268255
rect 201634 263824 201662 272251
rect 201826 271427 201854 278018
rect 201814 271421 201866 271427
rect 201814 271363 201866 271369
rect 202870 269941 202922 269947
rect 202870 269883 202922 269889
rect 202294 267869 202346 267875
rect 202294 267811 202346 267817
rect 201154 263796 201408 263824
rect 201634 263796 201888 263824
rect 202306 263810 202334 267811
rect 202882 263810 202910 269883
rect 202978 269503 203006 278018
rect 204022 272531 204074 272537
rect 204022 272473 204074 272479
rect 203542 272457 203594 272463
rect 203542 272399 203594 272405
rect 203350 270015 203402 270021
rect 203350 269957 203402 269963
rect 202966 269497 203018 269503
rect 202966 269439 203018 269445
rect 203362 263810 203390 269957
rect 203554 263824 203582 272399
rect 204034 263824 204062 272473
rect 204130 269429 204158 278018
rect 205174 271569 205226 271575
rect 205174 271511 205226 271517
rect 204694 270089 204746 270095
rect 204694 270031 204746 270037
rect 204118 269423 204170 269429
rect 204118 269365 204170 269371
rect 203554 263796 203808 263824
rect 204034 263796 204288 263824
rect 204706 263810 204734 270031
rect 205186 269947 205214 271511
rect 205378 271131 205406 278018
rect 206038 272679 206090 272685
rect 206038 272621 206090 272627
rect 205750 272605 205802 272611
rect 205750 272547 205802 272553
rect 205366 271125 205418 271131
rect 205366 271067 205418 271073
rect 205270 270163 205322 270169
rect 205270 270105 205322 270111
rect 205174 269941 205226 269947
rect 205174 269883 205226 269889
rect 205282 263810 205310 270105
rect 205762 263810 205790 272547
rect 205942 271347 205994 271353
rect 205942 271289 205994 271295
rect 205846 271199 205898 271205
rect 205846 271141 205898 271147
rect 205858 269799 205886 271141
rect 205954 269873 205982 271289
rect 205942 269867 205994 269873
rect 205942 269809 205994 269815
rect 205846 269793 205898 269799
rect 205846 269735 205898 269741
rect 206050 263824 206078 272621
rect 206422 270237 206474 270243
rect 206422 270179 206474 270185
rect 206434 263824 206462 270179
rect 206530 269577 206558 278018
rect 207478 273567 207530 273573
rect 207478 273509 207530 273515
rect 207382 273271 207434 273277
rect 207382 273213 207434 273219
rect 207286 273049 207338 273055
rect 207286 272991 207338 272997
rect 207094 272827 207146 272833
rect 207094 272769 207146 272775
rect 206518 269571 206570 269577
rect 206518 269513 206570 269519
rect 206050 263796 206208 263824
rect 206434 263796 206688 263824
rect 207106 263810 207134 272769
rect 207298 267875 207326 272991
rect 207394 268097 207422 273213
rect 207490 268319 207518 273509
rect 207682 272315 207710 278018
rect 207862 272753 207914 272759
rect 207862 272695 207914 272701
rect 207670 272309 207722 272315
rect 207670 272251 207722 272257
rect 207574 270311 207626 270317
rect 207574 270253 207626 270259
rect 207478 268313 207530 268319
rect 207478 268255 207530 268261
rect 207382 268091 207434 268097
rect 207382 268033 207434 268039
rect 207286 267869 207338 267875
rect 207286 267811 207338 267817
rect 207586 263810 207614 270253
rect 207874 263824 207902 272695
rect 208930 272463 208958 278018
rect 209590 273419 209642 273425
rect 209590 273361 209642 273367
rect 209014 272901 209066 272907
rect 209014 272843 209066 272849
rect 208918 272457 208970 272463
rect 208918 272399 208970 272405
rect 208342 270385 208394 270391
rect 208342 270327 208394 270333
rect 208354 263824 208382 270327
rect 207874 263796 208128 263824
rect 208354 263796 208608 263824
rect 209026 263810 209054 272843
rect 209602 268139 209630 273361
rect 209782 273345 209834 273351
rect 209782 273287 209834 273293
rect 209588 268130 209644 268139
rect 209588 268065 209644 268074
rect 209794 267875 209822 273287
rect 209878 273197 209930 273203
rect 209878 273139 209930 273145
rect 209890 268023 209918 273139
rect 209974 273123 210026 273129
rect 209974 273065 210026 273071
rect 209878 268017 209930 268023
rect 209878 267959 209930 267965
rect 209494 267869 209546 267875
rect 209494 267811 209546 267817
rect 209782 267869 209834 267875
rect 209782 267811 209834 267817
rect 209506 263810 209534 267811
rect 209986 263810 210014 273065
rect 210082 272537 210110 278018
rect 210166 272975 210218 272981
rect 210166 272917 210218 272923
rect 210070 272531 210122 272537
rect 210070 272473 210122 272479
rect 210178 267968 210206 272917
rect 211234 272611 211262 278018
rect 212482 272759 212510 278018
rect 212470 272753 212522 272759
rect 212470 272695 212522 272701
rect 213634 272685 213662 278018
rect 214786 272833 214814 278018
rect 216034 272981 216062 278018
rect 217186 273055 217214 278018
rect 218338 273129 218366 278018
rect 219586 273277 219614 278018
rect 219574 273271 219626 273277
rect 219574 273213 219626 273219
rect 220738 273203 220766 278018
rect 221494 273493 221546 273499
rect 221494 273435 221546 273441
rect 220726 273197 220778 273203
rect 220726 273139 220778 273145
rect 218326 273123 218378 273129
rect 218326 273065 218378 273071
rect 217174 273049 217226 273055
rect 217174 272991 217226 272997
rect 216022 272975 216074 272981
rect 216022 272917 216074 272923
rect 214774 272827 214826 272833
rect 214774 272769 214826 272775
rect 213622 272679 213674 272685
rect 213622 272621 213674 272627
rect 211222 272605 211274 272611
rect 211222 272547 211274 272553
rect 210646 272087 210698 272093
rect 210646 272029 210698 272035
rect 210550 272013 210602 272019
rect 210550 271955 210602 271961
rect 210454 271643 210506 271649
rect 210454 271585 210506 271591
rect 210358 271495 210410 271501
rect 210358 271437 210410 271443
rect 210262 271273 210314 271279
rect 210262 271215 210314 271221
rect 210274 270095 210302 271215
rect 210370 270169 210398 271437
rect 210358 270163 210410 270169
rect 210358 270105 210410 270111
rect 210262 270089 210314 270095
rect 210262 270031 210314 270037
rect 210466 270021 210494 271585
rect 210562 270243 210590 271955
rect 210550 270237 210602 270243
rect 210550 270179 210602 270185
rect 210454 270015 210506 270021
rect 210454 269957 210506 269963
rect 210178 267940 210302 267968
rect 210658 267949 210686 272029
rect 214966 270681 215018 270687
rect 214966 270623 215018 270629
rect 213814 270607 213866 270613
rect 213814 270549 213866 270555
rect 212662 270533 212714 270539
rect 212662 270475 212714 270481
rect 211894 270459 211946 270465
rect 211894 270401 211946 270407
rect 210742 268165 210794 268171
rect 210742 268107 210794 268113
rect 210274 263824 210302 267940
rect 210646 267943 210698 267949
rect 210646 267885 210698 267891
rect 210754 263824 210782 268107
rect 211414 268017 211466 268023
rect 211414 267959 211466 267965
rect 210274 263796 210528 263824
rect 210754 263796 211008 263824
rect 211426 263810 211454 267959
rect 211906 263810 211934 270401
rect 212470 268313 212522 268319
rect 212470 268255 212522 268261
rect 212482 267875 212510 268255
rect 212374 267869 212426 267875
rect 212374 267811 212426 267817
rect 212470 267869 212522 267875
rect 212470 267811 212522 267817
rect 212386 263810 212414 267811
rect 212674 263824 212702 270475
rect 213332 269906 213388 269915
rect 213332 269841 213388 269850
rect 212674 263796 212928 263824
rect 213346 263810 213374 269841
rect 213826 263810 213854 270549
rect 214486 269201 214538 269207
rect 214486 269143 214538 269149
rect 214292 268130 214348 268139
rect 214292 268065 214348 268074
rect 214306 263810 214334 268065
rect 214498 263824 214526 269143
rect 214978 263824 215006 270623
rect 220534 269645 220586 269651
rect 220534 269587 220586 269593
rect 216214 269127 216266 269133
rect 216214 269069 216266 269075
rect 215734 269053 215786 269059
rect 215734 268995 215786 269001
rect 214498 263796 214752 263824
rect 214978 263796 215232 263824
rect 215746 263810 215774 268995
rect 216226 263810 216254 269069
rect 216694 268979 216746 268985
rect 216694 268921 216746 268927
rect 216706 263810 216734 268921
rect 218134 268905 218186 268911
rect 218134 268847 218186 268853
rect 217366 268757 217418 268763
rect 217366 268699 217418 268705
rect 216886 268091 216938 268097
rect 216886 268033 216938 268039
rect 216898 263824 216926 268033
rect 217378 263824 217406 268699
rect 216898 263796 217152 263824
rect 217378 263796 217632 263824
rect 218146 263810 218174 268847
rect 219958 268831 220010 268837
rect 219958 268773 220010 268779
rect 219286 268683 219338 268689
rect 219286 268625 219338 268631
rect 218614 268239 218666 268245
rect 218614 268181 218666 268187
rect 218626 263810 218654 268181
rect 218902 267869 218954 267875
rect 218902 267811 218954 267817
rect 218914 263824 218942 267811
rect 219298 263824 219326 268625
rect 218914 263796 219072 263824
rect 219298 263796 219552 263824
rect 219970 263810 219998 268773
rect 220546 263810 220574 269587
rect 221206 268535 221258 268541
rect 221206 268477 221258 268483
rect 221014 267943 221066 267949
rect 221014 267885 221066 267891
rect 221026 263810 221054 267885
rect 221218 263824 221246 268477
rect 221506 268319 221534 273435
rect 221686 271939 221738 271945
rect 221686 271881 221738 271887
rect 221590 271717 221642 271723
rect 221590 271659 221642 271665
rect 221494 268313 221546 268319
rect 221494 268255 221546 268261
rect 221602 268097 221630 271659
rect 221590 268091 221642 268097
rect 221590 268033 221642 268039
rect 221698 268023 221726 271881
rect 221890 271057 221918 278018
rect 221878 271051 221930 271057
rect 221878 270993 221930 270999
rect 223042 270983 223070 278018
rect 223702 271421 223754 271427
rect 223702 271363 223754 271369
rect 223030 270977 223082 270983
rect 223030 270919 223082 270925
rect 222838 270237 222890 270243
rect 222838 270179 222890 270185
rect 222358 269719 222410 269725
rect 222358 269661 222410 269667
rect 221782 268609 221834 268615
rect 221782 268551 221834 268557
rect 221686 268017 221738 268023
rect 221686 267959 221738 267965
rect 221794 263824 221822 268551
rect 221218 263796 221472 263824
rect 221794 263796 221952 263824
rect 222370 263810 222398 269661
rect 222850 263810 222878 270179
rect 223414 268461 223466 268467
rect 223414 268403 223466 268409
rect 223426 263810 223454 268403
rect 223606 268387 223658 268393
rect 223606 268329 223658 268335
rect 223618 263824 223646 268329
rect 223714 268171 223742 271363
rect 224290 270909 224318 278018
rect 224374 272235 224426 272241
rect 224374 272177 224426 272183
rect 224278 270903 224330 270909
rect 224278 270845 224330 270851
rect 224086 269941 224138 269947
rect 224086 269883 224138 269889
rect 223702 268165 223754 268171
rect 223702 268107 223754 268113
rect 224098 263824 224126 269883
rect 224386 268245 224414 272177
rect 224470 272161 224522 272167
rect 224470 272103 224522 272109
rect 224374 268239 224426 268245
rect 224374 268181 224426 268187
rect 224482 267949 224510 272103
rect 224566 271791 224618 271797
rect 224566 271733 224618 271739
rect 224470 267943 224522 267949
rect 224470 267885 224522 267891
rect 224578 267875 224606 271733
rect 225442 270835 225470 278018
rect 225910 272753 225962 272759
rect 225910 272695 225962 272701
rect 225922 272241 225950 272695
rect 225910 272235 225962 272241
rect 225910 272177 225962 272183
rect 225430 270829 225482 270835
rect 225430 270771 225482 270777
rect 226594 270761 226622 278018
rect 227842 272167 227870 278018
rect 228994 273573 229022 278018
rect 228982 273567 229034 273573
rect 228982 273509 229034 273515
rect 227830 272161 227882 272167
rect 227830 272103 227882 272109
rect 230146 272093 230174 278018
rect 230134 272087 230186 272093
rect 230134 272029 230186 272035
rect 231394 272019 231422 278018
rect 232546 272389 232574 278018
rect 233698 272759 233726 278018
rect 233686 272753 233738 272759
rect 233686 272695 233738 272701
rect 234550 272531 234602 272537
rect 234550 272473 234602 272479
rect 234358 272457 234410 272463
rect 234358 272399 234410 272405
rect 232534 272383 232586 272389
rect 232534 272325 232586 272331
rect 233878 272309 233930 272315
rect 233878 272251 233930 272257
rect 231382 272013 231434 272019
rect 231382 271955 231434 271961
rect 227158 271865 227210 271871
rect 227158 271807 227210 271813
rect 226582 270755 226634 270761
rect 226582 270697 226634 270703
rect 225526 270163 225578 270169
rect 225526 270105 225578 270111
rect 224758 270015 224810 270021
rect 224758 269957 224810 269963
rect 224566 267869 224618 267875
rect 224566 267811 224618 267817
rect 223618 263796 223872 263824
rect 224098 263796 224352 263824
rect 224770 263810 224798 269957
rect 225238 269867 225290 269873
rect 225238 269809 225290 269815
rect 225250 263810 225278 269809
rect 225538 263824 225566 270105
rect 226678 270089 226730 270095
rect 226678 270031 226730 270037
rect 226006 269793 226058 269799
rect 226006 269735 226058 269741
rect 226018 263824 226046 269735
rect 225538 263796 225792 263824
rect 226018 263796 226272 263824
rect 226690 263810 226718 270031
rect 227170 263810 227198 271807
rect 232630 271125 232682 271131
rect 232630 271067 232682 271073
rect 231958 269497 232010 269503
rect 231958 269439 232010 269445
rect 230998 269349 231050 269355
rect 230998 269291 231050 269297
rect 229558 269275 229610 269281
rect 229558 269217 229610 269223
rect 227830 268313 227882 268319
rect 227830 268255 227882 268261
rect 227638 267869 227690 267875
rect 227638 267811 227690 267817
rect 227650 263810 227678 267811
rect 227842 263824 227870 268255
rect 229078 268017 229130 268023
rect 229078 267959 229130 267965
rect 228406 267943 228458 267949
rect 228406 267885 228458 267891
rect 228418 263824 228446 267885
rect 227842 263796 228096 263824
rect 228418 263796 228672 263824
rect 229090 263810 229118 267959
rect 229570 263810 229598 269217
rect 230038 268239 230090 268245
rect 230038 268181 230090 268187
rect 230050 263810 230078 268181
rect 230518 268091 230570 268097
rect 230518 268033 230570 268039
rect 230530 264120 230558 268033
rect 230482 264092 230558 264120
rect 230482 263810 230510 264092
rect 231010 263810 231038 269291
rect 231478 268165 231530 268171
rect 231478 268107 231530 268113
rect 231490 263810 231518 268107
rect 231970 263810 231998 269439
rect 232150 269423 232202 269429
rect 232150 269365 232202 269371
rect 232162 263824 232190 269365
rect 232642 263824 232670 271067
rect 233398 269571 233450 269577
rect 233398 269513 233450 269519
rect 232162 263796 232416 263824
rect 232642 263796 232896 263824
rect 233410 263810 233438 269513
rect 233890 263810 233918 272251
rect 234370 263810 234398 272399
rect 234562 263824 234590 272473
rect 234946 272463 234974 278018
rect 235030 272605 235082 272611
rect 235030 272547 235082 272553
rect 234934 272457 234986 272463
rect 234934 272399 234986 272405
rect 235042 263824 235070 272547
rect 236098 272315 236126 278018
rect 236950 272975 237002 272981
rect 236950 272917 237002 272923
rect 236470 272901 236522 272907
rect 236470 272843 236522 272849
rect 236278 272827 236330 272833
rect 236278 272769 236330 272775
rect 236086 272309 236138 272315
rect 236086 272251 236138 272257
rect 235702 272235 235754 272241
rect 235702 272177 235754 272183
rect 234562 263796 234816 263824
rect 235042 263796 235296 263824
rect 235714 263810 235742 272177
rect 236290 263810 236318 272769
rect 236482 263824 236510 272843
rect 236962 263824 236990 272917
rect 237250 271279 237278 278018
rect 238102 273123 238154 273129
rect 238102 273065 238154 273071
rect 237622 273049 237674 273055
rect 237622 272991 237674 272997
rect 237238 271273 237290 271279
rect 237238 271215 237290 271221
rect 236482 263796 236736 263824
rect 236962 263796 237216 263824
rect 237634 263810 237662 272991
rect 238114 263810 238142 273065
rect 238498 271205 238526 278018
rect 238678 273271 238730 273277
rect 238678 273213 238730 273219
rect 238486 271199 238538 271205
rect 238486 271141 238538 271147
rect 238690 263810 238718 273213
rect 239158 273197 239210 273203
rect 239158 273139 239210 273145
rect 239170 263824 239198 273139
rect 239350 271051 239402 271057
rect 239350 270993 239402 270999
rect 239542 271051 239594 271057
rect 239542 270993 239594 270999
rect 239136 263796 239198 263824
rect 239362 263824 239390 270993
rect 239554 270761 239582 270993
rect 239650 270761 239678 278018
rect 240802 271131 240830 278018
rect 240790 271125 240842 271131
rect 240790 271067 240842 271073
rect 241954 271057 241982 278018
rect 242422 273567 242474 273573
rect 242422 273509 242474 273515
rect 242134 272161 242186 272167
rect 242134 272103 242186 272109
rect 241270 271051 241322 271057
rect 241270 270993 241322 270999
rect 241942 271051 241994 271057
rect 241942 270993 241994 270999
rect 240022 270977 240074 270983
rect 240022 270919 240074 270925
rect 239542 270755 239594 270761
rect 239542 270697 239594 270703
rect 239638 270755 239690 270761
rect 239638 270697 239690 270703
rect 239362 263796 239616 263824
rect 240034 263810 240062 270919
rect 240502 270903 240554 270909
rect 240502 270845 240554 270851
rect 240514 263810 240542 270845
rect 241078 270829 241130 270835
rect 241078 270771 241130 270777
rect 241090 263810 241118 270771
rect 241282 263824 241310 270993
rect 242146 263824 242174 272103
rect 241282 263796 241536 263824
rect 242016 263796 242174 263824
rect 242434 263810 242462 273509
rect 242902 272087 242954 272093
rect 242902 272029 242954 272035
rect 242914 263810 242942 272029
rect 243094 272013 243146 272019
rect 243094 271955 243146 271961
rect 243106 263824 243134 271955
rect 243202 270983 243230 278018
rect 244054 272753 244106 272759
rect 244054 272695 244106 272701
rect 243670 272383 243722 272389
rect 243670 272325 243722 272331
rect 243190 270977 243242 270983
rect 243190 270919 243242 270925
rect 243682 263824 243710 272325
rect 244066 263824 244094 272695
rect 244354 270909 244382 278018
rect 244822 272457 244874 272463
rect 244822 272399 244874 272405
rect 244342 270903 244394 270909
rect 244342 270845 244394 270851
rect 243106 263796 243360 263824
rect 243682 263796 243936 263824
rect 244066 263796 244368 263824
rect 244834 263810 244862 272399
rect 245302 272309 245354 272315
rect 245302 272251 245354 272257
rect 245314 263810 245342 272251
rect 245506 270835 245534 278018
rect 245590 271273 245642 271279
rect 245590 271215 245642 271221
rect 245494 270829 245546 270835
rect 245494 270771 245546 270777
rect 245602 263824 245630 271215
rect 246070 271199 246122 271205
rect 246070 271141 246122 271147
rect 246082 263824 246110 271141
rect 246754 270761 246782 278018
rect 247222 271125 247274 271131
rect 247222 271067 247274 271073
rect 246454 270755 246506 270761
rect 246454 270697 246506 270703
rect 246742 270755 246794 270761
rect 246742 270697 246794 270703
rect 246466 263824 246494 270697
rect 245602 263796 245760 263824
rect 246082 263796 246336 263824
rect 246466 263796 246768 263824
rect 247234 263810 247262 271067
rect 247702 271051 247754 271057
rect 247702 270993 247754 270999
rect 247714 263810 247742 270993
rect 247906 268393 247934 278018
rect 247990 270977 248042 270983
rect 247990 270919 248042 270925
rect 247894 268387 247946 268393
rect 247894 268329 247946 268335
rect 248002 263824 248030 270919
rect 248662 270903 248714 270909
rect 248662 270845 248714 270851
rect 248002 263796 248160 263824
rect 248674 263810 248702 270845
rect 249058 269651 249086 278018
rect 250320 278004 250526 278032
rect 249142 270829 249194 270835
rect 249142 270771 249194 270777
rect 250498 270780 250526 278004
rect 249046 269645 249098 269651
rect 249046 269587 249098 269593
rect 249154 263810 249182 270771
rect 249622 270755 249674 270761
rect 250498 270752 250718 270780
rect 249622 270697 249674 270703
rect 249634 263810 249662 270697
rect 250294 269645 250346 269651
rect 250294 269587 250346 269593
rect 249814 268387 249866 268393
rect 249814 268329 249866 268335
rect 249826 263824 249854 268329
rect 250306 263824 250334 269587
rect 250690 263824 250718 270752
rect 251458 263824 251486 278018
rect 252322 278004 252624 278032
rect 252322 263824 252350 278004
rect 253366 269127 253418 269133
rect 253366 269069 253418 269075
rect 253174 268979 253226 268985
rect 253174 268921 253226 268927
rect 252694 268091 252746 268097
rect 252694 268033 252746 268039
rect 252706 263824 252734 268033
rect 253186 263824 253214 268921
rect 249826 263796 250080 263824
rect 250306 263796 250560 263824
rect 250690 263796 250992 263824
rect 251458 263796 251568 263824
rect 252048 263796 252350 263824
rect 252480 263796 252734 263824
rect 252960 263796 253214 263824
rect 253378 263810 253406 269069
rect 253762 268097 253790 278018
rect 253942 270459 253994 270465
rect 253942 270401 253994 270407
rect 253750 268091 253802 268097
rect 253750 268033 253802 268039
rect 253954 263810 253982 270401
rect 255010 268985 255038 278018
rect 255286 270311 255338 270317
rect 255286 270253 255338 270259
rect 254998 268979 255050 268985
rect 254998 268921 255050 268927
rect 254614 268683 254666 268689
rect 254614 268625 254666 268631
rect 254626 263824 254654 268625
rect 255094 268387 255146 268393
rect 255094 268329 255146 268335
rect 255106 263824 255134 268329
rect 254400 263796 254654 263824
rect 254880 263796 255134 263824
rect 255298 263810 255326 270253
rect 255766 269793 255818 269799
rect 255766 269735 255818 269741
rect 255778 263810 255806 269735
rect 256162 269133 256190 278018
rect 257314 270465 257342 278018
rect 257302 270459 257354 270465
rect 257302 270401 257354 270407
rect 256246 269941 256298 269947
rect 256246 269883 256298 269889
rect 256150 269127 256202 269133
rect 256150 269069 256202 269075
rect 256258 263810 256286 269883
rect 257014 269127 257066 269133
rect 257014 269069 257066 269075
rect 257026 263824 257054 269069
rect 258166 268831 258218 268837
rect 258166 268773 258218 268779
rect 257686 268757 257738 268763
rect 257686 268699 257738 268705
rect 257494 268239 257546 268245
rect 257494 268181 257546 268187
rect 257506 263824 257534 268181
rect 256800 263796 257054 263824
rect 257280 263796 257534 263824
rect 257698 263810 257726 268699
rect 258178 263810 258206 268773
rect 258562 268689 258590 278018
rect 258646 269423 258698 269429
rect 258646 269365 258698 269371
rect 258550 268683 258602 268689
rect 258550 268625 258602 268631
rect 258658 263810 258686 269365
rect 259414 268979 259466 268985
rect 259414 268921 259466 268927
rect 259426 263824 259454 268921
rect 259714 268393 259742 278018
rect 260866 270317 260894 278018
rect 260854 270311 260906 270317
rect 260854 270253 260906 270259
rect 262006 270311 262058 270317
rect 262006 270253 262058 270259
rect 261814 269867 261866 269873
rect 261814 269809 261866 269815
rect 259894 269645 259946 269651
rect 259894 269587 259946 269593
rect 259702 268387 259754 268393
rect 259702 268329 259754 268335
rect 259906 263824 259934 269587
rect 260566 269275 260618 269281
rect 260566 269217 260618 269223
rect 260086 268905 260138 268911
rect 260086 268847 260138 268853
rect 259200 263796 259454 263824
rect 259680 263796 259934 263824
rect 260098 263810 260126 268847
rect 260578 263810 260606 269217
rect 261238 268535 261290 268541
rect 261238 268477 261290 268483
rect 261250 263824 261278 268477
rect 261826 263824 261854 269809
rect 261024 263796 261278 263824
rect 261600 263796 261854 263824
rect 262018 263810 262046 270253
rect 262114 269799 262142 278018
rect 262966 270533 263018 270539
rect 262966 270475 263018 270481
rect 262486 270459 262538 270465
rect 262486 270401 262538 270407
rect 262102 269793 262154 269799
rect 262102 269735 262154 269741
rect 262498 263810 262526 270401
rect 262978 263810 263006 270475
rect 263266 269947 263294 278018
rect 263254 269941 263306 269947
rect 263254 269883 263306 269889
rect 264418 269133 264446 278018
rect 264886 270237 264938 270243
rect 264886 270179 264938 270185
rect 264694 270163 264746 270169
rect 264694 270105 264746 270111
rect 264406 269127 264458 269133
rect 264406 269069 264458 269075
rect 264118 268165 264170 268171
rect 264118 268107 264170 268113
rect 263638 267943 263690 267949
rect 263638 267885 263690 267891
rect 263650 263824 263678 267885
rect 264130 263824 264158 268107
rect 264706 263824 264734 270105
rect 263424 263796 263678 263824
rect 263904 263796 264158 263824
rect 264432 263796 264734 263824
rect 264898 263810 264926 270179
rect 265366 270089 265418 270095
rect 265366 270031 265418 270037
rect 265378 263810 265406 270031
rect 265666 268245 265694 278018
rect 266518 269941 266570 269947
rect 266518 269883 266570 269889
rect 266038 269127 266090 269133
rect 266038 269069 266090 269075
rect 265654 268239 265706 268245
rect 265654 268181 265706 268187
rect 266050 263824 266078 269069
rect 266530 263824 266558 269883
rect 266818 268763 266846 278018
rect 267094 270015 267146 270021
rect 267094 269957 267146 269963
rect 266806 268757 266858 268763
rect 266806 268699 266858 268705
rect 267106 263824 267134 269957
rect 267286 269793 267338 269799
rect 267286 269735 267338 269741
rect 265824 263796 266078 263824
rect 266304 263796 266558 263824
rect 266832 263796 267134 263824
rect 267298 263810 267326 269735
rect 267970 268837 267998 278018
rect 268630 269497 268682 269503
rect 268630 269439 268682 269445
rect 267958 268831 268010 268837
rect 267958 268773 268010 268779
rect 268438 268831 268490 268837
rect 268438 268773 268490 268779
rect 267718 264095 267770 264101
rect 267718 264037 267770 264043
rect 267730 263810 267758 264037
rect 268450 263824 268478 268773
rect 268224 263796 268478 263824
rect 268642 263810 268670 269439
rect 269122 269429 269150 278018
rect 270262 272605 270314 272611
rect 270262 272547 270314 272553
rect 269686 270681 269738 270687
rect 269686 270623 269738 270629
rect 269206 269571 269258 269577
rect 269206 269513 269258 269519
rect 269110 269423 269162 269429
rect 269110 269365 269162 269371
rect 269218 263810 269246 269513
rect 269698 263810 269726 270623
rect 270274 263824 270302 272547
rect 270370 268985 270398 278018
rect 271030 273567 271082 273573
rect 271030 273509 271082 273515
rect 270550 272531 270602 272537
rect 270550 272473 270602 272479
rect 270358 268979 270410 268985
rect 270358 268921 270410 268927
rect 270144 263796 270302 263824
rect 270562 263676 270590 272473
rect 271042 263810 271070 273509
rect 271522 269651 271550 278018
rect 272278 271939 272330 271945
rect 272278 271881 272330 271887
rect 271510 269645 271562 269651
rect 271510 269587 271562 269593
rect 271510 268683 271562 268689
rect 271510 268625 271562 268631
rect 271522 263810 271550 268625
rect 272290 263824 272318 271881
rect 272674 268911 272702 278018
rect 272758 272457 272810 272463
rect 272758 272399 272810 272405
rect 272662 268905 272714 268911
rect 272662 268847 272714 268853
rect 272770 263824 272798 272399
rect 273430 272383 273482 272389
rect 273430 272325 273482 272331
rect 272950 269423 273002 269429
rect 272950 269365 273002 269371
rect 272064 263796 272318 263824
rect 272544 263796 272798 263824
rect 272962 263810 272990 269365
rect 273442 263810 273470 272325
rect 273922 269281 273950 278018
rect 274198 272975 274250 272981
rect 274198 272917 274250 272923
rect 273910 269275 273962 269281
rect 273910 269217 273962 269223
rect 274210 263824 274238 272917
rect 274678 269349 274730 269355
rect 274678 269291 274730 269297
rect 274690 263824 274718 269291
rect 275074 268541 275102 278018
rect 275350 272309 275402 272315
rect 275350 272251 275402 272257
rect 275158 272235 275210 272241
rect 275158 272177 275210 272183
rect 275062 268535 275114 268541
rect 275062 268477 275114 268483
rect 275170 263824 275198 272177
rect 273936 263796 274238 263824
rect 274464 263796 274718 263824
rect 274944 263796 275198 263824
rect 275362 263810 275390 272251
rect 276226 269873 276254 278018
rect 277078 273493 277130 273499
rect 277078 273435 277130 273441
rect 276310 272161 276362 272167
rect 276310 272103 276362 272109
rect 276214 269867 276266 269873
rect 276214 269809 276266 269815
rect 275830 269275 275882 269281
rect 275830 269217 275882 269223
rect 275842 263810 275870 269217
rect 276322 263810 276350 272103
rect 276502 269645 276554 269651
rect 276502 269587 276554 269593
rect 276514 264101 276542 269587
rect 276502 264095 276554 264101
rect 276502 264037 276554 264043
rect 277090 263824 277118 273435
rect 277474 270317 277502 278018
rect 277750 273419 277802 273425
rect 277750 273361 277802 273367
rect 277462 270311 277514 270317
rect 277462 270253 277514 270259
rect 277558 268979 277610 268985
rect 277558 268921 277610 268927
rect 277570 263824 277598 268921
rect 276864 263796 277118 263824
rect 277344 263796 277598 263824
rect 277762 263810 277790 273361
rect 278230 273271 278282 273277
rect 278230 273213 278282 273219
rect 278242 263810 278270 273213
rect 278626 270465 278654 278018
rect 279670 273345 279722 273351
rect 279670 273287 279722 273293
rect 278614 270459 278666 270465
rect 278614 270401 278666 270407
rect 279286 270459 279338 270465
rect 279286 270401 279338 270407
rect 278902 270385 278954 270391
rect 278902 270327 278954 270333
rect 278914 263824 278942 270327
rect 279298 263824 279326 270401
rect 278688 263796 278942 263824
rect 279168 263796 279326 263824
rect 279682 263810 279710 273287
rect 279778 270539 279806 278018
rect 279766 270533 279818 270539
rect 279766 270475 279818 270481
rect 280150 270533 280202 270539
rect 280150 270475 280202 270481
rect 280162 263810 280190 270475
rect 280630 269941 280682 269947
rect 280630 269883 280682 269889
rect 280642 263810 280670 269883
rect 281026 267949 281054 278018
rect 281782 274825 281834 274831
rect 281782 274767 281834 274773
rect 281302 269127 281354 269133
rect 281302 269069 281354 269075
rect 281014 267943 281066 267949
rect 281014 267885 281066 267891
rect 281314 263824 281342 269069
rect 281794 263824 281822 274767
rect 282070 269053 282122 269059
rect 282070 268995 282122 269001
rect 281088 263796 281342 263824
rect 281568 263796 281822 263824
rect 282082 263810 282110 268995
rect 282178 268171 282206 278018
rect 283030 274899 283082 274905
rect 283030 274841 283082 274847
rect 282166 268165 282218 268171
rect 282166 268107 282218 268113
rect 282550 267943 282602 267949
rect 282550 267885 282602 267891
rect 282562 263810 282590 267885
rect 283042 263810 283070 274841
rect 283330 270169 283358 278018
rect 284470 274973 284522 274979
rect 284470 274915 284522 274921
rect 284374 270607 284426 270613
rect 284374 270549 284426 270555
rect 284278 270459 284330 270465
rect 284278 270401 284330 270407
rect 284290 270359 284318 270401
rect 284386 270391 284414 270549
rect 284374 270385 284426 270391
rect 284276 270350 284332 270359
rect 284374 270327 284426 270333
rect 284276 270285 284332 270294
rect 283702 270237 283754 270243
rect 283702 270179 283754 270185
rect 283318 270163 283370 270169
rect 283318 270105 283370 270111
rect 283714 263824 283742 270179
rect 284182 270163 284234 270169
rect 284182 270105 284234 270111
rect 284194 263824 284222 270105
rect 283488 263796 283742 263824
rect 283968 263796 284222 263824
rect 284482 263810 284510 274915
rect 284578 270317 284606 278018
rect 285622 273197 285674 273203
rect 285622 273139 285674 273145
rect 284950 273049 285002 273055
rect 284950 272991 285002 272997
rect 284662 270607 284714 270613
rect 284714 270567 284798 270595
rect 284662 270549 284714 270555
rect 284770 270465 284798 270567
rect 284758 270459 284810 270465
rect 284758 270401 284810 270407
rect 284854 270385 284906 270391
rect 284660 270350 284716 270359
rect 284566 270311 284618 270317
rect 284854 270327 284906 270333
rect 284660 270285 284662 270294
rect 284566 270253 284618 270259
rect 284714 270285 284716 270294
rect 284662 270253 284714 270259
rect 284866 269947 284894 270327
rect 284854 269941 284906 269947
rect 284854 269883 284906 269889
rect 284962 263810 284990 272991
rect 285634 263824 285662 273139
rect 285730 270095 285758 278018
rect 286102 276453 286154 276459
rect 286102 276395 286154 276401
rect 285718 270089 285770 270095
rect 285718 270031 285770 270037
rect 286114 263824 286142 276395
rect 286774 273123 286826 273129
rect 286774 273065 286826 273071
rect 286294 270089 286346 270095
rect 286294 270031 286346 270037
rect 285408 263796 285662 263824
rect 285888 263796 286142 263824
rect 286306 263810 286334 270031
rect 286786 263810 286814 273065
rect 286882 269207 286910 278018
rect 287350 276305 287402 276311
rect 287350 276247 287402 276253
rect 286870 269201 286922 269207
rect 286870 269143 286922 269149
rect 286966 269201 287018 269207
rect 286966 269143 287018 269149
rect 286978 268837 287006 269143
rect 286966 268831 287018 268837
rect 286966 268773 287018 268779
rect 287362 263810 287390 276247
rect 288034 269873 288062 278018
rect 288694 276379 288746 276385
rect 288694 276321 288746 276327
rect 288502 269941 288554 269947
rect 288502 269883 288554 269889
rect 288022 269867 288074 269873
rect 288022 269809 288074 269815
rect 287926 269719 287978 269725
rect 287926 269661 287978 269667
rect 287938 263824 287966 269661
rect 288514 263824 288542 269883
rect 287808 263796 287966 263824
rect 288288 263796 288542 263824
rect 288706 263810 288734 276321
rect 289282 270021 289310 278018
rect 290326 276157 290378 276163
rect 290326 276099 290378 276105
rect 289942 272901 289994 272907
rect 289942 272843 289994 272849
rect 289270 270015 289322 270021
rect 289270 269957 289322 269963
rect 289174 268831 289226 268837
rect 289174 268773 289226 268779
rect 289186 263810 289214 268773
rect 289954 263824 289982 272843
rect 290338 263824 290366 276099
rect 290434 269799 290462 278018
rect 290614 269867 290666 269873
rect 290614 269809 290666 269815
rect 290422 269793 290474 269799
rect 290422 269735 290474 269741
rect 289728 263796 289982 263824
rect 290208 263796 290366 263824
rect 290626 263810 290654 269809
rect 291094 269793 291146 269799
rect 291094 269735 291146 269741
rect 291106 263810 291134 269735
rect 291586 269651 291614 278018
rect 291862 276231 291914 276237
rect 291862 276173 291914 276179
rect 291574 269645 291626 269651
rect 291574 269587 291626 269593
rect 291874 263824 291902 276173
rect 292246 272827 292298 272833
rect 292246 272769 292298 272775
rect 292258 263824 292286 272769
rect 292726 272753 292778 272759
rect 292726 272695 292778 272701
rect 292738 263824 292766 272695
rect 292834 269207 292862 278018
rect 293986 276494 294014 278018
rect 293890 276466 294014 276494
rect 293014 276083 293066 276089
rect 293014 276025 293066 276031
rect 292822 269201 292874 269207
rect 292822 269143 292874 269149
rect 291600 263796 291902 263824
rect 292032 263796 292286 263824
rect 292608 263796 292766 263824
rect 293026 263810 293054 276025
rect 293494 269645 293546 269651
rect 293494 269587 293546 269593
rect 293506 263810 293534 269587
rect 293890 269503 293918 276466
rect 294646 276009 294698 276015
rect 294646 275951 294698 275957
rect 293974 270607 294026 270613
rect 293974 270549 294026 270555
rect 293878 269497 293930 269503
rect 293878 269439 293930 269445
rect 293986 263810 294014 270549
rect 294658 263824 294686 275951
rect 295138 269577 295166 278018
rect 295894 275861 295946 275867
rect 295894 275803 295946 275809
rect 295414 272679 295466 272685
rect 295414 272621 295466 272627
rect 295126 269571 295178 269577
rect 295126 269513 295178 269519
rect 295222 268757 295274 268763
rect 295222 268699 295274 268705
rect 295234 263824 295262 268699
rect 294432 263796 294686 263824
rect 295008 263796 295262 263824
rect 295426 263810 295454 272621
rect 295906 263810 295934 275803
rect 296386 270687 296414 278018
rect 297334 275935 297386 275941
rect 297334 275877 297386 275883
rect 296470 275787 296522 275793
rect 296470 275729 296522 275735
rect 296374 270681 296426 270687
rect 296374 270623 296426 270629
rect 296482 263824 296510 275729
rect 296566 270607 296618 270613
rect 296566 270549 296618 270555
rect 296578 268985 296606 270549
rect 297046 269571 297098 269577
rect 297046 269513 297098 269519
rect 296566 268979 296618 268985
rect 296566 268921 296618 268927
rect 297058 263824 297086 269513
rect 296352 263796 296510 263824
rect 296832 263796 297086 263824
rect 297346 263810 297374 275877
rect 297538 272611 297566 278018
rect 297814 275639 297866 275645
rect 297814 275581 297866 275587
rect 297526 272605 297578 272611
rect 297526 272547 297578 272553
rect 297826 263810 297854 275581
rect 298294 272605 298346 272611
rect 298294 272547 298346 272553
rect 298306 263810 298334 272547
rect 298690 272537 298718 278018
rect 298966 275713 299018 275719
rect 298966 275655 299018 275661
rect 298678 272531 298730 272537
rect 298678 272473 298730 272479
rect 298978 263824 299006 275655
rect 299158 275491 299210 275497
rect 299158 275433 299210 275439
rect 298752 263796 299006 263824
rect 299170 263676 299198 275433
rect 299938 273573 299966 278018
rect 301090 276494 301118 278018
rect 300994 276466 301118 276494
rect 301954 278004 302256 278032
rect 300214 275565 300266 275571
rect 300214 275507 300266 275513
rect 299926 273567 299978 273573
rect 299926 273509 299978 273515
rect 299446 272087 299498 272093
rect 299446 272029 299498 272035
rect 299350 271865 299402 271871
rect 299350 271807 299402 271813
rect 299362 267949 299390 271807
rect 299458 269059 299486 272029
rect 299638 269497 299690 269503
rect 299638 269439 299690 269445
rect 299446 269053 299498 269059
rect 299446 268995 299498 269001
rect 299350 267943 299402 267949
rect 299350 267885 299402 267891
rect 299650 263810 299678 269439
rect 300226 263810 300254 275507
rect 300694 268905 300746 268911
rect 300694 268847 300746 268853
rect 300706 263810 300734 268847
rect 300994 268689 301022 276466
rect 301366 272531 301418 272537
rect 301366 272473 301418 272479
rect 301078 271939 301130 271945
rect 301078 271881 301130 271887
rect 301090 269133 301118 271881
rect 301078 269127 301130 269133
rect 301078 269069 301130 269075
rect 300982 268683 301034 268689
rect 300982 268625 301034 268631
rect 301378 263824 301406 272473
rect 301954 272019 301982 278004
rect 303286 275417 303338 275423
rect 303286 275359 303338 275365
rect 301942 272013 301994 272019
rect 301942 271955 301994 271961
rect 302038 268979 302090 268985
rect 302038 268921 302090 268927
rect 301846 266981 301898 266987
rect 301846 266923 301898 266929
rect 301858 263824 301886 266923
rect 301152 263796 301406 263824
rect 301632 263796 301886 263824
rect 302050 263810 302078 268921
rect 302614 268165 302666 268171
rect 302614 268107 302666 268113
rect 302626 263810 302654 268107
rect 303298 263824 303326 275359
rect 303490 272463 303518 278018
rect 304438 275343 304490 275349
rect 304438 275285 304490 275291
rect 303478 272457 303530 272463
rect 303478 272399 303530 272405
rect 303958 272457 304010 272463
rect 303958 272399 304010 272405
rect 303766 269127 303818 269133
rect 303766 269069 303818 269075
rect 303778 263824 303806 269069
rect 303072 263796 303326 263824
rect 303552 263796 303806 263824
rect 303970 263810 303998 272399
rect 304450 263810 304478 275285
rect 304642 269429 304670 278018
rect 305794 272389 305822 278018
rect 306946 272981 306974 278018
rect 307318 275269 307370 275275
rect 307318 275211 307370 275217
rect 306934 272975 306986 272981
rect 306934 272917 306986 272923
rect 307030 272975 307082 272981
rect 307030 272917 307082 272923
rect 305782 272383 305834 272389
rect 305782 272325 305834 272331
rect 306838 272383 306890 272389
rect 306838 272325 306890 272331
rect 306646 272087 306698 272093
rect 306646 272029 306698 272035
rect 306658 271871 306686 272029
rect 306646 271865 306698 271871
rect 306646 271807 306698 271813
rect 304630 269423 304682 269429
rect 304630 269365 304682 269371
rect 306358 269201 306410 269207
rect 306358 269143 306410 269149
rect 305686 269053 305738 269059
rect 305686 268995 305738 269001
rect 305014 266833 305066 266839
rect 305014 266775 305066 266781
rect 305026 263810 305054 266775
rect 305698 263824 305726 268995
rect 306166 266907 306218 266913
rect 306166 266849 306218 266855
rect 306178 263824 306206 266849
rect 305472 263796 305726 263824
rect 305952 263796 306206 263824
rect 306370 263810 306398 269143
rect 306850 263810 306878 272325
rect 307042 268763 307070 272917
rect 307030 268757 307082 268763
rect 307030 268699 307082 268705
rect 307330 263810 307358 275211
rect 308194 269355 308222 278018
rect 308374 273567 308426 273573
rect 308374 273509 308426 273515
rect 308278 269423 308330 269429
rect 308278 269365 308330 269371
rect 308182 269349 308234 269355
rect 308182 269291 308234 269297
rect 308086 266685 308138 266691
rect 308086 266627 308138 266633
rect 308098 263824 308126 266627
rect 307872 263796 308126 263824
rect 308290 263810 308318 269365
rect 308386 268837 308414 273509
rect 309346 272241 309374 278018
rect 310390 275195 310442 275201
rect 310390 275137 310442 275143
rect 309334 272235 309386 272241
rect 309334 272177 309386 272183
rect 309910 272235 309962 272241
rect 309910 272177 309962 272183
rect 308374 268831 308426 268837
rect 308374 268773 308426 268779
rect 309238 268239 309290 268245
rect 309238 268181 309290 268187
rect 308758 266759 308810 266765
rect 308758 266701 308810 266707
rect 308770 263810 308798 266701
rect 309250 263810 309278 268181
rect 309922 263824 309950 272177
rect 310402 263824 310430 275137
rect 310498 272315 310526 278018
rect 311638 275047 311690 275053
rect 311638 274989 311690 274995
rect 310486 272309 310538 272315
rect 310486 272251 310538 272257
rect 311158 269349 311210 269355
rect 311158 269291 311210 269297
rect 310678 266611 310730 266617
rect 310678 266553 310730 266559
rect 309696 263796 309950 263824
rect 310272 263796 310430 263824
rect 310690 263810 310718 266553
rect 311170 263810 311198 269291
rect 311650 263810 311678 274989
rect 311746 269281 311774 278018
rect 312790 272235 312842 272241
rect 312790 272177 312842 272183
rect 311734 269275 311786 269281
rect 311734 269217 311786 269223
rect 312310 268313 312362 268319
rect 312310 268255 312362 268261
rect 312322 263824 312350 268255
rect 312802 263824 312830 272177
rect 312898 272167 312926 278018
rect 314050 273499 314078 278018
rect 314710 275121 314762 275127
rect 314710 275063 314762 275069
rect 314038 273493 314090 273499
rect 314038 273435 314090 273441
rect 312886 272161 312938 272167
rect 312886 272103 312938 272109
rect 314230 269275 314282 269281
rect 314230 269217 314282 269223
rect 313558 266537 313610 266543
rect 313558 266479 313610 266485
rect 313078 266463 313130 266469
rect 313078 266405 313130 266411
rect 312096 263796 312350 263824
rect 312672 263796 312830 263824
rect 313090 263810 313118 266405
rect 313570 263810 313598 266479
rect 314242 263824 314270 269217
rect 314722 263824 314750 275063
rect 314016 263796 314270 263824
rect 314496 263796 314750 263824
rect 314914 263810 314942 278245
rect 316630 278229 316682 278235
rect 316630 278171 316682 278177
rect 411862 278229 411914 278235
rect 411914 278177 412176 278180
rect 411862 278171 412176 278177
rect 315298 270613 315326 278018
rect 315958 274233 316010 274239
rect 315958 274175 316010 274181
rect 315478 272161 315530 272167
rect 315478 272103 315530 272109
rect 315286 270607 315338 270613
rect 315286 270549 315338 270555
rect 315490 263810 315518 272103
rect 315970 263810 315998 274175
rect 316450 273425 316478 278018
rect 316438 273419 316490 273425
rect 316438 273361 316490 273367
rect 316642 263824 316670 278171
rect 319510 278155 319562 278161
rect 411874 278152 412176 278171
rect 418978 278161 419280 278180
rect 418966 278155 419280 278161
rect 319510 278097 319562 278103
rect 419018 278152 419280 278155
rect 418966 278097 419018 278103
rect 317302 274159 317354 274165
rect 317302 274101 317354 274107
rect 317110 268387 317162 268393
rect 317110 268329 317162 268335
rect 317122 263824 317150 268329
rect 316416 263796 316670 263824
rect 316896 263796 317150 263824
rect 317314 263810 317342 274101
rect 317602 273277 317630 278018
rect 317878 277785 317930 277791
rect 317878 277727 317930 277733
rect 317590 273271 317642 273277
rect 317590 273213 317642 273219
rect 317890 263810 317918 277727
rect 318358 271273 318410 271279
rect 318358 271215 318410 271221
rect 318370 263810 318398 271215
rect 318850 270465 318878 278018
rect 318838 270459 318890 270465
rect 318838 270401 318890 270407
rect 319030 265501 319082 265507
rect 319030 265443 319082 265449
rect 319042 263824 319070 265443
rect 319522 263824 319550 278097
rect 320950 278081 321002 278087
rect 422518 278081 422570 278087
rect 320950 278023 321002 278029
rect 320002 270317 320030 278018
rect 320182 274307 320234 274313
rect 320182 274249 320234 274255
rect 319990 270311 320042 270317
rect 319990 270253 320042 270259
rect 319702 268461 319754 268467
rect 319702 268403 319754 268409
rect 318816 263796 319070 263824
rect 319296 263796 319550 263824
rect 319714 263810 319742 268403
rect 320194 263810 320222 274249
rect 320962 263824 320990 278023
rect 321154 273351 321182 278018
rect 322102 277859 322154 277865
rect 322102 277801 322154 277807
rect 321142 273345 321194 273351
rect 321142 273287 321194 273293
rect 321430 271347 321482 271353
rect 321430 271289 321482 271295
rect 321442 263824 321470 271289
rect 321622 265649 321674 265655
rect 321622 265591 321674 265597
rect 320736 263796 320990 263824
rect 321216 263796 321470 263824
rect 321634 263810 321662 265591
rect 322114 263810 322142 277801
rect 322402 270539 322430 278018
rect 323350 274381 323402 274387
rect 323350 274323 323402 274329
rect 322390 270533 322442 270539
rect 322390 270475 322442 270481
rect 322582 268535 322634 268541
rect 322582 268477 322634 268483
rect 322594 263810 322622 268477
rect 323362 263824 323390 274323
rect 323554 270391 323582 278018
rect 323830 277933 323882 277939
rect 323830 277875 323882 277881
rect 323542 270385 323594 270391
rect 323542 270327 323594 270333
rect 323842 263824 323870 277875
rect 324706 271945 324734 278018
rect 325858 274831 325886 278018
rect 326422 276527 326474 276533
rect 326422 276469 326474 276475
rect 325846 274825 325898 274831
rect 325846 274767 325898 274773
rect 325942 274455 325994 274461
rect 325942 274397 325994 274403
rect 324694 271939 324746 271945
rect 324694 271881 324746 271887
rect 324022 271421 324074 271427
rect 324022 271363 324074 271369
rect 323136 263796 323390 263824
rect 323616 263796 323870 263824
rect 324034 263810 324062 271363
rect 325750 268609 325802 268615
rect 325750 268551 325802 268557
rect 324502 265723 324554 265729
rect 324502 265665 324554 265671
rect 324514 263810 324542 265665
rect 324982 264095 325034 264101
rect 324982 264037 325034 264043
rect 324994 263810 325022 264037
rect 325762 263824 325790 268551
rect 325536 263796 325790 263824
rect 325954 263810 325982 274397
rect 326434 263810 326462 276469
rect 326806 274011 326858 274017
rect 326806 273953 326858 273959
rect 326818 268911 326846 273953
rect 327106 272019 327134 278018
rect 328258 272093 328286 278018
rect 329302 277711 329354 277717
rect 329302 277653 329354 277659
rect 328822 274529 328874 274535
rect 328822 274471 328874 274477
rect 328246 272087 328298 272093
rect 328246 272029 328298 272035
rect 327094 272013 327146 272019
rect 327094 271955 327146 271961
rect 326902 271495 326954 271501
rect 326902 271437 326954 271443
rect 326806 268905 326858 268911
rect 326806 268847 326858 268853
rect 326914 263810 326942 271437
rect 328342 268683 328394 268689
rect 328342 268625 328394 268631
rect 327574 265797 327626 265803
rect 327574 265739 327626 265745
rect 327586 263824 327614 265739
rect 328054 264761 328106 264767
rect 328054 264703 328106 264709
rect 328066 263824 328094 264703
rect 327360 263796 327614 263824
rect 327840 263796 328094 263824
rect 328354 263810 328382 268625
rect 328834 263810 328862 274471
rect 329314 263810 329342 277653
rect 329410 274905 329438 278018
rect 329398 274899 329450 274905
rect 329398 274841 329450 274847
rect 330454 274603 330506 274609
rect 330454 274545 330506 274551
rect 329974 271569 330026 271575
rect 329974 271511 330026 271517
rect 329986 263824 330014 271511
rect 330466 263824 330494 274545
rect 330658 270243 330686 278018
rect 331222 273715 331274 273721
rect 331222 273657 331274 273663
rect 330646 270237 330698 270243
rect 330646 270179 330698 270185
rect 331234 268985 331262 273657
rect 331810 270169 331838 278018
rect 332374 277637 332426 277643
rect 332374 277579 332426 277585
rect 331798 270163 331850 270169
rect 331798 270105 331850 270111
rect 331222 268979 331274 268985
rect 331222 268921 331274 268927
rect 331222 268757 331274 268763
rect 331222 268699 331274 268705
rect 331126 264687 331178 264693
rect 331126 264629 331178 264635
rect 331138 263824 331166 264629
rect 329760 263796 330014 263824
rect 330240 263796 330494 263824
rect 330768 263796 331166 263824
rect 331234 263810 331262 268699
rect 331894 265871 331946 265877
rect 331894 265813 331946 265819
rect 331906 263824 331934 265813
rect 332386 263824 332414 277579
rect 332962 274979 332990 278018
rect 332950 274973 333002 274979
rect 332950 274915 333002 274921
rect 333142 274677 333194 274683
rect 333142 274619 333194 274625
rect 332566 271643 332618 271649
rect 332566 271585 332618 271591
rect 331680 263796 331934 263824
rect 332160 263796 332414 263824
rect 332578 263810 332606 271585
rect 333154 263810 333182 274619
rect 334210 273055 334238 278018
rect 334966 277563 335018 277569
rect 334966 277505 335018 277511
rect 334294 273863 334346 273869
rect 334294 273805 334346 273811
rect 334198 273049 334250 273055
rect 334198 272991 334250 272997
rect 334102 270903 334154 270909
rect 334102 270845 334154 270851
rect 334114 270095 334142 270845
rect 334102 270089 334154 270095
rect 334102 270031 334154 270037
rect 334306 269133 334334 273805
rect 334294 269127 334346 269133
rect 334294 269069 334346 269075
rect 334294 268831 334346 268837
rect 334294 268773 334346 268779
rect 333622 268017 333674 268023
rect 333622 267959 333674 267965
rect 333634 263810 333662 267959
rect 334306 263824 334334 268773
rect 334774 265945 334826 265951
rect 334774 265887 334826 265893
rect 334786 263824 334814 265887
rect 334080 263796 334334 263824
rect 334560 263796 334814 263824
rect 334978 263810 335006 277505
rect 335362 273203 335390 278018
rect 336514 276459 336542 278018
rect 336502 276453 336554 276459
rect 336502 276395 336554 276401
rect 336022 274751 336074 274757
rect 336022 274693 336074 274699
rect 335350 273197 335402 273203
rect 335350 273139 335402 273145
rect 335446 271717 335498 271723
rect 335446 271659 335498 271665
rect 335458 263810 335486 271659
rect 336034 263810 336062 274693
rect 337762 270909 337790 278018
rect 337846 277489 337898 277495
rect 337846 277431 337898 277437
rect 337750 270903 337802 270909
rect 337750 270845 337802 270851
rect 336886 268905 336938 268911
rect 336886 268847 336938 268853
rect 336694 267943 336746 267949
rect 336694 267885 336746 267891
rect 336706 263824 336734 267885
rect 336480 263796 336734 263824
rect 336898 263824 336926 268847
rect 337366 266019 337418 266025
rect 337366 265961 337418 265967
rect 336898 263796 336960 263824
rect 337378 263810 337406 265961
rect 337858 263810 337886 277431
rect 338914 273129 338942 278018
rect 340066 276311 340094 278018
rect 341014 277415 341066 277421
rect 341014 277357 341066 277363
rect 340054 276305 340106 276311
rect 340054 276247 340106 276253
rect 339094 274825 339146 274831
rect 339094 274767 339146 274773
rect 338902 273123 338954 273129
rect 338902 273065 338954 273071
rect 338614 271791 338666 271797
rect 338614 271733 338666 271739
rect 337942 270755 337994 270761
rect 337942 270697 337994 270703
rect 337954 269947 337982 270697
rect 337942 269941 337994 269947
rect 337942 269883 337994 269889
rect 338626 263824 338654 271733
rect 339106 263824 339134 274767
rect 339766 268979 339818 268985
rect 339766 268921 339818 268927
rect 339286 267869 339338 267875
rect 339286 267811 339338 267817
rect 338400 263796 338654 263824
rect 338880 263796 339134 263824
rect 339298 263810 339326 267811
rect 339778 263810 339806 268921
rect 340246 266093 340298 266099
rect 340246 266035 340298 266041
rect 340258 263810 340286 266035
rect 341026 263824 341054 277357
rect 341314 270761 341342 278018
rect 341684 274494 341740 274503
rect 341684 274429 341740 274438
rect 341494 271865 341546 271871
rect 341494 271807 341546 271813
rect 341302 270755 341354 270761
rect 341302 270697 341354 270703
rect 341506 263824 341534 271807
rect 340800 263796 341054 263824
rect 341280 263796 341534 263824
rect 341698 263810 341726 274429
rect 342166 273937 342218 273943
rect 342166 273879 342218 273885
rect 342178 269207 342206 273879
rect 342466 270021 342494 278018
rect 343618 276385 343646 278018
rect 343894 277341 343946 277347
rect 343894 277283 343946 277289
rect 343606 276379 343658 276385
rect 343606 276321 343658 276327
rect 342742 270977 342794 270983
rect 342742 270919 342794 270925
rect 342454 270015 342506 270021
rect 342454 269957 342506 269963
rect 342754 269873 342782 270919
rect 342742 269867 342794 269873
rect 342742 269809 342794 269815
rect 342166 269201 342218 269207
rect 342166 269143 342218 269149
rect 342646 269127 342698 269133
rect 342646 269069 342698 269075
rect 342166 268091 342218 268097
rect 342166 268033 342218 268039
rect 342178 263810 342206 268033
rect 342658 263810 342686 269069
rect 343318 266167 343370 266173
rect 343318 266109 343370 266115
rect 343330 263824 343358 266109
rect 343906 263824 343934 277283
rect 344566 274899 344618 274905
rect 344566 274841 344618 274847
rect 344086 271939 344138 271945
rect 344086 271881 344138 271887
rect 343104 263796 343358 263824
rect 343632 263796 343934 263824
rect 344098 263810 344126 271881
rect 344578 263810 344606 274841
rect 344770 273573 344798 278018
rect 344758 273567 344810 273573
rect 344758 273509 344810 273515
rect 346018 272907 346046 278018
rect 347170 276163 347198 278018
rect 347158 276157 347210 276163
rect 347158 276099 347210 276105
rect 347636 274642 347692 274651
rect 347636 274577 347692 274586
rect 347062 273789 347114 273795
rect 347062 273731 347114 273737
rect 346006 272901 346058 272907
rect 346006 272843 346058 272849
rect 346966 272087 347018 272093
rect 346966 272029 347018 272035
rect 346486 272013 346538 272019
rect 346486 271955 346538 271961
rect 345430 270607 345482 270613
rect 345430 270549 345482 270555
rect 345238 269201 345290 269207
rect 345238 269143 345290 269149
rect 345250 263824 345278 269143
rect 345024 263796 345278 263824
rect 345442 263676 345470 270549
rect 346006 266241 346058 266247
rect 346006 266183 346058 266189
rect 346018 263810 346046 266183
rect 346498 263810 346526 271955
rect 346978 263810 347006 272029
rect 347074 268245 347102 273731
rect 347062 268239 347114 268245
rect 347062 268181 347114 268187
rect 347650 263824 347678 274577
rect 348322 270983 348350 278018
rect 348502 274085 348554 274091
rect 348502 274027 348554 274033
rect 348310 270977 348362 270983
rect 348310 270919 348362 270925
rect 348406 270533 348458 270539
rect 348406 270475 348458 270481
rect 348118 270459 348170 270465
rect 348118 270401 348170 270407
rect 348130 263824 348158 270401
rect 347424 263796 347678 263824
rect 347904 263796 348158 263824
rect 348418 263810 348446 270475
rect 348514 268319 348542 274027
rect 349462 273493 349514 273499
rect 349462 273435 349514 273441
rect 348502 268313 348554 268319
rect 348502 268255 348554 268261
rect 348886 266315 348938 266321
rect 348886 266257 348938 266263
rect 348898 263810 348926 266257
rect 349474 263824 349502 273435
rect 349570 269799 349598 278018
rect 350722 276237 350750 278018
rect 350710 276231 350762 276237
rect 350710 276173 350762 276179
rect 350228 274790 350284 274799
rect 350228 274725 350284 274734
rect 350038 273567 350090 273573
rect 350038 273509 350090 273515
rect 349558 269793 349610 269799
rect 349558 269735 349610 269741
rect 350050 263824 350078 273509
rect 349344 263796 349502 263824
rect 349824 263796 350078 263824
rect 350242 263810 350270 274725
rect 351874 272833 351902 278018
rect 352438 273419 352490 273425
rect 352438 273361 352490 273367
rect 351862 272827 351914 272833
rect 351862 272769 351914 272775
rect 351382 270829 351434 270835
rect 351382 270771 351434 270777
rect 350710 270385 350762 270391
rect 350710 270327 350762 270333
rect 350722 263810 350750 270327
rect 351286 270311 351338 270317
rect 351286 270253 351338 270259
rect 351298 263810 351326 270253
rect 351394 269651 351422 270771
rect 351382 269645 351434 269651
rect 351382 269587 351434 269593
rect 351382 268017 351434 268023
rect 351382 267959 351434 267965
rect 351394 264471 351422 267959
rect 351958 267795 352010 267801
rect 351958 267737 352010 267743
rect 351382 264465 351434 264471
rect 351382 264407 351434 264413
rect 351970 263824 351998 267737
rect 352450 263824 352478 273361
rect 352630 273345 352682 273351
rect 352630 273287 352682 273293
rect 351744 263796 351998 263824
rect 352224 263796 352478 263824
rect 352642 263810 352670 273287
rect 353122 272759 353150 278018
rect 354274 276089 354302 278018
rect 354262 276083 354314 276089
rect 354262 276025 354314 276031
rect 353396 274938 353452 274947
rect 353396 274873 353452 274882
rect 353110 272753 353162 272759
rect 353110 272695 353162 272701
rect 353410 263824 353438 274873
rect 355030 273197 355082 273203
rect 355030 273139 355082 273145
rect 354070 270237 354122 270243
rect 354070 270179 354122 270185
rect 353686 270163 353738 270169
rect 353686 270105 353738 270111
rect 353136 263796 353438 263824
rect 353698 263810 353726 270105
rect 354082 264120 354110 270179
rect 354262 267943 354314 267949
rect 354262 267885 354314 267891
rect 354274 264619 354302 267885
rect 354838 267721 354890 267727
rect 354838 267663 354890 267669
rect 354262 264613 354314 264619
rect 354262 264555 354314 264561
rect 354082 264092 354158 264120
rect 354130 263810 354158 264092
rect 354850 263824 354878 267663
rect 354624 263796 354878 263824
rect 355042 263810 355070 273139
rect 355426 270835 355454 278018
rect 356182 274973 356234 274979
rect 356182 274915 356234 274921
rect 355510 273271 355562 273277
rect 355510 273213 355562 273219
rect 355414 270829 355466 270835
rect 355414 270771 355466 270777
rect 355522 263810 355550 273213
rect 356194 263824 356222 274915
rect 356674 270687 356702 278018
rect 357826 276015 357854 278018
rect 357814 276009 357866 276015
rect 357814 275951 357866 275957
rect 358582 273123 358634 273129
rect 358582 273065 358634 273071
rect 357910 271199 357962 271205
rect 357910 271141 357962 271147
rect 356662 270681 356714 270687
rect 356662 270623 356714 270629
rect 356758 270089 356810 270095
rect 356758 270031 356810 270037
rect 356770 263824 356798 270031
rect 356950 270015 357002 270021
rect 356950 269957 357002 269963
rect 355968 263796 356222 263824
rect 356544 263796 356798 263824
rect 356962 263810 356990 269957
rect 357430 267647 357482 267653
rect 357430 267589 357482 267595
rect 357442 263810 357470 267589
rect 357922 263810 357950 271141
rect 358594 263824 358622 273065
rect 358978 272981 359006 278018
rect 359158 276453 359210 276459
rect 359158 276395 359210 276401
rect 358966 272975 359018 272981
rect 358966 272917 359018 272923
rect 359170 263824 359198 276395
rect 360226 272685 360254 278018
rect 361378 275867 361406 278018
rect 361750 276379 361802 276385
rect 361750 276321 361802 276327
rect 361366 275861 361418 275867
rect 361366 275803 361418 275809
rect 360982 273049 361034 273055
rect 360982 272991 361034 272997
rect 360214 272679 360266 272685
rect 360214 272621 360266 272627
rect 359830 269941 359882 269947
rect 359830 269883 359882 269889
rect 359350 269867 359402 269873
rect 359350 269809 359402 269815
rect 358368 263796 358622 263824
rect 358944 263796 359198 263824
rect 359362 263810 359390 269809
rect 359446 268091 359498 268097
rect 359446 268033 359498 268039
rect 359458 264841 359486 268033
rect 359446 264835 359498 264841
rect 359446 264777 359498 264783
rect 359842 263810 359870 269883
rect 360406 267869 360458 267875
rect 360406 267811 360458 267817
rect 360310 267573 360362 267579
rect 360310 267515 360362 267521
rect 360322 263810 360350 267515
rect 360418 264545 360446 267811
rect 360406 264539 360458 264545
rect 360406 264481 360458 264487
rect 360994 263824 361022 272991
rect 361270 272975 361322 272981
rect 361270 272917 361322 272923
rect 360768 263796 361022 263824
rect 361282 263810 361310 272917
rect 361762 263810 361790 276321
rect 362530 275793 362558 278018
rect 362518 275787 362570 275793
rect 362518 275729 362570 275735
rect 363574 272901 363626 272907
rect 363574 272843 363626 272849
rect 362806 269793 362858 269799
rect 362806 269735 362858 269741
rect 362230 269719 362282 269725
rect 362230 269661 362282 269667
rect 362242 263810 362270 269661
rect 362818 263824 362846 269735
rect 363382 267499 363434 267505
rect 363382 267441 363434 267447
rect 363394 263824 363422 267441
rect 362688 263796 362846 263824
rect 363168 263796 363422 263824
rect 363586 263810 363614 272843
rect 363682 269577 363710 278018
rect 364630 276305 364682 276311
rect 364630 276247 364682 276253
rect 364150 272827 364202 272833
rect 364150 272769 364202 272775
rect 363670 269571 363722 269577
rect 363670 269513 363722 269519
rect 364162 263810 364190 272769
rect 364642 263810 364670 276247
rect 364930 275941 364958 278018
rect 364918 275935 364970 275941
rect 364918 275877 364970 275883
rect 366082 275645 366110 278018
rect 366070 275639 366122 275645
rect 366070 275581 366122 275587
rect 366550 272753 366602 272759
rect 366550 272695 366602 272701
rect 365302 269645 365354 269651
rect 365302 269587 365354 269593
rect 365314 263824 365342 269587
rect 365686 269571 365738 269577
rect 365686 269513 365738 269519
rect 365698 263824 365726 269513
rect 365974 267425 366026 267431
rect 365974 267367 366026 267373
rect 365088 263796 365342 263824
rect 365568 263796 365726 263824
rect 365986 263810 366014 267367
rect 366562 263810 366590 272695
rect 367126 272679 367178 272685
rect 367126 272621 367178 272627
rect 367138 263824 367166 272621
rect 367234 272611 367262 278018
rect 367702 276231 367754 276237
rect 367702 276173 367754 276179
rect 367222 272605 367274 272611
rect 367222 272547 367274 272553
rect 367714 263824 367742 276173
rect 368482 275719 368510 278018
rect 368470 275713 368522 275719
rect 368470 275655 368522 275661
rect 369634 275497 369662 278018
rect 370294 276157 370346 276163
rect 370294 276099 370346 276105
rect 369622 275491 369674 275497
rect 369622 275433 369674 275439
rect 370100 271830 370156 271839
rect 370100 271765 370156 271774
rect 369620 271682 369676 271691
rect 369620 271617 369676 271626
rect 368372 269166 368428 269175
rect 368372 269101 368428 269110
rect 367892 269018 367948 269027
rect 367892 268953 367948 268962
rect 367008 263796 367166 263824
rect 367488 263796 367742 263824
rect 367906 263810 367934 268953
rect 368386 263810 368414 269101
rect 368950 267351 369002 267357
rect 368950 267293 369002 267299
rect 368962 263810 368990 267293
rect 369634 263824 369662 271617
rect 370114 263824 370142 271765
rect 369408 263796 369662 263824
rect 369888 263796 370142 263824
rect 370306 263810 370334 276099
rect 370786 269503 370814 278018
rect 371062 276083 371114 276089
rect 371062 276025 371114 276031
rect 370774 269497 370826 269503
rect 370774 269439 370826 269445
rect 371074 263824 371102 276025
rect 371926 276009 371978 276015
rect 371926 275951 371978 275957
rect 371254 270681 371306 270687
rect 371254 270623 371306 270629
rect 370800 263796 371102 263824
rect 371266 263810 371294 270623
rect 371938 263824 371966 275951
rect 372034 275571 372062 278018
rect 372022 275565 372074 275571
rect 372022 275507 372074 275513
rect 373186 274017 373214 278018
rect 373846 277267 373898 277273
rect 373846 277209 373898 277215
rect 373462 275935 373514 275941
rect 373462 275877 373514 275883
rect 373174 274011 373226 274017
rect 373174 273953 373226 273959
rect 372694 272605 372746 272611
rect 372694 272547 372746 272553
rect 372502 267277 372554 267283
rect 372502 267219 372554 267225
rect 372514 263824 372542 267219
rect 371808 263796 371966 263824
rect 372288 263796 372542 263824
rect 372706 263810 372734 272547
rect 373474 263824 373502 275877
rect 373858 263824 373886 277209
rect 374338 272537 374366 278018
rect 375298 278004 375600 278032
rect 375094 277193 375146 277199
rect 375094 277135 375146 277141
rect 374614 275861 374666 275867
rect 374614 275803 374666 275809
rect 374518 272753 374570 272759
rect 374518 272695 374570 272701
rect 374530 272611 374558 272695
rect 374518 272605 374570 272611
rect 374518 272547 374570 272553
rect 374326 272531 374378 272537
rect 374326 272473 374378 272479
rect 374324 270498 374380 270507
rect 374324 270433 374380 270442
rect 374338 263824 374366 270433
rect 373200 263796 373502 263824
rect 373632 263796 373886 263824
rect 374208 263796 374366 263824
rect 374626 263810 374654 275803
rect 374998 273123 375050 273129
rect 374998 273065 375050 273071
rect 374806 273049 374858 273055
rect 374806 272991 374858 272997
rect 374818 272907 374846 272991
rect 374806 272901 374858 272907
rect 374806 272843 374858 272849
rect 375010 271205 375038 273065
rect 374998 271199 375050 271205
rect 374998 271141 375050 271147
rect 375106 263810 375134 277135
rect 375298 266987 375326 278004
rect 376246 275713 376298 275719
rect 376246 275655 376298 275661
rect 375572 271978 375628 271987
rect 375572 271913 375628 271922
rect 375286 266981 375338 266987
rect 375286 266923 375338 266929
rect 375586 263810 375614 271913
rect 376258 263824 376286 275655
rect 376738 273721 376766 278018
rect 376822 277119 376874 277125
rect 376822 277061 376874 277067
rect 376726 273715 376778 273721
rect 376726 273657 376778 273663
rect 376834 263824 376862 277061
rect 377494 275787 377546 275793
rect 377494 275729 377546 275735
rect 377012 270350 377068 270359
rect 377012 270285 377068 270294
rect 376032 263796 376286 263824
rect 376608 263796 376862 263824
rect 377026 263810 377054 270285
rect 377506 263810 377534 275729
rect 377890 268171 377918 278018
rect 377974 277045 378026 277051
rect 377974 276987 378026 276993
rect 377878 268165 377930 268171
rect 377878 268107 377930 268113
rect 377986 263810 378014 276987
rect 379028 276122 379084 276131
rect 379028 276057 379084 276066
rect 378644 273310 378700 273319
rect 378644 273245 378700 273254
rect 378658 263824 378686 273245
rect 379042 263824 379070 276057
rect 379138 275423 379166 278018
rect 379414 276971 379466 276977
rect 379414 276913 379466 276919
rect 379126 275417 379178 275423
rect 379126 275359 379178 275365
rect 378432 263796 378686 263824
rect 378912 263796 379070 263824
rect 379426 263810 379454 276913
rect 380290 273869 380318 278018
rect 381046 276897 381098 276903
rect 381046 276839 381098 276845
rect 380566 275639 380618 275645
rect 380566 275581 380618 275587
rect 380278 273863 380330 273869
rect 380278 273805 380330 273811
rect 379894 269497 379946 269503
rect 379894 269439 379946 269445
rect 379906 263810 379934 269439
rect 380578 263824 380606 275581
rect 381058 263824 381086 276839
rect 381442 272463 381470 278018
rect 382294 276823 382346 276829
rect 382294 276765 382346 276771
rect 381814 275565 381866 275571
rect 381814 275507 381866 275513
rect 381430 272457 381482 272463
rect 381430 272399 381482 272405
rect 381526 272457 381578 272463
rect 381526 272399 381578 272405
rect 381538 263824 381566 272399
rect 380352 263796 380606 263824
rect 380832 263796 381086 263824
rect 381264 263796 381566 263824
rect 381826 263810 381854 275507
rect 382306 263810 382334 276765
rect 382594 275349 382622 278018
rect 383638 276749 383690 276755
rect 383638 276691 383690 276697
rect 383444 275974 383500 275983
rect 383444 275909 383500 275918
rect 382582 275343 382634 275349
rect 382582 275285 382634 275291
rect 382964 273162 383020 273171
rect 382964 273097 383020 273106
rect 382978 263824 383006 273097
rect 383458 263824 383486 275909
rect 382752 263796 383006 263824
rect 383232 263796 383486 263824
rect 383650 263810 383678 276691
rect 383842 266839 383870 278018
rect 384994 269059 385022 278018
rect 385366 276601 385418 276607
rect 385366 276543 385418 276549
rect 384982 269053 385034 269059
rect 384982 268995 385034 269001
rect 384118 268165 384170 268171
rect 384118 268107 384170 268113
rect 383830 266833 383882 266839
rect 383830 266775 383882 266781
rect 384130 263810 384158 268107
rect 384886 267203 384938 267209
rect 384886 267145 384938 267151
rect 384898 263824 384926 267145
rect 385378 263824 385406 276543
rect 385556 268870 385612 268879
rect 385556 268805 385612 268814
rect 384672 263796 384926 263824
rect 385152 263796 385406 263824
rect 385570 263810 385598 268805
rect 386038 267129 386090 267135
rect 386038 267071 386090 267077
rect 386050 263810 386078 267071
rect 386146 266913 386174 278018
rect 386518 276675 386570 276681
rect 386518 276617 386570 276623
rect 386134 266907 386186 266913
rect 386134 266849 386186 266855
rect 386530 263810 386558 276617
rect 387394 273943 387422 278018
rect 387382 273937 387434 273943
rect 387382 273879 387434 273885
rect 388546 272389 388574 278018
rect 388918 275491 388970 275497
rect 388918 275433 388970 275439
rect 388534 272383 388586 272389
rect 388534 272325 388586 272331
rect 387286 271199 387338 271205
rect 387286 271141 387338 271147
rect 387298 263824 387326 271141
rect 388436 270202 388492 270211
rect 388436 270137 388492 270146
rect 387766 267055 387818 267061
rect 387766 266997 387818 267003
rect 387778 263824 387806 266997
rect 387958 264021 388010 264027
rect 387958 263963 388010 263969
rect 387072 263796 387326 263824
rect 387552 263796 387806 263824
rect 387970 263810 387998 263963
rect 388450 263810 388478 270137
rect 388930 263810 388958 275433
rect 389590 275417 389642 275423
rect 389590 275359 389642 275365
rect 389602 263824 389630 275359
rect 389698 275275 389726 278018
rect 390356 275826 390412 275835
rect 390356 275761 390412 275770
rect 389686 275269 389738 275275
rect 389686 275211 389738 275217
rect 390164 273014 390220 273023
rect 390164 272949 390220 272958
rect 390178 263824 390206 272949
rect 389472 263796 389630 263824
rect 389952 263796 390206 263824
rect 390370 263810 390398 275761
rect 390946 266691 390974 278018
rect 391990 275343 392042 275349
rect 391990 275285 392042 275291
rect 391508 270054 391564 270063
rect 391508 269989 391564 269998
rect 390934 266685 390986 266691
rect 390934 266627 390986 266633
rect 390838 263947 390890 263953
rect 390838 263889 390890 263895
rect 390850 263810 390878 263889
rect 391522 263824 391550 269989
rect 392002 263824 392030 275285
rect 392098 269429 392126 278018
rect 392278 278007 392330 278013
rect 392278 277949 392330 277955
rect 392962 278004 393264 278032
rect 422570 278029 422832 278032
rect 422518 278023 422832 278029
rect 392086 269423 392138 269429
rect 392086 269365 392138 269371
rect 391296 263796 391550 263824
rect 391776 263796 392030 263824
rect 392290 263810 392318 277949
rect 392756 272866 392812 272875
rect 392756 272801 392812 272810
rect 392770 263810 392798 272801
rect 392962 266765 392990 278004
rect 394498 273795 394526 278018
rect 395156 276566 395212 276575
rect 395156 276501 395212 276510
rect 394486 273789 394538 273795
rect 394486 273731 394538 273737
rect 394390 269423 394442 269429
rect 394390 269365 394442 269371
rect 393238 266907 393290 266913
rect 393238 266849 393290 266855
rect 392950 266759 393002 266765
rect 392950 266701 393002 266707
rect 393250 263810 393278 266849
rect 393910 263873 393962 263879
rect 393696 263821 393910 263824
rect 394402 263824 394430 269365
rect 394678 266981 394730 266987
rect 394678 266923 394730 266929
rect 393696 263815 393962 263821
rect 393696 263796 393950 263815
rect 394176 263796 394430 263824
rect 394690 263810 394718 266923
rect 395170 263810 395198 276501
rect 395650 272315 395678 278018
rect 396310 275269 396362 275275
rect 396310 275211 396362 275217
rect 395638 272309 395690 272315
rect 395638 272251 395690 272257
rect 395926 272309 395978 272315
rect 395926 272251 395978 272257
rect 395938 263824 395966 272251
rect 396322 263824 396350 275211
rect 396802 275201 396830 278018
rect 396790 275195 396842 275201
rect 396790 275137 396842 275143
rect 397076 269906 397132 269915
rect 397076 269841 397132 269850
rect 395664 263796 395966 263824
rect 396096 263796 396350 263824
rect 396576 263805 396830 263824
rect 397090 263810 397118 269841
rect 397558 266833 397610 266839
rect 397558 266775 397610 266781
rect 397570 263810 397598 266775
rect 398050 266617 398078 278018
rect 398900 275678 398956 275687
rect 398900 275613 398956 275622
rect 398708 272718 398764 272727
rect 398708 272653 398764 272662
rect 398230 266759 398282 266765
rect 398230 266701 398282 266707
rect 398038 266611 398090 266617
rect 398038 266553 398090 266559
rect 398242 263824 398270 266701
rect 398722 263824 398750 272653
rect 396576 263799 396842 263805
rect 396576 263796 396790 263799
rect 398016 263796 398270 263824
rect 398496 263796 398750 263824
rect 398914 263810 398942 275613
rect 399202 269355 399230 278018
rect 400354 275053 400382 278018
rect 400342 275047 400394 275053
rect 400342 274989 400394 274995
rect 401506 274091 401534 278018
rect 402548 276714 402604 276723
rect 402548 276649 402604 276658
rect 401494 274085 401546 274091
rect 401494 274027 401546 274033
rect 401782 274085 401834 274091
rect 401782 274027 401834 274033
rect 399190 269349 399242 269355
rect 399190 269291 399242 269297
rect 399958 269349 400010 269355
rect 399958 269291 400010 269297
rect 399382 264169 399434 264175
rect 399382 264111 399434 264117
rect 399394 263810 399422 264111
rect 399970 263810 399998 269291
rect 401302 267869 401354 267875
rect 401302 267811 401354 267817
rect 400630 266685 400682 266691
rect 400630 266627 400682 266633
rect 400642 263824 400670 266627
rect 400416 263796 400670 263824
rect 401314 263810 401342 267811
rect 401794 263810 401822 274027
rect 402562 263824 402590 276649
rect 402754 272241 402782 278018
rect 402742 272235 402794 272241
rect 402742 272177 402794 272183
rect 402934 272235 402986 272241
rect 402934 272177 402986 272183
rect 402946 267875 402974 272177
rect 403028 269758 403084 269767
rect 403028 269693 403084 269702
rect 402934 267869 402986 267875
rect 402934 267811 402986 267817
rect 403042 263824 403070 269693
rect 403222 266611 403274 266617
rect 403222 266553 403274 266559
rect 402336 263796 402590 263824
rect 402816 263796 403070 263824
rect 403234 263810 403262 266553
rect 403906 266469 403934 278018
rect 404950 275195 405002 275201
rect 404950 275137 405002 275143
rect 404180 272570 404236 272579
rect 404180 272505 404236 272514
rect 403894 266463 403946 266469
rect 403894 266405 403946 266411
rect 404194 263810 404222 272505
rect 404962 263824 404990 275137
rect 405058 266543 405086 278018
rect 405428 276862 405484 276871
rect 405428 276797 405484 276806
rect 405046 266537 405098 266543
rect 405046 266479 405098 266485
rect 405442 263824 405470 276797
rect 405620 269610 405676 269619
rect 405620 269545 405676 269554
rect 404736 263796 404990 263824
rect 405216 263796 405470 263824
rect 405634 263810 405662 269545
rect 406306 269281 406334 278018
rect 407458 275127 407486 278018
rect 407828 275530 407884 275539
rect 407828 275465 407884 275474
rect 407734 275195 407786 275201
rect 407734 275137 407786 275143
rect 407446 275121 407498 275127
rect 407446 275063 407498 275069
rect 407746 274091 407774 275137
rect 407734 274085 407786 274091
rect 407734 274027 407786 274033
rect 407252 272422 407308 272431
rect 407252 272357 407308 272366
rect 407446 272383 407498 272389
rect 406294 269275 406346 269281
rect 406294 269217 406346 269223
rect 406582 269053 406634 269059
rect 406582 268995 406634 269001
rect 406102 266537 406154 266543
rect 406102 266479 406154 266485
rect 406114 263810 406142 266479
rect 406594 263810 406622 268995
rect 407266 263824 407294 272357
rect 407446 272325 407498 272331
rect 407458 271205 407486 272325
rect 407446 271199 407498 271205
rect 407446 271141 407498 271147
rect 407842 263824 407870 275465
rect 408406 275121 408458 275127
rect 408406 275063 408458 275069
rect 408418 269059 408446 275063
rect 409858 272167 409886 278018
rect 411010 274239 411038 278018
rect 410998 274233 411050 274239
rect 410998 274175 411050 274181
rect 410900 272274 410956 272283
rect 410900 272209 410956 272218
rect 409846 272161 409898 272167
rect 409846 272103 409898 272109
rect 408982 270755 409034 270761
rect 408982 270697 409034 270703
rect 408406 269053 408458 269059
rect 408406 268995 408458 269001
rect 408994 268393 409022 270697
rect 410420 269462 410476 269471
rect 410420 269397 410476 269406
rect 408982 268387 409034 268393
rect 408982 268329 409034 268335
rect 408502 268239 408554 268245
rect 408502 268181 408554 268187
rect 408022 265575 408074 265581
rect 408022 265517 408074 265523
rect 407040 263796 407294 263824
rect 407616 263796 407870 263824
rect 408034 263810 408062 265517
rect 408514 263810 408542 268181
rect 409942 267869 409994 267875
rect 409942 267811 409994 267817
rect 409174 266463 409226 266469
rect 409174 266405 409226 266411
rect 409186 263824 409214 266405
rect 408960 263796 409214 263824
rect 409954 263810 409982 267811
rect 410434 263810 410462 269397
rect 410914 263810 410942 272209
rect 411764 272126 411820 272135
rect 411764 272061 411820 272070
rect 411572 269314 411628 269323
rect 411572 269249 411628 269258
rect 410998 264169 411050 264175
rect 410998 264111 411050 264117
rect 396790 263741 396842 263747
rect 411010 263731 411038 264111
rect 411586 263824 411614 269249
rect 411360 263796 411614 263824
rect 411778 263824 411806 272061
rect 413410 270761 413438 278018
rect 414562 274165 414590 278018
rect 415714 277791 415742 278018
rect 415702 277785 415754 277791
rect 415702 277727 415754 277733
rect 414550 274159 414602 274165
rect 414550 274101 414602 274107
rect 413686 272161 413738 272167
rect 413686 272103 413738 272109
rect 413398 270755 413450 270761
rect 413398 270697 413450 270703
rect 413698 267875 413726 272103
rect 416962 271279 416990 278018
rect 416950 271273 417002 271279
rect 416950 271215 417002 271221
rect 413686 267869 413738 267875
rect 413686 267811 413738 267817
rect 418114 265507 418142 278018
rect 420514 268467 420542 278018
rect 421666 274313 421694 278018
rect 422530 278004 422832 278023
rect 421654 274307 421706 274313
rect 421654 274249 421706 274255
rect 423970 271353 423998 278018
rect 423958 271347 424010 271353
rect 423958 271289 424010 271295
rect 420502 268461 420554 268467
rect 420502 268403 420554 268409
rect 425218 265655 425246 278018
rect 426370 277865 426398 278018
rect 426358 277859 426410 277865
rect 426358 277801 426410 277807
rect 427522 268541 427550 278018
rect 428770 274387 428798 278018
rect 429634 278004 429936 278032
rect 429634 277939 429662 278004
rect 429622 277933 429674 277939
rect 429622 277875 429674 277881
rect 428758 274381 428810 274387
rect 428758 274323 428810 274329
rect 431074 271427 431102 278018
rect 431062 271421 431114 271427
rect 431062 271363 431114 271369
rect 427510 268535 427562 268541
rect 427510 268477 427562 268483
rect 432322 265729 432350 278018
rect 432310 265723 432362 265729
rect 432310 265665 432362 265671
rect 425206 265649 425258 265655
rect 425206 265591 425258 265597
rect 418102 265501 418154 265507
rect 418102 265443 418154 265449
rect 433474 264101 433502 278018
rect 434626 268615 434654 278018
rect 435874 274461 435902 278018
rect 437026 276533 437054 278018
rect 437014 276527 437066 276533
rect 437014 276469 437066 276475
rect 435862 274455 435914 274461
rect 435862 274397 435914 274403
rect 438178 271501 438206 278018
rect 438166 271495 438218 271501
rect 438166 271437 438218 271443
rect 434614 268609 434666 268615
rect 434614 268551 434666 268557
rect 439330 265803 439358 278018
rect 439318 265797 439370 265803
rect 439318 265739 439370 265745
rect 440578 264767 440606 278018
rect 441730 268689 441758 278018
rect 442882 274535 442910 278018
rect 444130 277717 444158 278018
rect 444118 277711 444170 277717
rect 444118 277653 444170 277659
rect 442870 274529 442922 274535
rect 442870 274471 442922 274477
rect 445282 271575 445310 278018
rect 446434 274609 446462 278018
rect 446422 274603 446474 274609
rect 446422 274545 446474 274551
rect 445270 271569 445322 271575
rect 445270 271511 445322 271517
rect 441718 268683 441770 268689
rect 441718 268625 441770 268631
rect 440566 264761 440618 264767
rect 440566 264703 440618 264709
rect 447682 264693 447710 278018
rect 448834 268763 448862 278018
rect 448822 268757 448874 268763
rect 448822 268699 448874 268705
rect 449986 265877 450014 278018
rect 451234 277643 451262 278018
rect 451222 277637 451274 277643
rect 451222 277579 451274 277585
rect 452386 271649 452414 278018
rect 453538 274683 453566 278018
rect 453526 274677 453578 274683
rect 453526 274619 453578 274625
rect 452374 271643 452426 271649
rect 452374 271585 452426 271591
rect 449974 265871 450026 265877
rect 449974 265813 450026 265819
rect 447670 264687 447722 264693
rect 447670 264629 447722 264635
rect 454786 264471 454814 278018
rect 455938 268837 455966 278018
rect 455926 268831 455978 268837
rect 455926 268773 455978 268779
rect 457090 265951 457118 278018
rect 458242 277569 458270 278018
rect 458230 277563 458282 277569
rect 458230 277505 458282 277511
rect 459490 271723 459518 278018
rect 460642 274757 460670 278018
rect 460630 274751 460682 274757
rect 460630 274693 460682 274699
rect 459478 271717 459530 271723
rect 459478 271659 459530 271665
rect 457078 265945 457130 265951
rect 457078 265887 457130 265893
rect 461794 264619 461822 278018
rect 463042 268911 463070 278018
rect 463030 268905 463082 268911
rect 463030 268847 463082 268853
rect 464194 266025 464222 278018
rect 465346 277495 465374 278018
rect 465334 277489 465386 277495
rect 465334 277431 465386 277437
rect 466594 271797 466622 278018
rect 467746 274831 467774 278018
rect 467734 274825 467786 274831
rect 467734 274767 467786 274773
rect 466582 271791 466634 271797
rect 466582 271733 466634 271739
rect 464182 266019 464234 266025
rect 464182 265961 464234 265967
rect 461782 264613 461834 264619
rect 461782 264555 461834 264561
rect 468898 264545 468926 278018
rect 470146 268985 470174 278018
rect 470134 268979 470186 268985
rect 470134 268921 470186 268927
rect 471298 266099 471326 278018
rect 472450 277421 472478 278018
rect 472438 277415 472490 277421
rect 472438 277357 472490 277363
rect 473698 271871 473726 278018
rect 474850 274503 474878 278018
rect 474836 274494 474892 274503
rect 474836 274429 474892 274438
rect 473686 271865 473738 271871
rect 473686 271807 473738 271813
rect 471286 266093 471338 266099
rect 471286 266035 471338 266041
rect 476002 264841 476030 278018
rect 477154 269133 477182 278018
rect 477142 269127 477194 269133
rect 477142 269069 477194 269075
rect 478402 266173 478430 278018
rect 479554 277347 479582 278018
rect 479542 277341 479594 277347
rect 479542 277283 479594 277289
rect 480706 271945 480734 278018
rect 481954 274905 481982 278018
rect 481942 274899 481994 274905
rect 481942 274841 481994 274847
rect 480694 271939 480746 271945
rect 480694 271881 480746 271887
rect 483106 269207 483134 278018
rect 484258 270613 484286 278018
rect 484246 270607 484298 270613
rect 484246 270549 484298 270555
rect 483094 269201 483146 269207
rect 483094 269143 483146 269149
rect 485506 266247 485534 278018
rect 486658 272019 486686 278018
rect 487810 272093 487838 278018
rect 489058 274651 489086 278018
rect 489044 274642 489100 274651
rect 489044 274577 489100 274586
rect 487798 272087 487850 272093
rect 487798 272029 487850 272035
rect 486646 272013 486698 272019
rect 486646 271955 486698 271961
rect 490210 270465 490238 278018
rect 491362 270539 491390 278018
rect 491350 270533 491402 270539
rect 491350 270475 491402 270481
rect 490198 270459 490250 270465
rect 490198 270401 490250 270407
rect 492610 266321 492638 278018
rect 493762 273499 493790 278018
rect 494914 273573 494942 278018
rect 496066 274799 496094 278018
rect 496052 274790 496108 274799
rect 496052 274725 496108 274734
rect 494902 273567 494954 273573
rect 494902 273509 494954 273515
rect 493750 273493 493802 273499
rect 493750 273435 493802 273441
rect 497314 270391 497342 278018
rect 497302 270385 497354 270391
rect 497302 270327 497354 270333
rect 498466 270317 498494 278018
rect 498454 270311 498506 270317
rect 498454 270253 498506 270259
rect 499618 267801 499646 278018
rect 500866 273425 500894 278018
rect 500854 273419 500906 273425
rect 500854 273361 500906 273367
rect 502018 273351 502046 278018
rect 503170 274947 503198 278018
rect 503156 274938 503212 274947
rect 503156 274873 503212 274882
rect 502006 273345 502058 273351
rect 502006 273287 502058 273293
rect 504418 270169 504446 278018
rect 505570 270243 505598 278018
rect 505558 270237 505610 270243
rect 505558 270179 505610 270185
rect 504406 270163 504458 270169
rect 504406 270105 504458 270111
rect 499606 267795 499658 267801
rect 499606 267737 499658 267743
rect 506722 267727 506750 278018
rect 507970 273203 507998 278018
rect 509122 273277 509150 278018
rect 510274 274979 510302 278018
rect 510262 274973 510314 274979
rect 510262 274915 510314 274921
rect 509110 273271 509162 273277
rect 509110 273213 509162 273219
rect 509206 273271 509258 273277
rect 509206 273213 509258 273219
rect 507958 273197 508010 273203
rect 507958 273139 508010 273145
rect 508246 273197 508298 273203
rect 508246 273139 508298 273145
rect 506710 267721 506762 267727
rect 506710 267663 506762 267669
rect 492598 266315 492650 266321
rect 492598 266257 492650 266263
rect 485494 266241 485546 266247
rect 485494 266183 485546 266189
rect 478390 266167 478442 266173
rect 478390 266109 478442 266115
rect 508258 265581 508286 273139
rect 509218 270687 509246 273213
rect 509206 270681 509258 270687
rect 509206 270623 509258 270629
rect 511522 270095 511550 278018
rect 511510 270089 511562 270095
rect 511510 270031 511562 270037
rect 512674 270021 512702 278018
rect 512662 270015 512714 270021
rect 512662 269957 512714 269963
rect 513826 267653 513854 278018
rect 514978 273129 515006 278018
rect 514966 273123 515018 273129
rect 514966 273065 515018 273071
rect 516226 273055 516254 278018
rect 517378 276459 517406 278018
rect 517366 276453 517418 276459
rect 517366 276395 517418 276401
rect 516214 273049 516266 273055
rect 516214 272991 516266 272997
rect 516310 273049 516362 273055
rect 516310 272991 516362 272997
rect 516322 268171 516350 272991
rect 518530 269873 518558 278018
rect 519778 269947 519806 278018
rect 519766 269941 519818 269947
rect 519766 269883 519818 269889
rect 518518 269867 518570 269873
rect 518518 269809 518570 269815
rect 516310 268165 516362 268171
rect 516310 268107 516362 268113
rect 513814 267647 513866 267653
rect 513814 267589 513866 267595
rect 520930 267579 520958 278018
rect 521300 276862 521356 276871
rect 521300 276797 521356 276806
rect 521314 273573 521342 276797
rect 521302 273567 521354 273573
rect 521302 273509 521354 273515
rect 522082 272907 522110 278018
rect 523330 272981 523358 278018
rect 524482 276385 524510 278018
rect 524470 276379 524522 276385
rect 524470 276321 524522 276327
rect 523318 272975 523370 272981
rect 523318 272917 523370 272923
rect 522070 272901 522122 272907
rect 522070 272843 522122 272849
rect 523030 272901 523082 272907
rect 523030 272843 523082 272849
rect 523042 268879 523070 272843
rect 525634 269725 525662 278018
rect 526882 269799 526910 278018
rect 526870 269793 526922 269799
rect 526870 269735 526922 269741
rect 525622 269719 525674 269725
rect 525622 269661 525674 269667
rect 523028 268870 523084 268879
rect 523028 268805 523084 268814
rect 520918 267573 520970 267579
rect 520918 267515 520970 267521
rect 528034 267505 528062 278018
rect 529186 272833 529214 278018
rect 529844 276714 529900 276723
rect 529844 276649 529900 276658
rect 529858 273499 529886 276649
rect 529846 273493 529898 273499
rect 529846 273435 529898 273441
rect 529174 272827 529226 272833
rect 529174 272769 529226 272775
rect 530434 272759 530462 278018
rect 531586 276311 531614 278018
rect 531574 276305 531626 276311
rect 531574 276247 531626 276253
rect 530422 272753 530474 272759
rect 530422 272695 530474 272701
rect 532738 269651 532766 278018
rect 532726 269645 532778 269651
rect 532726 269587 532778 269593
rect 533890 269577 533918 278018
rect 533878 269571 533930 269577
rect 533878 269513 533930 269519
rect 528022 267499 528074 267505
rect 528022 267441 528074 267447
rect 535138 267431 535166 278018
rect 536290 272611 536318 278018
rect 537442 272685 537470 278018
rect 538690 276237 538718 278018
rect 538678 276231 538730 276237
rect 538678 276173 538730 276179
rect 537430 272679 537482 272685
rect 537430 272621 537482 272627
rect 536278 272605 536330 272611
rect 536278 272547 536330 272553
rect 539842 269027 539870 278018
rect 540994 269175 541022 278018
rect 540980 269166 541036 269175
rect 540980 269101 541036 269110
rect 539828 269018 539884 269027
rect 539828 268953 539884 268962
rect 535126 267425 535178 267431
rect 535126 267367 535178 267373
rect 542242 267357 542270 278018
rect 543394 271691 543422 278018
rect 544546 271839 544574 278018
rect 545794 276163 545822 278018
rect 545782 276157 545834 276163
rect 545782 276099 545834 276105
rect 546946 276089 546974 278018
rect 546934 276083 546986 276089
rect 546934 276025 546986 276031
rect 548098 273277 548126 278018
rect 549346 276015 549374 278018
rect 549334 276009 549386 276015
rect 549334 275951 549386 275957
rect 548086 273271 548138 273277
rect 548086 273213 548138 273219
rect 544532 271830 544588 271839
rect 544532 271765 544588 271774
rect 543380 271682 543436 271691
rect 543380 271617 543436 271626
rect 542230 267351 542282 267357
rect 542230 267293 542282 267299
rect 550498 267283 550526 278018
rect 551650 272537 551678 278018
rect 552802 275941 552830 278018
rect 554050 277273 554078 278018
rect 554038 277267 554090 277273
rect 554038 277209 554090 277215
rect 552790 275935 552842 275941
rect 552790 275877 552842 275883
rect 551638 272531 551690 272537
rect 551638 272473 551690 272479
rect 555202 270507 555230 278018
rect 556354 275867 556382 278018
rect 557602 277199 557630 278018
rect 557590 277193 557642 277199
rect 557590 277135 557642 277141
rect 556342 275861 556394 275867
rect 556342 275803 556394 275809
rect 558754 271987 558782 278018
rect 559906 275719 559934 278018
rect 561154 277125 561182 278018
rect 561142 277119 561194 277125
rect 561142 277061 561194 277067
rect 559894 275713 559946 275719
rect 559894 275655 559946 275661
rect 558740 271978 558796 271987
rect 558740 271913 558796 271922
rect 555188 270498 555244 270507
rect 555188 270433 555244 270442
rect 562306 270359 562334 278018
rect 563458 275793 563486 278018
rect 564706 277051 564734 278018
rect 564694 277045 564746 277051
rect 564694 276987 564746 276993
rect 563446 275787 563498 275793
rect 563446 275729 563498 275735
rect 565858 273319 565886 278018
rect 567010 276131 567038 278018
rect 568258 276977 568286 278018
rect 568246 276971 568298 276977
rect 568246 276913 568298 276919
rect 566996 276122 567052 276131
rect 566996 276057 567052 276066
rect 565844 273310 565900 273319
rect 565844 273245 565900 273254
rect 562292 270350 562348 270359
rect 562292 270285 562348 270294
rect 569410 269503 569438 278018
rect 570562 275645 570590 278018
rect 571714 276903 571742 278018
rect 571702 276897 571754 276903
rect 571702 276839 571754 276845
rect 570550 275639 570602 275645
rect 570550 275581 570602 275587
rect 572962 272463 572990 278018
rect 574114 275571 574142 278018
rect 575266 276829 575294 278018
rect 575254 276823 575306 276829
rect 575254 276765 575306 276771
rect 574102 275565 574154 275571
rect 574102 275507 574154 275513
rect 576514 273171 576542 278018
rect 577666 275983 577694 278018
rect 578818 276755 578846 278018
rect 578806 276749 578858 276755
rect 578806 276691 578858 276697
rect 577652 275974 577708 275983
rect 577652 275909 577708 275918
rect 576500 273162 576556 273171
rect 576500 273097 576556 273106
rect 580066 273055 580094 278018
rect 580054 273049 580106 273055
rect 580054 272991 580106 272997
rect 572950 272457 573002 272463
rect 572950 272399 573002 272405
rect 569398 269497 569450 269503
rect 569398 269439 569450 269445
rect 550486 267277 550538 267283
rect 550486 267219 550538 267225
rect 581218 267209 581246 278018
rect 582370 276607 582398 278018
rect 582358 276601 582410 276607
rect 582358 276543 582410 276549
rect 583618 272907 583646 278018
rect 583606 272901 583658 272907
rect 583606 272843 583658 272849
rect 581206 267203 581258 267209
rect 581206 267145 581258 267151
rect 584770 267135 584798 278018
rect 585922 276681 585950 278018
rect 585910 276675 585962 276681
rect 585910 276617 585962 276623
rect 587170 272389 587198 278018
rect 587158 272383 587210 272389
rect 587158 272325 587210 272331
rect 584758 267129 584810 267135
rect 584758 267071 584810 267077
rect 588322 267061 588350 278018
rect 588310 267055 588362 267061
rect 588310 266997 588362 267003
rect 508246 265575 508298 265581
rect 508246 265517 508298 265523
rect 475990 264835 476042 264841
rect 475990 264777 476042 264783
rect 468886 264539 468938 264545
rect 468886 264481 468938 264487
rect 454774 264465 454826 264471
rect 454774 264407 454826 264413
rect 433462 264095 433514 264101
rect 433462 264037 433514 264043
rect 589474 264027 589502 278018
rect 590626 270211 590654 278018
rect 591874 275497 591902 278018
rect 591862 275491 591914 275497
rect 591862 275433 591914 275439
rect 593026 275423 593054 278018
rect 593014 275417 593066 275423
rect 593014 275359 593066 275365
rect 594178 273023 594206 278018
rect 595426 275835 595454 278018
rect 595412 275826 595468 275835
rect 595412 275761 595468 275770
rect 594164 273014 594220 273023
rect 594164 272949 594220 272958
rect 590612 270202 590668 270211
rect 590612 270137 590668 270146
rect 589462 264021 589514 264027
rect 589462 263963 589514 263969
rect 596578 263953 596606 278018
rect 597730 270063 597758 278018
rect 598978 275349 599006 278018
rect 599842 278013 600144 278032
rect 599830 278007 600144 278013
rect 599882 278004 600144 278007
rect 599830 277949 599882 277955
rect 598966 275343 599018 275349
rect 598966 275285 599018 275291
rect 601282 272875 601310 278018
rect 601268 272866 601324 272875
rect 601268 272801 601324 272810
rect 597716 270054 597772 270063
rect 597716 269989 597772 269998
rect 602530 266913 602558 278018
rect 602518 266907 602570 266913
rect 602518 266849 602570 266855
rect 596566 263947 596618 263953
rect 596566 263889 596618 263895
rect 603682 263879 603710 278018
rect 604834 269429 604862 278018
rect 604822 269423 604874 269429
rect 604822 269365 604874 269371
rect 606082 266987 606110 278018
rect 607234 276575 607262 278018
rect 607220 276566 607276 276575
rect 607220 276501 607276 276510
rect 608386 272315 608414 278018
rect 609538 275275 609566 278018
rect 609526 275269 609578 275275
rect 609526 275211 609578 275217
rect 608374 272309 608426 272315
rect 608374 272251 608426 272257
rect 606070 266981 606122 266987
rect 606070 266923 606122 266929
rect 603670 263873 603722 263879
rect 411778 263796 411840 263824
rect 603670 263815 603722 263821
rect 610786 263805 610814 278018
rect 611938 269915 611966 278018
rect 611924 269906 611980 269915
rect 611924 269841 611980 269850
rect 613090 266839 613118 278018
rect 613078 266833 613130 266839
rect 613078 266775 613130 266781
rect 614338 266765 614366 278018
rect 615490 272727 615518 278018
rect 616642 275687 616670 278018
rect 616628 275678 616684 275687
rect 616628 275613 616684 275622
rect 615476 272718 615532 272727
rect 615476 272653 615532 272662
rect 614326 266759 614378 266765
rect 614326 266701 614378 266707
rect 610774 263799 610826 263805
rect 610774 263741 610826 263747
rect 617890 263731 617918 278018
rect 619042 269355 619070 278018
rect 619030 269349 619082 269355
rect 619030 269291 619082 269297
rect 620194 266691 620222 278018
rect 620182 266685 620234 266691
rect 620182 266627 620234 266633
rect 401110 263725 401162 263731
rect 270562 263648 270624 263676
rect 299170 263648 299232 263676
rect 345442 263648 345504 263676
rect 400896 263673 401110 263676
rect 410998 263725 411050 263731
rect 400896 263667 401162 263673
rect 400896 263648 401150 263667
rect 403728 263657 404030 263676
rect 410998 263667 411050 263673
rect 617878 263725 617930 263731
rect 617878 263667 617930 263673
rect 621442 263657 621470 278018
rect 622594 272241 622622 278018
rect 623746 275201 623774 278018
rect 623734 275195 623786 275201
rect 623734 275137 623786 275143
rect 624994 273499 625022 278018
rect 624982 273493 625034 273499
rect 624982 273435 625034 273441
rect 622582 272235 622634 272241
rect 622582 272177 622634 272183
rect 626146 269767 626174 278018
rect 626132 269758 626188 269767
rect 626132 269693 626188 269702
rect 627298 266617 627326 278018
rect 627286 266611 627338 266617
rect 627286 266553 627338 266559
rect 403728 263651 404042 263657
rect 403728 263648 403990 263651
rect 403990 263593 404042 263599
rect 621430 263651 621482 263657
rect 621430 263593 621482 263599
rect 628450 263583 628478 278018
rect 629698 272579 629726 278018
rect 630850 275053 630878 278018
rect 630838 275047 630890 275053
rect 630838 274989 630890 274995
rect 632002 273573 632030 278018
rect 631990 273567 632042 273573
rect 631990 273509 632042 273515
rect 629684 272570 629740 272579
rect 629684 272505 629740 272514
rect 633250 269619 633278 278018
rect 633236 269610 633292 269619
rect 633236 269545 633292 269554
rect 634402 266543 634430 278018
rect 635554 275127 635582 278018
rect 635542 275121 635594 275127
rect 635542 275063 635594 275069
rect 636802 272431 636830 278018
rect 637954 275539 637982 278018
rect 637940 275530 637996 275539
rect 637940 275465 637996 275474
rect 639106 273203 639134 278018
rect 639094 273197 639146 273203
rect 639094 273139 639146 273145
rect 636788 272422 636844 272431
rect 636788 272357 636844 272366
rect 640354 268245 640382 278018
rect 640342 268239 640394 268245
rect 640342 268181 640394 268187
rect 634390 266537 634442 266543
rect 634390 266479 634442 266485
rect 641506 266469 641534 278018
rect 641494 266463 641546 266469
rect 641494 266405 641546 266411
rect 409654 263577 409706 263583
rect 409440 263525 409654 263528
rect 409440 263519 409706 263525
rect 628438 263577 628490 263583
rect 628438 263519 628490 263525
rect 409440 263500 409694 263519
rect 642658 263509 642686 278018
rect 643906 272167 643934 278018
rect 643894 272161 643946 272167
rect 643894 272103 643946 272109
rect 645058 269471 645086 278018
rect 646210 272283 646238 278018
rect 646484 275382 646540 275391
rect 646484 275317 646540 275326
rect 646196 272274 646252 272283
rect 646196 272209 646252 272218
rect 645044 269462 645100 269471
rect 645044 269397 645100 269406
rect 642646 263503 642698 263509
rect 642646 263445 642698 263451
rect 420404 262210 420460 262219
rect 420404 262145 420406 262154
rect 420458 262145 420460 262154
rect 606166 262171 606218 262177
rect 420406 262113 420458 262119
rect 606166 262113 606218 262119
rect 187222 260691 187274 260697
rect 187222 260633 187274 260639
rect 189718 260691 189770 260697
rect 189718 260633 189770 260639
rect 186262 255141 186314 255147
rect 186262 255083 186314 255089
rect 186070 255067 186122 255073
rect 186070 255009 186122 255015
rect 185974 254919 186026 254925
rect 185974 254861 186026 254867
rect 185782 246705 185834 246711
rect 185782 246647 185834 246653
rect 185590 242857 185642 242863
rect 185590 242799 185642 242805
rect 185602 220335 185630 242799
rect 185686 242709 185738 242715
rect 185686 242651 185738 242657
rect 185588 220326 185644 220335
rect 185588 220261 185644 220270
rect 185492 198274 185548 198283
rect 185492 198209 185548 198218
rect 184244 197682 184300 197691
rect 184244 197617 184300 197626
rect 183094 195867 183146 195873
rect 183094 195809 183146 195815
rect 182998 149765 183050 149771
rect 182998 149707 183050 149713
rect 183106 143999 183134 195809
rect 184534 195793 184586 195799
rect 184534 195735 184586 195741
rect 184438 195719 184490 195725
rect 184438 195661 184490 195667
rect 184342 195645 184394 195651
rect 184342 195587 184394 195593
rect 184354 195323 184382 195587
rect 184340 195314 184396 195323
rect 184340 195249 184396 195258
rect 184450 194435 184478 195661
rect 184436 194426 184492 194435
rect 184436 194361 184492 194370
rect 184546 193843 184574 195735
rect 184532 193834 184588 193843
rect 184532 193769 184588 193778
rect 184630 192981 184682 192987
rect 184436 192946 184492 192955
rect 184630 192923 184682 192929
rect 184436 192881 184492 192890
rect 184534 192907 184586 192913
rect 184342 192833 184394 192839
rect 184342 192775 184394 192781
rect 184354 192363 184382 192775
rect 184450 192765 184478 192881
rect 184534 192849 184586 192855
rect 184438 192759 184490 192765
rect 184438 192701 184490 192707
rect 184340 192354 184396 192363
rect 184340 192289 184396 192298
rect 184546 191475 184574 192849
rect 184532 191466 184588 191475
rect 184532 191401 184588 191410
rect 184642 190735 184670 192923
rect 184628 190726 184684 190735
rect 184628 190661 184684 190670
rect 184534 190095 184586 190101
rect 184534 190037 184586 190043
rect 184342 190021 184394 190027
rect 184340 189986 184342 189995
rect 184394 189986 184396 189995
rect 184340 189921 184396 189930
rect 184438 189947 184490 189953
rect 184438 189889 184490 189895
rect 184342 189873 184394 189879
rect 184342 189815 184394 189821
rect 184354 188515 184382 189815
rect 184340 188506 184396 188515
rect 184340 188441 184396 188450
rect 184450 187627 184478 189889
rect 184546 189255 184574 190037
rect 184532 189246 184588 189255
rect 184532 189181 184588 189190
rect 184436 187618 184492 187627
rect 184436 187553 184492 187562
rect 184438 187209 184490 187215
rect 184438 187151 184490 187157
rect 184342 187061 184394 187067
rect 184342 187003 184394 187009
rect 184354 186887 184382 187003
rect 184340 186878 184396 186887
rect 184340 186813 184396 186822
rect 184450 186147 184478 187151
rect 184534 187135 184586 187141
rect 184534 187077 184586 187083
rect 184436 186138 184492 186147
rect 184436 186073 184492 186082
rect 184546 184667 184574 187077
rect 184630 186987 184682 186993
rect 184630 186929 184682 186935
rect 184642 185407 184670 186929
rect 184628 185398 184684 185407
rect 184628 185333 184684 185342
rect 184532 184658 184588 184667
rect 184532 184593 184588 184602
rect 184342 184323 184394 184329
rect 184342 184265 184394 184271
rect 184354 183927 184382 184265
rect 184438 184249 184490 184255
rect 184438 184191 184490 184197
rect 184340 183918 184396 183927
rect 184340 183853 184396 183862
rect 184450 181559 184478 184191
rect 184436 181550 184492 181559
rect 184436 181485 184492 181494
rect 184630 181437 184682 181443
rect 184630 181379 184682 181385
rect 184342 181363 184394 181369
rect 184342 181305 184394 181311
rect 184354 180819 184382 181305
rect 184438 181289 184490 181295
rect 184438 181231 184490 181237
rect 184340 180810 184396 180819
rect 184340 180745 184396 180754
rect 184450 180079 184478 181231
rect 184534 181215 184586 181221
rect 184534 181157 184586 181163
rect 184436 180070 184492 180079
rect 184436 180005 184492 180014
rect 184546 178599 184574 181157
rect 184642 179339 184670 181379
rect 185302 180105 185354 180111
rect 185302 180047 185354 180053
rect 184628 179330 184684 179339
rect 184628 179265 184684 179274
rect 184532 178590 184588 178599
rect 184438 178551 184490 178557
rect 184532 178525 184588 178534
rect 184438 178493 184490 178499
rect 184342 178403 184394 178409
rect 184342 178345 184394 178351
rect 184354 177119 184382 178345
rect 184450 177711 184478 178493
rect 184534 178477 184586 178483
rect 184534 178419 184586 178425
rect 184436 177702 184492 177711
rect 184436 177637 184492 177646
rect 184340 177110 184396 177119
rect 184340 177045 184396 177054
rect 184546 176231 184574 178419
rect 184532 176222 184588 176231
rect 184532 176157 184588 176166
rect 184438 175665 184490 175671
rect 184340 175630 184396 175639
rect 184438 175607 184490 175613
rect 184340 175565 184342 175574
rect 184394 175565 184396 175574
rect 184342 175533 184394 175539
rect 184450 174011 184478 175607
rect 184436 174002 184492 174011
rect 184436 173937 184492 173946
rect 184630 172779 184682 172785
rect 184630 172721 184682 172727
rect 184438 172705 184490 172711
rect 184438 172647 184490 172653
rect 184342 172631 184394 172637
rect 184342 172573 184394 172579
rect 184354 172531 184382 172573
rect 184340 172522 184396 172531
rect 184340 172457 184396 172466
rect 184450 171791 184478 172647
rect 184534 172557 184586 172563
rect 184534 172499 184586 172505
rect 184436 171782 184492 171791
rect 184436 171717 184492 171726
rect 184546 170311 184574 172499
rect 184642 170903 184670 172721
rect 184628 170894 184684 170903
rect 184628 170829 184684 170838
rect 184532 170302 184588 170311
rect 184532 170237 184588 170246
rect 184438 169893 184490 169899
rect 184438 169835 184490 169841
rect 184342 169745 184394 169751
rect 184342 169687 184394 169693
rect 184354 168683 184382 169687
rect 184450 169423 184478 169835
rect 184630 169819 184682 169825
rect 184630 169761 184682 169767
rect 184534 169671 184586 169677
rect 184534 169613 184586 169619
rect 184436 169414 184492 169423
rect 184436 169349 184492 169358
rect 184340 168674 184396 168683
rect 184340 168609 184396 168618
rect 184546 167203 184574 169613
rect 184642 167943 184670 169761
rect 184628 167934 184684 167943
rect 184628 167869 184684 167878
rect 184532 167194 184588 167203
rect 184532 167129 184588 167138
rect 184342 167007 184394 167013
rect 184342 166949 184394 166955
rect 184354 166463 184382 166949
rect 184438 166933 184490 166939
rect 184438 166875 184490 166881
rect 184340 166454 184396 166463
rect 184340 166389 184396 166398
rect 184450 165723 184478 166875
rect 184534 166859 184586 166865
rect 184534 166801 184586 166807
rect 184436 165714 184492 165723
rect 184436 165649 184492 165658
rect 184546 164835 184574 166801
rect 185314 165626 185342 180047
rect 185698 175694 185726 242651
rect 185794 182447 185822 246647
rect 185878 242783 185930 242789
rect 185878 242725 185930 242731
rect 185890 195854 185918 242725
rect 185986 204351 186014 254861
rect 186082 212047 186110 255009
rect 186166 246335 186218 246341
rect 186166 246277 186218 246283
rect 186068 212038 186124 212047
rect 186068 211973 186124 211982
rect 185972 204342 186028 204351
rect 185972 204277 186028 204286
rect 186178 202871 186206 246277
rect 186274 215007 186302 255083
rect 186454 254993 186506 254999
rect 186454 254935 186506 254941
rect 186358 246631 186410 246637
rect 186358 246573 186410 246579
rect 186260 214998 186316 215007
rect 186260 214933 186316 214942
rect 186370 207311 186398 246573
rect 186466 213527 186494 254935
rect 186646 252033 186698 252039
rect 186646 251975 186698 251981
rect 186550 246557 186602 246563
rect 186550 246499 186602 246505
rect 186452 213518 186508 213527
rect 186452 213453 186508 213462
rect 186356 207302 186412 207311
rect 186356 207237 186412 207246
rect 186562 205979 186590 246499
rect 186658 210567 186686 251975
rect 186742 246483 186794 246489
rect 186742 246425 186794 246431
rect 186644 210558 186700 210567
rect 186644 210493 186700 210502
rect 186754 209087 186782 246425
rect 186838 246409 186890 246415
rect 186838 246351 186890 246357
rect 186850 218115 186878 246351
rect 187030 246261 187082 246267
rect 187030 246203 187082 246209
rect 186934 244929 186986 244935
rect 186934 244871 186986 244877
rect 186946 221075 186974 244871
rect 186932 221066 186988 221075
rect 186932 221001 186988 221010
rect 186836 218106 186892 218115
rect 186836 218041 186892 218050
rect 187042 216487 187070 246203
rect 187124 243414 187180 243423
rect 187124 243349 187180 243358
rect 187138 227545 187166 243349
rect 187126 227539 187178 227545
rect 187126 227481 187178 227487
rect 187138 226139 187166 227481
rect 187126 226133 187178 226139
rect 187126 226075 187178 226081
rect 187028 216478 187084 216487
rect 187028 216413 187084 216422
rect 186740 209078 186796 209087
rect 186740 209013 186796 209022
rect 186548 205970 186604 205979
rect 186548 205905 186604 205914
rect 186164 202862 186220 202871
rect 186164 202797 186220 202806
rect 185974 201565 186026 201571
rect 185974 201507 186026 201513
rect 185986 199763 186014 201507
rect 185972 199754 186028 199763
rect 185972 199689 186028 199698
rect 187234 199171 187262 260633
rect 420404 259842 420460 259851
rect 420404 259777 420460 259786
rect 191540 259398 191596 259407
rect 191540 259333 191596 259342
rect 190196 251702 190252 251711
rect 190196 251637 190252 251646
rect 190210 228581 190238 251637
rect 190198 228575 190250 228581
rect 190198 228517 190250 228523
rect 190774 227539 190826 227545
rect 190774 227481 190826 227487
rect 190786 221792 190814 227481
rect 190786 221764 190862 221792
rect 190834 221482 190862 221764
rect 191554 221482 191582 259333
rect 420418 259291 420446 259777
rect 420406 259285 420458 259291
rect 420406 259227 420458 259233
rect 420404 257030 420460 257039
rect 420404 256965 420460 256974
rect 420418 256405 420446 256965
rect 420406 256399 420458 256405
rect 420406 256341 420458 256347
rect 420404 255254 420460 255263
rect 420404 255189 420460 255198
rect 420418 253519 420446 255189
rect 420406 253513 420458 253519
rect 420406 253455 420458 253461
rect 603286 253513 603338 253519
rect 603286 253455 603338 253461
rect 420404 252886 420460 252895
rect 420404 252821 420460 252830
rect 420418 250633 420446 252821
rect 420406 250627 420458 250633
rect 420406 250569 420458 250575
rect 420308 250518 420364 250527
rect 420308 250453 420364 250462
rect 420322 247821 420350 250453
rect 420404 248150 420460 248159
rect 420404 248085 420460 248094
rect 420310 247815 420362 247821
rect 420310 247757 420362 247763
rect 420418 247747 420446 248085
rect 420406 247741 420458 247747
rect 420406 247683 420458 247689
rect 420404 245338 420460 245347
rect 420404 245273 420460 245282
rect 420418 244861 420446 245273
rect 420406 244855 420458 244861
rect 420406 244797 420458 244803
rect 420404 243562 420460 243571
rect 420404 243497 420460 243506
rect 420418 241975 420446 243497
rect 420406 241969 420458 241975
rect 420406 241911 420458 241917
rect 600406 241969 600458 241975
rect 600406 241911 600458 241917
rect 420404 241194 420460 241203
rect 420404 241129 420460 241138
rect 412148 240158 412204 240167
rect 412148 240093 412204 240102
rect 412052 240010 412108 240019
rect 380640 239977 380894 239996
rect 380640 239971 380906 239977
rect 380640 239968 380854 239971
rect 412052 239945 412054 239954
rect 380854 239913 380906 239919
rect 412106 239945 412108 239954
rect 412054 239913 412106 239919
rect 412162 239903 412190 240093
rect 409558 239897 409610 239903
rect 409344 239845 409558 239848
rect 409344 239839 409610 239845
rect 412150 239897 412202 239903
rect 412150 239839 412202 239845
rect 357142 239823 357194 239829
rect 409344 239820 409598 239839
rect 357142 239765 357194 239771
rect 192418 233317 192446 239686
rect 192768 239672 192926 239700
rect 192898 233539 192926 239672
rect 193138 239404 193166 239686
rect 193282 239672 193488 239700
rect 193138 239376 193214 239404
rect 193186 236174 193214 239376
rect 193090 236146 193214 236174
rect 192886 233533 192938 233539
rect 192886 233475 192938 233481
rect 192406 233311 192458 233317
rect 192406 233253 192458 233259
rect 192310 228575 192362 228581
rect 192310 228517 192362 228523
rect 192322 221482 192350 228517
rect 193090 221792 193118 236146
rect 193282 233391 193310 239672
rect 193858 233465 193886 239686
rect 194242 233613 194270 239686
rect 194626 236174 194654 239686
rect 194976 239672 195230 239700
rect 195360 239672 195614 239700
rect 194626 236146 194750 236174
rect 194230 233607 194282 233613
rect 194230 233549 194282 233555
rect 193846 233459 193898 233465
rect 193846 233401 193898 233407
rect 193270 233385 193322 233391
rect 193270 233327 193322 233333
rect 194614 233385 194666 233391
rect 194614 233327 194666 233333
rect 193750 233311 193802 233317
rect 193750 233253 193802 233259
rect 193042 221764 193118 221792
rect 193042 221482 193070 221764
rect 193762 221482 193790 233253
rect 194626 221482 194654 233327
rect 194722 233317 194750 236146
rect 195202 233391 195230 239672
rect 195586 233539 195614 239672
rect 195682 233687 195710 239686
rect 195670 233681 195722 233687
rect 195670 233623 195722 233629
rect 195286 233533 195338 233539
rect 195286 233475 195338 233481
rect 195574 233533 195626 233539
rect 195574 233475 195626 233481
rect 195190 233385 195242 233391
rect 195190 233327 195242 233333
rect 194710 233311 194762 233317
rect 194710 233253 194762 233259
rect 195298 221792 195326 233475
rect 196162 233317 196190 239686
rect 196546 233761 196574 239686
rect 196930 233835 196958 239686
rect 197280 239672 197534 239700
rect 197664 239672 197918 239700
rect 197506 233909 197534 239672
rect 197494 233903 197546 233909
rect 197494 233845 197546 233851
rect 196918 233829 196970 233835
rect 196918 233771 196970 233777
rect 196534 233755 196586 233761
rect 196534 233697 196586 233703
rect 196822 233459 196874 233465
rect 196822 233401 196874 233407
rect 196054 233311 196106 233317
rect 196054 233253 196106 233259
rect 196150 233311 196202 233317
rect 196150 233253 196202 233259
rect 195298 221764 195374 221792
rect 195346 221482 195374 221764
rect 196066 221482 196094 233253
rect 196834 221482 196862 233401
rect 197890 233391 197918 239672
rect 197986 233465 198014 239686
rect 198370 233983 198398 239686
rect 198754 234057 198782 239686
rect 198742 234051 198794 234057
rect 198742 233993 198794 233999
rect 198358 233977 198410 233983
rect 198358 233919 198410 233925
rect 199138 233613 199166 239686
rect 199488 239672 199742 239700
rect 199968 239672 200222 239700
rect 198358 233607 198410 233613
rect 198358 233549 198410 233555
rect 199126 233607 199178 233613
rect 199126 233549 199178 233555
rect 197974 233459 198026 233465
rect 197974 233401 198026 233407
rect 197494 233385 197546 233391
rect 197494 233327 197546 233333
rect 197878 233385 197930 233391
rect 197878 233327 197930 233333
rect 197506 221792 197534 233327
rect 197506 221764 197582 221792
rect 197554 221482 197582 221764
rect 198370 221482 198398 233549
rect 199714 233317 199742 239672
rect 200194 234131 200222 239672
rect 200290 234205 200318 239686
rect 200278 234199 200330 234205
rect 200278 234141 200330 234147
rect 200182 234125 200234 234131
rect 200182 234067 200234 234073
rect 200566 233755 200618 233761
rect 200566 233697 200618 233703
rect 199798 233533 199850 233539
rect 199798 233475 199850 233481
rect 199126 233311 199178 233317
rect 199126 233253 199178 233259
rect 199702 233311 199754 233317
rect 199702 233253 199754 233259
rect 199138 221482 199166 233253
rect 199810 221792 199838 233475
rect 199810 221764 199886 221792
rect 199858 221482 199886 221764
rect 200578 221482 200606 233697
rect 200674 233539 200702 239686
rect 201058 233761 201086 239686
rect 201408 239672 201566 239700
rect 201792 239672 202046 239700
rect 202176 239672 202430 239700
rect 201538 234279 201566 239672
rect 202018 234575 202046 239672
rect 202006 234569 202058 234575
rect 202006 234511 202058 234517
rect 201526 234273 201578 234279
rect 201526 234215 201578 234221
rect 201046 233755 201098 233761
rect 201046 233697 201098 233703
rect 201334 233681 201386 233687
rect 201334 233623 201386 233629
rect 200662 233533 200714 233539
rect 200662 233475 200714 233481
rect 201346 221482 201374 233623
rect 202402 233391 202430 239672
rect 202498 233687 202526 239686
rect 202882 234649 202910 239686
rect 202870 234643 202922 234649
rect 202870 234585 202922 234591
rect 203266 234353 203294 239686
rect 203712 239672 203966 239700
rect 204096 239672 204254 239700
rect 203254 234347 203306 234353
rect 203254 234289 203306 234295
rect 202870 233829 202922 233835
rect 202870 233771 202922 233777
rect 202486 233681 202538 233687
rect 202486 233623 202538 233629
rect 202102 233385 202154 233391
rect 202102 233327 202154 233333
rect 202390 233385 202442 233391
rect 202390 233327 202442 233333
rect 202114 221792 202142 233327
rect 202114 221764 202190 221792
rect 202162 221482 202190 221764
rect 202882 221482 202910 233771
rect 203938 233465 203966 239672
rect 204226 233835 204254 239672
rect 204418 239672 204480 239700
rect 204418 234871 204446 239672
rect 204406 234865 204458 234871
rect 204406 234807 204458 234813
rect 204802 234797 204830 239686
rect 204790 234791 204842 234797
rect 204790 234733 204842 234739
rect 205186 233909 205214 239686
rect 204310 233903 204362 233909
rect 204310 233845 204362 233851
rect 205174 233903 205226 233909
rect 205174 233845 205226 233851
rect 204214 233829 204266 233835
rect 204214 233771 204266 233777
rect 203638 233459 203690 233465
rect 203638 233401 203690 233407
rect 203926 233459 203978 233465
rect 203926 233401 203978 233407
rect 203650 221482 203678 233401
rect 204322 221792 204350 233845
rect 205570 233613 205598 239686
rect 205920 239672 206174 239700
rect 206304 239672 206558 239700
rect 206688 239672 206942 239700
rect 206146 234501 206174 239672
rect 206530 234723 206558 239672
rect 206518 234717 206570 234723
rect 206518 234659 206570 234665
rect 206134 234495 206186 234501
rect 206134 234437 206186 234443
rect 206914 234353 206942 239672
rect 207010 234427 207038 239686
rect 207490 235093 207518 239686
rect 207478 235087 207530 235093
rect 207478 235029 207530 235035
rect 206998 234421 207050 234427
rect 206998 234363 207050 234369
rect 206806 234347 206858 234353
rect 206806 234289 206858 234295
rect 206902 234347 206954 234353
rect 206902 234289 206954 234295
rect 206818 233983 206846 234289
rect 207874 234057 207902 239686
rect 208224 239672 208478 239700
rect 208608 239672 208862 239700
rect 208450 236055 208478 239672
rect 208438 236049 208490 236055
rect 208438 235991 208490 235997
rect 208834 235833 208862 239672
rect 208930 235907 208958 239686
rect 208918 235901 208970 235907
rect 208918 235843 208970 235849
rect 208822 235827 208874 235833
rect 208822 235769 208874 235775
rect 209314 235315 209342 239686
rect 209698 235981 209726 239686
rect 209686 235975 209738 235981
rect 209686 235917 209738 235923
rect 210082 235611 210110 239686
rect 210432 239672 210686 239700
rect 210816 239672 211070 239700
rect 210658 235685 210686 239672
rect 210646 235679 210698 235685
rect 210646 235621 210698 235627
rect 210070 235605 210122 235611
rect 210070 235547 210122 235553
rect 209302 235309 209354 235315
rect 209302 235251 209354 235257
rect 211042 235019 211070 239672
rect 211234 235759 211262 239686
rect 211222 235753 211274 235759
rect 211222 235695 211274 235701
rect 211618 235167 211646 239686
rect 212002 235463 212030 239686
rect 211990 235457 212042 235463
rect 211990 235399 212042 235405
rect 211606 235161 211658 235167
rect 211606 235103 211658 235109
rect 211030 235013 211082 235019
rect 211030 234955 211082 234961
rect 210166 234865 210218 234871
rect 210166 234807 210218 234813
rect 208822 234125 208874 234131
rect 208822 234067 208874 234073
rect 207382 234051 207434 234057
rect 207382 233993 207434 233999
rect 207862 234051 207914 234057
rect 207862 233993 207914 233999
rect 205942 233977 205994 233983
rect 205942 233919 205994 233925
rect 206806 233977 206858 233983
rect 206806 233919 206858 233925
rect 205078 233607 205130 233613
rect 205078 233549 205130 233555
rect 205558 233607 205610 233613
rect 205558 233549 205610 233555
rect 204322 221764 204398 221792
rect 204370 221482 204398 221764
rect 205090 221482 205118 233549
rect 205954 221496 205982 233919
rect 206614 233311 206666 233317
rect 206614 233253 206666 233259
rect 205920 221468 205982 221496
rect 206626 221496 206654 233253
rect 206626 221468 206688 221496
rect 207394 221482 207422 233993
rect 208150 233533 208202 233539
rect 208150 233475 208202 233481
rect 208162 221496 208190 233475
rect 208128 221468 208190 221496
rect 208834 221496 208862 234067
rect 210178 233761 210206 234807
rect 210454 234791 210506 234797
rect 210454 234733 210506 234739
rect 210466 234205 210494 234733
rect 211990 234495 212042 234501
rect 211990 234437 212042 234443
rect 212002 234279 212030 234437
rect 211894 234273 211946 234279
rect 211894 234215 211946 234221
rect 211990 234273 212042 234279
rect 211990 234215 212042 234221
rect 210358 234199 210410 234205
rect 210358 234141 210410 234147
rect 210454 234199 210506 234205
rect 210454 234141 210506 234147
rect 209686 233755 209738 233761
rect 209686 233697 209738 233703
rect 210166 233755 210218 233761
rect 210166 233697 210218 233703
rect 208834 221468 208896 221496
rect 209698 221482 209726 233697
rect 210370 221681 210398 234141
rect 211126 233385 211178 233391
rect 211126 233327 211178 233333
rect 210370 221653 210446 221681
rect 210418 221482 210446 221653
rect 211138 221482 211166 233327
rect 211906 221482 211934 234215
rect 212386 225991 212414 239686
rect 212736 239672 212990 239700
rect 212962 235537 212990 239672
rect 213058 239672 213120 239700
rect 212950 235531 213002 235537
rect 212950 235473 213002 235479
rect 212566 233681 212618 233687
rect 212566 233623 212618 233629
rect 212374 225985 212426 225991
rect 212374 225927 212426 225933
rect 212578 221681 212606 233623
rect 213058 227027 213086 239672
rect 213442 234945 213470 239686
rect 213430 234939 213482 234945
rect 213430 234881 213482 234887
rect 213430 234569 213482 234575
rect 213430 234511 213482 234517
rect 213046 227021 213098 227027
rect 213046 226963 213098 226969
rect 212578 221653 212654 221681
rect 212626 221482 212654 221653
rect 213442 221482 213470 234511
rect 213826 226361 213854 239686
rect 214210 235389 214238 239686
rect 214198 235383 214250 235389
rect 214198 235325 214250 235331
rect 214198 233459 214250 233465
rect 214198 233401 214250 233407
rect 213814 226355 213866 226361
rect 213814 226297 213866 226303
rect 214210 221482 214238 233401
rect 214594 226065 214622 239686
rect 215040 239672 215294 239700
rect 215424 239672 215678 239700
rect 214870 234643 214922 234649
rect 214870 234585 214922 234591
rect 214582 226059 214634 226065
rect 214582 226001 214634 226007
rect 214882 221681 214910 234585
rect 215266 229025 215294 239672
rect 215542 233829 215594 233835
rect 215542 233771 215594 233777
rect 215254 229019 215306 229025
rect 215254 228961 215306 228967
rect 215554 226084 215582 233771
rect 215650 226213 215678 239672
rect 215746 227471 215774 239686
rect 216144 239672 216446 239700
rect 215734 227465 215786 227471
rect 215734 227407 215786 227413
rect 216418 226287 216446 239672
rect 216514 236174 216542 239686
rect 216864 239672 217118 239700
rect 217248 239672 217502 239700
rect 217632 239672 217886 239700
rect 216514 236146 216638 236174
rect 216502 233977 216554 233983
rect 216502 233919 216554 233925
rect 216406 226281 216458 226287
rect 216406 226223 216458 226229
rect 215638 226207 215690 226213
rect 215638 226149 215690 226155
rect 215554 226056 215678 226084
rect 214882 221653 214958 221681
rect 214930 221482 214958 221653
rect 215650 221482 215678 226056
rect 216514 221482 216542 233919
rect 216610 232799 216638 236146
rect 216598 232793 216650 232799
rect 216598 232735 216650 232741
rect 217090 227397 217118 239672
rect 217174 233903 217226 233909
rect 217174 233845 217226 233851
rect 217078 227391 217130 227397
rect 217078 227333 217130 227339
rect 217186 221792 217214 233845
rect 217474 227545 217502 239672
rect 217462 227539 217514 227545
rect 217462 227481 217514 227487
rect 217858 227249 217886 239672
rect 217954 236174 217982 239686
rect 217954 236146 218078 236174
rect 217942 233755 217994 233761
rect 217942 233697 217994 233703
rect 217846 227243 217898 227249
rect 217846 227185 217898 227191
rect 217186 221764 217262 221792
rect 217234 221482 217262 221764
rect 217954 221482 217982 233697
rect 218050 232577 218078 236146
rect 218038 232571 218090 232577
rect 218038 232513 218090 232519
rect 218338 226139 218366 239686
rect 218710 233533 218762 233539
rect 218710 233475 218762 233481
rect 218326 226133 218378 226139
rect 218326 226075 218378 226081
rect 218722 221482 218750 233475
rect 218818 225917 218846 239686
rect 219168 239672 219422 239700
rect 219552 239672 219806 239700
rect 219936 239672 220190 239700
rect 219394 236174 219422 239672
rect 219394 236146 219518 236174
rect 219382 234199 219434 234205
rect 219382 234141 219434 234147
rect 218806 225911 218858 225917
rect 218806 225853 218858 225859
rect 219394 221792 219422 234141
rect 219490 227323 219518 236146
rect 219778 232651 219806 239672
rect 219766 232645 219818 232651
rect 219766 232587 219818 232593
rect 220162 229765 220190 239672
rect 220258 236174 220286 239686
rect 220258 236146 220382 236174
rect 220246 234347 220298 234353
rect 220246 234289 220298 234295
rect 220150 229759 220202 229765
rect 220150 229701 220202 229707
rect 219478 227317 219530 227323
rect 219478 227259 219530 227265
rect 219394 221764 219470 221792
rect 219442 221482 219470 221764
rect 220258 221482 220286 234289
rect 220354 227175 220382 236146
rect 220642 235389 220670 239686
rect 221026 236174 221054 239686
rect 221376 239672 221630 239700
rect 221026 236146 221150 236174
rect 220534 235383 220586 235389
rect 220534 235325 220586 235331
rect 220630 235383 220682 235389
rect 220630 235325 220682 235331
rect 220546 234945 220574 235325
rect 220534 234939 220586 234945
rect 220534 234881 220586 234887
rect 221014 234273 221066 234279
rect 221014 234215 221066 234221
rect 220342 227169 220394 227175
rect 220342 227111 220394 227117
rect 221026 221482 221054 234215
rect 221122 232503 221150 236146
rect 221110 232497 221162 232503
rect 221110 232439 221162 232445
rect 221602 229617 221630 239672
rect 221746 239404 221774 239686
rect 222144 239672 222302 239700
rect 221698 239376 221774 239404
rect 221590 229611 221642 229617
rect 221590 229553 221642 229559
rect 221698 226953 221726 239376
rect 222274 234649 222302 239672
rect 222454 234717 222506 234723
rect 222454 234659 222506 234665
rect 222262 234643 222314 234649
rect 222262 234585 222314 234591
rect 221782 234421 221834 234427
rect 221782 234363 221834 234369
rect 221686 226947 221738 226953
rect 221686 226889 221738 226895
rect 221794 221792 221822 234363
rect 221746 221764 221822 221792
rect 221746 221482 221774 221764
rect 222466 221482 222494 234659
rect 222562 232429 222590 239686
rect 222550 232423 222602 232429
rect 222550 232365 222602 232371
rect 222946 232355 222974 239686
rect 223222 236049 223274 236055
rect 223222 235991 223274 235997
rect 222934 232349 222986 232355
rect 222934 232291 222986 232297
rect 223234 221482 223262 235991
rect 223330 226805 223358 239686
rect 223680 239672 223934 239700
rect 224064 239672 224318 239700
rect 223906 235167 223934 239672
rect 223894 235161 223946 235167
rect 223894 235103 223946 235109
rect 223990 235087 224042 235093
rect 223990 235029 224042 235035
rect 223318 226799 223370 226805
rect 223318 226741 223370 226747
rect 224002 221792 224030 235029
rect 224290 232281 224318 239672
rect 224278 232275 224330 232281
rect 224278 232217 224330 232223
rect 224386 228507 224414 239686
rect 224770 236174 224798 239686
rect 224770 236146 224894 236174
rect 224758 235827 224810 235833
rect 224758 235769 224810 235775
rect 224374 228501 224426 228507
rect 224374 228443 224426 228449
rect 224002 221764 224078 221792
rect 224050 221482 224078 221764
rect 224770 221482 224798 235769
rect 224866 226879 224894 236146
rect 225154 234723 225182 239686
rect 225538 234871 225566 239686
rect 225984 239672 226238 239700
rect 226368 239672 226622 239700
rect 226210 236174 226238 239672
rect 226210 236146 226334 236174
rect 226198 235975 226250 235981
rect 226198 235917 226250 235923
rect 225526 234865 225578 234871
rect 225526 234807 225578 234813
rect 225142 234717 225194 234723
rect 225142 234659 225194 234665
rect 225526 234125 225578 234131
rect 225526 234067 225578 234073
rect 224854 226873 224906 226879
rect 224854 226815 224906 226821
rect 225538 221482 225566 234067
rect 226210 221792 226238 235917
rect 226306 232207 226334 236146
rect 226294 232201 226346 232207
rect 226294 232143 226346 232149
rect 226594 226657 226622 239672
rect 226690 233391 226718 239686
rect 226966 235901 227018 235907
rect 226966 235843 227018 235849
rect 226678 233385 226730 233391
rect 226678 233327 226730 233333
rect 226582 226651 226634 226657
rect 226582 226593 226634 226599
rect 226210 221764 226286 221792
rect 226258 221482 226286 221764
rect 226978 221482 227006 235843
rect 227074 232133 227102 239686
rect 227062 232127 227114 232133
rect 227062 232069 227114 232075
rect 227458 229913 227486 239686
rect 227856 239672 227966 239700
rect 228192 239672 228446 239700
rect 228576 239672 228830 239700
rect 227830 235605 227882 235611
rect 227830 235547 227882 235553
rect 227446 229907 227498 229913
rect 227446 229849 227498 229855
rect 227842 221482 227870 235547
rect 227938 226731 227966 239672
rect 228418 233613 228446 239672
rect 228502 235309 228554 235315
rect 228502 235251 228554 235257
rect 228406 233607 228458 233613
rect 228406 233549 228458 233555
rect 227926 226725 227978 226731
rect 227926 226667 227978 226673
rect 228514 221792 228542 235251
rect 228802 228581 228830 239672
rect 228898 229469 228926 239686
rect 229296 239672 229598 239700
rect 229270 235753 229322 235759
rect 229270 235695 229322 235701
rect 228886 229463 228938 229469
rect 228886 229405 228938 229411
rect 228790 228575 228842 228581
rect 228790 228517 228842 228523
rect 228514 221764 228590 221792
rect 228562 221482 228590 221764
rect 229282 221482 229310 235695
rect 229570 226583 229598 239672
rect 229762 235315 229790 239686
rect 230112 239672 230366 239700
rect 230496 239672 230654 239700
rect 230880 239672 231134 239700
rect 230038 235679 230090 235685
rect 230038 235621 230090 235627
rect 229750 235309 229802 235315
rect 229750 235251 229802 235257
rect 229558 226577 229610 226583
rect 229558 226519 229610 226525
rect 230050 221482 230078 235621
rect 230338 229395 230366 239672
rect 230326 229389 230378 229395
rect 230326 229331 230378 229337
rect 230626 228655 230654 239672
rect 230710 235235 230762 235241
rect 230710 235177 230762 235183
rect 230614 228649 230666 228655
rect 230614 228591 230666 228597
rect 230722 221792 230750 235177
rect 231106 225769 231134 239672
rect 231202 235759 231230 239686
rect 231600 239672 231902 239700
rect 231190 235753 231242 235759
rect 231190 235695 231242 235701
rect 231574 235013 231626 235019
rect 231574 234955 231626 234961
rect 231094 225763 231146 225769
rect 231094 225705 231146 225711
rect 230722 221764 230798 221792
rect 230770 221482 230798 221764
rect 231586 221482 231614 234955
rect 231874 228729 231902 239672
rect 231970 229247 231998 239686
rect 232320 239672 232574 239700
rect 232704 239672 232958 239700
rect 233088 239672 233246 239700
rect 232342 235531 232394 235537
rect 232342 235473 232394 235479
rect 231958 229241 232010 229247
rect 231958 229183 232010 229189
rect 231862 228723 231914 228729
rect 231862 228665 231914 228671
rect 232354 221482 232382 235473
rect 232546 226435 232574 239672
rect 232930 235241 232958 239672
rect 233014 235457 233066 235463
rect 233014 235399 233066 235405
rect 232918 235235 232970 235241
rect 232918 235177 232970 235183
rect 232534 226429 232586 226435
rect 232534 226371 232586 226377
rect 233026 221792 233054 235399
rect 233218 231911 233246 239672
rect 233206 231905 233258 231911
rect 233206 231847 233258 231853
rect 233506 229321 233534 239686
rect 233890 232059 233918 239686
rect 234274 235907 234302 239686
rect 234624 239672 234878 239700
rect 235008 239672 235262 239700
rect 235392 239672 235646 239700
rect 234262 235901 234314 235907
rect 234262 235843 234314 235849
rect 233878 232053 233930 232059
rect 233878 231995 233930 232001
rect 234850 231985 234878 239672
rect 234838 231979 234890 231985
rect 234838 231921 234890 231927
rect 233494 229315 233546 229321
rect 233494 229257 233546 229263
rect 235234 229173 235262 239672
rect 235318 234939 235370 234945
rect 235318 234881 235370 234887
rect 235222 229167 235274 229173
rect 235222 229109 235274 229115
rect 233782 227021 233834 227027
rect 233782 226963 233834 226969
rect 233026 221764 233102 221792
rect 233074 221482 233102 221764
rect 233794 221482 233822 226963
rect 234550 225985 234602 225991
rect 234550 225927 234602 225933
rect 234562 221482 234590 225927
rect 235330 221496 235358 234881
rect 235618 234501 235646 239672
rect 235714 234945 235742 239686
rect 236002 239672 236112 239700
rect 235702 234939 235754 234945
rect 235702 234881 235754 234887
rect 235606 234495 235658 234501
rect 235606 234437 235658 234443
rect 236002 231837 236030 239672
rect 236482 235611 236510 239686
rect 236832 239672 237086 239700
rect 237312 239672 237566 239700
rect 236470 235605 236522 235611
rect 236470 235547 236522 235553
rect 236086 234791 236138 234797
rect 236086 234733 236138 234739
rect 235990 231831 236042 231837
rect 235990 231773 236042 231779
rect 235330 221468 235392 221496
rect 236098 221482 236126 234733
rect 237058 234427 237086 239672
rect 237538 235833 237566 239672
rect 237526 235827 237578 235833
rect 237526 235769 237578 235775
rect 237046 234421 237098 234427
rect 237046 234363 237098 234369
rect 237634 232725 237662 239686
rect 238018 235537 238046 239686
rect 238006 235531 238058 235537
rect 238006 235473 238058 235479
rect 238102 233607 238154 233613
rect 238102 233549 238154 233555
rect 237622 232719 237674 232725
rect 237622 232661 237674 232667
rect 238114 227027 238142 233549
rect 238402 229099 238430 239686
rect 238390 229093 238442 229099
rect 238390 229035 238442 229041
rect 238390 227465 238442 227471
rect 238390 227407 238442 227413
rect 238102 227021 238154 227027
rect 238102 226963 238154 226969
rect 237526 226355 237578 226361
rect 237526 226297 237578 226303
rect 236854 226059 236906 226065
rect 236854 226001 236906 226007
rect 236866 221496 236894 226001
rect 236832 221468 236894 221496
rect 237538 221496 237566 226297
rect 237538 221468 237600 221496
rect 238402 221482 238430 227407
rect 238786 227101 238814 239686
rect 239136 239672 239390 239700
rect 239520 239672 239774 239700
rect 239362 235685 239390 239672
rect 239350 235679 239402 235685
rect 239350 235621 239402 235627
rect 238966 233385 239018 233391
rect 238966 233327 239018 233333
rect 238774 227095 238826 227101
rect 238774 227037 238826 227043
rect 238978 226065 239006 233327
rect 239062 229019 239114 229025
rect 239062 228961 239114 228967
rect 238966 226059 239018 226065
rect 238966 226001 239018 226007
rect 239074 221792 239102 228961
rect 239746 228877 239774 239672
rect 239842 234353 239870 239686
rect 240226 234649 240254 239686
rect 240214 234643 240266 234649
rect 240214 234585 240266 234591
rect 239830 234347 239882 234353
rect 239830 234289 239882 234295
rect 240610 233539 240638 239686
rect 240598 233533 240650 233539
rect 240598 233475 240650 233481
rect 241090 229025 241118 239686
rect 241440 239672 241694 239700
rect 241078 229019 241130 229025
rect 241078 228961 241130 228967
rect 239734 228871 239786 228877
rect 239734 228813 239786 228819
rect 241666 228803 241694 239672
rect 241762 239672 241824 239700
rect 241654 228797 241706 228803
rect 241654 228739 241706 228745
rect 241270 227539 241322 227545
rect 241270 227481 241322 227487
rect 239830 226281 239882 226287
rect 239830 226223 239882 226229
rect 239074 221764 239150 221792
rect 239122 221482 239150 221764
rect 239842 221482 239870 226223
rect 240598 226207 240650 226213
rect 240598 226149 240650 226155
rect 240610 221482 240638 226149
rect 241282 221792 241310 227481
rect 241762 226361 241790 239672
rect 242146 235463 242174 239686
rect 242134 235457 242186 235463
rect 242134 235399 242186 235405
rect 241846 235383 241898 235389
rect 241846 235325 241898 235331
rect 241750 226355 241802 226361
rect 241750 226297 241802 226303
rect 241858 225621 241886 235325
rect 242134 232793 242186 232799
rect 242134 232735 242186 232741
rect 241846 225615 241898 225621
rect 241846 225557 241898 225563
rect 241282 221764 241358 221792
rect 241330 221482 241358 221764
rect 242146 221482 242174 232735
rect 242530 228951 242558 239686
rect 242914 234279 242942 239686
rect 243298 235981 243326 239686
rect 243648 239672 243902 239700
rect 244032 239672 244286 239700
rect 243286 235975 243338 235981
rect 243286 235917 243338 235923
rect 243874 235019 243902 239672
rect 243862 235013 243914 235019
rect 243862 234955 243914 234961
rect 243958 234569 244010 234575
rect 243958 234511 244010 234517
rect 242902 234273 242954 234279
rect 242902 234215 242954 234221
rect 242518 228945 242570 228951
rect 242518 228887 242570 228893
rect 243574 227391 243626 227397
rect 243574 227333 243626 227339
rect 242902 227243 242954 227249
rect 242902 227185 242954 227191
rect 242914 221482 242942 227185
rect 243586 221792 243614 227333
rect 243970 225177 243998 234511
rect 244258 229691 244286 239672
rect 244354 234131 244382 239686
rect 244848 239672 245054 239700
rect 244726 235161 244778 235167
rect 244726 235103 244778 235109
rect 244342 234125 244394 234131
rect 244342 234067 244394 234073
rect 244246 229685 244298 229691
rect 244246 229627 244298 229633
rect 244738 227545 244766 235103
rect 244726 227539 244778 227545
rect 244726 227481 244778 227487
rect 245026 226287 245054 239672
rect 245110 232571 245162 232577
rect 245110 232513 245162 232519
rect 245014 226281 245066 226287
rect 245014 226223 245066 226229
rect 244342 225911 244394 225917
rect 244342 225853 244394 225859
rect 243958 225171 244010 225177
rect 243958 225113 244010 225119
rect 243586 221764 243662 221792
rect 243634 221482 243662 221764
rect 244354 221482 244382 225853
rect 245122 221482 245150 232513
rect 245218 231319 245246 239686
rect 245568 239672 245822 239700
rect 245952 239672 246206 239700
rect 246336 239672 246590 239700
rect 245206 231313 245258 231319
rect 245206 231255 245258 231261
rect 245794 230357 245822 239672
rect 246178 230431 246206 239672
rect 246166 230425 246218 230431
rect 246166 230367 246218 230373
rect 245782 230351 245834 230357
rect 245782 230293 245834 230299
rect 245878 227317 245930 227323
rect 245878 227259 245930 227265
rect 245890 221792 245918 227259
rect 246562 226213 246590 239672
rect 246658 235093 246686 239686
rect 246646 235087 246698 235093
rect 246646 235029 246698 235035
rect 247042 230209 247070 239686
rect 247426 234057 247454 239686
rect 247776 239672 248030 239700
rect 248160 239672 248414 239700
rect 248640 239672 248798 239700
rect 248002 236055 248030 239672
rect 247990 236049 248042 236055
rect 247990 235991 248042 235997
rect 247702 234717 247754 234723
rect 247702 234659 247754 234665
rect 247414 234051 247466 234057
rect 247414 233993 247466 233999
rect 247030 230203 247082 230209
rect 247030 230145 247082 230151
rect 247414 227169 247466 227175
rect 247414 227111 247466 227117
rect 246550 226207 246602 226213
rect 246550 226149 246602 226155
rect 246646 226133 246698 226139
rect 246646 226075 246698 226081
rect 245890 221764 245966 221792
rect 245938 221482 245966 221764
rect 246658 221482 246686 226075
rect 247426 221482 247454 227111
rect 247714 226509 247742 234659
rect 248086 232645 248138 232651
rect 248086 232587 248138 232593
rect 247702 226503 247754 226509
rect 247702 226445 247754 226451
rect 248098 221792 248126 232587
rect 248386 231541 248414 239672
rect 248374 231535 248426 231541
rect 248374 231477 248426 231483
rect 248770 230135 248798 239672
rect 248962 230283 248990 239686
rect 248950 230277 249002 230283
rect 248950 230219 249002 230225
rect 248758 230129 248810 230135
rect 248758 230071 248810 230077
rect 249346 227397 249374 239686
rect 249730 235389 249758 239686
rect 250080 239672 250238 239700
rect 249718 235383 249770 235389
rect 249718 235325 249770 235331
rect 249718 229759 249770 229765
rect 249718 229701 249770 229707
rect 249334 227391 249386 227397
rect 249334 227333 249386 227339
rect 248854 225615 248906 225621
rect 248854 225557 248906 225563
rect 248098 221764 248174 221792
rect 248146 221482 248174 221764
rect 248866 221482 248894 225557
rect 249730 221482 249758 229701
rect 250210 227841 250238 239672
rect 250450 239404 250478 239686
rect 250848 239672 251102 239700
rect 250450 239376 250526 239404
rect 250498 234501 250526 239376
rect 251074 236129 251102 239672
rect 251062 236123 251114 236129
rect 251062 236065 251114 236071
rect 251170 234723 251198 239686
rect 251158 234717 251210 234723
rect 251158 234659 251210 234665
rect 250582 234569 250634 234575
rect 250582 234511 250634 234517
rect 250486 234495 250538 234501
rect 250486 234437 250538 234443
rect 250594 228137 250622 234511
rect 251158 232497 251210 232503
rect 251158 232439 251210 232445
rect 250582 228131 250634 228137
rect 250582 228073 250634 228079
rect 250198 227835 250250 227841
rect 250198 227777 250250 227783
rect 250390 226947 250442 226953
rect 250390 226889 250442 226895
rect 250402 221792 250430 226889
rect 250402 221764 250478 221792
rect 250450 221482 250478 221764
rect 251170 221482 251198 232439
rect 251554 229987 251582 239686
rect 251938 230061 251966 239686
rect 252384 239672 252638 239700
rect 252768 239672 253022 239700
rect 252610 236174 252638 239672
rect 252610 236146 252734 236174
rect 251926 230055 251978 230061
rect 251926 229997 251978 230003
rect 251542 229981 251594 229987
rect 251542 229923 251594 229929
rect 252598 229611 252650 229617
rect 252598 229553 252650 229559
rect 252118 227095 252170 227101
rect 252118 227037 252170 227043
rect 252130 226361 252158 227037
rect 252118 226355 252170 226361
rect 252118 226297 252170 226303
rect 251926 225171 251978 225177
rect 251926 225113 251978 225119
rect 251938 221482 251966 225113
rect 252610 221792 252638 229553
rect 252706 225103 252734 236146
rect 252994 231097 253022 239672
rect 252982 231091 253034 231097
rect 252982 231033 253034 231039
rect 253090 229765 253118 239686
rect 253474 233835 253502 239686
rect 253558 235309 253610 235315
rect 253558 235251 253610 235257
rect 253462 233829 253514 233835
rect 253462 233771 253514 233777
rect 253078 229759 253130 229765
rect 253078 229701 253130 229707
rect 253570 226953 253598 235251
rect 253858 233317 253886 239686
rect 254242 234797 254270 239686
rect 254592 239672 254846 239700
rect 254976 239672 255230 239700
rect 254230 234791 254282 234797
rect 254230 234733 254282 234739
rect 253846 233311 253898 233317
rect 253846 233253 253898 233259
rect 254230 232423 254282 232429
rect 254230 232365 254282 232371
rect 253558 226947 253610 226953
rect 253558 226889 253610 226895
rect 253462 226799 253514 226805
rect 253462 226741 253514 226747
rect 252694 225097 252746 225103
rect 252694 225039 252746 225045
rect 252610 221764 252686 221792
rect 252658 221482 252686 221764
rect 253474 221482 253502 226741
rect 254242 221482 254270 232365
rect 254818 229839 254846 239672
rect 254806 229833 254858 229839
rect 254806 229775 254858 229781
rect 255202 229617 255230 239672
rect 255298 234575 255326 239686
rect 255286 234569 255338 234575
rect 255286 234511 255338 234517
rect 255670 232349 255722 232355
rect 255670 232291 255722 232297
rect 255190 229611 255242 229617
rect 255190 229553 255242 229559
rect 254902 227539 254954 227545
rect 254902 227481 254954 227487
rect 254914 221792 254942 227481
rect 254914 221764 254990 221792
rect 254962 221482 254990 221764
rect 255682 221482 255710 232291
rect 255778 231615 255806 239686
rect 255766 231609 255818 231615
rect 255766 231551 255818 231557
rect 256162 231171 256190 239686
rect 256546 234205 256574 239686
rect 256896 239672 257150 239700
rect 257280 239672 257534 239700
rect 256534 234199 256586 234205
rect 256534 234141 256586 234147
rect 256246 233311 256298 233317
rect 256246 233253 256298 233259
rect 256150 231165 256202 231171
rect 256150 231107 256202 231113
rect 256258 227471 256286 233253
rect 256246 227465 256298 227471
rect 256246 227407 256298 227413
rect 256438 226873 256490 226879
rect 256438 226815 256490 226821
rect 256450 221482 256478 226815
rect 257122 226805 257150 239672
rect 257506 235315 257534 239672
rect 257494 235309 257546 235315
rect 257494 235251 257546 235257
rect 257206 232275 257258 232281
rect 257206 232217 257258 232223
rect 257110 226799 257162 226805
rect 257110 226741 257162 226747
rect 257218 221792 257246 232217
rect 257602 231689 257630 239686
rect 257986 233317 258014 239686
rect 258370 233909 258398 239686
rect 258358 233903 258410 233909
rect 258358 233845 258410 233851
rect 257974 233311 258026 233317
rect 257974 233253 258026 233259
rect 258754 233243 258782 239686
rect 259104 239672 259166 239700
rect 259584 239672 259838 239700
rect 259030 235753 259082 235759
rect 259030 235695 259082 235701
rect 258934 234421 258986 234427
rect 258934 234363 258986 234369
rect 258742 233237 258794 233243
rect 258742 233179 258794 233185
rect 257590 231683 257642 231689
rect 257590 231625 257642 231631
rect 258742 228501 258794 228507
rect 258742 228443 258794 228449
rect 257974 226503 258026 226509
rect 257974 226445 258026 226451
rect 257218 221764 257294 221792
rect 257266 221482 257294 221764
rect 257986 221482 258014 226445
rect 258754 221482 258782 228443
rect 258946 227989 258974 234363
rect 258934 227983 258986 227989
rect 258934 227925 258986 227931
rect 259042 225473 259070 235695
rect 259138 231763 259166 239672
rect 259810 233983 259838 239672
rect 259798 233977 259850 233983
rect 259798 233919 259850 233925
rect 259906 233613 259934 239686
rect 260290 234871 260318 239686
rect 260182 234865 260234 234871
rect 260182 234807 260234 234813
rect 260278 234865 260330 234871
rect 260278 234807 260330 234813
rect 259894 233607 259946 233613
rect 259894 233549 259946 233555
rect 259126 231757 259178 231763
rect 259126 231699 259178 231705
rect 259414 226651 259466 226657
rect 259414 226593 259466 226599
rect 259030 225467 259082 225473
rect 259030 225409 259082 225415
rect 259426 221792 259454 226593
rect 259426 221764 259502 221792
rect 259474 221482 259502 221764
rect 260194 221482 260222 234807
rect 260674 233169 260702 239686
rect 261024 239672 261278 239700
rect 261408 239672 261662 239700
rect 261792 239672 261950 239700
rect 260950 234347 261002 234353
rect 260950 234289 261002 234295
rect 260662 233163 260714 233169
rect 260662 233105 260714 233111
rect 260962 228063 260990 234289
rect 261250 234279 261278 239672
rect 261142 234273 261194 234279
rect 261142 234215 261194 234221
rect 261238 234273 261290 234279
rect 261238 234215 261290 234221
rect 261154 228285 261182 234215
rect 261634 233391 261662 239672
rect 261622 233385 261674 233391
rect 261622 233327 261674 233333
rect 261718 232201 261770 232207
rect 261718 232143 261770 232149
rect 261142 228279 261194 228285
rect 261142 228221 261194 228227
rect 260950 228057 261002 228063
rect 260950 227999 261002 228005
rect 261046 226059 261098 226065
rect 261046 226001 261098 226007
rect 261058 221482 261086 226001
rect 261730 221792 261758 232143
rect 261922 223697 261950 239672
rect 262006 235161 262058 235167
rect 262006 235103 262058 235109
rect 262018 225917 262046 235103
rect 262114 233095 262142 239686
rect 262498 234427 262526 239686
rect 262882 235759 262910 239686
rect 263328 239672 263582 239700
rect 263712 239672 263966 239700
rect 264096 239672 264350 239700
rect 262870 235753 262922 235759
rect 262870 235695 262922 235701
rect 262486 234421 262538 234427
rect 262486 234363 262538 234369
rect 262102 233089 262154 233095
rect 262102 233031 262154 233037
rect 263254 232127 263306 232133
rect 263254 232069 263306 232075
rect 262486 226725 262538 226731
rect 262486 226667 262538 226673
rect 262006 225911 262058 225917
rect 262006 225853 262058 225859
rect 261910 223691 261962 223697
rect 261910 223633 261962 223639
rect 261730 221764 261806 221792
rect 261778 221482 261806 221764
rect 262498 221482 262526 226667
rect 263266 221482 263294 232069
rect 263554 223771 263582 239672
rect 263830 234643 263882 234649
rect 263830 234585 263882 234591
rect 263842 227175 263870 234585
rect 263938 232873 263966 239672
rect 263926 232867 263978 232873
rect 263926 232809 263978 232815
rect 264322 229543 264350 239672
rect 264418 233465 264446 239686
rect 264706 239672 264816 239700
rect 264706 236174 264734 239672
rect 264610 236146 264734 236174
rect 264406 233459 264458 233465
rect 264406 233401 264458 233407
rect 264310 229537 264362 229543
rect 264310 229479 264362 229485
rect 263830 227169 263882 227175
rect 263830 227111 263882 227117
rect 264022 227021 264074 227027
rect 264022 226963 264074 226969
rect 263542 223765 263594 223771
rect 263542 223707 263594 223713
rect 264034 221496 264062 226963
rect 264610 223475 264638 236146
rect 264694 235901 264746 235907
rect 264694 235843 264746 235849
rect 264706 225399 264734 235843
rect 265078 234939 265130 234945
rect 265078 234881 265130 234887
rect 264886 234125 264938 234131
rect 264886 234067 264938 234073
rect 264790 229907 264842 229913
rect 264790 229849 264842 229855
rect 264694 225393 264746 225399
rect 264694 225335 264746 225341
rect 264598 223469 264650 223475
rect 264598 223411 264650 223417
rect 264034 221468 264096 221496
rect 264802 221482 264830 229849
rect 264898 228433 264926 234067
rect 264886 228427 264938 228433
rect 264886 228369 264938 228375
rect 265090 225695 265118 234881
rect 265186 232799 265214 239686
rect 265536 239672 265790 239700
rect 265920 239672 266174 239700
rect 266304 239672 266462 239700
rect 265762 233021 265790 239672
rect 266146 235167 266174 239672
rect 266134 235161 266186 235167
rect 266134 235103 266186 235109
rect 266326 234051 266378 234057
rect 266326 233993 266378 233999
rect 265750 233015 265802 233021
rect 265750 232957 265802 232963
rect 265174 232793 265226 232799
rect 265174 232735 265226 232741
rect 266338 228581 266366 233993
rect 266230 228575 266282 228581
rect 266230 228517 266282 228523
rect 266326 228575 266378 228581
rect 266326 228517 266378 228523
rect 265558 226577 265610 226583
rect 265558 226519 265610 226525
rect 265078 225689 265130 225695
rect 265078 225631 265130 225637
rect 265570 221496 265598 226519
rect 265536 221468 265598 221496
rect 266242 221496 266270 228517
rect 266434 223623 266462 239672
rect 266626 232651 266654 239686
rect 267106 234057 267134 239686
rect 267490 234649 267518 239686
rect 267840 239672 268094 239700
rect 268224 239672 268478 239700
rect 267478 234643 267530 234649
rect 267478 234585 267530 234591
rect 267958 234495 268010 234501
rect 267958 234437 268010 234443
rect 267094 234051 267146 234057
rect 267094 233993 267146 233999
rect 267766 233607 267818 233613
rect 267766 233549 267818 233555
rect 266614 232645 266666 232651
rect 266614 232587 266666 232593
rect 266998 226947 267050 226953
rect 266998 226889 267050 226895
rect 266422 223617 266474 223623
rect 266422 223559 266474 223565
rect 266242 221468 266304 221496
rect 267010 221482 267038 226889
rect 267778 225991 267806 233549
rect 267862 229463 267914 229469
rect 267862 229405 267914 229411
rect 267766 225985 267818 225991
rect 267766 225927 267818 225933
rect 267874 221792 267902 229405
rect 267970 228359 267998 234437
rect 267958 228353 268010 228359
rect 267958 228295 268010 228301
rect 268066 223549 268094 239672
rect 268150 235827 268202 235833
rect 268150 235769 268202 235775
rect 268162 226509 268190 235769
rect 268450 232577 268478 239672
rect 268546 234131 268574 239686
rect 268930 234945 268958 239686
rect 269314 236174 269342 239686
rect 269314 236146 269438 236174
rect 268918 234939 268970 234945
rect 268918 234881 268970 234887
rect 268534 234125 268586 234131
rect 268534 234067 268586 234073
rect 269014 233385 269066 233391
rect 269014 233327 269066 233333
rect 268438 232571 268490 232577
rect 268438 232513 268490 232519
rect 268150 226503 268202 226509
rect 268150 226445 268202 226451
rect 269026 225843 269054 233327
rect 269110 233311 269162 233317
rect 269110 233253 269162 233259
rect 269122 228211 269150 233253
rect 269302 229389 269354 229395
rect 269302 229331 269354 229337
rect 269110 228205 269162 228211
rect 269110 228147 269162 228153
rect 269014 225837 269066 225843
rect 269014 225779 269066 225785
rect 268534 225763 268586 225769
rect 268534 225705 268586 225711
rect 268054 223543 268106 223549
rect 268054 223485 268106 223491
rect 267826 221764 267902 221792
rect 267826 221482 267854 221764
rect 268546 221482 268574 225705
rect 269314 221482 269342 229331
rect 269410 223327 269438 236146
rect 269698 232503 269726 239686
rect 270048 239672 270302 239700
rect 270274 233317 270302 239672
rect 270418 239404 270446 239686
rect 270418 239376 270494 239404
rect 270466 233391 270494 239376
rect 270850 236174 270878 239686
rect 270850 236146 270974 236174
rect 270838 233829 270890 233835
rect 270838 233771 270890 233777
rect 270454 233385 270506 233391
rect 270454 233327 270506 233333
rect 270262 233311 270314 233317
rect 270262 233253 270314 233259
rect 269686 232497 269738 232503
rect 269686 232439 269738 232445
rect 270742 228649 270794 228655
rect 270742 228591 270794 228597
rect 269974 225467 270026 225473
rect 269974 225409 270026 225415
rect 269398 223321 269450 223327
rect 269398 223263 269450 223269
rect 269986 221792 270014 225409
rect 269986 221764 270062 221792
rect 270034 221482 270062 221764
rect 270754 221482 270782 228591
rect 270850 228507 270878 233771
rect 270838 228501 270890 228507
rect 270838 228443 270890 228449
rect 270946 223401 270974 236146
rect 271030 235975 271082 235981
rect 271030 235917 271082 235923
rect 271042 226583 271070 235917
rect 271234 232429 271262 239686
rect 271618 234353 271646 239686
rect 271606 234347 271658 234353
rect 271606 234289 271658 234295
rect 271798 233459 271850 233465
rect 271798 233401 271850 233407
rect 271222 232423 271274 232429
rect 271222 232365 271274 232371
rect 271030 226577 271082 226583
rect 271030 226519 271082 226525
rect 271606 226429 271658 226435
rect 271606 226371 271658 226377
rect 270934 223395 270986 223401
rect 270934 223337 270986 223343
rect 271618 221482 271646 226371
rect 271810 226065 271838 233401
rect 272002 227249 272030 239686
rect 272352 239672 272606 239700
rect 272736 239672 272990 239700
rect 272278 228723 272330 228729
rect 272278 228665 272330 228671
rect 271990 227243 272042 227249
rect 271990 227185 272042 227191
rect 271798 226059 271850 226065
rect 271798 226001 271850 226007
rect 272290 221792 272318 228665
rect 272578 223253 272606 239672
rect 272962 232207 272990 239672
rect 273058 234501 273086 239686
rect 273046 234495 273098 234501
rect 273046 234437 273098 234443
rect 272950 232201 273002 232207
rect 272950 232143 273002 232149
rect 273442 226953 273470 239686
rect 273840 239672 274142 239700
rect 273622 236123 273674 236129
rect 273622 236065 273674 236071
rect 273526 233311 273578 233317
rect 273526 233253 273578 233259
rect 273538 229395 273566 233253
rect 273526 229389 273578 229395
rect 273526 229331 273578 229337
rect 273430 226947 273482 226953
rect 273430 226889 273482 226895
rect 273238 226799 273290 226805
rect 273238 226741 273290 226747
rect 273250 225991 273278 226741
rect 273238 225985 273290 225991
rect 273238 225927 273290 225933
rect 273046 225911 273098 225917
rect 273046 225853 273098 225859
rect 272566 223247 272618 223253
rect 272566 223189 272618 223195
rect 272290 221764 272366 221792
rect 272338 221482 272366 221764
rect 273058 221482 273086 225853
rect 273634 225473 273662 236065
rect 273814 229241 273866 229247
rect 273814 229183 273866 229189
rect 273622 225467 273674 225473
rect 273622 225409 273674 225415
rect 273826 221482 273854 229183
rect 274114 222365 274142 239672
rect 274210 232281 274238 239686
rect 274656 239672 274910 239700
rect 275040 239672 275294 239700
rect 274882 232355 274910 239672
rect 275062 233385 275114 233391
rect 275062 233327 275114 233333
rect 274870 232349 274922 232355
rect 274870 232291 274922 232297
rect 274198 232275 274250 232281
rect 274198 232217 274250 232223
rect 274486 232053 274538 232059
rect 274486 231995 274538 232001
rect 274102 222359 274154 222365
rect 274102 222301 274154 222307
rect 274498 221792 274526 231995
rect 275074 227323 275102 233327
rect 275062 227317 275114 227323
rect 275062 227259 275114 227265
rect 275266 227101 275294 239672
rect 275362 237757 275390 239686
rect 275350 237751 275402 237757
rect 275350 237693 275402 237699
rect 275746 232059 275774 239686
rect 276130 236055 276158 239686
rect 276480 239672 276734 239700
rect 276864 239672 277118 239700
rect 277248 239672 277502 239700
rect 276118 236049 276170 236055
rect 276118 235991 276170 235997
rect 276214 235975 276266 235981
rect 276214 235917 276266 235923
rect 275734 232053 275786 232059
rect 275734 231995 275786 232001
rect 275350 231905 275402 231911
rect 275350 231847 275402 231853
rect 275254 227095 275306 227101
rect 275254 227037 275306 227043
rect 274498 221764 274574 221792
rect 274546 221482 274574 221764
rect 275362 221482 275390 231847
rect 276226 225399 276254 235917
rect 276706 227027 276734 239672
rect 277090 237683 277118 239672
rect 277078 237677 277130 237683
rect 277078 237619 277130 237625
rect 277474 232133 277502 239672
rect 277570 236129 277598 239686
rect 277558 236123 277610 236129
rect 277558 236065 277610 236071
rect 277462 232127 277514 232133
rect 277462 232069 277514 232075
rect 276790 229315 276842 229321
rect 276790 229257 276842 229263
rect 276694 227021 276746 227027
rect 276694 226963 276746 226969
rect 276118 225393 276170 225399
rect 276118 225335 276170 225341
rect 276214 225393 276266 225399
rect 276214 225335 276266 225341
rect 276130 221482 276158 225335
rect 276802 221792 276830 229257
rect 277558 228131 277610 228137
rect 277558 228073 277610 228079
rect 276802 221764 276878 221792
rect 276850 221482 276878 221764
rect 277570 221482 277598 228073
rect 277954 224881 277982 239686
rect 278434 236795 278462 239686
rect 278784 239672 279038 239700
rect 279168 239672 279326 239700
rect 279552 239672 279806 239700
rect 278422 236789 278474 236795
rect 278422 236731 278474 236737
rect 278038 234569 278090 234575
rect 278038 234511 278090 234517
rect 278050 227397 278078 234511
rect 278326 231979 278378 231985
rect 278326 231921 278378 231927
rect 278038 227391 278090 227397
rect 278038 227333 278090 227339
rect 277942 224875 277994 224881
rect 277942 224817 277994 224823
rect 278338 221482 278366 231921
rect 279010 231911 279038 239672
rect 279298 235907 279326 239672
rect 279286 235901 279338 235907
rect 279286 235843 279338 235849
rect 279286 234199 279338 234205
rect 279286 234141 279338 234147
rect 279190 233903 279242 233909
rect 279190 233845 279242 233851
rect 278998 231905 279050 231911
rect 278998 231847 279050 231853
rect 279202 225769 279230 233845
rect 279298 227693 279326 234141
rect 279286 227687 279338 227693
rect 279286 227629 279338 227635
rect 279286 227391 279338 227397
rect 279286 227333 279338 227339
rect 279190 225763 279242 225769
rect 279190 225705 279242 225711
rect 279298 225695 279326 227333
rect 279778 226805 279806 239672
rect 279874 236869 279902 239686
rect 279862 236863 279914 236869
rect 279862 236805 279914 236811
rect 280258 231985 280286 239686
rect 280642 235981 280670 239686
rect 280992 239672 281246 239700
rect 281376 239672 281630 239700
rect 281760 239672 282014 239700
rect 281218 236174 281246 239672
rect 281218 236146 281342 236174
rect 280630 235975 280682 235981
rect 280630 235917 280682 235923
rect 281206 233977 281258 233983
rect 281206 233919 281258 233925
rect 280246 231979 280298 231985
rect 280246 231921 280298 231927
rect 279862 229167 279914 229173
rect 279862 229109 279914 229115
rect 279766 226799 279818 226805
rect 279766 226741 279818 226747
rect 279094 225689 279146 225695
rect 279094 225631 279146 225637
rect 279286 225689 279338 225695
rect 279286 225631 279338 225637
rect 279106 221792 279134 225631
rect 279106 221764 279182 221792
rect 279154 221482 279182 221764
rect 279874 221482 279902 229109
rect 280630 227983 280682 227989
rect 280630 227925 280682 227931
rect 280642 221482 280670 227925
rect 281218 227767 281246 233919
rect 281314 232947 281342 236146
rect 281302 232941 281354 232947
rect 281302 232883 281354 232889
rect 281302 231831 281354 231837
rect 281302 231773 281354 231779
rect 281206 227761 281258 227767
rect 281206 227703 281258 227709
rect 281314 221792 281342 231773
rect 281602 222439 281630 239672
rect 281986 231837 282014 239672
rect 281974 231831 282026 231837
rect 281974 231773 282026 231779
rect 282178 228729 282206 239686
rect 282358 234643 282410 234649
rect 282358 234585 282410 234591
rect 282166 228723 282218 228729
rect 282166 228665 282218 228671
rect 282070 226503 282122 226509
rect 282070 226445 282122 226451
rect 281590 222433 281642 222439
rect 281590 222375 281642 222381
rect 281314 221764 281390 221792
rect 281362 221482 281390 221764
rect 282082 221482 282110 226445
rect 282370 225251 282398 234585
rect 282562 226731 282590 239686
rect 282960 239672 283070 239700
rect 283296 239672 283550 239700
rect 283680 239672 283934 239700
rect 282934 235605 282986 235611
rect 282934 235547 282986 235553
rect 282550 226725 282602 226731
rect 282550 226667 282602 226673
rect 282358 225245 282410 225251
rect 282358 225187 282410 225193
rect 282946 221482 282974 235547
rect 283042 222513 283070 239672
rect 283522 229469 283550 239672
rect 283906 234575 283934 239672
rect 283894 234569 283946 234575
rect 283894 234511 283946 234517
rect 284002 234205 284030 239686
rect 284400 239672 284702 239700
rect 283990 234199 284042 234205
rect 283990 234141 284042 234147
rect 284374 232719 284426 232725
rect 284374 232661 284426 232667
rect 283510 229463 283562 229469
rect 283510 229405 283562 229411
rect 283606 229093 283658 229099
rect 283606 229035 283658 229041
rect 283030 222507 283082 222513
rect 283030 222449 283082 222455
rect 283618 221792 283646 229035
rect 283618 221764 283694 221792
rect 283666 221482 283694 221764
rect 284386 221482 284414 232661
rect 284674 226435 284702 239672
rect 284770 229321 284798 239686
rect 285154 233835 285182 239686
rect 285504 239672 285758 239700
rect 285984 239672 286238 239700
rect 285142 233829 285194 233835
rect 285142 233771 285194 233777
rect 284758 229315 284810 229321
rect 284758 229257 284810 229263
rect 285730 226657 285758 239672
rect 285910 235531 285962 235537
rect 285910 235473 285962 235479
rect 285718 226651 285770 226657
rect 285718 226593 285770 226599
rect 284662 226429 284714 226435
rect 284662 226371 284714 226377
rect 285142 226355 285194 226361
rect 285142 226297 285194 226303
rect 285154 221482 285182 226297
rect 285922 221792 285950 235473
rect 286210 222735 286238 239672
rect 286306 229247 286334 239686
rect 286690 234649 286718 239686
rect 287074 235685 287102 239686
rect 287062 235679 287114 235685
rect 287062 235621 287114 235627
rect 287350 235605 287402 235611
rect 287350 235547 287402 235553
rect 286678 234643 286730 234649
rect 286678 234585 286730 234591
rect 286294 229241 286346 229247
rect 286294 229183 286346 229189
rect 287362 228304 287390 235547
rect 287458 233465 287486 239686
rect 287808 239672 287966 239700
rect 288192 239672 288446 239700
rect 287446 233459 287498 233465
rect 287446 233401 287498 233407
rect 287938 229173 287966 239672
rect 288022 234273 288074 234279
rect 288022 234215 288074 234221
rect 287926 229167 287978 229173
rect 287926 229109 287978 229115
rect 287362 228276 287486 228304
rect 286678 228057 286730 228063
rect 286678 227999 286730 228005
rect 286198 222729 286250 222735
rect 286198 222671 286250 222677
rect 285922 221764 285998 221792
rect 285970 221482 285998 221764
rect 286690 221482 286718 227999
rect 287458 221482 287486 228276
rect 288034 227619 288062 234215
rect 288418 233391 288446 239672
rect 288406 233385 288458 233391
rect 288406 233327 288458 233333
rect 288022 227613 288074 227619
rect 288022 227555 288074 227561
rect 288118 227169 288170 227175
rect 288118 227111 288170 227117
rect 288130 221792 288158 227111
rect 288514 226509 288542 239686
rect 288898 235241 288926 239686
rect 288886 235235 288938 235241
rect 288886 235177 288938 235183
rect 288982 232941 289034 232947
rect 288982 232883 289034 232889
rect 288886 228871 288938 228877
rect 288886 228813 288938 228819
rect 288502 226503 288554 226509
rect 288502 226445 288554 226451
rect 288130 221764 288206 221792
rect 288178 221482 288206 221764
rect 288898 221482 288926 228813
rect 288994 227175 289022 232883
rect 289378 228729 289406 239686
rect 289728 239672 289982 239700
rect 290112 239672 290366 239700
rect 290496 239672 290750 239700
rect 289954 232947 289982 239672
rect 290338 235833 290366 239672
rect 290326 235827 290378 235833
rect 290326 235769 290378 235775
rect 290422 233533 290474 233539
rect 290422 233475 290474 233481
rect 289942 232941 289994 232947
rect 289942 232883 289994 232889
rect 289366 228723 289418 228729
rect 289366 228665 289418 228671
rect 289750 228649 289802 228655
rect 289750 228591 289802 228597
rect 288982 227169 289034 227175
rect 288982 227111 289034 227117
rect 289762 221482 289790 228591
rect 290434 221792 290462 233475
rect 290722 230801 290750 239672
rect 290818 231467 290846 239686
rect 290902 234421 290954 234427
rect 290902 234363 290954 234369
rect 290806 231461 290858 231467
rect 290806 231403 290858 231409
rect 290710 230795 290762 230801
rect 290710 230737 290762 230743
rect 290914 229913 290942 234363
rect 290998 234051 291050 234057
rect 290998 233993 291050 233999
rect 290902 229907 290954 229913
rect 290902 229849 290954 229855
rect 291010 228137 291038 233993
rect 291202 229099 291230 239686
rect 291190 229093 291242 229099
rect 291190 229035 291242 229041
rect 290998 228131 291050 228137
rect 290998 228073 291050 228079
rect 291586 226361 291614 239686
rect 291936 239672 292190 239700
rect 292320 239672 292574 239700
rect 292704 239672 292958 239700
rect 292162 229067 292190 239672
rect 292546 231393 292574 239672
rect 292930 234427 292958 239672
rect 292918 234421 292970 234427
rect 292918 234363 292970 234369
rect 292534 231387 292586 231393
rect 292534 231329 292586 231335
rect 292148 229058 292204 229067
rect 291958 229019 292010 229025
rect 292148 228993 292204 229002
rect 291958 228961 292010 228967
rect 291574 226355 291626 226361
rect 291574 226297 291626 226303
rect 291190 226281 291242 226287
rect 291190 226223 291242 226229
rect 290434 221764 290510 221792
rect 290482 221482 290510 221764
rect 291202 221482 291230 226223
rect 291970 221482 291998 228961
rect 293122 228919 293150 239686
rect 293398 235457 293450 235463
rect 293398 235399 293450 235405
rect 293108 228910 293164 228919
rect 293108 228845 293164 228854
rect 292630 228279 292682 228285
rect 292630 228221 292682 228227
rect 292642 221792 292670 228221
rect 293410 228156 293438 235399
rect 293506 231245 293534 239686
rect 293782 234125 293834 234131
rect 293782 234067 293834 234073
rect 293494 231239 293546 231245
rect 293494 231181 293546 231187
rect 293410 228128 293534 228156
rect 292642 221764 292718 221792
rect 292690 221482 292718 221764
rect 293506 221482 293534 228128
rect 293794 227989 293822 234067
rect 293890 228655 293918 239686
rect 294240 239672 294494 239700
rect 294624 239672 294878 239700
rect 295008 239672 295262 239700
rect 294466 233761 294494 239672
rect 294850 235463 294878 239672
rect 294838 235457 294890 235463
rect 294838 235399 294890 235405
rect 295234 234279 295262 239672
rect 295222 234273 295274 234279
rect 295222 234215 295274 234221
rect 294454 233755 294506 233761
rect 294454 233697 294506 233703
rect 295330 232725 295358 239686
rect 295714 234131 295742 239686
rect 295702 234125 295754 234131
rect 295702 234067 295754 234073
rect 296098 233909 296126 239686
rect 296448 239672 296606 239700
rect 296928 239672 297182 239700
rect 296470 235013 296522 235019
rect 296470 234955 296522 234961
rect 296086 233903 296138 233909
rect 296086 233845 296138 233851
rect 295318 232719 295370 232725
rect 295318 232661 295370 232667
rect 294166 229315 294218 229321
rect 294166 229257 294218 229263
rect 293974 229241 294026 229247
rect 293974 229183 294026 229189
rect 293986 229099 294014 229183
rect 293974 229093 294026 229099
rect 293974 229035 294026 229041
rect 294178 228877 294206 229257
rect 294934 228945 294986 228951
rect 294934 228887 294986 228893
rect 294166 228871 294218 228877
rect 294166 228813 294218 228819
rect 293878 228649 293930 228655
rect 293878 228591 293930 228597
rect 293782 227983 293834 227989
rect 293782 227925 293834 227931
rect 294262 226577 294314 226583
rect 294262 226519 294314 226525
rect 294274 221496 294302 226519
rect 294240 221468 294302 221496
rect 294946 221496 294974 228887
rect 295798 228649 295850 228655
rect 295798 228591 295850 228597
rect 295810 228433 295838 228591
rect 295702 228427 295754 228433
rect 295702 228369 295754 228375
rect 295798 228427 295850 228433
rect 295798 228369 295850 228375
rect 294946 221468 295008 221496
rect 295714 221482 295742 228369
rect 296482 221496 296510 234955
rect 296578 229215 296606 239672
rect 297154 233317 297182 239672
rect 297250 233539 297278 239686
rect 297238 233533 297290 233539
rect 297238 233475 297290 233481
rect 297142 233311 297194 233317
rect 297142 233253 297194 233259
rect 297334 230795 297386 230801
rect 297334 230737 297386 230743
rect 296564 229206 296620 229215
rect 296564 229141 296620 229150
rect 297346 226583 297374 230737
rect 297334 226577 297386 226583
rect 297334 226519 297386 226525
rect 297634 226287 297662 239686
rect 298018 235019 298046 239686
rect 298416 239672 298622 239700
rect 298752 239672 299006 239700
rect 299136 239672 299390 239700
rect 298006 235013 298058 235019
rect 298006 234955 298058 234961
rect 298594 229691 298622 239672
rect 298978 236943 299006 239672
rect 298966 236937 299018 236943
rect 298966 236879 299018 236885
rect 299254 235087 299306 235093
rect 299254 235029 299306 235035
rect 299266 230505 299294 235029
rect 299362 234691 299390 239672
rect 299458 234987 299486 239686
rect 299842 235537 299870 239686
rect 299830 235531 299882 235537
rect 299830 235473 299882 235479
rect 299444 234978 299500 234987
rect 299444 234913 299500 234922
rect 299348 234682 299404 234691
rect 299348 234617 299404 234626
rect 300226 231319 300254 239686
rect 299446 231313 299498 231319
rect 299446 231255 299498 231261
rect 300214 231313 300266 231319
rect 300214 231255 300266 231261
rect 299254 230499 299306 230505
rect 299254 230441 299306 230447
rect 298678 230425 298730 230431
rect 298678 230367 298730 230373
rect 298006 229685 298058 229691
rect 298006 229627 298058 229633
rect 298582 229685 298634 229691
rect 298582 229627 298634 229633
rect 297622 226281 297674 226287
rect 297622 226223 297674 226229
rect 297238 226207 297290 226213
rect 297238 226149 297290 226155
rect 296448 221468 296510 221496
rect 297250 221482 297278 226149
rect 298018 221482 298046 229627
rect 298690 221792 298718 230367
rect 298690 221764 298766 221792
rect 298738 221482 298766 221764
rect 299458 221482 299486 231255
rect 300706 226139 300734 239686
rect 301056 239672 301310 239700
rect 301440 239672 301694 239700
rect 301776 239672 302078 239700
rect 300982 230351 301034 230357
rect 300982 230293 301034 230299
rect 300214 226133 300266 226139
rect 300214 226075 300266 226081
rect 300694 226133 300746 226139
rect 300694 226075 300746 226081
rect 300226 221482 300254 226075
rect 300994 221792 301022 230293
rect 301282 226213 301310 239672
rect 301666 234057 301694 239672
rect 301654 234051 301706 234057
rect 301654 233993 301706 233999
rect 301750 228575 301802 228581
rect 301750 228517 301802 228523
rect 301270 226207 301322 226213
rect 301270 226149 301322 226155
rect 300994 221764 301070 221792
rect 301042 221482 301070 221764
rect 301762 221482 301790 228517
rect 302050 222587 302078 239672
rect 302146 236174 302174 239686
rect 302544 239672 302846 239700
rect 302146 236146 302270 236174
rect 302134 234347 302186 234353
rect 302134 234289 302186 234295
rect 302146 227915 302174 234289
rect 302134 227909 302186 227915
rect 302134 227851 302186 227857
rect 302242 225325 302270 236146
rect 302326 235383 302378 235389
rect 302326 235325 302378 235331
rect 302338 230653 302366 235325
rect 302326 230647 302378 230653
rect 302326 230589 302378 230595
rect 302518 230499 302570 230505
rect 302518 230441 302570 230447
rect 302230 225319 302282 225325
rect 302230 225261 302282 225267
rect 302038 222581 302090 222587
rect 302038 222523 302090 222529
rect 302530 221482 302558 230441
rect 302818 222661 302846 239672
rect 302914 233613 302942 239686
rect 303264 239672 303518 239700
rect 303648 239672 303902 239700
rect 303984 239672 304286 239700
rect 302902 233607 302954 233613
rect 302902 233549 302954 233555
rect 303490 228581 303518 239672
rect 303478 228575 303530 228581
rect 303478 228517 303530 228523
rect 303874 225399 303902 239672
rect 304150 234717 304202 234723
rect 304150 234659 304202 234665
rect 304162 230505 304190 234659
rect 304150 230499 304202 230505
rect 304150 230441 304202 230447
rect 303958 230203 304010 230209
rect 303958 230145 304010 230151
rect 303190 225393 303242 225399
rect 303190 225335 303242 225341
rect 303862 225393 303914 225399
rect 303862 225335 303914 225341
rect 302806 222655 302858 222661
rect 302806 222597 302858 222603
rect 303202 221792 303230 225335
rect 303202 221764 303278 221792
rect 303250 221482 303278 221764
rect 303970 221482 303998 230145
rect 304258 222883 304286 239672
rect 304450 228803 304478 239686
rect 304834 235389 304862 239686
rect 305184 239672 305246 239700
rect 305568 239672 305822 239700
rect 305952 239672 306206 239700
rect 305014 235753 305066 235759
rect 305014 235695 305066 235701
rect 304822 235383 304874 235389
rect 304822 235325 304874 235331
rect 304822 230277 304874 230283
rect 304822 230219 304874 230225
rect 304438 228797 304490 228803
rect 304438 228739 304490 228745
rect 304246 222877 304298 222883
rect 304246 222819 304298 222825
rect 304834 221482 304862 230219
rect 305026 225177 305054 235695
rect 305110 234495 305162 234501
rect 305110 234437 305162 234443
rect 305122 228063 305150 234437
rect 305218 233983 305246 239672
rect 305794 237017 305822 239672
rect 305782 237011 305834 237017
rect 305782 236953 305834 236959
rect 305206 233977 305258 233983
rect 305206 233919 305258 233925
rect 305494 231535 305546 231541
rect 305494 231477 305546 231483
rect 305110 228057 305162 228063
rect 305110 227999 305162 228005
rect 305014 225171 305066 225177
rect 305014 225113 305066 225119
rect 305506 221792 305534 231477
rect 306178 228729 306206 239672
rect 306274 233687 306302 239686
rect 306262 233681 306314 233687
rect 306262 233623 306314 233629
rect 306166 228723 306218 228729
rect 306166 228665 306218 228671
rect 306262 227539 306314 227545
rect 306262 227481 306314 227487
rect 305506 221764 305582 221792
rect 305554 221482 305582 221764
rect 306274 221482 306302 227481
rect 306658 225473 306686 239686
rect 307056 239672 307262 239700
rect 307392 239672 307646 239700
rect 307776 239672 308030 239700
rect 308256 239672 308510 239700
rect 306742 234791 306794 234797
rect 306742 234733 306794 234739
rect 306754 230579 306782 234733
rect 306742 230573 306794 230579
rect 306742 230515 306794 230521
rect 307030 230129 307082 230135
rect 307030 230071 307082 230077
rect 306646 225467 306698 225473
rect 306646 225409 306698 225415
rect 307042 221482 307070 230071
rect 307234 222957 307262 239672
rect 307618 231139 307646 239672
rect 307604 231130 307660 231139
rect 307604 231065 307660 231074
rect 307702 228353 307754 228359
rect 307702 228295 307754 228301
rect 307222 222951 307274 222957
rect 307222 222893 307274 222899
rect 307714 221792 307742 228295
rect 308002 222809 308030 239672
rect 308182 235309 308234 235315
rect 308182 235251 308234 235257
rect 308194 231023 308222 235251
rect 308482 234353 308510 239672
rect 308578 237165 308606 239686
rect 308566 237159 308618 237165
rect 308566 237101 308618 237107
rect 308470 234347 308522 234353
rect 308470 234289 308522 234295
rect 308182 231017 308234 231023
rect 308182 230959 308234 230965
rect 308566 230647 308618 230653
rect 308566 230589 308618 230595
rect 307990 222803 308042 222809
rect 307990 222745 308042 222751
rect 307714 221764 307790 221792
rect 307762 221482 307790 221764
rect 308578 221482 308606 230589
rect 308962 228951 308990 239686
rect 309346 235093 309374 239686
rect 309696 239672 309950 239700
rect 310080 239672 310334 239700
rect 310464 239672 310718 239700
rect 309334 235087 309386 235093
rect 309334 235029 309386 235035
rect 308950 228945 309002 228951
rect 308950 228887 309002 228893
rect 309334 225615 309386 225621
rect 309334 225557 309386 225563
rect 309346 221482 309374 225557
rect 309922 225547 309950 239672
rect 310198 236049 310250 236055
rect 310198 235991 310250 235997
rect 310210 228063 310238 235991
rect 310102 228057 310154 228063
rect 310102 227999 310154 228005
rect 310198 228057 310250 228063
rect 310198 227999 310250 228005
rect 310114 227841 310142 227999
rect 310006 227835 310058 227841
rect 310006 227777 310058 227783
rect 310102 227835 310154 227841
rect 310102 227777 310154 227783
rect 309910 225541 309962 225547
rect 309910 225483 309962 225489
rect 310018 221792 310046 227777
rect 310306 223105 310334 239672
rect 310690 228877 310718 239672
rect 310786 237091 310814 239686
rect 310774 237085 310826 237091
rect 310774 237027 310826 237033
rect 311170 235611 311198 239686
rect 311554 237239 311582 239686
rect 312000 239672 312254 239700
rect 312384 239672 312638 239700
rect 311542 237233 311594 237239
rect 311542 237175 311594 237181
rect 311158 235605 311210 235611
rect 311158 235547 311210 235553
rect 311158 234421 311210 234427
rect 311158 234363 311210 234369
rect 311062 233385 311114 233391
rect 311062 233327 311114 233333
rect 310774 230055 310826 230061
rect 310774 229997 310826 230003
rect 310678 228871 310730 228877
rect 310678 228813 310730 228819
rect 310294 223099 310346 223105
rect 310294 223041 310346 223047
rect 310018 221764 310094 221792
rect 310066 221482 310094 221764
rect 310786 221482 310814 229997
rect 311074 228285 311102 233327
rect 311170 228359 311198 234363
rect 311350 234199 311402 234205
rect 311350 234141 311402 234147
rect 311254 233459 311306 233465
rect 311254 233401 311306 233407
rect 311158 228353 311210 228359
rect 311158 228295 311210 228301
rect 311062 228279 311114 228285
rect 311062 228221 311114 228227
rect 311266 227397 311294 233401
rect 311362 227545 311390 234141
rect 312226 231541 312254 239672
rect 312214 231535 312266 231541
rect 312214 231477 312266 231483
rect 311638 230499 311690 230505
rect 311638 230441 311690 230447
rect 311350 227539 311402 227545
rect 311350 227481 311402 227487
rect 311254 227391 311306 227397
rect 311254 227333 311306 227339
rect 311650 221482 311678 230441
rect 312310 225097 312362 225103
rect 312310 225039 312362 225045
rect 312322 221792 312350 225039
rect 312610 223031 312638 239672
rect 312706 234427 312734 239686
rect 313104 239672 313406 239700
rect 312694 234421 312746 234427
rect 312694 234363 312746 234369
rect 313078 229981 313130 229987
rect 313078 229923 313130 229929
rect 312598 223025 312650 223031
rect 312598 222967 312650 222973
rect 312322 221764 312398 221792
rect 312370 221482 312398 221764
rect 313090 221482 313118 229923
rect 313378 223179 313406 239672
rect 313474 230209 313502 239686
rect 313858 236055 313886 239686
rect 314208 239672 314462 239700
rect 314592 239672 314846 239700
rect 313942 236123 313994 236129
rect 313942 236065 313994 236071
rect 313846 236049 313898 236055
rect 313846 235991 313898 235997
rect 313954 230801 313982 236065
rect 314434 234501 314462 239672
rect 314818 237313 314846 239672
rect 314806 237307 314858 237313
rect 314806 237249 314858 237255
rect 314422 234495 314474 234501
rect 314422 234437 314474 234443
rect 314518 231091 314570 231097
rect 314518 231033 314570 231039
rect 313942 230795 313994 230801
rect 313942 230737 313994 230743
rect 313462 230203 313514 230209
rect 313462 230145 313514 230151
rect 313846 228501 313898 228507
rect 313846 228443 313898 228449
rect 313366 223173 313418 223179
rect 313366 223115 313418 223121
rect 313858 221482 313886 228443
rect 314530 221792 314558 231033
rect 314914 230357 314942 239686
rect 315298 234723 315326 239686
rect 315286 234717 315338 234723
rect 315286 234659 315338 234665
rect 314902 230351 314954 230357
rect 314902 230293 314954 230299
rect 315382 227465 315434 227471
rect 315382 227407 315434 227413
rect 314530 221764 314606 221792
rect 314578 221482 314606 221764
rect 315394 221482 315422 227407
rect 315778 225621 315806 239686
rect 316176 239672 316382 239700
rect 316512 239672 316766 239700
rect 316896 239672 317150 239700
rect 316150 229759 316202 229765
rect 316150 229701 316202 229707
rect 315766 225615 315818 225621
rect 315766 225557 315818 225563
rect 316162 221482 316190 229701
rect 316354 224659 316382 239672
rect 316738 231287 316766 239672
rect 317122 237387 317150 239672
rect 317110 237381 317162 237387
rect 317110 237323 317162 237329
rect 317218 235759 317246 239686
rect 317602 237461 317630 239686
rect 317590 237455 317642 237461
rect 317590 237397 317642 237403
rect 317206 235753 317258 235759
rect 317206 235695 317258 235701
rect 317878 233311 317930 233317
rect 317878 233253 317930 233259
rect 316724 231278 316780 231287
rect 316724 231213 316780 231222
rect 317590 230573 317642 230579
rect 317590 230515 317642 230521
rect 316822 229611 316874 229617
rect 316822 229553 316874 229559
rect 316342 224653 316394 224659
rect 316342 224595 316394 224601
rect 316834 221792 316862 229553
rect 316834 221764 316910 221792
rect 316882 221482 316910 221764
rect 317602 221482 317630 230515
rect 317890 228507 317918 233253
rect 317986 230283 318014 239686
rect 318262 235901 318314 235907
rect 318262 235843 318314 235849
rect 318274 230727 318302 235843
rect 318370 234205 318398 239686
rect 318720 239672 318974 239700
rect 319200 239672 319454 239700
rect 318454 235679 318506 235685
rect 318454 235621 318506 235627
rect 318358 234199 318410 234205
rect 318358 234141 318410 234147
rect 318262 230721 318314 230727
rect 318262 230663 318314 230669
rect 317974 230277 318026 230283
rect 317974 230219 318026 230225
rect 317878 228501 317930 228507
rect 317878 228443 317930 228449
rect 318466 227471 318494 235621
rect 318454 227465 318506 227471
rect 318454 227407 318506 227413
rect 318358 225689 318410 225695
rect 318358 225631 318410 225637
rect 318370 221482 318398 225631
rect 318946 225367 318974 239672
rect 319126 229833 319178 229839
rect 319126 229775 319178 229781
rect 318932 225358 318988 225367
rect 318932 225293 318988 225302
rect 319138 221792 319166 229775
rect 319426 224585 319454 239672
rect 319522 231435 319550 239686
rect 319906 233317 319934 239686
rect 320290 233465 320318 239686
rect 320640 239672 320894 239700
rect 321024 239672 321278 239700
rect 321408 239672 321662 239700
rect 320866 237535 320894 239672
rect 320854 237529 320906 237535
rect 320854 237471 320906 237477
rect 320278 233459 320330 233465
rect 320278 233401 320330 233407
rect 319894 233311 319946 233317
rect 319894 233253 319946 233259
rect 320662 231609 320714 231615
rect 320662 231551 320714 231557
rect 319508 231426 319564 231435
rect 319508 231361 319564 231370
rect 319894 227687 319946 227693
rect 319894 227629 319946 227635
rect 319414 224579 319466 224585
rect 319414 224521 319466 224527
rect 319138 221764 319214 221792
rect 319186 221482 319214 221764
rect 319906 221482 319934 227629
rect 320674 221482 320702 231551
rect 321250 227693 321278 239672
rect 321634 234797 321662 239672
rect 321622 234791 321674 234797
rect 321622 234733 321674 234739
rect 321238 227687 321290 227693
rect 321238 227629 321290 227635
rect 321334 225985 321386 225991
rect 321334 225927 321386 225933
rect 321346 221792 321374 225927
rect 321730 225695 321758 239686
rect 322128 239672 322334 239700
rect 322006 235975 322058 235981
rect 322006 235917 322058 235923
rect 322018 230505 322046 235917
rect 322198 234569 322250 234575
rect 322198 234511 322250 234517
rect 322102 231165 322154 231171
rect 322102 231107 322154 231113
rect 322006 230499 322058 230505
rect 322006 230441 322058 230447
rect 321718 225689 321770 225695
rect 321718 225631 321770 225637
rect 321346 221764 321422 221792
rect 321394 221482 321422 221764
rect 322114 221482 322142 231107
rect 322210 230653 322238 234511
rect 322198 230647 322250 230653
rect 322198 230589 322250 230595
rect 322306 224437 322334 239672
rect 322498 231583 322526 239686
rect 322944 239672 323198 239700
rect 323328 239672 323582 239700
rect 323712 239672 323966 239700
rect 323170 236174 323198 239672
rect 323170 236146 323294 236174
rect 323158 234865 323210 234871
rect 323158 234807 323210 234813
rect 322484 231574 322540 231583
rect 322484 231509 322540 231518
rect 323170 230949 323198 234807
rect 323158 230943 323210 230949
rect 323158 230885 323210 230891
rect 322966 228205 323018 228211
rect 322966 228147 323018 228153
rect 322294 224431 322346 224437
rect 322294 224373 322346 224379
rect 322978 221496 323006 228147
rect 323266 224511 323294 236146
rect 323554 234575 323582 239672
rect 323938 238941 323966 239672
rect 323926 238935 323978 238941
rect 323926 238877 323978 238883
rect 323542 234569 323594 234575
rect 323542 234511 323594 234517
rect 323638 231017 323690 231023
rect 323638 230959 323690 230965
rect 323254 224505 323306 224511
rect 323254 224447 323306 224453
rect 322944 221468 323006 221496
rect 323650 221496 323678 230959
rect 324034 230431 324062 239686
rect 324418 239015 324446 239686
rect 324406 239009 324458 239015
rect 324406 238951 324458 238957
rect 324118 235161 324170 235167
rect 324118 235103 324170 235109
rect 324022 230425 324074 230431
rect 324022 230367 324074 230373
rect 324130 226879 324158 235103
rect 324802 233391 324830 239686
rect 325152 239672 325214 239700
rect 325536 239672 325790 239700
rect 325920 239672 326174 239700
rect 325186 236174 325214 239672
rect 325762 236174 325790 239672
rect 325186 236146 325310 236174
rect 325762 236146 325886 236174
rect 324790 233385 324842 233391
rect 324790 233327 324842 233333
rect 325174 231683 325226 231689
rect 325174 231625 325226 231631
rect 324118 226873 324170 226879
rect 324118 226815 324170 226821
rect 324406 225763 324458 225769
rect 324406 225705 324458 225711
rect 323650 221468 323712 221496
rect 324418 221482 324446 225705
rect 325186 221496 325214 231625
rect 325282 224363 325310 236146
rect 325750 234643 325802 234649
rect 325750 234585 325802 234591
rect 325366 233829 325418 233835
rect 325366 233771 325418 233777
rect 325378 230579 325406 233771
rect 325762 230875 325790 234585
rect 325750 230869 325802 230875
rect 325750 230811 325802 230817
rect 325366 230573 325418 230579
rect 325366 230515 325418 230521
rect 325858 230135 325886 236146
rect 326146 236129 326174 239672
rect 326134 236123 326186 236129
rect 326134 236065 326186 236071
rect 326242 235907 326270 239686
rect 326722 238867 326750 239686
rect 326710 238861 326762 238867
rect 326710 238803 326762 238809
rect 326230 235901 326282 235907
rect 326230 235843 326282 235849
rect 326710 233237 326762 233243
rect 326710 233179 326762 233185
rect 325846 230129 325898 230135
rect 325846 230071 325898 230077
rect 325846 227761 325898 227767
rect 325846 227703 325898 227709
rect 325270 224357 325322 224363
rect 325270 224299 325322 224305
rect 325152 221468 325214 221496
rect 325858 221496 325886 227703
rect 325858 221468 325920 221496
rect 326722 221482 326750 233179
rect 327106 231615 327134 239686
rect 327456 239672 327710 239700
rect 327840 239672 328094 239700
rect 327682 234871 327710 239672
rect 327670 234865 327722 234871
rect 327670 234807 327722 234813
rect 327286 233385 327338 233391
rect 327286 233327 327338 233333
rect 327094 231609 327146 231615
rect 327094 231551 327146 231557
rect 327298 225515 327326 233327
rect 327382 225911 327434 225917
rect 327382 225853 327434 225859
rect 327284 225506 327340 225515
rect 327284 225441 327340 225450
rect 327394 221792 327422 225853
rect 328066 225663 328094 239672
rect 328162 236174 328190 239686
rect 328162 236146 328286 236174
rect 328150 231757 328202 231763
rect 328150 231699 328202 231705
rect 328052 225654 328108 225663
rect 328052 225589 328108 225598
rect 327394 221764 327470 221792
rect 327442 221482 327470 221764
rect 328162 221482 328190 231699
rect 328258 224141 328286 236146
rect 328342 233533 328394 233539
rect 328342 233475 328394 233481
rect 328354 231023 328382 233475
rect 328342 231017 328394 231023
rect 328342 230959 328394 230965
rect 328546 230061 328574 239686
rect 328930 238793 328958 239686
rect 328918 238787 328970 238793
rect 328918 238729 328970 238735
rect 329314 234649 329342 239686
rect 329664 239672 329918 239700
rect 330048 239672 330302 239700
rect 330480 239672 330782 239700
rect 329890 238719 329918 239672
rect 329878 238713 329930 238719
rect 329878 238655 329930 238661
rect 329302 234643 329354 234649
rect 329302 234585 329354 234591
rect 330274 231731 330302 239672
rect 330260 231722 330316 231731
rect 330260 231657 330316 231666
rect 329590 230943 329642 230949
rect 329590 230885 329642 230891
rect 328534 230055 328586 230061
rect 328534 229997 328586 230003
rect 328918 227613 328970 227619
rect 328918 227555 328970 227561
rect 328246 224135 328298 224141
rect 328246 224077 328298 224083
rect 328930 221482 328958 227555
rect 329602 221792 329630 230885
rect 330454 225837 330506 225843
rect 330454 225779 330506 225785
rect 329602 221764 329678 221792
rect 329650 221482 329678 221764
rect 330466 221482 330494 225779
rect 330754 224215 330782 239672
rect 330850 225811 330878 239686
rect 331248 239672 331550 239700
rect 331414 234939 331466 234945
rect 331414 234881 331466 234887
rect 331222 233755 331274 233761
rect 331222 233697 331274 233703
rect 331234 230949 331262 233697
rect 331318 233163 331370 233169
rect 331318 233105 331370 233111
rect 331222 230943 331274 230949
rect 331222 230885 331274 230891
rect 331330 226972 331358 233105
rect 331234 226944 331358 226972
rect 330836 225802 330892 225811
rect 330836 225737 330892 225746
rect 330742 224209 330794 224215
rect 330742 224151 330794 224157
rect 331234 221482 331262 226944
rect 331426 225917 331454 234881
rect 331414 225911 331466 225917
rect 331414 225853 331466 225859
rect 331522 224289 331550 239672
rect 331618 229987 331646 239686
rect 331968 239672 332222 239700
rect 332352 239672 332606 239700
rect 332194 235167 332222 239672
rect 332182 235161 332234 235167
rect 332182 235103 332234 235109
rect 332578 234099 332606 239672
rect 332674 238645 332702 239686
rect 332662 238639 332714 238645
rect 332662 238581 332714 238587
rect 332564 234090 332620 234099
rect 332564 234025 332620 234034
rect 331606 229981 331658 229987
rect 331606 229923 331658 229929
rect 331894 229907 331946 229913
rect 331894 229849 331946 229855
rect 331510 224283 331562 224289
rect 331510 224225 331562 224231
rect 331906 221792 331934 229849
rect 333058 228179 333086 239686
rect 333442 234945 333470 239686
rect 333430 234939 333482 234945
rect 333430 234881 333482 234887
rect 333826 231879 333854 239686
rect 334272 239672 334526 239700
rect 334656 239672 334910 239700
rect 334294 239527 334346 239533
rect 334294 239469 334346 239475
rect 334306 236129 334334 239469
rect 334294 236123 334346 236129
rect 334294 236065 334346 236071
rect 334102 235827 334154 235833
rect 334102 235769 334154 235775
rect 333812 231870 333868 231879
rect 333812 231805 333868 231814
rect 333044 228170 333100 228179
rect 333044 228105 333100 228114
rect 333526 225171 333578 225177
rect 333526 225113 333578 225119
rect 332662 223691 332714 223697
rect 332662 223633 332714 223639
rect 331906 221764 331982 221792
rect 331954 221482 331982 221764
rect 332674 221482 332702 223633
rect 333538 221482 333566 225113
rect 334114 224807 334142 235769
rect 334198 233089 334250 233095
rect 334198 233031 334250 233037
rect 334102 224801 334154 224807
rect 334102 224743 334154 224749
rect 334210 221792 334238 233031
rect 334498 224067 334526 239672
rect 334882 231689 334910 239672
rect 334978 235315 335006 239686
rect 334966 235309 335018 235315
rect 334966 235251 335018 235257
rect 335362 233391 335390 239686
rect 335746 238571 335774 239686
rect 336096 239672 336350 239700
rect 336480 239672 336734 239700
rect 335734 238565 335786 238571
rect 335734 238507 335786 238513
rect 335350 233385 335402 233391
rect 335350 233327 335402 233333
rect 334870 231683 334922 231689
rect 334870 231625 334922 231631
rect 336322 229839 336350 239672
rect 336706 238497 336734 239672
rect 336850 239404 336878 239686
rect 336850 239376 336926 239404
rect 336694 238491 336746 238497
rect 336694 238433 336746 238439
rect 336310 229833 336362 229839
rect 336310 229775 336362 229781
rect 334966 229537 335018 229543
rect 334966 229479 335018 229485
rect 334486 224061 334538 224067
rect 334486 224003 334538 224009
rect 334210 221764 334286 221792
rect 334258 221482 334286 221764
rect 334978 221482 335006 229479
rect 336898 227439 336926 239376
rect 336884 227430 336940 227439
rect 336884 227365 336940 227374
rect 336406 226059 336458 226065
rect 336406 226001 336458 226007
rect 335734 223765 335786 223771
rect 335734 223707 335786 223713
rect 335746 221482 335774 223707
rect 336418 221792 336446 226001
rect 337186 223993 337214 239686
rect 337366 233607 337418 233613
rect 337366 233549 337418 233555
rect 337270 232867 337322 232873
rect 337270 232809 337322 232815
rect 337174 223987 337226 223993
rect 337174 223929 337226 223935
rect 336418 221764 336494 221792
rect 336466 221482 336494 221764
rect 337282 221482 337310 232809
rect 337378 231171 337406 233549
rect 337570 231763 337598 239686
rect 338050 233761 338078 239686
rect 338400 239672 338654 239700
rect 338784 239672 339038 239700
rect 339168 239672 339422 239700
rect 338038 233755 338090 233761
rect 338038 233697 338090 233703
rect 338626 233539 338654 239672
rect 339010 238423 339038 239672
rect 338998 238417 339050 238423
rect 338998 238359 339050 238365
rect 338902 235457 338954 235463
rect 338902 235399 338954 235405
rect 338614 233533 338666 233539
rect 338614 233475 338666 233481
rect 338038 233015 338090 233021
rect 338038 232957 338090 232963
rect 337558 231757 337610 231763
rect 337558 231699 337610 231705
rect 337366 231165 337418 231171
rect 337366 231107 337418 231113
rect 338050 221482 338078 232957
rect 338914 225769 338942 235399
rect 339094 233903 339146 233909
rect 339094 233845 339146 233851
rect 338902 225763 338954 225769
rect 338902 225705 338954 225711
rect 339106 225177 339134 233845
rect 339394 228327 339422 239672
rect 339490 235463 339518 239686
rect 339888 239672 340190 239700
rect 340272 239672 340478 239700
rect 340608 239672 340862 239700
rect 340992 239672 341246 239700
rect 341376 239672 341630 239700
rect 339478 235457 339530 235463
rect 339478 235399 339530 235405
rect 339380 228318 339436 228327
rect 339380 228253 339436 228262
rect 339478 226873 339530 226879
rect 339478 226815 339530 226821
rect 339094 225171 339146 225177
rect 339094 225113 339146 225119
rect 338710 223469 338762 223475
rect 338710 223411 338762 223417
rect 338722 221792 338750 223411
rect 338722 221764 338798 221792
rect 338770 221482 338798 221764
rect 339490 221482 339518 226815
rect 340162 225959 340190 239672
rect 340246 232793 340298 232799
rect 340246 232735 340298 232741
rect 340148 225950 340204 225959
rect 340148 225885 340204 225894
rect 340258 221482 340286 232735
rect 340450 223919 340478 239672
rect 340834 233243 340862 239672
rect 341218 236129 341246 239672
rect 341206 236123 341258 236129
rect 341206 236065 341258 236071
rect 341602 234247 341630 239672
rect 341794 238349 341822 239686
rect 341782 238343 341834 238349
rect 341782 238285 341834 238291
rect 341588 234238 341644 234247
rect 341588 234173 341644 234182
rect 341206 234125 341258 234131
rect 341206 234067 341258 234073
rect 340822 233237 340874 233243
rect 340822 233179 340874 233185
rect 341218 228137 341246 234067
rect 342178 228475 342206 239686
rect 342562 235727 342590 239686
rect 342912 239672 343166 239700
rect 343296 239672 343550 239700
rect 342548 235718 342604 235727
rect 342548 235653 342604 235662
rect 342164 228466 342220 228475
rect 342164 228401 342220 228410
rect 341014 228131 341066 228137
rect 341014 228073 341066 228079
rect 341206 228131 341258 228137
rect 341206 228073 341258 228079
rect 340438 223913 340490 223919
rect 340438 223855 340490 223861
rect 341026 221792 341054 228073
rect 343138 227291 343166 239672
rect 343522 235833 343550 239672
rect 343510 235827 343562 235833
rect 343510 235769 343562 235775
rect 343222 232645 343274 232651
rect 343222 232587 343274 232593
rect 343124 227282 343180 227291
rect 343124 227217 343180 227226
rect 342550 225245 342602 225251
rect 342550 225187 342602 225193
rect 341782 223617 341834 223623
rect 341782 223559 341834 223565
rect 341026 221764 341102 221792
rect 341074 221482 341102 221764
rect 341794 221482 341822 223559
rect 342562 221482 342590 225187
rect 343234 221792 343262 232587
rect 343618 223845 343646 239686
rect 344002 233211 344030 239686
rect 344386 234057 344414 239686
rect 344086 234051 344138 234057
rect 344086 233993 344138 233999
rect 344374 234051 344426 234057
rect 344374 233993 344426 233999
rect 343988 233202 344044 233211
rect 343988 233137 344044 233146
rect 344098 228211 344126 233993
rect 344470 233681 344522 233687
rect 344470 233623 344522 233629
rect 344482 231097 344510 233623
rect 344470 231091 344522 231097
rect 344470 231033 344522 231039
rect 344086 228205 344138 228211
rect 344086 228147 344138 228153
rect 343990 227983 344042 227989
rect 343990 227925 344042 227931
rect 343606 223839 343658 223845
rect 343606 223781 343658 223787
rect 343234 221764 343310 221792
rect 343282 221482 343310 221764
rect 344002 221482 344030 227925
rect 344770 227143 344798 239686
rect 345120 239672 345374 239700
rect 345346 238275 345374 239672
rect 345442 239672 345600 239700
rect 345334 238269 345386 238275
rect 345334 238211 345386 238217
rect 345442 228623 345470 239672
rect 345718 235235 345770 235241
rect 345718 235177 345770 235183
rect 345428 228614 345484 228623
rect 345428 228549 345484 228558
rect 344756 227134 344812 227143
rect 344756 227069 344812 227078
rect 345526 225911 345578 225917
rect 345526 225853 345578 225859
rect 344854 223543 344906 223549
rect 344854 223485 344906 223491
rect 344866 221482 344894 223485
rect 345538 221792 345566 225853
rect 345730 225843 345758 235177
rect 345922 234131 345950 239686
rect 346320 239672 346622 239700
rect 345910 234125 345962 234131
rect 345910 234067 345962 234073
rect 346294 232571 346346 232577
rect 346294 232513 346346 232519
rect 345718 225837 345770 225843
rect 345718 225779 345770 225785
rect 345538 221764 345614 221792
rect 345586 221482 345614 221764
rect 346306 221482 346334 232513
rect 346594 223771 346622 239672
rect 346690 238201 346718 239686
rect 346678 238195 346730 238201
rect 346678 238137 346730 238143
rect 347074 233169 347102 239686
rect 347424 239672 347678 239700
rect 347808 239672 348062 239700
rect 347650 234839 347678 239672
rect 347636 234830 347692 234839
rect 347636 234765 347692 234774
rect 347062 233163 347114 233169
rect 347062 233105 347114 233111
rect 346774 232571 346826 232577
rect 346774 232513 346826 232519
rect 346786 232355 346814 232513
rect 346966 232423 347018 232429
rect 346966 232365 347018 232371
rect 346774 232349 346826 232355
rect 346774 232291 346826 232297
rect 346978 232059 347006 232365
rect 346966 232053 347018 232059
rect 346966 231995 347018 232001
rect 346966 230425 347018 230431
rect 346966 230367 347018 230373
rect 346978 230061 347006 230367
rect 346966 230055 347018 230061
rect 346966 229997 347018 230003
rect 347062 229389 347114 229395
rect 347062 229331 347114 229337
rect 346582 223765 346634 223771
rect 346582 223707 346634 223713
rect 347074 221482 347102 229331
rect 348034 223549 348062 239672
rect 348130 223623 348158 239686
rect 348514 229765 348542 239686
rect 348694 234273 348746 234279
rect 348694 234215 348746 234221
rect 348502 229759 348554 229765
rect 348502 229701 348554 229707
rect 348598 227317 348650 227323
rect 348598 227259 348650 227265
rect 348118 223617 348170 223623
rect 348118 223559 348170 223565
rect 348022 223543 348074 223549
rect 348022 223485 348074 223491
rect 347734 223321 347786 223327
rect 347734 223263 347786 223269
rect 347746 221792 347774 223263
rect 347746 221764 347822 221792
rect 347794 221482 347822 221764
rect 348610 221482 348638 227259
rect 348706 225103 348734 234215
rect 348898 233613 348926 239686
rect 349344 239672 349598 239700
rect 349728 239672 349982 239700
rect 350112 239672 350366 239700
rect 348886 233607 348938 233613
rect 348886 233549 348938 233555
rect 349366 232497 349418 232503
rect 349366 232439 349418 232445
rect 348694 225097 348746 225103
rect 348694 225039 348746 225045
rect 349378 221482 349406 232439
rect 349570 223697 349598 239672
rect 349954 238127 349982 239672
rect 349942 238121 349994 238127
rect 349942 238063 349994 238069
rect 350338 233095 350366 239672
rect 350434 239163 350462 239686
rect 350832 239672 351134 239700
rect 350422 239157 350474 239163
rect 350422 239099 350474 239105
rect 350326 233089 350378 233095
rect 350326 233031 350378 233037
rect 350038 227909 350090 227915
rect 350038 227851 350090 227857
rect 349558 223691 349610 223697
rect 349558 223633 349610 223639
rect 350050 221792 350078 227851
rect 351106 223401 351134 239672
rect 350806 223395 350858 223401
rect 350806 223337 350858 223343
rect 351094 223395 351146 223401
rect 351094 223337 351146 223343
rect 350050 221764 350126 221792
rect 350098 221482 350126 221764
rect 350818 221482 350846 223337
rect 351202 223327 351230 239686
rect 351552 239672 351806 239700
rect 351936 239672 352190 239700
rect 352320 239672 352574 239700
rect 351382 233977 351434 233983
rect 351382 233919 351434 233925
rect 351394 225251 351422 233919
rect 351778 229617 351806 239672
rect 352162 234279 352190 239672
rect 352150 234273 352202 234279
rect 352150 234215 352202 234221
rect 352342 232349 352394 232355
rect 352342 232291 352394 232297
rect 351766 229611 351818 229617
rect 351766 229553 351818 229559
rect 351574 227243 351626 227249
rect 351574 227185 351626 227191
rect 351382 225245 351434 225251
rect 351382 225187 351434 225193
rect 351190 223321 351242 223327
rect 351190 223263 351242 223269
rect 351586 221482 351614 227185
rect 352354 221496 352382 232291
rect 352546 223475 352574 239672
rect 352738 237979 352766 239686
rect 352726 237973 352778 237979
rect 352726 237915 352778 237921
rect 353122 233021 353150 239686
rect 353506 238053 353534 239686
rect 353856 239672 354014 239700
rect 353494 238047 353546 238053
rect 353494 237989 353546 237995
rect 353110 233015 353162 233021
rect 353110 232957 353162 232963
rect 353110 227835 353162 227841
rect 353110 227777 353162 227783
rect 352534 223469 352586 223475
rect 352534 223411 352586 223417
rect 352354 221468 352416 221496
rect 353122 221482 353150 227777
rect 353986 223253 354014 239672
rect 354082 239672 354240 239700
rect 354624 239672 354878 239700
rect 354082 224627 354110 239672
rect 354262 235531 354314 235537
rect 354262 235473 354314 235479
rect 354274 232059 354302 235473
rect 354262 232053 354314 232059
rect 354262 231995 354314 232001
rect 354850 229543 354878 239672
rect 354946 233835 354974 239686
rect 355344 239672 355646 239700
rect 354934 233829 354986 233835
rect 354934 233771 354986 233777
rect 355318 232201 355370 232207
rect 355318 232143 355370 232149
rect 354838 229537 354890 229543
rect 354838 229479 354890 229485
rect 354550 226873 354602 226879
rect 354550 226815 354602 226821
rect 354068 224618 354124 224627
rect 354068 224553 354124 224562
rect 353878 223247 353930 223253
rect 353878 223189 353930 223195
rect 353974 223247 354026 223253
rect 353974 223189 354026 223195
rect 353890 221496 353918 223189
rect 353856 221468 353918 221496
rect 354562 221496 354590 226815
rect 354562 221468 354624 221496
rect 355330 221482 355358 232143
rect 355618 222703 355646 239672
rect 355714 237905 355742 239686
rect 356064 239672 356318 239700
rect 356544 239672 356798 239700
rect 355702 237899 355754 237905
rect 355702 237841 355754 237847
rect 355892 234978 355948 234987
rect 355892 234913 355948 234922
rect 355906 226879 355934 234913
rect 356290 232873 356318 239672
rect 356770 234987 356798 239672
rect 356866 236171 356894 239686
rect 356852 236162 356908 236171
rect 356852 236097 356908 236106
rect 357154 236055 357182 239765
rect 377302 239749 377354 239755
rect 357142 236049 357194 236055
rect 357142 235991 357194 235997
rect 356756 234978 356812 234987
rect 356756 234913 356812 234922
rect 356278 232867 356330 232873
rect 356278 232809 356330 232815
rect 356086 232571 356138 232577
rect 356086 232513 356138 232519
rect 355894 226873 355946 226879
rect 355894 226815 355946 226821
rect 355604 222694 355660 222703
rect 355604 222629 355660 222638
rect 356098 221792 356126 232513
rect 357250 224479 357278 239686
rect 357526 237751 357578 237757
rect 357526 237693 357578 237699
rect 357538 228063 357566 237693
rect 357634 229395 357662 239686
rect 358018 235685 358046 239686
rect 358368 239672 358622 239700
rect 358752 239672 359006 239700
rect 358006 235679 358058 235685
rect 358006 235621 358058 235627
rect 358294 232275 358346 232281
rect 358294 232217 358346 232223
rect 357622 229389 357674 229395
rect 357622 229331 357674 229337
rect 357526 228057 357578 228063
rect 357526 227999 357578 228005
rect 357622 227021 357674 227027
rect 357622 226963 357674 226969
rect 357236 224470 357292 224479
rect 357236 224405 357292 224414
rect 356854 222359 356906 222365
rect 356854 222301 356906 222307
rect 356098 221764 356174 221792
rect 356146 221482 356174 221764
rect 356866 221482 356894 222301
rect 357634 221482 357662 226963
rect 358306 221792 358334 232217
rect 358594 222999 358622 239672
rect 358978 230103 359006 239672
rect 359074 232799 359102 239686
rect 359062 232793 359114 232799
rect 359062 232735 359114 232741
rect 358964 230094 359020 230103
rect 358964 230029 359020 230038
rect 359158 227983 359210 227989
rect 359158 227925 359210 227931
rect 358580 222990 358636 222999
rect 358580 222925 358636 222934
rect 358306 221764 358382 221792
rect 358354 221482 358382 221764
rect 359170 221482 359198 227925
rect 359458 222851 359486 239686
rect 359842 236174 359870 239686
rect 359746 236146 359870 236174
rect 359746 224035 359774 236146
rect 359828 229058 359884 229067
rect 359828 228993 359884 229002
rect 359842 227101 359870 228993
rect 359926 228057 359978 228063
rect 359926 227999 359978 228005
rect 359830 227095 359882 227101
rect 359830 227037 359882 227043
rect 359732 224026 359788 224035
rect 359732 223961 359788 223970
rect 359444 222842 359500 222851
rect 359444 222777 359500 222786
rect 359938 221482 359966 227999
rect 360322 224331 360350 239686
rect 360672 239672 360830 239700
rect 361056 239672 361310 239700
rect 360802 228771 360830 239672
rect 361282 233983 361310 239672
rect 361378 236174 361406 239686
rect 361762 237757 361790 239686
rect 361750 237751 361802 237757
rect 361750 237693 361802 237699
rect 361378 236146 361502 236174
rect 361270 233977 361322 233983
rect 361270 233919 361322 233925
rect 361366 232423 361418 232429
rect 361366 232365 361418 232371
rect 360788 228762 360844 228771
rect 360788 228697 360844 228706
rect 360598 226947 360650 226953
rect 360598 226889 360650 226895
rect 360308 224322 360364 224331
rect 360308 224257 360364 224266
rect 360610 221792 360638 226889
rect 360610 221764 360686 221792
rect 360658 221482 360686 221764
rect 361378 221482 361406 232365
rect 361474 224183 361502 236146
rect 362146 232651 362174 239686
rect 362326 235383 362378 235389
rect 362326 235325 362378 235331
rect 362134 232645 362186 232651
rect 362134 232587 362186 232593
rect 362338 230801 362366 235325
rect 362530 235019 362558 239686
rect 362880 239672 363134 239700
rect 363264 239672 363518 239700
rect 363106 237831 363134 239672
rect 363094 237825 363146 237831
rect 363094 237767 363146 237773
rect 362422 235013 362474 235019
rect 362422 234955 362474 234961
rect 362518 235013 362570 235019
rect 362518 234955 362570 234961
rect 362134 230795 362186 230801
rect 362134 230737 362186 230743
rect 362326 230795 362378 230801
rect 362326 230737 362378 230743
rect 361460 224174 361516 224183
rect 361460 224109 361516 224118
rect 362146 221482 362174 230737
rect 362434 224733 362462 234955
rect 363490 233687 363518 239672
rect 363478 233681 363530 233687
rect 363478 233623 363530 233629
rect 363586 230251 363614 239686
rect 363670 237677 363722 237683
rect 363670 237619 363722 237625
rect 363572 230242 363628 230251
rect 363572 230177 363628 230186
rect 362804 229206 362860 229215
rect 362804 229141 362860 229150
rect 362818 224955 362846 229141
rect 363682 227268 363710 237619
rect 364066 233803 364094 239686
rect 364450 237683 364478 239686
rect 364800 239672 365054 239700
rect 365184 239672 365438 239700
rect 365568 239672 365726 239700
rect 364438 237677 364490 237683
rect 364438 237619 364490 237625
rect 364052 233794 364108 233803
rect 364052 233729 364108 233738
rect 363766 233681 363818 233687
rect 363766 233623 363818 233629
rect 363010 227240 363710 227268
rect 362806 224949 362858 224955
rect 362806 224891 362858 224897
rect 362422 224727 362474 224733
rect 362422 224669 362474 224675
rect 363010 221792 363038 227240
rect 363670 224875 363722 224881
rect 363670 224817 363722 224823
rect 362962 221764 363038 221792
rect 362962 221482 362990 221764
rect 363682 221482 363710 224817
rect 363778 223887 363806 233623
rect 365026 232503 365054 239672
rect 365410 232577 365438 239672
rect 365698 233359 365726 239672
rect 365890 237609 365918 239686
rect 365878 237603 365930 237609
rect 365878 237545 365930 237551
rect 365684 233350 365740 233359
rect 365684 233285 365740 233294
rect 365398 232571 365450 232577
rect 365398 232513 365450 232519
rect 365014 232497 365066 232503
rect 365014 232439 365066 232445
rect 366274 232355 366302 239686
rect 366262 232349 366314 232355
rect 366262 232291 366314 232297
rect 364438 232127 364490 232133
rect 364438 232069 364490 232075
rect 363764 223878 363820 223887
rect 363764 223813 363820 223822
rect 364450 221482 364478 232069
rect 365590 231239 365642 231245
rect 365590 231181 365642 231187
rect 365110 230721 365162 230727
rect 365110 230663 365162 230669
rect 365122 221792 365150 230663
rect 365602 227249 365630 231181
rect 366658 229955 366686 239686
rect 367008 239672 367262 239700
rect 367392 239672 367646 239700
rect 367872 239672 368126 239700
rect 366742 236789 366794 236795
rect 366742 236731 366794 236737
rect 366644 229946 366700 229955
rect 366644 229881 366700 229890
rect 365684 228910 365740 228919
rect 365684 228845 365740 228854
rect 365590 227243 365642 227249
rect 365590 227185 365642 227191
rect 365698 227027 365726 228845
rect 366754 228600 366782 236731
rect 367234 235579 367262 239672
rect 367220 235570 367276 235579
rect 367220 235505 367276 235514
rect 367126 232053 367178 232059
rect 367126 231995 367178 232001
rect 367138 230727 367166 231995
rect 367414 231905 367466 231911
rect 367414 231847 367466 231853
rect 367126 230721 367178 230727
rect 367126 230663 367178 230669
rect 365890 228572 366782 228600
rect 365686 227021 365738 227027
rect 365686 226963 365738 226969
rect 365122 221764 365198 221792
rect 365170 221482 365198 221764
rect 365890 221482 365918 228572
rect 367126 227243 367178 227249
rect 367126 227185 367178 227191
rect 367030 226947 367082 226953
rect 367030 226889 367082 226895
rect 366838 226873 366890 226879
rect 367042 226824 367070 226889
rect 367138 226879 367166 227185
rect 366890 226821 367070 226824
rect 366838 226815 367070 226821
rect 367126 226873 367178 226879
rect 367126 226815 367178 226821
rect 366742 226799 366794 226805
rect 366850 226796 367070 226815
rect 366742 226741 366794 226747
rect 366754 221482 366782 226741
rect 367426 221792 367454 231847
rect 367618 223739 367646 239672
rect 368098 232133 368126 239672
rect 368194 232429 368222 239686
rect 368578 239089 368606 239686
rect 368566 239083 368618 239089
rect 368566 239025 368618 239031
rect 368962 236467 368990 239686
rect 369312 239672 369566 239700
rect 369696 239672 369950 239700
rect 370080 239672 370334 239700
rect 368948 236458 369004 236467
rect 368948 236393 369004 236402
rect 368182 232423 368234 232429
rect 368182 232365 368234 232371
rect 369538 232281 369566 239672
rect 369526 232275 369578 232281
rect 369526 232217 369578 232223
rect 368086 232127 368138 232133
rect 368086 232069 368138 232075
rect 368660 231870 368716 231879
rect 368660 231805 368716 231814
rect 368182 230499 368234 230505
rect 368182 230441 368234 230447
rect 367604 223730 367660 223739
rect 367604 223665 367660 223674
rect 367426 221764 367502 221792
rect 367474 221482 367502 221764
rect 368194 221482 368222 230441
rect 368674 225219 368702 231805
rect 369922 230431 369950 239672
rect 370306 233909 370334 239672
rect 370402 236763 370430 239686
rect 370486 236863 370538 236869
rect 370486 236805 370538 236811
rect 370388 236754 370444 236763
rect 370388 236689 370444 236698
rect 370294 233903 370346 233909
rect 370294 233845 370346 233851
rect 370390 231979 370442 231985
rect 370390 231921 370442 231927
rect 369910 230425 369962 230431
rect 369910 230367 369962 230373
rect 368854 229463 368906 229469
rect 368854 229405 368906 229411
rect 368660 225210 368716 225219
rect 368660 225145 368716 225154
rect 368866 225029 368894 229405
rect 368950 228057 369002 228063
rect 368950 227999 369002 228005
rect 368854 225023 368906 225029
rect 368854 224965 368906 224971
rect 368962 221482 368990 227999
rect 370402 227534 370430 231921
rect 370498 228063 370526 236805
rect 370582 235087 370634 235093
rect 370582 235029 370634 235035
rect 370594 228063 370622 235029
rect 370786 232915 370814 239686
rect 371170 233063 371198 239686
rect 371616 239672 371870 239700
rect 372000 239672 372254 239700
rect 371842 236055 371870 239672
rect 372226 237059 372254 239672
rect 372212 237050 372268 237059
rect 372212 236985 372268 236994
rect 371830 236049 371882 236055
rect 371830 235991 371882 235997
rect 371638 234199 371690 234205
rect 371638 234141 371690 234147
rect 371156 233054 371212 233063
rect 371156 232989 371212 232998
rect 370772 232906 370828 232915
rect 370772 232841 370828 232850
rect 371254 229315 371306 229321
rect 371254 229257 371306 229263
rect 370486 228057 370538 228063
rect 370486 227999 370538 228005
rect 370582 228057 370634 228063
rect 370582 227999 370634 228005
rect 370402 227506 370526 227534
rect 369622 227169 369674 227175
rect 369622 227111 369674 227117
rect 369634 221792 369662 227111
rect 369634 221764 369710 221792
rect 369682 221482 369710 221764
rect 370498 221482 370526 227506
rect 371266 221482 371294 229257
rect 371542 229241 371594 229247
rect 371542 229183 371594 229189
rect 371554 224881 371582 229183
rect 371542 224875 371594 224881
rect 371542 224817 371594 224823
rect 371650 222365 371678 234141
rect 372322 232059 372350 239686
rect 372706 232207 372734 239686
rect 372694 232201 372746 232207
rect 372694 232143 372746 232149
rect 372310 232053 372362 232059
rect 372310 231995 372362 232001
rect 373090 229807 373118 239686
rect 373474 236911 373502 239686
rect 373824 239672 374078 239700
rect 373460 236902 373516 236911
rect 373460 236837 373516 236846
rect 374050 232767 374078 239672
rect 374194 239404 374222 239686
rect 374422 239601 374474 239607
rect 374422 239543 374474 239549
rect 374194 239376 374270 239404
rect 374036 232758 374092 232767
rect 374036 232693 374092 232702
rect 373462 231831 373514 231837
rect 373462 231773 373514 231779
rect 373076 229798 373132 229807
rect 373076 229733 373132 229742
rect 372694 226725 372746 226731
rect 372694 226667 372746 226673
rect 371926 222433 371978 222439
rect 371926 222375 371978 222381
rect 371638 222359 371690 222365
rect 371638 222301 371690 222307
rect 371938 221792 371966 222375
rect 371938 221764 372014 221792
rect 371986 221482 372014 221764
rect 372706 221482 372734 226667
rect 373474 221482 373502 231773
rect 374134 230647 374186 230653
rect 374134 230589 374186 230595
rect 374146 227534 374174 230589
rect 374242 229321 374270 239376
rect 374434 236129 374462 239543
rect 374422 236123 374474 236129
rect 374422 236065 374474 236071
rect 374530 231985 374558 239686
rect 374914 236319 374942 239686
rect 374900 236310 374956 236319
rect 374900 236245 374956 236254
rect 375394 232619 375422 239686
rect 375380 232610 375436 232619
rect 375380 232545 375436 232554
rect 374518 231979 374570 231985
rect 374518 231921 374570 231927
rect 375778 231911 375806 239686
rect 376128 239672 376382 239700
rect 376512 239672 376766 239700
rect 377302 239691 377354 239697
rect 376354 236129 376382 239672
rect 376342 236123 376394 236129
rect 376342 236065 376394 236071
rect 375766 231905 375818 231911
rect 375766 231847 375818 231853
rect 374614 231461 374666 231467
rect 374614 231403 374666 231409
rect 374230 229315 374282 229321
rect 374230 229257 374282 229263
rect 374422 229167 374474 229173
rect 374422 229109 374474 229115
rect 374146 227506 374270 227534
rect 374242 221792 374270 227506
rect 374326 225985 374378 225991
rect 374326 225927 374378 225933
rect 374338 224807 374366 225927
rect 374434 225843 374462 229109
rect 374518 229093 374570 229099
rect 374518 229035 374570 229041
rect 374422 225837 374474 225843
rect 374422 225779 374474 225785
rect 374530 224807 374558 229035
rect 374626 226731 374654 231403
rect 375766 227539 375818 227545
rect 375766 227481 375818 227487
rect 374614 226725 374666 226731
rect 374614 226667 374666 226673
rect 374326 224801 374378 224807
rect 374326 224743 374378 224749
rect 374518 224801 374570 224807
rect 374518 224743 374570 224749
rect 374998 222507 375050 222513
rect 374998 222449 375050 222455
rect 374242 221764 374318 221792
rect 374290 221482 374318 221764
rect 375010 221482 375038 222449
rect 375778 221482 375806 227481
rect 376438 225023 376490 225029
rect 376438 224965 376490 224971
rect 376450 221792 376478 224965
rect 376738 223443 376766 239672
rect 376834 229099 376862 239686
rect 377110 230573 377162 230579
rect 377110 230515 377162 230521
rect 376822 229093 376874 229099
rect 376822 229035 376874 229041
rect 377122 227534 377150 230515
rect 377218 229173 377246 239686
rect 377314 233317 377342 239691
rect 377302 233311 377354 233317
rect 377302 233253 377354 233259
rect 377206 229167 377258 229173
rect 377206 229109 377258 229115
rect 377122 227506 377246 227534
rect 376724 223434 376780 223443
rect 376724 223369 376780 223378
rect 376450 221764 376526 221792
rect 376498 221482 376526 221764
rect 377218 221482 377246 227506
rect 377602 223591 377630 239686
rect 378000 239672 378206 239700
rect 378336 239672 378590 239700
rect 378720 239672 378974 239700
rect 378178 236425 378206 239672
rect 378166 236419 378218 236425
rect 378166 236361 378218 236367
rect 378562 234205 378590 239672
rect 378550 234199 378602 234205
rect 378550 234141 378602 234147
rect 378946 231837 378974 239672
rect 379138 234543 379166 239686
rect 379522 236615 379550 239686
rect 379508 236606 379564 236615
rect 379508 236541 379564 236550
rect 379124 234534 379180 234543
rect 379124 234469 379180 234478
rect 378934 231831 378986 231837
rect 378934 231773 378986 231779
rect 379906 229659 379934 239686
rect 380256 239672 380510 239700
rect 381024 239672 381278 239700
rect 380084 233350 380140 233359
rect 380482 233317 380510 239672
rect 380084 233285 380140 233294
rect 380470 233311 380522 233317
rect 379990 231387 380042 231393
rect 379990 231329 380042 231335
rect 379892 229650 379948 229659
rect 379892 229585 379948 229594
rect 378742 226651 378794 226657
rect 378742 226593 378794 226599
rect 378070 226429 378122 226435
rect 378070 226371 378122 226377
rect 377588 223582 377644 223591
rect 377588 223517 377644 223526
rect 378082 221482 378110 226371
rect 378646 225023 378698 225029
rect 378646 224965 378698 224971
rect 378658 224733 378686 224965
rect 378646 224727 378698 224733
rect 378646 224669 378698 224675
rect 378754 221792 378782 226593
rect 380002 226065 380030 231329
rect 380098 229469 380126 233285
rect 380470 233253 380522 233259
rect 380278 230869 380330 230875
rect 380278 230811 380330 230817
rect 380086 229463 380138 229469
rect 380086 229405 380138 229411
rect 380086 228649 380138 228655
rect 380086 228591 380138 228597
rect 379990 226059 380042 226065
rect 379990 226001 380042 226007
rect 380098 224881 380126 228591
rect 379510 224875 379562 224881
rect 379510 224817 379562 224823
rect 380086 224875 380138 224881
rect 380086 224817 380138 224823
rect 378754 221764 378830 221792
rect 378802 221482 378830 221764
rect 379522 221482 379550 224817
rect 380290 221482 380318 230811
rect 381250 223295 381278 239672
rect 381346 229511 381374 239686
rect 381730 232471 381758 239686
rect 382114 234395 382142 239686
rect 382560 239672 382622 239700
rect 382390 236789 382442 236795
rect 382390 236731 382442 236737
rect 382402 236615 382430 236731
rect 382594 236615 382622 239672
rect 382690 239672 382944 239700
rect 383328 239672 383582 239700
rect 382388 236606 382444 236615
rect 382388 236541 382444 236550
rect 382580 236606 382636 236615
rect 382580 236541 382636 236550
rect 382100 234386 382156 234395
rect 382100 234321 382156 234330
rect 381716 232462 381772 232471
rect 381716 232397 381772 232406
rect 382690 232175 382718 239672
rect 382966 233311 383018 233317
rect 382966 233253 383018 233259
rect 382774 232941 382826 232947
rect 382774 232883 382826 232889
rect 382676 232166 382732 232175
rect 382676 232101 382732 232110
rect 381332 229502 381388 229511
rect 381332 229437 381388 229446
rect 381814 227465 381866 227471
rect 381814 227407 381866 227413
rect 381236 223286 381292 223295
rect 381236 223221 381292 223230
rect 381046 222729 381098 222735
rect 381046 222671 381098 222677
rect 381058 221496 381086 222671
rect 381058 221468 381120 221496
rect 381826 221482 381854 227407
rect 382678 226429 382730 226435
rect 382678 226371 382730 226377
rect 382690 225917 382718 226371
rect 382678 225911 382730 225917
rect 382678 225853 382730 225859
rect 382582 224801 382634 224807
rect 382582 224743 382634 224749
rect 382594 221496 382622 224743
rect 382786 224733 382814 232883
rect 382978 229025 383006 233253
rect 383554 229363 383582 239672
rect 383650 233687 383678 239686
rect 384048 239672 384350 239700
rect 383638 233681 383690 233687
rect 383638 233623 383690 233629
rect 383540 229354 383596 229363
rect 383540 229289 383596 229298
rect 382870 229019 382922 229025
rect 382870 228961 382922 228967
rect 382966 229019 383018 229025
rect 382966 228961 383018 228967
rect 382882 225917 382910 228961
rect 382966 228427 383018 228433
rect 382966 228369 383018 228375
rect 382978 226657 383006 228369
rect 383254 228279 383306 228285
rect 383254 228221 383306 228227
rect 382966 226651 383018 226657
rect 382966 226593 383018 226599
rect 382870 225911 382922 225917
rect 382870 225853 382922 225859
rect 382774 224727 382826 224733
rect 382774 224669 382826 224675
rect 382560 221468 382622 221496
rect 383266 221496 383294 228221
rect 384022 227391 384074 227397
rect 384022 227333 384074 227339
rect 383266 221468 383328 221496
rect 384034 221482 384062 227333
rect 384322 223147 384350 239672
rect 384418 229215 384446 239686
rect 384768 239672 385022 239700
rect 385152 239672 385310 239700
rect 384994 232323 385022 239672
rect 384980 232314 385036 232323
rect 384980 232249 385036 232258
rect 385282 232027 385310 239672
rect 385366 239675 385418 239681
rect 385536 239672 385790 239700
rect 385366 239617 385418 239623
rect 385378 235167 385406 239617
rect 385366 235161 385418 235167
rect 385366 235103 385418 235109
rect 385268 232018 385324 232027
rect 385268 231953 385324 231962
rect 384404 229206 384460 229215
rect 384404 229141 384460 229150
rect 385762 226509 385790 239672
rect 385858 236023 385886 239686
rect 386352 239672 386654 239700
rect 385844 236014 385900 236023
rect 385844 235949 385900 235958
rect 386134 233755 386186 233761
rect 386134 233697 386186 233703
rect 385846 231313 385898 231319
rect 385846 231255 385898 231261
rect 384790 226503 384842 226509
rect 384790 226445 384842 226451
rect 385750 226503 385802 226509
rect 385750 226445 385802 226451
rect 384308 223138 384364 223147
rect 384308 223073 384364 223082
rect 384802 221792 384830 226445
rect 385558 225837 385610 225843
rect 385558 225779 385610 225785
rect 384802 221764 384878 221792
rect 384850 221482 384878 221764
rect 385570 221482 385598 225779
rect 385858 224807 385886 231255
rect 385846 224801 385898 224807
rect 385846 224743 385898 224749
rect 386146 222439 386174 233697
rect 386626 226805 386654 239672
rect 386722 235981 386750 239686
rect 387072 239672 387326 239700
rect 387456 239672 387710 239700
rect 386996 237050 387052 237059
rect 386996 236985 387052 236994
rect 387010 236869 387038 236985
rect 386998 236863 387050 236869
rect 386998 236805 387050 236811
rect 387092 236606 387148 236615
rect 387092 236541 387148 236550
rect 387190 236567 387242 236573
rect 387106 236351 387134 236541
rect 387190 236509 387242 236515
rect 387202 236467 387230 236509
rect 387188 236458 387244 236467
rect 387188 236393 387244 236402
rect 387094 236345 387146 236351
rect 387094 236287 387146 236293
rect 387298 236174 387326 239672
rect 387476 237050 387532 237059
rect 387476 236985 387532 236994
rect 387490 236467 387518 236985
rect 387574 236863 387626 236869
rect 387574 236805 387626 236811
rect 387586 236763 387614 236805
rect 387572 236754 387628 236763
rect 387572 236689 387628 236698
rect 387476 236458 387532 236467
rect 387476 236393 387532 236402
rect 387478 236345 387530 236351
rect 387476 236310 387478 236319
rect 387530 236310 387532 236319
rect 387476 236245 387532 236254
rect 387298 236146 387422 236174
rect 386710 235975 386762 235981
rect 386710 235917 386762 235923
rect 387286 234791 387338 234797
rect 387286 234733 387338 234739
rect 387298 230875 387326 234733
rect 387286 230869 387338 230875
rect 387286 230811 387338 230817
rect 387286 230425 387338 230431
rect 387286 230367 387338 230373
rect 387298 229321 387326 230367
rect 387286 229315 387338 229321
rect 387286 229257 387338 229263
rect 386614 226799 386666 226805
rect 386614 226741 386666 226747
rect 386998 226429 387050 226435
rect 386998 226371 387050 226377
rect 386422 225911 386474 225917
rect 386422 225853 386474 225859
rect 386434 224733 386462 225853
rect 386326 224727 386378 224733
rect 386326 224669 386378 224675
rect 386422 224727 386474 224733
rect 386422 224669 386474 224675
rect 386134 222433 386186 222439
rect 386134 222375 386186 222381
rect 386338 221482 386366 224669
rect 387010 221792 387038 226371
rect 387394 225917 387422 236146
rect 387682 235167 387710 239672
rect 387670 235161 387722 235167
rect 387670 235103 387722 235109
rect 387778 227619 387806 239686
rect 387860 237050 387916 237059
rect 387860 236985 387916 236994
rect 387874 236573 387902 236985
rect 387862 236567 387914 236573
rect 387862 236509 387914 236515
rect 387766 227613 387818 227619
rect 387766 227555 387818 227561
rect 388162 225991 388190 239686
rect 388546 227471 388574 239686
rect 388930 227545 388958 239686
rect 389280 239672 389534 239700
rect 389664 239672 389918 239700
rect 388918 227539 388970 227545
rect 388918 227481 388970 227487
rect 388534 227465 388586 227471
rect 388534 227407 388586 227413
rect 388726 226799 388778 226805
rect 388726 226741 388778 226747
rect 387766 225985 387818 225991
rect 387766 225927 387818 225933
rect 388150 225985 388202 225991
rect 388150 225927 388202 225933
rect 388738 225936 388766 226741
rect 387382 225911 387434 225917
rect 387382 225853 387434 225859
rect 387010 221764 387086 221792
rect 387058 221482 387086 221764
rect 387778 221482 387806 225927
rect 388738 225908 388862 225936
rect 388834 225843 388862 225908
rect 388822 225837 388874 225843
rect 388822 225779 388874 225785
rect 388630 224875 388682 224881
rect 388630 224817 388682 224823
rect 388642 221482 388670 224817
rect 389506 224733 389534 239672
rect 389890 235875 389918 239672
rect 389876 235866 389932 235875
rect 389876 235801 389932 235810
rect 390082 227323 390110 239686
rect 390466 227397 390494 239686
rect 390742 236345 390794 236351
rect 390742 236287 390794 236293
rect 390754 235727 390782 236287
rect 390740 235718 390796 235727
rect 390740 235653 390796 235662
rect 390454 227391 390506 227397
rect 390454 227333 390506 227339
rect 390070 227317 390122 227323
rect 390070 227259 390122 227265
rect 390850 227249 390878 239686
rect 390838 227243 390890 227249
rect 390838 227185 390890 227191
rect 391234 226847 391262 239686
rect 391584 239672 391646 239700
rect 391968 239672 392222 239700
rect 391618 226995 391646 239672
rect 391702 235309 391754 235315
rect 391702 235251 391754 235257
rect 391714 228433 391742 235251
rect 392194 235241 392222 239672
rect 392182 235235 392234 235241
rect 392182 235177 392234 235183
rect 391702 228427 391754 228433
rect 391702 228369 391754 228375
rect 391604 226986 391660 226995
rect 391604 226921 391660 226930
rect 391220 226838 391276 226847
rect 391220 226773 391276 226782
rect 391510 226725 391562 226731
rect 391510 226667 391562 226673
rect 390070 226577 390122 226583
rect 390070 226519 390122 226525
rect 389302 224727 389354 224733
rect 389302 224669 389354 224675
rect 389494 224727 389546 224733
rect 389494 224669 389546 224675
rect 389314 221792 389342 224669
rect 389314 221764 389390 221792
rect 389362 221482 389390 221764
rect 390082 221482 390110 226519
rect 390838 226355 390890 226361
rect 390838 226297 390890 226303
rect 390850 221482 390878 226297
rect 391522 221792 391550 226667
rect 392290 224807 392318 239686
rect 392470 234865 392522 234871
rect 392470 234807 392522 234813
rect 392482 228359 392510 234807
rect 392374 228353 392426 228359
rect 392374 228295 392426 228301
rect 392470 228353 392522 228359
rect 392470 228295 392522 228301
rect 392278 224801 392330 224807
rect 392278 224743 392330 224749
rect 391522 221764 391598 221792
rect 391570 221482 391598 221764
rect 392386 221482 392414 228295
rect 392674 227175 392702 239686
rect 393058 235727 393086 239686
rect 393044 235718 393100 235727
rect 393044 235653 393100 235662
rect 393442 235389 393470 239686
rect 393888 239672 394142 239700
rect 394272 239672 394526 239700
rect 394608 239672 394910 239700
rect 393430 235383 393482 235389
rect 393430 235325 393482 235331
rect 392662 227169 392714 227175
rect 392662 227111 392714 227117
rect 393142 227095 393194 227101
rect 393142 227037 393194 227043
rect 393154 221482 393182 227037
rect 393814 227021 393866 227027
rect 393814 226963 393866 226969
rect 393826 221792 393854 226963
rect 394114 226699 394142 239672
rect 394100 226690 394156 226699
rect 394100 226625 394156 226634
rect 394498 226551 394526 239672
rect 394678 239453 394730 239459
rect 394678 239395 394730 239401
rect 394582 236271 394634 236277
rect 394582 236213 394634 236219
rect 394594 233613 394622 236213
rect 394690 235019 394718 239395
rect 394882 235093 394910 239672
rect 394978 235537 395006 239686
rect 395376 239672 395582 239700
rect 395712 239672 395966 239700
rect 396096 239672 396350 239700
rect 396480 239672 396734 239700
rect 394966 235531 395018 235537
rect 394966 235473 395018 235479
rect 395062 235457 395114 235463
rect 395062 235399 395114 235405
rect 394870 235087 394922 235093
rect 394870 235029 394922 235035
rect 394678 235013 394730 235019
rect 394678 234955 394730 234961
rect 394774 234939 394826 234945
rect 394774 234881 394826 234887
rect 394678 234717 394730 234723
rect 394678 234659 394730 234665
rect 394582 233607 394634 233613
rect 394582 233549 394634 233555
rect 394690 228285 394718 234659
rect 394786 231245 394814 234881
rect 394870 234051 394922 234057
rect 394870 233993 394922 233999
rect 394774 231239 394826 231245
rect 394774 231181 394826 231187
rect 394678 228279 394730 228285
rect 394678 228221 394730 228227
rect 394484 226542 394540 226551
rect 394484 226477 394540 226486
rect 394774 226503 394826 226509
rect 394774 226445 394826 226451
rect 394582 226059 394634 226065
rect 394582 226001 394634 226007
rect 394678 226059 394730 226065
rect 394678 226001 394730 226007
rect 393826 221764 393902 221792
rect 393874 221482 393902 221764
rect 394594 221482 394622 226001
rect 394690 225917 394718 226001
rect 394786 225917 394814 226445
rect 394678 225911 394730 225917
rect 394678 225853 394730 225859
rect 394774 225911 394826 225917
rect 394774 225853 394826 225859
rect 394882 222513 394910 233993
rect 395074 231319 395102 235399
rect 395062 231313 395114 231319
rect 395062 231255 395114 231261
rect 395350 230943 395402 230949
rect 395350 230885 395402 230891
rect 394870 222507 394922 222513
rect 394870 222449 394922 222455
rect 395362 221482 395390 230885
rect 395554 226805 395582 239672
rect 395938 233317 395966 239672
rect 396322 235315 396350 239672
rect 396310 235309 396362 235315
rect 396310 235251 396362 235257
rect 396706 234057 396734 239672
rect 396802 235463 396830 239686
rect 397078 236715 397130 236721
rect 397078 236657 397130 236663
rect 397090 236319 397118 236657
rect 397076 236310 397132 236319
rect 397076 236245 397132 236254
rect 396790 235457 396842 235463
rect 396790 235399 396842 235405
rect 396694 234051 396746 234057
rect 396694 233993 396746 233999
rect 395926 233311 395978 233317
rect 395926 233253 395978 233259
rect 396406 227613 396458 227619
rect 396406 227555 396458 227561
rect 396418 227323 396446 227555
rect 396406 227317 396458 227323
rect 396406 227259 396458 227265
rect 396118 226873 396170 226879
rect 396118 226815 396170 226821
rect 395542 226799 395594 226805
rect 395542 226741 395594 226747
rect 396130 221792 396158 226815
rect 397186 226731 397214 239686
rect 397460 236754 397516 236763
rect 397460 236689 397516 236698
rect 397474 236647 397502 236689
rect 397462 236641 397514 236647
rect 397462 236583 397514 236589
rect 397462 236493 397514 236499
rect 397462 236435 397514 236441
rect 397366 236419 397418 236425
rect 397366 236361 397418 236367
rect 397378 236319 397406 236361
rect 397364 236310 397420 236319
rect 397364 236245 397420 236254
rect 397474 235579 397502 236435
rect 397460 235570 397516 235579
rect 397460 235505 397516 235514
rect 397366 232719 397418 232725
rect 397366 232661 397418 232667
rect 397378 232596 397406 232661
rect 397378 232568 397502 232596
rect 397474 226805 397502 232568
rect 397666 227101 397694 239686
rect 398016 239672 398270 239700
rect 398400 239672 398654 239700
rect 398784 239672 399038 239700
rect 399120 239672 399422 239700
rect 397942 239379 397994 239385
rect 397942 239321 397994 239327
rect 397748 237050 397804 237059
rect 397748 236985 397804 236994
rect 397762 236721 397790 236985
rect 397844 236902 397900 236911
rect 397844 236837 397846 236846
rect 397898 236837 397900 236846
rect 397846 236805 397898 236811
rect 397750 236715 397802 236721
rect 397750 236657 397802 236663
rect 397954 236499 397982 239321
rect 398036 236902 398092 236911
rect 398036 236837 398092 236846
rect 398050 236795 398078 236837
rect 398038 236789 398090 236795
rect 398038 236731 398090 236737
rect 397942 236493 397994 236499
rect 397942 236435 397994 236441
rect 398242 234279 398270 239672
rect 398626 234945 398654 239672
rect 399010 235019 399038 239672
rect 398998 235013 399050 235019
rect 398998 234955 399050 234961
rect 398614 234939 398666 234945
rect 398614 234881 398666 234887
rect 398134 234273 398186 234279
rect 398134 234215 398186 234221
rect 398230 234273 398282 234279
rect 398230 234215 398282 234221
rect 398146 233761 398174 234215
rect 399190 234199 399242 234205
rect 399190 234141 399242 234147
rect 398134 233755 398186 233761
rect 398134 233697 398186 233703
rect 399202 232725 399230 234141
rect 399190 232719 399242 232725
rect 399190 232661 399242 232667
rect 398326 228131 398378 228137
rect 398326 228073 398378 228079
rect 397654 227095 397706 227101
rect 397654 227037 397706 227043
rect 397462 226799 397514 226805
rect 397462 226741 397514 226747
rect 397174 226725 397226 226731
rect 397174 226667 397226 226673
rect 397654 226651 397706 226657
rect 397654 226593 397706 226599
rect 396886 225763 396938 225769
rect 396886 225705 396938 225711
rect 396130 221764 396206 221792
rect 396178 221482 396206 221764
rect 396898 221482 396926 225705
rect 397666 221482 397694 226593
rect 398338 221792 398366 228073
rect 399394 225103 399422 239672
rect 399490 228919 399518 239686
rect 399874 235579 399902 239686
rect 400224 239672 400286 239700
rect 400608 239672 400862 239700
rect 400992 239672 401246 239700
rect 399860 235570 399916 235579
rect 399860 235505 399916 235514
rect 400150 234125 400202 234131
rect 400150 234067 400202 234073
rect 400162 231393 400190 234067
rect 400258 233951 400286 239672
rect 400342 236197 400394 236203
rect 400342 236139 400394 236145
rect 400354 235685 400382 236139
rect 400342 235679 400394 235685
rect 400342 235621 400394 235627
rect 400244 233942 400300 233951
rect 400244 233877 400300 233886
rect 400246 233311 400298 233317
rect 400246 233253 400298 233259
rect 400150 231387 400202 231393
rect 400150 231329 400202 231335
rect 400258 229067 400286 233253
rect 400244 229058 400300 229067
rect 400244 228993 400300 229002
rect 399476 228910 399532 228919
rect 399476 228845 399532 228854
rect 400630 226799 400682 226805
rect 400630 226741 400682 226747
rect 399958 225171 400010 225177
rect 399958 225113 400010 225119
rect 399094 225097 399146 225103
rect 399094 225039 399146 225045
rect 399382 225097 399434 225103
rect 399382 225039 399434 225045
rect 398338 221764 398414 221792
rect 398386 221482 398414 221764
rect 399106 221482 399134 225039
rect 399970 221482 399998 225113
rect 400642 221792 400670 226741
rect 400834 226657 400862 239672
rect 401218 233317 401246 239672
rect 401410 235431 401438 239686
rect 401396 235422 401452 235431
rect 401396 235357 401452 235366
rect 401794 234131 401822 239686
rect 402192 239672 402398 239700
rect 402528 239672 402686 239700
rect 401782 234125 401834 234131
rect 401782 234067 401834 234073
rect 401206 233311 401258 233317
rect 401206 233253 401258 233259
rect 401398 231017 401450 231023
rect 401398 230959 401450 230965
rect 400822 226651 400874 226657
rect 400822 226593 400874 226599
rect 400642 221764 400718 221792
rect 400690 221482 400718 221764
rect 401410 221482 401438 230959
rect 402370 226583 402398 239672
rect 402358 226577 402410 226583
rect 402358 226519 402410 226525
rect 402658 226509 402686 239672
rect 402754 239672 402912 239700
rect 403248 239672 403550 239700
rect 402754 235283 402782 239672
rect 402740 235274 402796 235283
rect 402740 235209 402796 235218
rect 403124 234978 403180 234987
rect 403124 234913 403180 234922
rect 403030 233755 403082 233761
rect 403030 233697 403082 233703
rect 402646 226503 402698 226509
rect 402646 226445 402698 226451
rect 402838 226281 402890 226287
rect 402838 226223 402890 226229
rect 402166 224949 402218 224955
rect 402166 224891 402218 224897
rect 402178 221482 402206 224891
rect 402850 221792 402878 226223
rect 403042 222735 403070 233697
rect 403138 231467 403166 234913
rect 403522 234205 403550 239672
rect 403618 234871 403646 239686
rect 404002 234987 404030 239686
rect 403988 234978 404044 234987
rect 403988 234913 404044 234922
rect 403606 234865 403658 234871
rect 403606 234807 403658 234813
rect 403510 234199 403562 234205
rect 403510 234141 403562 234147
rect 403126 231461 403178 231467
rect 403126 231403 403178 231409
rect 403702 228501 403754 228507
rect 403702 228443 403754 228449
rect 403030 222729 403082 222735
rect 403030 222671 403082 222677
rect 402850 221764 402926 221792
rect 402898 221482 402926 221764
rect 403714 221482 403742 228443
rect 404386 226403 404414 239686
rect 404736 239672 404990 239700
rect 405216 239672 405470 239700
rect 404470 236937 404522 236943
rect 404470 236879 404522 236885
rect 404372 226394 404428 226403
rect 404372 226329 404428 226338
rect 404482 221482 404510 236879
rect 404962 226435 404990 239672
rect 405442 235135 405470 239672
rect 405428 235126 405484 235135
rect 405428 235061 405484 235070
rect 405538 234839 405566 239686
rect 405826 239672 405936 239700
rect 405622 235975 405674 235981
rect 405622 235917 405674 235923
rect 405634 235611 405662 235917
rect 405622 235605 405674 235611
rect 405622 235547 405674 235553
rect 405332 234830 405388 234839
rect 405332 234765 405388 234774
rect 405524 234830 405580 234839
rect 405524 234765 405580 234774
rect 405346 228507 405374 234765
rect 405716 234682 405772 234691
rect 405716 234617 405772 234626
rect 405334 228501 405386 228507
rect 405334 228443 405386 228449
rect 404950 226429 405002 226435
rect 404950 226371 405002 226377
rect 405730 226084 405758 234617
rect 405826 226255 405854 239672
rect 406006 239305 406058 239311
rect 406006 239247 406058 239253
rect 405910 236937 405962 236943
rect 405910 236879 405962 236885
rect 405922 233803 405950 236879
rect 406018 236055 406046 239247
rect 406306 236055 406334 239686
rect 406484 236162 406540 236171
rect 406484 236097 406540 236106
rect 406006 236049 406058 236055
rect 406006 235991 406058 235997
rect 406294 236049 406346 236055
rect 406294 235991 406346 235997
rect 406006 234273 406058 234279
rect 406006 234215 406058 234221
rect 405908 233794 405964 233803
rect 405908 233729 405964 233738
rect 406018 231879 406046 234215
rect 406004 231870 406060 231879
rect 406004 231805 406060 231814
rect 405812 226246 405868 226255
rect 405812 226181 405868 226190
rect 405730 226056 405950 226084
rect 405142 225023 405194 225029
rect 405142 224965 405194 224971
rect 405154 221792 405182 224965
rect 405154 221764 405230 221792
rect 405202 221482 405230 221764
rect 405922 221482 405950 226056
rect 406498 222555 406526 236097
rect 406690 234797 406718 239686
rect 407040 239672 407294 239700
rect 407424 239672 407678 239700
rect 406678 234791 406730 234797
rect 406678 234733 406730 234739
rect 407266 234279 407294 239672
rect 407444 236754 407500 236763
rect 407444 236689 407500 236698
rect 407458 236319 407486 236689
rect 407444 236310 407500 236319
rect 407444 236245 407500 236254
rect 407446 234421 407498 234427
rect 407446 234363 407498 234369
rect 407254 234273 407306 234279
rect 407254 234215 407306 234221
rect 407458 233835 407486 234363
rect 407350 233829 407402 233835
rect 407350 233771 407402 233777
rect 407446 233829 407498 233835
rect 407446 233771 407498 233777
rect 406774 229685 406826 229691
rect 406774 229627 406826 229633
rect 406484 222546 406540 222555
rect 406484 222481 406540 222490
rect 406786 221482 406814 229627
rect 407362 228655 407390 233771
rect 407350 228649 407402 228655
rect 407350 228591 407402 228597
rect 407446 227317 407498 227323
rect 407446 227259 407498 227265
rect 407458 227101 407486 227259
rect 407350 227095 407402 227101
rect 407350 227037 407402 227043
rect 407446 227095 407498 227101
rect 407446 227037 407498 227043
rect 407362 226805 407390 227037
rect 407350 226799 407402 226805
rect 407350 226741 407402 226747
rect 407650 226107 407678 239672
rect 407746 226361 407774 239686
rect 408130 234723 408158 239686
rect 408118 234717 408170 234723
rect 408514 234691 408542 239686
rect 408960 239672 409214 239700
rect 409728 239672 409982 239700
rect 409186 235685 409214 239672
rect 409954 236171 409982 239672
rect 409940 236162 409996 236171
rect 410050 236129 410078 239686
rect 409940 236097 409996 236106
rect 410038 236123 410090 236129
rect 410038 236065 410090 236071
rect 408982 235679 409034 235685
rect 408982 235621 409034 235627
rect 409174 235679 409226 235685
rect 409174 235621 409226 235627
rect 408118 234659 408170 234665
rect 408500 234682 408556 234691
rect 408500 234617 408556 234626
rect 408994 233761 409022 235621
rect 409844 234534 409900 234543
rect 409844 234469 409900 234478
rect 408982 233755 409034 233761
rect 408982 233697 409034 233703
rect 408118 233681 408170 233687
rect 408118 233623 408170 233629
rect 408130 230399 408158 233623
rect 408886 233311 408938 233317
rect 408886 233253 408938 233259
rect 408116 230390 408172 230399
rect 408116 230325 408172 230334
rect 408214 226947 408266 226953
rect 408214 226889 408266 226895
rect 407734 226355 407786 226361
rect 407734 226297 407786 226303
rect 407636 226098 407692 226107
rect 407636 226033 407692 226042
rect 407446 224875 407498 224881
rect 407446 224817 407498 224823
rect 407458 221792 407486 224817
rect 407458 221764 407534 221792
rect 407506 221482 407534 221764
rect 408226 221482 408254 226889
rect 408898 225769 408926 233253
rect 409654 230721 409706 230727
rect 409654 230663 409706 230669
rect 408982 226133 409034 226139
rect 408982 226075 409034 226081
rect 408886 225763 408938 225769
rect 408886 225705 408938 225711
rect 408994 221482 409022 226075
rect 409666 221792 409694 230663
rect 409858 229691 409886 234469
rect 410036 234386 410092 234395
rect 410036 234321 410092 234330
rect 410050 232947 410078 234321
rect 410038 232941 410090 232947
rect 410038 232883 410090 232889
rect 409846 229685 409898 229691
rect 409846 229627 409898 229633
rect 410434 226287 410462 239686
rect 410710 236419 410762 236425
rect 410710 236361 410762 236367
rect 410722 235759 410750 236361
rect 410710 235753 410762 235759
rect 410710 235695 410762 235701
rect 410818 234395 410846 239686
rect 411168 239672 411422 239700
rect 411552 239672 411710 239700
rect 411936 239672 412190 239700
rect 411394 234543 411422 239672
rect 411380 234534 411436 234543
rect 411380 234469 411436 234478
rect 410804 234386 410860 234395
rect 410804 234321 410860 234330
rect 410614 233755 410666 233761
rect 410614 233697 410666 233703
rect 410422 226281 410474 226287
rect 410422 226223 410474 226229
rect 410626 222587 410654 233697
rect 411286 226207 411338 226213
rect 411286 226149 411338 226155
rect 410518 222581 410570 222587
rect 410518 222523 410570 222529
rect 410614 222581 410666 222587
rect 410614 222523 410666 222529
rect 409666 221764 409742 221792
rect 409714 221482 409742 221764
rect 410530 221482 410558 222523
rect 411298 221496 411326 226149
rect 411682 226139 411710 239672
rect 411862 235753 411914 235759
rect 411862 235695 411914 235701
rect 411874 235611 411902 235695
rect 412162 235611 412190 239672
rect 420418 239237 420446 241129
rect 569012 240010 569068 240019
rect 569012 239945 569068 239954
rect 434614 239823 434666 239829
rect 434614 239765 434666 239771
rect 420406 239231 420458 239237
rect 420406 239173 420458 239179
rect 413396 238974 413452 238983
rect 413396 238909 413452 238918
rect 413410 236647 413438 238909
rect 414068 238826 414124 238835
rect 414068 238761 414124 238770
rect 413684 238678 413740 238687
rect 413602 238636 413684 238664
rect 413602 236869 413630 238636
rect 413684 238613 413740 238622
rect 413972 238382 414028 238391
rect 413698 238340 413972 238368
rect 413590 236863 413642 236869
rect 413590 236805 413642 236811
rect 413398 236641 413450 236647
rect 413398 236583 413450 236589
rect 413698 236319 413726 238340
rect 413972 238317 414028 238326
rect 414082 237480 414110 238761
rect 415220 238234 415276 238243
rect 415220 238169 415276 238178
rect 414452 238086 414508 238095
rect 414452 238021 414508 238030
rect 413794 237452 414110 237480
rect 413684 236310 413740 236319
rect 413684 236245 413740 236254
rect 413794 236148 413822 237452
rect 414466 236943 414494 238021
rect 414454 236937 414506 236943
rect 414454 236879 414506 236885
rect 415234 236319 415262 238169
rect 432406 237233 432458 237239
rect 432406 237175 432458 237181
rect 426358 237159 426410 237165
rect 426358 237101 426410 237107
rect 420310 237011 420362 237017
rect 420310 236953 420362 236959
rect 415220 236310 415276 236319
rect 415220 236245 415276 236254
rect 415412 236310 415468 236319
rect 415412 236245 415468 236254
rect 413698 236120 413822 236148
rect 413876 236162 413932 236171
rect 413698 235759 413726 236120
rect 413876 236097 413932 236106
rect 413890 235981 413918 236097
rect 415426 236055 415454 236245
rect 415414 236049 415466 236055
rect 415414 235991 415466 235997
rect 413878 235975 413930 235981
rect 413878 235917 413930 235923
rect 413686 235753 413738 235759
rect 413686 235695 413738 235701
rect 411862 235605 411914 235611
rect 411862 235547 411914 235553
rect 412150 235605 412202 235611
rect 412150 235547 412202 235553
rect 414742 234347 414794 234353
rect 414742 234289 414794 234295
rect 414754 231171 414782 234289
rect 414742 231165 414794 231171
rect 414742 231107 414794 231113
rect 415702 231017 415754 231023
rect 415702 230959 415754 230965
rect 413494 228575 413546 228581
rect 413494 228517 413546 228523
rect 412726 228205 412778 228211
rect 412726 228147 412778 228153
rect 411670 226133 411722 226139
rect 411670 226075 411722 226081
rect 411958 225319 412010 225325
rect 411958 225261 412010 225267
rect 411264 221468 411326 221496
rect 411970 221496 411998 225261
rect 411970 221468 412032 221496
rect 412738 221482 412766 228147
rect 413506 221496 413534 228517
rect 415030 225393 415082 225399
rect 415030 225335 415082 225341
rect 414262 222655 414314 222661
rect 414262 222597 414314 222603
rect 413472 221468 413534 221496
rect 414274 221482 414302 222597
rect 415042 221482 415070 225335
rect 415714 221792 415742 230959
rect 419542 230943 419594 230949
rect 419542 230885 419594 230891
rect 416470 230795 416522 230801
rect 416470 230737 416522 230743
rect 415714 221764 415790 221792
rect 415762 221482 415790 221764
rect 416482 221482 416510 230737
rect 418774 228797 418826 228803
rect 418774 228739 418826 228745
rect 418006 225245 418058 225251
rect 418006 225187 418058 225193
rect 417238 222877 417290 222883
rect 417238 222819 417290 222825
rect 417250 221482 417278 222819
rect 418018 221792 418046 225187
rect 418018 221764 418094 221792
rect 418066 221482 418094 221764
rect 418786 221482 418814 228739
rect 419554 221482 419582 230885
rect 420322 221792 420350 236953
rect 426166 234495 426218 234501
rect 426166 234437 426218 234443
rect 423286 233829 423338 233835
rect 423286 233771 423338 233777
rect 421846 228723 421898 228729
rect 421846 228665 421898 228671
rect 420982 225467 421034 225473
rect 420982 225409 421034 225415
rect 420274 221764 420350 221792
rect 420274 221482 420302 221764
rect 420994 221482 421022 225409
rect 421858 221482 421886 228665
rect 423298 227619 423326 233771
rect 424054 231165 424106 231171
rect 424054 231107 424106 231113
rect 424724 231130 424780 231139
rect 423286 227613 423338 227619
rect 423286 227555 423338 227561
rect 423286 222951 423338 222957
rect 423286 222893 423338 222899
rect 422518 222803 422570 222809
rect 422518 222745 422570 222751
rect 422530 221792 422558 222745
rect 422530 221764 422606 221792
rect 422578 221482 422606 221764
rect 423298 221482 423326 222893
rect 424066 221482 424094 231107
rect 424724 231065 424780 231074
rect 424738 221792 424766 231065
rect 426178 230505 426206 234437
rect 426166 230499 426218 230505
rect 426166 230441 426218 230447
rect 425590 228057 425642 228063
rect 425590 227999 425642 228005
rect 424738 221764 424814 221792
rect 424786 221482 424814 221764
rect 425602 221482 425630 227999
rect 426370 221482 426398 237101
rect 428662 237085 428714 237091
rect 428662 237027 428714 237033
rect 427894 233903 427946 233909
rect 427894 233845 427946 233851
rect 427906 228951 427934 233845
rect 427798 228945 427850 228951
rect 427798 228887 427850 228893
rect 427894 228945 427946 228951
rect 427894 228887 427946 228893
rect 427030 225541 427082 225547
rect 427030 225483 427082 225489
rect 427042 221792 427070 225483
rect 427042 221764 427118 221792
rect 427090 221482 427118 221764
rect 427810 221482 427838 228887
rect 428674 221482 428702 237027
rect 432022 233977 432074 233983
rect 432022 233919 432074 233925
rect 432034 228877 432062 233919
rect 430870 228871 430922 228877
rect 430870 228813 430922 228819
rect 432022 228871 432074 228877
rect 432022 228813 432074 228819
rect 429334 223099 429386 223105
rect 429334 223041 429386 223047
rect 429346 221792 429374 223041
rect 430102 222581 430154 222587
rect 430102 222523 430154 222529
rect 429346 221764 429422 221792
rect 429394 221482 429422 221764
rect 430114 221482 430142 222523
rect 430882 221482 430910 228813
rect 431542 223025 431594 223031
rect 431542 222967 431594 222973
rect 431554 221792 431582 222967
rect 431554 221764 431630 221792
rect 431602 221482 431630 221764
rect 432418 221482 432446 237175
rect 433846 231535 433898 231541
rect 433846 231477 433898 231483
rect 433174 227613 433226 227619
rect 433174 227555 433226 227561
rect 433186 221482 433214 227555
rect 433858 221792 433886 231477
rect 433858 221764 433934 221792
rect 433906 221482 433934 221764
rect 434626 221482 434654 239765
rect 446710 239749 446762 239755
rect 446710 239691 446762 239697
rect 444502 237455 444554 237461
rect 444502 237397 444554 237403
rect 440662 237381 440714 237387
rect 440662 237323 440714 237329
rect 438358 237307 438410 237313
rect 438358 237249 438410 237255
rect 434902 234569 434954 234575
rect 434902 234511 434954 234517
rect 434914 230431 434942 234511
rect 436150 230499 436202 230505
rect 436150 230441 436202 230447
rect 434902 230425 434954 230431
rect 434902 230367 434954 230373
rect 435382 223173 435434 223179
rect 435382 223115 435434 223121
rect 435394 221482 435422 223115
rect 436162 221792 436190 230441
rect 436918 230203 436970 230209
rect 436918 230145 436970 230151
rect 436162 221764 436238 221792
rect 436210 221482 436238 221764
rect 436930 221482 436958 230145
rect 437686 228279 437738 228285
rect 437686 228221 437738 228227
rect 437698 221482 437726 228221
rect 438370 221792 438398 237249
rect 439990 230351 440042 230357
rect 439990 230293 440042 230299
rect 439126 225615 439178 225621
rect 439126 225557 439178 225563
rect 438370 221764 438446 221792
rect 438418 221482 438446 221764
rect 439138 221482 439166 225557
rect 440002 221496 440030 230293
rect 439968 221468 440030 221496
rect 440674 221496 440702 237323
rect 442198 236419 442250 236425
rect 442198 236361 442250 236367
rect 441430 224653 441482 224659
rect 441430 224595 441482 224601
rect 440674 221468 440736 221496
rect 441442 221482 441470 224595
rect 442210 221496 442238 236361
rect 442868 231278 442924 231287
rect 442868 231213 442924 231222
rect 442176 221468 442238 221496
rect 442882 221496 442910 231213
rect 443734 222359 443786 222365
rect 443734 222301 443786 222307
rect 442882 221468 442944 221496
rect 443746 221482 443774 222301
rect 444514 221792 444542 237397
rect 445942 230277 445994 230283
rect 445942 230219 445994 230225
rect 445172 225358 445228 225367
rect 445172 225293 445228 225302
rect 444466 221764 444542 221792
rect 444466 221482 444494 221764
rect 445186 221482 445214 225293
rect 445954 221482 445982 230219
rect 446722 221792 446750 239691
rect 470902 239675 470954 239681
rect 470902 239617 470954 239623
rect 458806 239527 458858 239533
rect 458806 239469 458858 239475
rect 455158 239009 455210 239015
rect 455158 238951 455210 238957
rect 455062 238935 455114 238941
rect 455062 238877 455114 238883
rect 450454 237529 450506 237535
rect 450454 237471 450506 237477
rect 449302 234643 449354 234649
rect 449302 234585 449354 234591
rect 448246 233459 448298 233465
rect 448246 233401 448298 233407
rect 447478 224579 447530 224585
rect 447478 224521 447530 224527
rect 446674 221764 446750 221792
rect 446674 221482 446702 221764
rect 447490 221482 447518 224521
rect 448258 221482 448286 233401
rect 448916 231426 448972 231435
rect 448916 231361 448972 231370
rect 448930 221792 448958 231361
rect 449314 230209 449342 234585
rect 449686 230869 449738 230875
rect 449686 230811 449738 230817
rect 449302 230203 449354 230209
rect 449302 230145 449354 230151
rect 448930 221764 449006 221792
rect 448978 221482 449006 221764
rect 449698 221482 449726 230811
rect 450466 221482 450494 237471
rect 454294 230425 454346 230431
rect 454294 230367 454346 230373
rect 451990 227687 452042 227693
rect 451990 227629 452042 227635
rect 451222 225689 451274 225695
rect 451222 225631 451274 225637
rect 451234 221792 451262 225631
rect 451234 221764 451310 221792
rect 451282 221482 451310 221764
rect 452002 221482 452030 227629
rect 452758 224505 452810 224511
rect 452758 224447 452810 224453
rect 452770 221482 452798 224447
rect 453430 224431 453482 224437
rect 453430 224373 453482 224379
rect 453442 221792 453470 224373
rect 453442 221764 453518 221792
rect 453490 221482 453518 221764
rect 454306 221482 454334 230367
rect 455074 228581 455102 238877
rect 455170 236174 455198 238951
rect 455170 236146 455774 236174
rect 455156 231574 455212 231583
rect 455156 231509 455212 231518
rect 455062 228575 455114 228581
rect 455062 228517 455114 228523
rect 455170 226232 455198 231509
rect 455074 226204 455198 226232
rect 455074 221482 455102 226204
rect 455746 221792 455774 236146
rect 458038 230055 458090 230061
rect 458038 229997 458090 230003
rect 456502 228575 456554 228581
rect 456502 228517 456554 228523
rect 455746 221764 455822 221792
rect 455794 221482 455822 221764
rect 456514 221482 456542 228517
rect 457268 225506 457324 225515
rect 457268 225441 457324 225450
rect 457282 221482 457310 225441
rect 458050 221792 458078 229997
rect 458050 221764 458126 221792
rect 458098 221482 458126 221764
rect 458818 221482 458846 239469
rect 462550 238861 462602 238867
rect 462550 238803 462602 238809
rect 460246 235901 460298 235907
rect 460246 235843 460298 235849
rect 459574 224357 459626 224363
rect 459574 224299 459626 224305
rect 459586 221482 459614 224299
rect 460258 221792 460286 235843
rect 461014 230129 461066 230135
rect 461014 230071 461066 230077
rect 460258 221764 460334 221792
rect 460306 221482 460334 221764
rect 461026 221482 461054 230071
rect 461878 228353 461930 228359
rect 461878 228295 461930 228301
rect 461890 221482 461918 228295
rect 462562 221792 462590 238803
rect 464758 238787 464810 238793
rect 464758 238729 464810 238735
rect 463606 233385 463658 233391
rect 463606 233327 463658 233333
rect 463618 230135 463646 233327
rect 464086 231609 464138 231615
rect 464086 231551 464138 231557
rect 463606 230129 463658 230135
rect 463606 230071 463658 230077
rect 463316 225654 463372 225663
rect 463316 225589 463372 225598
rect 462562 221764 462638 221792
rect 462610 221482 462638 221764
rect 463330 221482 463358 225589
rect 464098 221482 464126 231551
rect 464770 221792 464798 238729
rect 468598 238713 468650 238719
rect 468598 238655 468650 238661
rect 466486 233533 466538 233539
rect 466486 233475 466538 233481
rect 466390 230203 466442 230209
rect 466390 230145 466442 230151
rect 465622 224135 465674 224141
rect 465622 224077 465674 224083
rect 464770 221764 464846 221792
rect 464818 221482 464846 221764
rect 465634 221482 465662 224077
rect 466402 221482 466430 230145
rect 466498 230061 466526 233475
rect 466486 230055 466538 230061
rect 466486 229997 466538 230003
rect 467062 229981 467114 229987
rect 467062 229923 467114 229929
rect 467074 221792 467102 229923
rect 467830 224209 467882 224215
rect 467830 224151 467882 224157
rect 467074 221764 467150 221792
rect 467122 221482 467150 221764
rect 467842 221482 467870 224151
rect 468610 221482 468638 238655
rect 470132 231722 470188 231731
rect 470132 231657 470188 231666
rect 469364 225802 469420 225811
rect 469364 225737 469420 225746
rect 469378 221496 469406 225737
rect 469378 221468 469440 221496
rect 470146 221482 470174 231657
rect 470914 221496 470942 239617
rect 488278 239601 488330 239607
rect 488278 239543 488330 239549
rect 474646 238639 474698 238645
rect 474646 238581 474698 238587
rect 472340 234090 472396 234099
rect 472340 234025 472396 234034
rect 471574 224283 471626 224289
rect 471574 224225 471626 224231
rect 470880 221468 470942 221496
rect 471586 221496 471614 224225
rect 471586 221468 471648 221496
rect 472354 221482 472382 234025
rect 473878 231239 473930 231245
rect 473878 231181 473930 231187
rect 473110 229907 473162 229913
rect 473110 229849 473162 229855
rect 473122 221792 473150 229849
rect 473122 221764 473198 221792
rect 473170 221482 473198 221764
rect 473890 221482 473918 231181
rect 474658 221482 474686 238581
rect 480694 238565 480746 238571
rect 480694 238507 480746 238513
rect 478102 238491 478154 238497
rect 478102 238433 478154 238439
rect 475222 234051 475274 234057
rect 475222 233993 475274 233999
rect 475234 229987 475262 233993
rect 475222 229981 475274 229987
rect 475222 229923 475274 229929
rect 476950 228427 477002 228433
rect 476950 228369 477002 228375
rect 476180 228170 476236 228179
rect 476180 228105 476236 228114
rect 475316 225210 475372 225219
rect 475316 225145 475372 225154
rect 475330 221792 475358 225145
rect 475330 221764 475406 221792
rect 475378 221482 475406 221764
rect 476194 221482 476222 228105
rect 476962 221482 476990 228369
rect 477622 224061 477674 224067
rect 477622 224003 477674 224009
rect 477634 221792 477662 224003
rect 477634 221764 477710 221792
rect 478114 221773 478142 238433
rect 479158 231683 479210 231689
rect 479158 231625 479210 231631
rect 478390 230129 478442 230135
rect 478390 230071 478442 230077
rect 477682 221482 477710 221764
rect 478102 221767 478154 221773
rect 478102 221709 478154 221715
rect 478402 221482 478430 230071
rect 479170 221482 479198 231625
rect 479974 221767 480026 221773
rect 479974 221709 480026 221715
rect 479986 221482 480014 221709
rect 480706 221482 480734 238507
rect 486742 238417 486794 238423
rect 486742 238359 486794 238365
rect 484630 234125 484682 234131
rect 484630 234067 484682 234073
rect 480884 233942 480940 233951
rect 480884 233877 480940 233886
rect 480898 229913 480926 233877
rect 484438 230055 484490 230061
rect 484438 229997 484490 230003
rect 480886 229907 480938 229913
rect 480886 229849 480938 229855
rect 482134 229833 482186 229839
rect 482134 229775 482186 229781
rect 481460 227430 481516 227439
rect 481460 227365 481516 227374
rect 481474 221482 481502 227365
rect 482146 221792 482174 229775
rect 483766 223987 483818 223993
rect 483766 223929 483818 223935
rect 482902 222433 482954 222439
rect 482902 222375 482954 222381
rect 482146 221764 482222 221792
rect 482194 221482 482222 221764
rect 482914 221482 482942 222375
rect 483778 221482 483806 223929
rect 484450 221792 484478 229997
rect 484642 229839 484670 234067
rect 485206 231757 485258 231763
rect 485206 231699 485258 231705
rect 484630 229833 484682 229839
rect 484630 229775 484682 229781
rect 484450 221764 484526 221792
rect 484498 221482 484526 221764
rect 485218 221482 485246 231699
rect 485974 231313 486026 231319
rect 485974 231255 486026 231261
rect 485986 221482 486014 231255
rect 486754 221792 486782 238359
rect 488290 236174 488318 239543
rect 532822 239453 532874 239459
rect 532822 239395 532874 239401
rect 508630 239157 508682 239163
rect 508630 239099 508682 239105
rect 492790 238343 492842 238349
rect 492790 238285 492842 238291
rect 492022 236345 492074 236351
rect 492022 236287 492074 236293
rect 488290 236146 488990 236174
rect 488276 228318 488332 228327
rect 488276 228253 488332 228262
rect 487508 225950 487564 225959
rect 487508 225885 487564 225894
rect 486706 221764 486782 221792
rect 486706 221482 486734 221764
rect 487522 221482 487550 225885
rect 488290 221482 488318 228253
rect 488962 221792 488990 236146
rect 490484 234238 490540 234247
rect 490484 234173 490540 234182
rect 489718 223913 489770 223919
rect 489718 223855 489770 223861
rect 488962 221764 489038 221792
rect 489010 221482 489038 221764
rect 489730 221482 489758 223855
rect 490498 221482 490526 234173
rect 491254 233237 491306 233243
rect 491254 233179 491306 233185
rect 491266 221792 491294 233179
rect 491266 221764 491342 221792
rect 491314 221482 491342 221764
rect 492034 221482 492062 236287
rect 492802 221482 492830 238285
rect 500278 238269 500330 238275
rect 500278 238211 500330 238217
rect 495766 235827 495818 235833
rect 495766 235769 495818 235775
rect 495382 234199 495434 234205
rect 495382 234141 495434 234147
rect 495394 233243 495422 234141
rect 495382 233237 495434 233243
rect 495092 233202 495148 233211
rect 495382 233179 495434 233185
rect 495092 233137 495148 233146
rect 494228 228466 494284 228475
rect 494228 228401 494284 228410
rect 493460 227282 493516 227291
rect 493460 227217 493516 227226
rect 493474 221792 493502 227217
rect 493474 221764 493550 221792
rect 493522 221482 493550 221764
rect 494242 221482 494270 228401
rect 495106 221482 495134 233137
rect 495778 221792 495806 235769
rect 499606 231387 499658 231393
rect 499606 231329 499658 231335
rect 497972 228614 498028 228623
rect 497972 228549 498028 228558
rect 497302 223839 497354 223845
rect 497302 223781 497354 223787
rect 496534 222507 496586 222513
rect 496534 222449 496586 222455
rect 495778 221764 495854 221792
rect 495826 221482 495854 221764
rect 496546 221482 496574 222449
rect 497314 221482 497342 223781
rect 497986 221792 498014 228549
rect 498836 227134 498892 227143
rect 498836 227069 498892 227078
rect 497986 221764 498062 221792
rect 498034 221482 498062 221764
rect 498850 221482 498878 227069
rect 499618 221496 499646 231329
rect 499584 221468 499646 221496
rect 500290 221496 500318 238211
rect 503350 238195 503402 238201
rect 503350 238137 503402 238143
rect 501046 233163 501098 233169
rect 501046 233105 501098 233111
rect 500290 221468 500352 221496
rect 501058 221482 501086 233105
rect 502582 228501 502634 228507
rect 502582 228443 502634 228449
rect 501814 223765 501866 223771
rect 501814 223707 501866 223713
rect 501826 221792 501854 223707
rect 501826 221764 501902 221792
rect 501874 221482 501902 221764
rect 502594 221482 502622 228443
rect 503362 221482 503390 238137
rect 505654 236271 505706 236277
rect 505654 236213 505706 236219
rect 503926 234273 503978 234279
rect 503926 234215 503978 234221
rect 503938 230061 503966 234215
rect 503926 230055 503978 230061
rect 503926 229997 503978 230003
rect 504022 229759 504074 229765
rect 504022 229701 504074 229707
rect 504034 221792 504062 229701
rect 504790 223543 504842 223549
rect 504790 223485 504842 223491
rect 504034 221764 504110 221792
rect 504082 221482 504110 221764
rect 504802 221482 504830 223485
rect 505666 221482 505694 236213
rect 507094 233089 507146 233095
rect 507094 233031 507146 233037
rect 506326 223617 506378 223623
rect 506326 223559 506378 223565
rect 506338 221792 506366 223559
rect 506338 221764 506414 221792
rect 506386 221482 506414 221764
rect 507106 221482 507134 233031
rect 507862 223691 507914 223697
rect 507862 223633 507914 223639
rect 507874 221482 507902 223633
rect 508642 221792 508670 239099
rect 509398 238121 509450 238127
rect 509398 238063 509450 238069
rect 508594 221764 508670 221792
rect 508594 221482 508622 221764
rect 509410 221482 509438 238063
rect 514678 238047 514730 238053
rect 514678 237989 514730 237995
rect 512758 237973 512810 237979
rect 512758 237915 512810 237921
rect 510166 229611 510218 229617
rect 510166 229553 510218 229559
rect 510178 221482 510206 229553
rect 510838 223395 510890 223401
rect 510838 223337 510890 223343
rect 510850 221792 510878 223337
rect 512374 223321 512426 223327
rect 512374 223263 512426 223269
rect 511606 222729 511658 222735
rect 511606 222671 511658 222677
rect 510850 221764 510926 221792
rect 510898 221482 510926 221764
rect 511618 221482 511646 222671
rect 512386 221482 512414 223263
rect 512770 221773 512798 237915
rect 513142 233015 513194 233021
rect 513142 232957 513194 232963
rect 513154 221792 513182 232957
rect 513910 223469 513962 223475
rect 513910 223411 513962 223417
rect 512758 221767 512810 221773
rect 513154 221764 513230 221792
rect 512758 221709 512810 221715
rect 513202 221482 513230 221764
rect 513922 221482 513950 223411
rect 514690 221482 514718 237989
rect 522166 237899 522218 237905
rect 522166 237841 522218 237847
rect 522178 236174 522206 237841
rect 521506 236146 522206 236174
rect 523798 236197 523850 236203
rect 519190 232867 519242 232873
rect 519190 232809 519242 232815
rect 516118 229537 516170 229543
rect 516118 229479 516170 229485
rect 515398 221767 515450 221773
rect 515398 221709 515450 221715
rect 515410 221482 515438 221709
rect 516130 221482 516158 229479
rect 517654 228649 517706 228655
rect 517654 228591 517706 228597
rect 516982 223247 517034 223253
rect 516982 223189 517034 223195
rect 516994 221482 517022 223189
rect 517666 221792 517694 228591
rect 518420 224618 518476 224627
rect 518420 224553 518476 224562
rect 517666 221764 517742 221792
rect 517714 221482 517742 221764
rect 518434 221482 518462 224553
rect 519202 221482 519230 232809
rect 520726 231461 520778 231467
rect 520726 231403 520778 231409
rect 519860 222694 519916 222703
rect 519860 222629 519916 222638
rect 519874 221792 519902 222629
rect 519874 221764 519950 221792
rect 519922 221482 519950 221764
rect 520738 221482 520766 231403
rect 521506 221482 521534 236146
rect 523798 236139 523850 236145
rect 522166 229389 522218 229395
rect 522166 229331 522218 229337
rect 522178 221792 522206 229331
rect 522932 222546 522988 222555
rect 522932 222481 522988 222490
rect 522178 221764 522254 221792
rect 522226 221482 522254 221764
rect 522946 221482 522974 222481
rect 523810 221482 523838 236139
rect 525238 232793 525290 232799
rect 525238 232735 525290 232741
rect 524468 224470 524524 224479
rect 524468 224405 524524 224414
rect 524482 221792 524510 224405
rect 524482 221764 524558 221792
rect 524530 221482 524558 221764
rect 525250 221482 525278 232735
rect 531286 232645 531338 232651
rect 531286 232587 531338 232593
rect 527540 230094 527596 230103
rect 527540 230029 527596 230038
rect 526004 222990 526060 222999
rect 526004 222925 526060 222934
rect 526018 221482 526046 222925
rect 526676 222842 526732 222851
rect 526676 222777 526732 222786
rect 526690 221792 526718 222777
rect 526690 221764 526766 221792
rect 526738 221482 526766 221764
rect 527554 221482 527582 230029
rect 529750 228871 529802 228877
rect 529750 228813 529802 228819
rect 528308 228762 528364 228771
rect 528308 228697 528364 228706
rect 528322 221496 528350 228697
rect 528980 224026 529036 224035
rect 528980 223961 529036 223970
rect 528288 221468 528350 221496
rect 528994 221496 529022 223961
rect 528994 221468 529056 221496
rect 529762 221482 529790 228813
rect 530516 224322 530572 224331
rect 530516 224257 530572 224266
rect 530530 221496 530558 224257
rect 530496 221468 530558 221496
rect 531298 221482 531326 232587
rect 532052 224174 532108 224183
rect 532052 224109 532108 224118
rect 532066 221482 532094 224109
rect 532834 221792 532862 239395
rect 541462 239379 541514 239385
rect 541462 239321 541514 239327
rect 538004 238086 538060 238095
rect 538004 238021 538060 238030
rect 535126 237825 535178 237831
rect 535126 237767 535178 237773
rect 533494 237751 533546 237757
rect 533494 237693 533546 237699
rect 532786 221764 532862 221792
rect 532786 221482 532814 221764
rect 533506 221482 533534 237693
rect 534260 230242 534316 230251
rect 534260 230177 534316 230186
rect 534274 221482 534302 230177
rect 535138 221792 535166 237767
rect 535798 237677 535850 237683
rect 535798 237619 535850 237625
rect 535810 228581 535838 237619
rect 538018 236174 538046 238021
rect 541078 237603 541130 237609
rect 541078 237545 541130 237551
rect 537922 236146 538046 236174
rect 537238 232571 537290 232577
rect 537238 232513 537290 232519
rect 535798 228575 535850 228581
rect 535798 228517 535850 228523
rect 535798 228427 535850 228433
rect 535798 228369 535850 228375
rect 535090 221764 535166 221792
rect 535090 221482 535118 221764
rect 535810 221482 535838 228369
rect 536564 223878 536620 223887
rect 536564 223813 536620 223822
rect 536578 221482 536606 223813
rect 537250 221792 537278 232513
rect 537922 228433 537950 236146
rect 539542 232497 539594 232503
rect 539542 232439 539594 232445
rect 538870 229463 538922 229469
rect 538870 229405 538922 229411
rect 538006 228575 538058 228581
rect 538006 228517 538058 228523
rect 537910 228427 537962 228433
rect 537910 228369 537962 228375
rect 537250 221764 537326 221792
rect 537298 221482 537326 221764
rect 538018 221482 538046 228517
rect 538882 221482 538910 229405
rect 539554 221792 539582 232439
rect 540308 229946 540364 229955
rect 540308 229881 540364 229890
rect 539554 221764 539630 221792
rect 539602 221482 539630 221764
rect 540322 221482 540350 229881
rect 541090 221482 541118 237545
rect 541474 236174 541502 239321
rect 550870 239305 550922 239311
rect 550870 239247 550922 239253
rect 544822 239083 544874 239089
rect 544822 239025 544874 239031
rect 544340 238382 544396 238391
rect 544340 238317 544396 238326
rect 541474 236146 541790 236174
rect 541762 221792 541790 236146
rect 543382 232423 543434 232429
rect 543382 232365 543434 232371
rect 542614 232349 542666 232355
rect 542614 232291 542666 232297
rect 541762 221764 541838 221792
rect 541810 221482 541838 221764
rect 542626 221482 542654 232291
rect 543394 221482 543422 232365
rect 544354 228581 544382 238317
rect 544342 228575 544394 228581
rect 544342 228517 544394 228523
rect 544052 223730 544108 223739
rect 544052 223665 544108 223674
rect 544066 221792 544094 223665
rect 544066 221764 544142 221792
rect 544114 221482 544142 221764
rect 544834 221482 544862 239025
rect 550196 238678 550252 238687
rect 550196 238613 550252 238622
rect 549428 233054 549484 233063
rect 549428 232989 549484 232998
rect 548566 232275 548618 232281
rect 548566 232217 548618 232223
rect 545590 232127 545642 232133
rect 545590 232069 545642 232075
rect 545602 221482 545630 232069
rect 546358 229315 546410 229321
rect 546358 229257 546410 229263
rect 546370 221792 546398 229257
rect 547894 228945 547946 228951
rect 547894 228887 547946 228893
rect 547126 228575 547178 228581
rect 547126 228517 547178 228523
rect 546370 221764 546446 221792
rect 546418 221482 546446 221764
rect 547138 221482 547166 228517
rect 547906 221482 547934 228887
rect 548578 221792 548606 232217
rect 548578 221764 548654 221792
rect 548626 221482 548654 221764
rect 549442 221482 549470 232989
rect 550210 221482 550238 238613
rect 550882 221792 550910 239247
rect 555380 238974 555436 238983
rect 555380 238909 555436 238918
rect 551636 232906 551692 232915
rect 551636 232841 551692 232850
rect 550882 221764 550958 221792
rect 550930 221482 550958 221764
rect 551650 221482 551678 232841
rect 552406 232201 552458 232207
rect 552406 232143 552458 232149
rect 552418 221482 552446 232143
rect 554710 232053 554762 232059
rect 554710 231995 554762 232001
rect 553940 229798 553996 229807
rect 553940 229733 553996 229742
rect 553270 224209 553322 224215
rect 553270 224151 553322 224157
rect 553282 221681 553310 224151
rect 553234 221653 553310 221681
rect 553234 221482 553262 221653
rect 553954 221482 553982 229733
rect 554722 221482 554750 231995
rect 555286 229241 555338 229247
rect 555286 229183 555338 229189
rect 555298 221792 555326 229183
rect 555394 224215 555422 238909
rect 559892 238234 559948 238243
rect 559892 238169 559948 238178
rect 559220 236606 559276 236615
rect 559220 236541 559276 236550
rect 558452 236458 558508 236467
rect 558452 236393 558508 236402
rect 557684 232758 557740 232767
rect 557684 232693 557740 232702
rect 557014 231979 557066 231985
rect 557014 231921 557066 231927
rect 556150 228575 556202 228581
rect 556150 228517 556202 228523
rect 555382 224209 555434 224215
rect 555382 224151 555434 224157
rect 555298 221764 555470 221792
rect 555442 221482 555470 221764
rect 556162 221482 556190 228517
rect 557026 221496 557054 231921
rect 556992 221468 557054 221496
rect 557698 221496 557726 232693
rect 558358 231905 558410 231911
rect 558358 231847 558410 231853
rect 558370 227534 558398 231847
rect 558466 228581 558494 236393
rect 558454 228575 558506 228581
rect 558454 228517 558506 228523
rect 558370 227506 558494 227534
rect 557698 221468 557760 221496
rect 558466 221482 558494 227506
rect 559234 221496 559262 236541
rect 559200 221468 559262 221496
rect 559906 221496 559934 238169
rect 567476 236902 567532 236911
rect 567476 236837 567532 236846
rect 565268 236754 565324 236763
rect 565268 236689 565324 236698
rect 560756 232610 560812 232619
rect 560756 232545 560812 232554
rect 559906 221468 559968 221496
rect 560770 221482 560798 232545
rect 564502 231831 564554 231837
rect 564502 231773 564554 231779
rect 561430 229167 561482 229173
rect 561430 229109 561482 229115
rect 561442 221792 561470 229109
rect 563638 229093 563690 229099
rect 563638 229035 563690 229041
rect 562964 223582 563020 223591
rect 562964 223517 563020 223526
rect 562196 223434 562252 223443
rect 562196 223369 562252 223378
rect 561442 221764 561518 221792
rect 561490 221482 561518 221764
rect 562210 221482 562238 223369
rect 562978 221482 563006 223517
rect 563650 221792 563678 229035
rect 563650 221764 563726 221792
rect 563698 221482 563726 221764
rect 564514 221482 564542 231773
rect 565282 221482 565310 236689
rect 567490 236174 567518 236837
rect 567490 236146 568286 236174
rect 566710 232719 566762 232725
rect 566710 232661 566762 232667
rect 565942 229685 565994 229691
rect 565942 229627 565994 229633
rect 565954 221792 565982 229627
rect 565954 221764 566030 221792
rect 566002 221482 566030 221764
rect 566722 221482 566750 232661
rect 567382 229019 567434 229025
rect 567382 228961 567434 228967
rect 567394 227534 567422 228961
rect 567394 227506 567518 227534
rect 567490 221482 567518 227506
rect 568258 221792 568286 236146
rect 568258 221764 568334 221792
rect 568306 221482 568334 221764
rect 569026 221482 569054 239945
rect 599158 239231 599210 239237
rect 599158 239173 599210 239179
rect 581780 238826 581836 238835
rect 581780 238761 581836 238770
rect 573140 237050 573196 237059
rect 573140 236985 573196 236994
rect 573154 236174 573182 236985
rect 573154 236146 574334 236174
rect 572086 232941 572138 232947
rect 572086 232883 572138 232889
rect 570452 232462 570508 232471
rect 570452 232397 570508 232406
rect 569780 229650 569836 229659
rect 569780 229585 569836 229594
rect 569794 221482 569822 229585
rect 570466 221681 570494 232397
rect 571316 223286 571372 223295
rect 571316 223221 571372 223230
rect 570466 221653 570542 221681
rect 570514 221482 570542 221653
rect 571330 221482 571358 223221
rect 572098 221482 572126 232883
rect 572756 229502 572812 229511
rect 572756 229437 572812 229446
rect 572770 221681 572798 229437
rect 573524 229354 573580 229363
rect 573524 229289 573580 229298
rect 572770 221653 572846 221681
rect 572818 221482 572846 221653
rect 573538 221482 573566 229289
rect 574306 221482 574334 236146
rect 580340 236014 580396 236023
rect 580340 235949 580396 235958
rect 576596 232314 576652 232323
rect 576596 232249 576652 232258
rect 575828 232166 575884 232175
rect 575828 232101 575884 232110
rect 575060 230390 575116 230399
rect 575060 230325 575116 230334
rect 575074 221792 575102 230325
rect 575074 221764 575150 221792
rect 575122 221482 575150 221764
rect 575842 221482 575870 232101
rect 576610 221482 576638 232249
rect 578036 232018 578092 232027
rect 578036 231953 578092 231962
rect 577268 223138 577324 223147
rect 577268 223073 577324 223082
rect 577282 221792 577310 223073
rect 577282 221764 577358 221792
rect 577330 221482 577358 221764
rect 578050 221482 578078 231953
rect 578900 229206 578956 229215
rect 578900 229141 578956 229150
rect 578914 221482 578942 229141
rect 579574 225911 579626 225917
rect 579574 225853 579626 225859
rect 579586 221792 579614 225853
rect 579586 221764 579662 221792
rect 579634 221482 579662 221764
rect 580354 221482 580382 235949
rect 581110 225837 581162 225843
rect 581110 225779 581162 225785
rect 581122 221482 581150 225779
rect 581794 221792 581822 238761
rect 590420 236162 590476 236171
rect 584566 236123 584618 236129
rect 590420 236097 590476 236106
rect 584566 236065 584618 236071
rect 583414 235161 583466 235167
rect 583414 235103 583466 235109
rect 582646 226059 582698 226065
rect 582646 226001 582698 226007
rect 581794 221764 581870 221792
rect 581842 221482 581870 221764
rect 582658 221482 582686 226001
rect 583426 221482 583454 235103
rect 584086 227095 584138 227101
rect 584086 227037 584138 227043
rect 584098 221792 584126 227037
rect 584578 226065 584606 236065
rect 587924 235866 587980 235875
rect 587924 235801 587980 235810
rect 587350 235531 587402 235537
rect 587350 235473 587402 235479
rect 587062 235383 587114 235389
rect 587062 235325 587114 235331
rect 586390 227539 586442 227545
rect 586390 227481 586442 227487
rect 585622 227465 585674 227471
rect 585622 227407 585674 227413
rect 584566 226059 584618 226065
rect 584566 226001 584618 226007
rect 584854 225985 584906 225991
rect 584854 225927 584906 225933
rect 584098 221764 584174 221792
rect 584146 221482 584174 221764
rect 584866 221482 584894 225927
rect 585634 221482 585662 227407
rect 586402 221496 586430 227481
rect 587074 226065 587102 235325
rect 587254 235235 587306 235241
rect 587254 235177 587306 235183
rect 587062 226059 587114 226065
rect 587062 226001 587114 226007
rect 587266 225695 587294 235177
rect 587362 226953 587390 235473
rect 587638 235309 587690 235315
rect 587638 235251 587690 235257
rect 587444 234386 587500 234395
rect 587444 234321 587500 234330
rect 587458 227323 587486 234321
rect 587650 227471 587678 235251
rect 587638 227465 587690 227471
rect 587638 227407 587690 227413
rect 587446 227317 587498 227323
rect 587446 227259 587498 227265
rect 587350 226947 587402 226953
rect 587350 226889 587402 226895
rect 587254 225689 587306 225695
rect 587254 225631 587306 225637
rect 587158 224727 587210 224733
rect 587158 224669 587210 224675
rect 586402 221468 586464 221496
rect 587170 221482 587198 224669
rect 587938 221496 587966 235801
rect 588886 235679 588938 235685
rect 588886 235621 588938 235627
rect 588406 235457 588458 235463
rect 588406 235399 588458 235405
rect 588418 225843 588446 235399
rect 588898 227249 588926 235621
rect 590434 227397 590462 236097
rect 591476 235718 591532 235727
rect 591476 235653 591532 235662
rect 590518 235605 590570 235611
rect 590518 235547 590570 235553
rect 589366 227391 589418 227397
rect 589366 227333 589418 227339
rect 590422 227391 590474 227397
rect 590422 227333 590474 227339
rect 588598 227243 588650 227249
rect 588598 227185 588650 227191
rect 588886 227243 588938 227249
rect 588886 227185 588938 227191
rect 588406 225837 588458 225843
rect 588406 225779 588458 225785
rect 587904 221468 587966 221496
rect 588610 221496 588638 227185
rect 588610 221468 588672 221496
rect 589378 221482 589406 227333
rect 590134 227169 590186 227175
rect 590134 227111 590186 227117
rect 590146 221792 590174 227111
rect 590530 227101 590558 235547
rect 590900 234534 590956 234543
rect 590900 234469 590956 234478
rect 590914 227175 590942 234469
rect 591490 227545 591518 235653
rect 596086 235087 596138 235093
rect 596086 235029 596138 235035
rect 591478 227539 591530 227545
rect 591478 227481 591530 227487
rect 594646 227539 594698 227545
rect 594646 227481 594698 227487
rect 590902 227169 590954 227175
rect 590902 227111 590954 227117
rect 590518 227095 590570 227101
rect 590518 227037 590570 227043
rect 593974 227021 594026 227027
rect 591668 226986 591724 226995
rect 593974 226963 594026 226969
rect 591668 226921 591724 226930
rect 590900 226838 590956 226847
rect 590900 226773 590956 226782
rect 590146 221764 590222 221792
rect 590194 221482 590222 221764
rect 590914 221482 590942 226773
rect 591682 221482 591710 226921
rect 592342 225689 592394 225695
rect 592342 225631 592394 225637
rect 592354 221792 592382 225631
rect 593110 224801 593162 224807
rect 593110 224743 593162 224749
rect 592354 221764 592430 221792
rect 592402 221482 592430 221764
rect 593122 221482 593150 224743
rect 593986 221482 594014 226963
rect 594658 221792 594686 227481
rect 595414 226059 595466 226065
rect 595414 226001 595466 226007
rect 594658 221764 594734 221792
rect 594706 221482 594734 221764
rect 595426 221482 595454 226001
rect 596098 224733 596126 235029
rect 599170 227027 599198 239173
rect 599924 229058 599980 229067
rect 599924 228993 599980 229002
rect 599158 227021 599210 227027
rect 599158 226963 599210 226969
rect 598486 226947 598538 226953
rect 598486 226889 598538 226895
rect 596180 226690 596236 226699
rect 596180 226625 596236 226634
rect 596086 224727 596138 224733
rect 596086 224669 596138 224675
rect 596194 221482 596222 226625
rect 596948 226542 597004 226551
rect 596948 226477 597004 226486
rect 596962 221792 596990 226477
rect 597718 224727 597770 224733
rect 597718 224669 597770 224675
rect 596962 221764 597038 221792
rect 597010 221482 597038 221764
rect 597730 221482 597758 224669
rect 598498 221482 598526 226889
rect 599158 226873 599210 226879
rect 599158 226815 599210 226821
rect 599170 221792 599198 226815
rect 599170 221764 599246 221792
rect 599218 221482 599246 221764
rect 599938 221482 599966 228993
rect 600418 226879 600446 241911
rect 601462 229981 601514 229987
rect 601462 229923 601514 229929
rect 600790 227465 600842 227471
rect 600790 227407 600842 227413
rect 600406 226873 600458 226879
rect 600406 226815 600458 226821
rect 600802 221482 600830 227407
rect 601474 221792 601502 229923
rect 603298 226731 603326 253455
rect 603382 250627 603434 250633
rect 603382 250569 603434 250575
rect 603394 226805 603422 250569
rect 603478 247815 603530 247821
rect 603478 247757 603530 247763
rect 603382 226799 603434 226805
rect 603382 226741 603434 226747
rect 602998 226725 603050 226731
rect 602998 226667 603050 226673
rect 603286 226725 603338 226731
rect 603286 226667 603338 226673
rect 602230 225837 602282 225843
rect 602230 225779 602282 225785
rect 601474 221764 601550 221792
rect 601522 221482 601550 221764
rect 602242 221482 602270 225779
rect 603010 221482 603038 226667
rect 603490 225991 603518 247757
rect 605974 235013 606026 235019
rect 605974 234955 606026 234961
rect 605302 234939 605354 234945
rect 605302 234881 605354 234887
rect 604532 231870 604588 231879
rect 604532 231805 604588 231814
rect 603670 226651 603722 226657
rect 603670 226593 603722 226599
rect 603478 225985 603530 225991
rect 603478 225927 603530 225933
rect 603682 221792 603710 226593
rect 603682 221764 603758 221792
rect 603730 221482 603758 221764
rect 604546 221482 604574 231805
rect 605314 221482 605342 234881
rect 605986 221792 606014 234955
rect 606178 226657 606206 262113
rect 606262 259285 606314 259291
rect 606262 259227 606314 259233
rect 606274 227545 606302 259227
rect 606358 256399 606410 256405
rect 606358 256341 606410 256347
rect 606262 227539 606314 227545
rect 606262 227481 606314 227487
rect 606370 227027 606398 256341
rect 629206 247741 629258 247747
rect 629206 247683 629258 247689
rect 627188 240158 627244 240167
rect 627188 240093 627244 240102
rect 621140 236310 621196 236319
rect 621140 236245 621196 236254
rect 608276 235570 608332 235579
rect 608276 235505 608332 235514
rect 607508 228910 607564 228919
rect 607508 228845 607564 228854
rect 606358 227021 606410 227027
rect 606358 226963 606410 226969
rect 606166 226651 606218 226657
rect 606166 226593 606218 226599
rect 606742 225171 606794 225177
rect 606742 225113 606794 225119
rect 605986 221764 606062 221792
rect 606034 221482 606062 221764
rect 606754 221482 606782 225113
rect 607522 221482 607550 228845
rect 608290 221792 608318 235505
rect 611252 235422 611308 235431
rect 611252 235357 611308 235366
rect 609046 229907 609098 229913
rect 609046 229849 609098 229855
rect 608290 221764 608366 221792
rect 608338 221482 608366 221764
rect 609058 221482 609086 229849
rect 609814 226577 609866 226583
rect 609814 226519 609866 226525
rect 609826 221482 609854 226519
rect 610486 225763 610538 225769
rect 610486 225705 610538 225711
rect 610498 221792 610526 225705
rect 610498 221764 610574 221792
rect 610546 221482 610574 221764
rect 611266 221482 611294 235357
rect 614324 235274 614380 235283
rect 614324 235209 614380 235218
rect 612118 229833 612170 229839
rect 612118 229775 612170 229781
rect 612130 221482 612158 229775
rect 612790 226503 612842 226509
rect 612790 226445 612842 226451
rect 612802 221792 612830 226445
rect 613558 226429 613610 226435
rect 613558 226371 613610 226377
rect 612802 221764 612878 221792
rect 612850 221482 612878 221764
rect 613570 221482 613598 226371
rect 614338 221482 614366 235209
rect 618836 235126 618892 235135
rect 618836 235061 618892 235070
rect 616628 234978 616684 234987
rect 616628 234913 616684 234922
rect 615862 234865 615914 234871
rect 615862 234807 615914 234813
rect 614998 233237 615050 233243
rect 614998 233179 615050 233185
rect 615010 221792 615038 233179
rect 615010 221764 615086 221792
rect 615058 221482 615086 221764
rect 615874 221482 615902 234807
rect 616642 221496 616670 234913
rect 617300 226394 617356 226403
rect 617300 226329 617356 226338
rect 618070 226355 618122 226361
rect 616608 221468 616670 221496
rect 617314 221496 617342 226329
rect 618070 226297 618122 226303
rect 617314 221468 617376 221496
rect 618082 221482 618110 226297
rect 618850 221792 618878 235061
rect 619604 234830 619660 234839
rect 619604 234765 619660 234774
rect 618850 221764 618926 221792
rect 618898 221482 618926 221764
rect 619618 221482 619646 234765
rect 620372 226246 620428 226255
rect 620372 226181 620428 226190
rect 620386 221482 620414 226181
rect 621154 221792 621182 236245
rect 621814 234791 621866 234797
rect 621814 234733 621866 234739
rect 621106 221764 621182 221792
rect 621106 221482 621134 221764
rect 621826 221482 621854 234733
rect 624886 234717 624938 234723
rect 624886 234659 624938 234665
rect 625556 234682 625612 234691
rect 622678 230055 622730 230061
rect 622678 229997 622730 230003
rect 622690 221482 622718 229997
rect 624118 226281 624170 226287
rect 624118 226223 624170 226229
rect 623348 226098 623404 226107
rect 623348 226033 623404 226042
rect 623362 221792 623390 226033
rect 623362 221764 623438 221792
rect 623410 221482 623438 221764
rect 624130 221482 624158 226223
rect 624898 221482 624926 234659
rect 625556 234617 625612 234626
rect 625570 221792 625598 234617
rect 626422 227243 626474 227249
rect 626422 227185 626474 227191
rect 625570 221764 625646 221792
rect 625618 221482 625646 221764
rect 626434 221482 626462 227185
rect 627202 221482 627230 240093
rect 627862 227391 627914 227397
rect 627862 227333 627914 227339
rect 627874 221792 627902 227333
rect 629218 226435 629246 247683
rect 629302 244855 629354 244861
rect 629302 244797 629354 244803
rect 629314 227545 629342 244797
rect 629302 227539 629354 227545
rect 629302 227481 629354 227487
rect 634006 227539 634058 227545
rect 634006 227481 634058 227487
rect 630166 227317 630218 227323
rect 630166 227259 630218 227265
rect 629206 226429 629258 226435
rect 629206 226371 629258 226377
rect 629398 226207 629450 226213
rect 629398 226149 629450 226155
rect 628630 226059 628682 226065
rect 628630 226001 628682 226007
rect 627874 221764 627950 221792
rect 627922 221482 627950 221764
rect 628642 221482 628670 226001
rect 629410 221482 629438 226149
rect 630178 221792 630206 227259
rect 630934 227169 630986 227175
rect 630934 227111 630986 227117
rect 630178 221764 630254 221792
rect 630226 221482 630254 221764
rect 630946 221482 630974 227111
rect 632374 227095 632426 227101
rect 632374 227037 632426 227043
rect 631702 226133 631754 226139
rect 631702 226075 631754 226081
rect 631714 221482 631742 226075
rect 632386 221792 632414 227037
rect 633142 226947 633194 226953
rect 633142 226889 633194 226895
rect 632386 221764 632462 221792
rect 632434 221482 632462 221764
rect 633154 221482 633182 226889
rect 634018 221482 634046 227481
rect 639190 227465 639242 227471
rect 639190 227407 639242 227413
rect 638518 227021 638570 227027
rect 638518 226963 638570 226969
rect 634678 226873 634730 226879
rect 634678 226815 634730 226821
rect 634690 221792 634718 226815
rect 636886 226799 636938 226805
rect 636886 226741 636938 226747
rect 635446 226429 635498 226435
rect 635446 226371 635498 226377
rect 634690 221764 634766 221792
rect 634738 221482 634766 221764
rect 635458 221482 635486 226371
rect 636214 225985 636266 225991
rect 636214 225927 636266 225933
rect 636226 221482 636254 225927
rect 636898 221792 636926 226741
rect 637750 226725 637802 226731
rect 637750 226667 637802 226673
rect 636898 221764 636974 221792
rect 636946 221482 636974 221764
rect 637762 221482 637790 226667
rect 638530 221482 638558 226963
rect 639202 221792 639230 227407
rect 639958 226651 640010 226657
rect 639958 226593 640010 226599
rect 639202 221764 639278 221792
rect 639250 221482 639278 221764
rect 639970 221482 639998 226593
rect 640148 212334 640204 212343
rect 640148 212269 640204 212278
rect 640162 211603 640190 212269
rect 640148 211594 640204 211603
rect 640148 211529 640204 211538
rect 190292 201382 190348 201391
rect 190292 201317 190348 201326
rect 190306 200577 190334 201317
rect 640148 200938 640204 200947
rect 640148 200873 640204 200882
rect 190292 200568 190348 200577
rect 190292 200503 190348 200512
rect 640162 200207 640190 200873
rect 640148 200198 640204 200207
rect 640148 200133 640204 200142
rect 187220 199162 187276 199171
rect 187220 199097 187276 199106
rect 185974 198605 186026 198611
rect 185974 198547 186026 198553
rect 185986 196803 186014 198547
rect 186070 198531 186122 198537
rect 186070 198473 186122 198479
rect 185972 196794 186028 196803
rect 185972 196729 186028 196738
rect 186082 196063 186110 198473
rect 186068 196054 186124 196063
rect 186068 195989 186124 195998
rect 185890 195826 186302 195854
rect 186070 185803 186122 185809
rect 186070 185745 186122 185751
rect 185974 182991 186026 182997
rect 185974 182933 186026 182939
rect 185780 182438 185836 182447
rect 185780 182373 185836 182382
rect 185602 175666 185726 175694
rect 185602 173271 185630 175666
rect 185588 173262 185644 173271
rect 185588 173197 185644 173206
rect 185314 165598 185822 165626
rect 184532 164826 184588 164835
rect 184532 164761 184588 164770
rect 184534 164121 184586 164127
rect 184340 164086 184396 164095
rect 184534 164063 184586 164069
rect 184340 164021 184342 164030
rect 184394 164021 184396 164030
rect 184342 163989 184394 163995
rect 184438 163973 184490 163979
rect 184438 163915 184490 163921
rect 184342 163899 184394 163905
rect 184342 163841 184394 163847
rect 184354 162615 184382 163841
rect 184340 162606 184396 162615
rect 184340 162541 184396 162550
rect 184450 161875 184478 163915
rect 184546 163355 184574 164063
rect 184532 163346 184588 163355
rect 184532 163281 184588 163290
rect 184436 161866 184492 161875
rect 184436 161801 184492 161810
rect 184438 161235 184490 161241
rect 184438 161177 184490 161183
rect 184342 161013 184394 161019
rect 184450 160987 184478 161177
rect 184534 161161 184586 161167
rect 184534 161103 184586 161109
rect 184342 160955 184394 160961
rect 184436 160978 184492 160987
rect 184354 159507 184382 160955
rect 184436 160913 184492 160922
rect 184546 160395 184574 161103
rect 184630 161087 184682 161093
rect 184630 161029 184682 161035
rect 184532 160386 184588 160395
rect 184532 160321 184588 160330
rect 184340 159498 184396 159507
rect 184340 159433 184396 159442
rect 184642 158915 184670 161029
rect 184628 158906 184684 158915
rect 184628 158841 184684 158850
rect 184342 158423 184394 158429
rect 184342 158365 184394 158371
rect 184354 158027 184382 158365
rect 184438 158349 184490 158355
rect 184438 158291 184490 158297
rect 184340 158018 184396 158027
rect 184340 157953 184396 157962
rect 184450 157435 184478 158291
rect 184534 158275 184586 158281
rect 184534 158217 184586 158223
rect 184436 157426 184492 157435
rect 184436 157361 184492 157370
rect 184546 156547 184574 158217
rect 184630 158201 184682 158207
rect 184630 158143 184682 158149
rect 184532 156538 184588 156547
rect 184532 156473 184588 156482
rect 184642 155659 184670 158143
rect 184628 155650 184684 155659
rect 184628 155585 184684 155594
rect 184534 155537 184586 155543
rect 184534 155479 184586 155485
rect 184438 155389 184490 155395
rect 184438 155331 184490 155337
rect 184342 155315 184394 155321
rect 184342 155257 184394 155263
rect 184354 155067 184382 155257
rect 184340 155058 184396 155067
rect 184340 154993 184396 155002
rect 184450 154179 184478 155331
rect 184436 154170 184492 154179
rect 184436 154105 184492 154114
rect 184546 153587 184574 155479
rect 184630 155463 184682 155469
rect 184630 155405 184682 155411
rect 184532 153578 184588 153587
rect 184532 153513 184588 153522
rect 184642 152699 184670 155405
rect 184628 152690 184684 152699
rect 184534 152651 184586 152657
rect 184628 152625 184684 152634
rect 184534 152593 184586 152599
rect 184342 152577 184394 152583
rect 184342 152519 184394 152525
rect 184354 151959 184382 152519
rect 184438 152503 184490 152509
rect 184438 152445 184490 152451
rect 184340 151950 184396 151959
rect 184340 151885 184396 151894
rect 184450 151219 184478 152445
rect 184436 151210 184492 151219
rect 184436 151145 184492 151154
rect 184546 150479 184574 152593
rect 184532 150470 184588 150479
rect 184532 150405 184588 150414
rect 184340 149730 184396 149739
rect 184340 149665 184396 149674
rect 184438 149691 184490 149697
rect 184354 149549 184382 149665
rect 184438 149633 184490 149639
rect 184342 149543 184394 149549
rect 184342 149485 184394 149491
rect 184450 148999 184478 149633
rect 184534 149617 184586 149623
rect 184534 149559 184586 149565
rect 184436 148990 184492 148999
rect 184436 148925 184492 148934
rect 184546 147371 184574 149559
rect 184532 147362 184588 147371
rect 184532 147297 184588 147306
rect 184534 146879 184586 146885
rect 184534 146821 184586 146827
rect 184438 146805 184490 146811
rect 184438 146747 184490 146753
rect 184342 146731 184394 146737
rect 184342 146673 184394 146679
rect 184354 145891 184382 146673
rect 184340 145882 184396 145891
rect 184340 145817 184396 145826
rect 184450 145151 184478 146747
rect 184436 145142 184492 145151
rect 184436 145077 184492 145086
rect 184546 144411 184574 146821
rect 184630 146657 184682 146663
rect 184628 146622 184630 146631
rect 184682 146622 184684 146631
rect 184628 146557 184684 146566
rect 184532 144402 184588 144411
rect 184532 144337 184588 144346
rect 183094 143993 183146 143999
rect 183094 143935 183146 143941
rect 184630 143993 184682 143999
rect 184630 143935 184682 143941
rect 184438 143919 184490 143925
rect 184438 143861 184490 143867
rect 184342 143845 184394 143851
rect 184342 143787 184394 143793
rect 184354 143671 184382 143787
rect 184340 143662 184396 143671
rect 184340 143597 184396 143606
rect 184450 142783 184478 143861
rect 184534 143771 184586 143777
rect 184534 143713 184586 143719
rect 184436 142774 184492 142783
rect 184436 142709 184492 142718
rect 184546 141303 184574 143713
rect 184642 142191 184670 143935
rect 184628 142182 184684 142191
rect 184628 142117 184684 142126
rect 184532 141294 184588 141303
rect 184532 141229 184588 141238
rect 184534 141107 184586 141113
rect 184534 141049 184586 141055
rect 184438 141033 184490 141039
rect 184438 140975 184490 140981
rect 184342 140959 184394 140965
rect 184342 140901 184394 140907
rect 184354 140563 184382 140901
rect 184340 140554 184396 140563
rect 184340 140489 184396 140498
rect 184450 139823 184478 140975
rect 184436 139814 184492 139823
rect 184436 139749 184492 139758
rect 184546 138935 184574 141049
rect 184532 138926 184588 138935
rect 184532 138861 184588 138870
rect 184438 135335 184490 135341
rect 184438 135277 184490 135283
rect 184342 135261 184394 135267
rect 184342 135203 184394 135209
rect 184354 134495 184382 135203
rect 184340 134486 184396 134495
rect 184340 134421 184396 134430
rect 184450 133015 184478 135277
rect 185794 135235 185822 165598
rect 185986 137455 186014 182933
rect 186082 138343 186110 185745
rect 186166 182917 186218 182923
rect 186166 182859 186218 182865
rect 186068 138334 186124 138343
rect 186068 138269 186124 138278
rect 185972 137446 186028 137455
rect 185972 137381 186028 137390
rect 186178 136863 186206 182859
rect 186274 174751 186302 195826
rect 640244 185694 640300 185703
rect 640244 185629 640300 185638
rect 640258 184963 640286 185629
rect 640244 184954 640300 184963
rect 640244 184889 640300 184898
rect 186742 184175 186794 184181
rect 186742 184117 186794 184123
rect 186754 183187 186782 184117
rect 186740 183178 186796 183187
rect 186740 183113 186796 183122
rect 645142 183139 645194 183145
rect 645142 183081 645194 183087
rect 645154 183039 645182 183081
rect 645140 183030 645196 183039
rect 645140 182965 645196 182974
rect 186454 180031 186506 180037
rect 186454 179973 186506 179979
rect 186260 174742 186316 174751
rect 186260 174677 186316 174686
rect 186262 174259 186314 174265
rect 186262 174201 186314 174207
rect 186164 136854 186220 136863
rect 186164 136789 186220 136798
rect 185780 135226 185836 135235
rect 185780 135161 185836 135170
rect 184726 134373 184778 134379
rect 184726 134315 184778 134321
rect 184436 133006 184492 133015
rect 184436 132941 184492 132950
rect 182998 132523 183050 132529
rect 182998 132465 183050 132471
rect 182902 112247 182954 112253
rect 182902 112189 182954 112195
rect 183010 106555 183038 132465
rect 184630 132449 184682 132455
rect 184630 132391 184682 132397
rect 184534 132375 184586 132381
rect 184534 132317 184586 132323
rect 184438 132301 184490 132307
rect 184340 132266 184396 132275
rect 184438 132243 184490 132249
rect 184340 132201 184342 132210
rect 184394 132201 184396 132210
rect 184342 132169 184394 132175
rect 184450 131535 184478 132243
rect 184436 131526 184492 131535
rect 184436 131461 184492 131470
rect 184546 130647 184574 132317
rect 184532 130638 184588 130647
rect 184532 130573 184588 130582
rect 184642 129907 184670 132391
rect 184628 129898 184684 129907
rect 184628 129833 184684 129842
rect 184438 129489 184490 129495
rect 184438 129431 184490 129437
rect 184342 129341 184394 129347
rect 184342 129283 184394 129289
rect 184354 128427 184382 129283
rect 184340 128418 184396 128427
rect 184340 128353 184396 128362
rect 184450 127687 184478 129431
rect 184534 129415 184586 129421
rect 184534 129357 184586 129363
rect 184436 127678 184492 127687
rect 184436 127613 184492 127622
rect 184546 126947 184574 129357
rect 184532 126938 184588 126947
rect 184532 126873 184588 126882
rect 184438 126677 184490 126683
rect 184438 126619 184490 126625
rect 184342 126529 184394 126535
rect 184342 126471 184394 126477
rect 184354 125467 184382 126471
rect 184450 126059 184478 126619
rect 184534 126603 184586 126609
rect 184534 126545 184586 126551
rect 184436 126050 184492 126059
rect 184436 125985 184492 125994
rect 184340 125458 184396 125467
rect 184340 125393 184396 125402
rect 184546 124579 184574 126545
rect 184532 124570 184588 124579
rect 184532 124505 184588 124514
rect 184534 123865 184586 123871
rect 184340 123830 184396 123839
rect 184534 123807 184586 123813
rect 184340 123765 184342 123774
rect 184394 123765 184396 123774
rect 184342 123733 184394 123739
rect 184438 123717 184490 123723
rect 184438 123659 184490 123665
rect 184342 123643 184394 123649
rect 184342 123585 184394 123591
rect 184354 122211 184382 123585
rect 184450 123099 184478 123659
rect 184436 123090 184492 123099
rect 184436 123025 184492 123034
rect 184340 122202 184396 122211
rect 184340 122137 184396 122146
rect 184546 121619 184574 123807
rect 184532 121610 184588 121619
rect 184532 121545 184588 121554
rect 184342 120979 184394 120985
rect 184342 120921 184394 120927
rect 184354 120731 184382 120921
rect 184438 120905 184490 120911
rect 184438 120847 184490 120853
rect 184340 120722 184396 120731
rect 184340 120657 184396 120666
rect 184450 120139 184478 120847
rect 184534 120831 184586 120837
rect 184534 120773 184586 120779
rect 184436 120130 184492 120139
rect 184436 120065 184492 120074
rect 184546 119251 184574 120773
rect 184532 119242 184588 119251
rect 184532 119177 184588 119186
rect 184738 118659 184766 134315
rect 186274 133755 186302 174201
rect 186466 135975 186494 179973
rect 645142 179439 645194 179445
rect 645142 179381 645194 179387
rect 645154 179339 645182 179381
rect 645140 179330 645196 179339
rect 645140 179265 645196 179274
rect 645142 174925 645194 174931
rect 645140 174890 645142 174899
rect 645194 174890 645196 174899
rect 645140 174825 645196 174834
rect 645142 171077 645194 171083
rect 645140 171042 645142 171051
rect 645194 171042 645196 171051
rect 645140 170977 645196 170986
rect 645142 168265 645194 168271
rect 645142 168207 645194 168213
rect 645154 167795 645182 168207
rect 645140 167786 645196 167795
rect 645140 167721 645196 167730
rect 645142 163381 645194 163387
rect 645140 163346 645142 163355
rect 645194 163346 645196 163355
rect 645140 163281 645196 163290
rect 645142 159755 645194 159761
rect 645142 159697 645194 159703
rect 645154 159507 645182 159697
rect 645140 159498 645196 159507
rect 645140 159433 645196 159442
rect 645142 156055 645194 156061
rect 645142 155997 645194 156003
rect 645154 155511 645182 155997
rect 645140 155502 645196 155511
rect 645140 155437 645196 155446
rect 645142 152577 645194 152583
rect 645140 152542 645142 152551
rect 645194 152542 645196 152551
rect 645140 152477 645196 152486
rect 186742 149765 186794 149771
rect 186742 149707 186794 149713
rect 186754 148111 186782 149707
rect 645142 148211 645194 148217
rect 645142 148153 645194 148159
rect 645154 148111 645182 148153
rect 186740 148102 186796 148111
rect 186740 148037 186796 148046
rect 645140 148102 645196 148111
rect 645140 148037 645196 148046
rect 186452 135966 186508 135975
rect 186452 135901 186508 135910
rect 186260 133746 186316 133755
rect 186260 133681 186316 133690
rect 185686 129637 185738 129643
rect 185686 129579 185738 129585
rect 645718 129637 645770 129643
rect 645718 129579 645770 129585
rect 184724 118650 184780 118659
rect 184724 118585 184780 118594
rect 184630 118093 184682 118099
rect 184630 118035 184682 118041
rect 184534 118019 184586 118025
rect 184534 117961 184586 117967
rect 184438 117945 184490 117951
rect 184438 117887 184490 117893
rect 184342 117871 184394 117877
rect 184342 117813 184394 117819
rect 184354 117771 184382 117813
rect 184340 117762 184396 117771
rect 184340 117697 184396 117706
rect 184450 117031 184478 117887
rect 184436 117022 184492 117031
rect 184436 116957 184492 116966
rect 184546 116291 184574 117961
rect 184532 116282 184588 116291
rect 184532 116217 184588 116226
rect 184642 115403 184670 118035
rect 184628 115394 184684 115403
rect 184628 115329 184684 115338
rect 184534 115207 184586 115213
rect 184534 115149 184586 115155
rect 184438 115133 184490 115139
rect 184438 115075 184490 115081
rect 184342 115059 184394 115065
rect 184342 115001 184394 115007
rect 184354 114811 184382 115001
rect 184340 114802 184396 114811
rect 184340 114737 184396 114746
rect 184450 113923 184478 115075
rect 184436 113914 184492 113923
rect 184436 113849 184492 113858
rect 184546 113183 184574 115149
rect 184630 114393 184682 114399
rect 184630 114335 184682 114341
rect 184532 113174 184588 113183
rect 184532 113109 184588 113118
rect 184642 112443 184670 114335
rect 184628 112434 184684 112443
rect 184628 112369 184684 112378
rect 184342 112321 184394 112327
rect 184342 112263 184394 112269
rect 184354 111703 184382 112263
rect 184534 112247 184586 112253
rect 184534 112189 184586 112195
rect 184438 112173 184490 112179
rect 184438 112115 184490 112121
rect 184340 111694 184396 111703
rect 184340 111629 184396 111638
rect 184450 110963 184478 112115
rect 184436 110954 184492 110963
rect 184436 110889 184492 110898
rect 184546 110223 184574 112189
rect 184532 110214 184588 110223
rect 184532 110149 184588 110158
rect 184438 109435 184490 109441
rect 184438 109377 184490 109383
rect 184342 109361 184394 109367
rect 184340 109326 184342 109335
rect 184394 109326 184396 109335
rect 184340 109261 184396 109270
rect 184450 107115 184478 109377
rect 185698 108743 185726 129579
rect 186742 129563 186794 129569
rect 186742 129505 186794 129511
rect 186754 129167 186782 129505
rect 186740 129158 186796 129167
rect 186740 129093 186796 129102
rect 645730 129019 645758 129579
rect 645716 129010 645772 129019
rect 645716 128945 645772 128954
rect 646498 126905 646526 275317
rect 647362 269323 647390 278018
rect 648610 272135 648638 278018
rect 648596 272126 648652 272135
rect 648596 272061 648652 272070
rect 647348 269314 647404 269323
rect 647348 269249 647404 269258
rect 646580 267094 646636 267103
rect 646580 267029 646636 267038
rect 646486 126899 646538 126905
rect 646486 126841 646538 126847
rect 186166 122459 186218 122465
rect 186166 122401 186218 122407
rect 185684 108734 185740 108743
rect 185684 108669 185740 108678
rect 186178 107855 186206 122401
rect 646498 122063 646526 126841
rect 646594 126831 646622 267029
rect 646678 253513 646730 253519
rect 646678 253455 646730 253461
rect 646690 144263 646718 253455
rect 646774 207411 646826 207417
rect 646774 207353 646826 207359
rect 646676 144254 646732 144263
rect 646676 144189 646732 144198
rect 646786 141007 646814 207353
rect 649378 183145 649406 861106
rect 655126 792085 655178 792091
rect 655126 792027 655178 792033
rect 654358 780541 654410 780547
rect 654358 780483 654410 780489
rect 654370 773559 654398 780483
rect 655138 775927 655166 792027
rect 656566 783427 656618 783433
rect 656566 783369 656618 783375
rect 655412 778286 655468 778295
rect 655412 778221 655468 778230
rect 655220 777694 655276 777703
rect 655220 777629 655276 777638
rect 655124 775918 655180 775927
rect 655124 775853 655180 775862
rect 654356 773550 654412 773559
rect 654356 773485 654412 773494
rect 654070 737473 654122 737479
rect 654070 737415 654122 737421
rect 654082 728567 654110 737415
rect 654166 737399 654218 737405
rect 654166 737341 654218 737347
rect 654178 730195 654206 737341
rect 655124 734478 655180 734487
rect 655124 734413 655180 734422
rect 654164 730186 654220 730195
rect 654164 730121 654220 730130
rect 654068 728558 654124 728567
rect 654068 728493 654124 728502
rect 654742 702841 654794 702847
rect 654742 702783 654794 702789
rect 649462 702767 649514 702773
rect 649462 702709 649514 702715
rect 649366 183139 649418 183145
rect 649366 183081 649418 183087
rect 649474 179445 649502 702709
rect 654166 694183 654218 694189
rect 654166 694125 654218 694131
rect 654070 691297 654122 691303
rect 654070 691239 654122 691245
rect 654082 684611 654110 691239
rect 654178 685351 654206 694125
rect 654754 686979 654782 702783
rect 654740 686970 654796 686979
rect 654740 686905 654796 686914
rect 654164 685342 654220 685351
rect 654164 685277 654220 685286
rect 654068 684602 654124 684611
rect 654068 684537 654124 684546
rect 655138 668215 655166 734413
rect 655234 714465 655262 777629
rect 655316 731666 655372 731675
rect 655316 731601 655372 731610
rect 655222 714459 655274 714465
rect 655222 714401 655274 714407
rect 655220 689486 655276 689495
rect 655220 689421 655276 689430
rect 655126 668209 655178 668215
rect 655126 668151 655178 668157
rect 652246 666803 652298 666809
rect 652246 666745 652298 666751
rect 649750 666729 649802 666735
rect 649750 666671 649802 666677
rect 649558 656739 649610 656745
rect 649558 656681 649610 656687
rect 649462 179439 649514 179445
rect 649462 179381 649514 179387
rect 649570 174931 649598 656681
rect 649654 610637 649706 610643
rect 649654 610579 649706 610585
rect 649558 174925 649610 174931
rect 649558 174867 649610 174873
rect 649666 171083 649694 610579
rect 649762 263551 649790 666671
rect 649846 564535 649898 564541
rect 649846 564477 649898 564483
rect 649748 263542 649804 263551
rect 649748 263477 649804 263486
rect 649654 171077 649706 171083
rect 649654 171019 649706 171025
rect 649858 168271 649886 564477
rect 649942 521319 649994 521325
rect 649942 521261 649994 521267
rect 649846 168265 649898 168271
rect 649846 168207 649898 168213
rect 647062 164343 647114 164349
rect 647062 164285 647114 164291
rect 646966 164269 647018 164275
rect 646966 164211 647018 164217
rect 646870 164195 646922 164201
rect 646870 164137 646922 164143
rect 646772 140998 646828 141007
rect 646772 140933 646828 140942
rect 646582 126825 646634 126831
rect 646582 126767 646634 126773
rect 646594 123839 646622 126767
rect 646882 125763 646910 164137
rect 646978 127687 647006 164211
rect 647074 134791 647102 164285
rect 649954 163387 649982 521261
rect 650038 478177 650090 478183
rect 650038 478119 650090 478125
rect 649942 163381 649994 163387
rect 649942 163323 649994 163329
rect 650050 159761 650078 478119
rect 650134 388859 650186 388865
rect 650134 388801 650186 388807
rect 650038 159755 650090 159761
rect 650038 159697 650090 159703
rect 650146 156061 650174 388801
rect 650230 345865 650282 345871
rect 650230 345807 650282 345813
rect 650134 156055 650186 156061
rect 650134 155997 650186 156003
rect 650242 152583 650270 345807
rect 650326 299615 650378 299621
rect 650326 299557 650378 299563
rect 650230 152577 650282 152583
rect 650230 152519 650282 152525
rect 650338 148217 650366 299557
rect 652258 266955 652286 666745
rect 654166 656813 654218 656819
rect 654166 656755 654218 656761
rect 654178 640655 654206 656755
rect 655124 642422 655180 642431
rect 655124 642357 655180 642366
rect 654164 640646 654220 640655
rect 654164 640581 654220 640590
rect 653974 602053 654026 602059
rect 653974 601995 654026 602001
rect 653986 594183 654014 601995
rect 653972 594174 654028 594183
rect 653972 594109 654028 594118
rect 655138 576381 655166 642357
rect 655234 622409 655262 689421
rect 655330 668437 655358 731601
rect 655426 714613 655454 778221
rect 655604 776066 655660 776075
rect 655604 776001 655660 776010
rect 655508 732702 655564 732711
rect 655508 732637 655564 732646
rect 655414 714607 655466 714613
rect 655414 714549 655466 714555
rect 655412 687118 655468 687127
rect 655412 687053 655468 687062
rect 655318 668431 655370 668437
rect 655318 668373 655370 668379
rect 655316 643014 655372 643023
rect 655316 642949 655372 642958
rect 655222 622403 655274 622409
rect 655222 622345 655274 622351
rect 655220 597874 655276 597883
rect 655220 597809 655276 597818
rect 655126 576375 655178 576381
rect 655126 576317 655178 576323
rect 654166 555877 654218 555883
rect 654166 555819 654218 555825
rect 654178 548599 654206 555819
rect 655124 553326 655180 553335
rect 655124 553261 655180 553270
rect 654164 548590 654220 548599
rect 654164 548525 654220 548534
rect 655138 489801 655166 553261
rect 655234 533165 655262 597809
rect 655330 576529 655358 642949
rect 655426 622557 655454 687053
rect 655522 668585 655550 732637
rect 655618 714761 655646 776001
rect 656578 774743 656606 783369
rect 656564 774734 656620 774743
rect 656564 774669 656620 774678
rect 655702 748869 655754 748875
rect 655702 748811 655754 748817
rect 655714 731379 655742 748811
rect 655700 731370 655756 731379
rect 655700 731305 655756 731314
rect 655606 714755 655658 714761
rect 655606 714697 655658 714703
rect 669718 713127 669770 713133
rect 669718 713069 669770 713075
rect 669526 711943 669578 711949
rect 669526 711885 669578 711891
rect 655604 688450 655660 688459
rect 655604 688385 655660 688394
rect 655510 668579 655562 668585
rect 655510 668521 655562 668527
rect 655508 640794 655564 640803
rect 655508 640729 655564 640738
rect 655414 622551 655466 622557
rect 655414 622493 655466 622499
rect 655412 596690 655468 596699
rect 655412 596625 655468 596634
rect 655318 576523 655370 576529
rect 655318 576465 655370 576471
rect 655316 550958 655372 550967
rect 655316 550893 655372 550902
rect 655222 533159 655274 533165
rect 655222 533101 655274 533107
rect 655330 489949 655358 550893
rect 655426 533313 655454 596625
rect 655522 576677 655550 640729
rect 655618 624999 655646 688385
rect 655798 648229 655850 648235
rect 655798 648171 655850 648177
rect 655810 639175 655838 648171
rect 655990 645195 656042 645201
rect 655990 645137 656042 645143
rect 655796 639166 655852 639175
rect 655796 639101 655852 639110
rect 656002 638287 656030 645137
rect 655988 638278 656044 638287
rect 655988 638213 656044 638222
rect 655606 624993 655658 624999
rect 655606 624935 655658 624941
rect 655798 613523 655850 613529
rect 655798 613465 655850 613471
rect 655604 595506 655660 595515
rect 655604 595441 655660 595450
rect 655510 576671 655562 576677
rect 655510 576613 655562 576619
rect 655508 552142 655564 552151
rect 655508 552077 655564 552086
rect 655414 533307 655466 533313
rect 655414 533249 655466 533255
rect 655522 490097 655550 552077
rect 655618 533461 655646 595441
rect 655810 595367 655838 613465
rect 656566 602127 656618 602133
rect 656566 602069 656618 602075
rect 655796 595358 655852 595367
rect 655796 595293 655852 595302
rect 656578 592999 656606 602069
rect 656564 592990 656620 592999
rect 656564 592925 656620 592934
rect 655702 567495 655754 567501
rect 655702 567437 655754 567443
rect 655714 550819 655742 567437
rect 656566 558837 656618 558843
rect 656566 558779 656618 558785
rect 655700 550810 655756 550819
rect 655700 550745 655756 550754
rect 656578 549783 656606 558779
rect 656564 549774 656620 549783
rect 656564 549709 656620 549718
rect 655606 533455 655658 533461
rect 655606 533397 655658 533403
rect 655510 490091 655562 490097
rect 655510 490033 655562 490039
rect 655318 489943 655370 489949
rect 655318 489885 655370 489891
rect 655126 489795 655178 489801
rect 655126 489737 655178 489743
rect 655510 400551 655562 400557
rect 655510 400493 655562 400499
rect 655318 400477 655370 400483
rect 655318 400419 655370 400425
rect 655126 400403 655178 400409
rect 655126 400345 655178 400351
rect 655138 373367 655166 400345
rect 655330 374403 655358 400419
rect 655316 374394 655372 374403
rect 655316 374329 655372 374338
rect 655124 373358 655180 373367
rect 655124 373293 655180 373302
rect 655522 372183 655550 400493
rect 656566 381607 656618 381613
rect 656566 381549 656618 381555
rect 655508 372174 655564 372183
rect 655508 372109 655564 372118
rect 656578 370999 656606 381549
rect 656564 370990 656620 370999
rect 656564 370925 656620 370934
rect 655318 357335 655370 357341
rect 655318 357277 655370 357283
rect 655222 357261 655274 357267
rect 655222 357203 655274 357209
rect 655126 357187 655178 357193
rect 655126 357129 655178 357135
rect 654166 328327 654218 328333
rect 654166 328269 654218 328275
rect 654178 326303 654206 328269
rect 655138 327487 655166 357129
rect 655234 329855 655262 357203
rect 655220 329846 655276 329855
rect 655220 329781 655276 329790
rect 655330 328079 655358 357277
rect 667798 340685 667850 340691
rect 667798 340627 667850 340633
rect 667810 328333 667838 340627
rect 667798 328327 667850 328333
rect 667798 328269 667850 328275
rect 655316 328070 655372 328079
rect 655316 328005 655372 328014
rect 655124 327478 655180 327487
rect 655124 327413 655180 327422
rect 654164 326294 654220 326303
rect 654164 326229 654220 326238
rect 654262 311233 654314 311239
rect 654262 311175 654314 311181
rect 654166 311159 654218 311165
rect 654166 311101 654218 311107
rect 654070 311085 654122 311091
rect 654070 311027 654122 311033
rect 654082 302179 654110 311027
rect 654178 303363 654206 311101
rect 654164 303354 654220 303363
rect 654164 303289 654220 303298
rect 654068 302170 654124 302179
rect 654068 302105 654124 302114
rect 654274 300995 654302 311175
rect 654260 300986 654316 300995
rect 654260 300921 654316 300930
rect 656564 298766 656620 298775
rect 656564 298701 656620 298710
rect 656276 297582 656332 297591
rect 656276 297517 656332 297526
rect 656084 296842 656140 296851
rect 656084 296777 656140 296786
rect 655892 294030 655948 294039
rect 655892 293965 655948 293974
rect 655796 292846 655852 292855
rect 655796 292781 655852 292790
rect 655604 289294 655660 289303
rect 655604 289229 655660 289238
rect 655412 288110 655468 288119
rect 655412 288045 655468 288054
rect 653780 284558 653836 284567
rect 653780 284493 653836 284502
rect 653794 284303 653822 284493
rect 653782 284297 653834 284303
rect 653782 284239 653834 284245
rect 655124 283374 655180 283383
rect 655124 283309 655180 283318
rect 654164 279822 654220 279831
rect 654164 279757 654220 279766
rect 654178 279493 654206 279757
rect 654166 279487 654218 279493
rect 654166 279429 654218 279435
rect 652244 266946 652300 266955
rect 652244 266881 652300 266890
rect 650326 148211 650378 148217
rect 650326 148153 650378 148159
rect 647060 134782 647116 134791
rect 647060 134717 647116 134726
rect 647828 130934 647884 130943
rect 647828 130869 647884 130878
rect 646964 127678 647020 127687
rect 646964 127613 647020 127622
rect 646868 125754 646924 125763
rect 646868 125689 646924 125698
rect 646580 123830 646636 123839
rect 646580 123765 646636 123774
rect 646484 122054 646540 122063
rect 646484 121989 646540 121998
rect 647842 118395 647870 130869
rect 655138 129865 655166 283309
rect 655316 282338 655372 282347
rect 655316 282273 655372 282282
rect 655220 281006 655276 281015
rect 655220 280941 655276 280950
rect 655234 130013 655262 280941
rect 655330 130161 655358 282273
rect 655426 175893 655454 288045
rect 655508 285742 655564 285751
rect 655508 285677 655564 285686
rect 655522 176041 655550 285677
rect 655618 201571 655646 289229
rect 655700 286926 655756 286935
rect 655700 286861 655756 286870
rect 655606 201565 655658 201571
rect 655606 201507 655658 201513
rect 655714 176189 655742 286861
rect 655810 219109 655838 292781
rect 655906 247673 655934 293965
rect 655988 290922 656044 290931
rect 655988 290857 656044 290866
rect 655894 247667 655946 247673
rect 655894 247609 655946 247615
rect 656002 219257 656030 290857
rect 656098 265137 656126 296777
rect 656180 291662 656236 291671
rect 656180 291597 656236 291606
rect 656086 265131 656138 265137
rect 656086 265073 656138 265079
rect 656194 221847 656222 291597
rect 656290 265285 656318 297517
rect 656372 295214 656428 295223
rect 656372 295149 656428 295158
rect 656386 290464 656414 295149
rect 656578 290889 656606 298701
rect 656566 290883 656618 290889
rect 656566 290825 656618 290831
rect 656386 290436 656606 290464
rect 656578 265433 656606 290436
rect 658006 284297 658058 284303
rect 658006 284239 658058 284245
rect 656566 265427 656618 265433
rect 656566 265369 656618 265375
rect 656278 265279 656330 265285
rect 656278 265221 656330 265227
rect 656182 221841 656234 221847
rect 656182 221783 656234 221789
rect 655990 219251 656042 219257
rect 655990 219193 656042 219199
rect 655798 219103 655850 219109
rect 655798 219045 655850 219051
rect 655702 176183 655754 176189
rect 655702 176125 655754 176131
rect 655510 176035 655562 176041
rect 655510 175977 655562 175983
rect 655414 175887 655466 175893
rect 655414 175829 655466 175835
rect 658018 155543 658046 284239
rect 663766 279487 663818 279493
rect 663766 279429 663818 279435
rect 658006 155537 658058 155543
rect 658006 155479 658058 155485
rect 655318 130155 655370 130161
rect 655318 130097 655370 130103
rect 655222 130007 655274 130013
rect 655222 129949 655274 129955
rect 655126 129859 655178 129865
rect 655126 129801 655178 129807
rect 647924 119538 647980 119547
rect 647924 119473 647980 119482
rect 647830 118389 647882 118395
rect 647830 118331 647882 118337
rect 647938 118247 647966 119473
rect 647926 118241 647978 118247
rect 647926 118183 647978 118189
rect 645238 118167 645290 118173
rect 645238 118109 645290 118115
rect 645250 117623 645278 118109
rect 645236 117614 645292 117623
rect 645236 117549 645292 117558
rect 647924 115690 647980 115699
rect 647924 115625 647980 115634
rect 647938 115287 647966 115625
rect 647926 115281 647978 115287
rect 647926 115223 647978 115229
rect 663778 115213 663806 279429
rect 669538 275495 669566 711885
rect 669622 623143 669674 623149
rect 669622 623085 669674 623091
rect 669524 275486 669580 275495
rect 669524 275421 669580 275430
rect 669634 264915 669662 623085
rect 669730 275643 669758 713069
rect 670678 712683 670730 712689
rect 670678 712625 670730 712631
rect 670582 711573 670634 711579
rect 670582 711515 670634 711521
rect 670594 666809 670622 711515
rect 670690 668067 670718 712625
rect 670882 711949 670910 890373
rect 670978 713133 671006 891409
rect 673654 737917 673706 737923
rect 673654 737859 673706 737865
rect 673462 733773 673514 733779
rect 673462 733715 673514 733721
rect 670966 713127 671018 713133
rect 670966 713069 671018 713075
rect 670870 711943 670922 711949
rect 670870 711885 670922 711891
rect 670774 699881 670826 699887
rect 670774 699823 670826 699829
rect 670786 669251 670814 699823
rect 670774 669245 670826 669251
rect 670774 669187 670826 669193
rect 670678 668061 670730 668067
rect 670678 668003 670730 668009
rect 670582 666803 670634 666809
rect 670582 666745 670634 666751
rect 670690 666735 670718 668003
rect 670870 667691 670922 667697
rect 670870 667633 670922 667639
rect 670678 666729 670730 666735
rect 670678 666671 670730 666677
rect 670882 623149 670910 667633
rect 670966 666359 671018 666365
rect 670966 666301 671018 666307
rect 670870 623143 670922 623149
rect 670870 623085 670922 623091
rect 670774 622477 670826 622483
rect 670774 622419 670826 622425
rect 669814 620035 669866 620041
rect 669814 619977 669866 619983
rect 669716 275634 669772 275643
rect 669716 275569 669772 275578
rect 669826 264989 669854 619977
rect 670786 575937 670814 622419
rect 670978 621965 671006 666301
rect 673474 659927 673502 733715
rect 673558 688781 673610 688787
rect 673558 688723 673610 688729
rect 673462 659921 673514 659927
rect 673462 659863 673514 659869
rect 673078 644603 673130 644609
rect 673078 644545 673130 644551
rect 672790 623439 672842 623445
rect 672790 623381 672842 623387
rect 670966 621959 671018 621965
rect 670966 621901 671018 621907
rect 670870 621367 670922 621373
rect 670870 621309 670922 621315
rect 670774 575931 670826 575937
rect 670774 575873 670826 575879
rect 669910 573267 669962 573273
rect 669910 573209 669962 573215
rect 669922 277907 669950 573209
rect 670786 573199 670814 575873
rect 670882 574975 670910 621309
rect 670978 620041 671006 621901
rect 670966 620035 671018 620041
rect 670966 619977 671018 619983
rect 672802 590367 672830 623381
rect 672886 598427 672938 598433
rect 672886 598369 672938 598375
rect 672790 590361 672842 590367
rect 672790 590303 672842 590309
rect 672790 576227 672842 576233
rect 672790 576169 672842 576175
rect 672598 575487 672650 575493
rect 672598 575429 672650 575435
rect 670870 574969 670922 574975
rect 670870 574911 670922 574917
rect 670882 573273 670910 574911
rect 670870 573267 670922 573273
rect 670870 573209 670922 573215
rect 670102 573193 670154 573199
rect 670102 573135 670154 573141
rect 670774 573193 670826 573199
rect 670774 573135 670826 573141
rect 670004 354710 670060 354719
rect 670004 354645 670060 354654
rect 669908 277898 669964 277907
rect 669908 277833 669964 277842
rect 670018 273615 670046 354645
rect 670114 277463 670142 573135
rect 672610 532721 672638 575429
rect 672694 574155 672746 574161
rect 672694 574097 672746 574103
rect 672598 532715 672650 532721
rect 672598 532657 672650 532663
rect 672406 531531 672458 531537
rect 672406 531473 672458 531479
rect 670294 488167 670346 488173
rect 670294 488109 670346 488115
rect 670196 356042 670252 356051
rect 670196 355977 670252 355986
rect 670100 277454 670156 277463
rect 670100 277389 670156 277398
rect 670210 277227 670238 355977
rect 670306 277611 670334 488109
rect 670486 487131 670538 487137
rect 670486 487073 670538 487079
rect 670388 308978 670444 308987
rect 670388 308913 670444 308922
rect 670292 277602 670348 277611
rect 670292 277537 670348 277546
rect 670196 277218 670252 277227
rect 670196 277153 670252 277162
rect 670402 277079 670430 308913
rect 670498 277759 670526 487073
rect 670966 434961 671018 434967
rect 670966 434903 671018 434909
rect 670978 399077 671006 434903
rect 670966 399071 671018 399077
rect 670966 399013 671018 399019
rect 670978 377294 671006 399013
rect 670690 377266 671006 377294
rect 670690 278055 670718 377266
rect 672418 278647 672446 531473
rect 672502 486835 672554 486841
rect 672502 486777 672554 486783
rect 672514 434967 672542 486777
rect 672502 434961 672554 434967
rect 672502 434903 672554 434909
rect 672502 400329 672554 400335
rect 672502 400271 672554 400277
rect 672404 278638 672460 278647
rect 672404 278573 672460 278582
rect 670676 278046 670732 278055
rect 670676 277981 670732 277990
rect 670484 277750 670540 277759
rect 670484 277685 670540 277694
rect 670388 277070 670444 277079
rect 670388 277005 670444 277014
rect 670004 273606 670060 273615
rect 670004 273541 670060 273550
rect 672514 273467 672542 400271
rect 672610 278203 672638 532657
rect 672706 531537 672734 574097
rect 672802 547225 672830 576169
rect 672790 547219 672842 547225
rect 672790 547161 672842 547167
rect 672694 531531 672746 531537
rect 672694 531473 672746 531479
rect 672898 524507 672926 598369
rect 672982 596577 673034 596583
rect 672982 596519 673034 596525
rect 672994 526357 673022 596519
rect 673090 568019 673118 644545
rect 673270 643937 673322 643943
rect 673270 643879 673322 643885
rect 673174 643419 673226 643425
rect 673174 643361 673226 643367
rect 673078 568013 673130 568019
rect 673078 567955 673130 567961
rect 673186 567723 673214 643361
rect 673282 569203 673310 643879
rect 673366 642309 673418 642315
rect 673366 642251 673418 642257
rect 673378 569573 673406 642251
rect 673570 614491 673598 688723
rect 673666 660667 673694 737859
rect 673858 722975 673886 892371
rect 676052 891506 676108 891515
rect 676052 891441 676054 891450
rect 676106 891441 676108 891450
rect 676054 891409 676106 891415
rect 676052 890470 676108 890479
rect 676052 890405 676054 890414
rect 676106 890405 676108 890414
rect 676054 890373 676106 890379
rect 680180 890174 680236 890183
rect 680180 890109 680236 890118
rect 676244 889286 676300 889295
rect 676244 889221 676300 889230
rect 676258 887921 676286 889221
rect 679988 888694 680044 888703
rect 679988 888629 680044 888638
rect 674038 887915 674090 887921
rect 674038 887857 674090 887863
rect 676246 887915 676298 887921
rect 676246 887857 676298 887863
rect 674050 876303 674078 887857
rect 676244 887806 676300 887815
rect 676244 887741 676300 887750
rect 676052 887436 676108 887445
rect 676052 887371 676108 887380
rect 676066 887181 676094 887371
rect 674230 887175 674282 887181
rect 674230 887117 674282 887123
rect 676054 887175 676106 887181
rect 676054 887117 676106 887123
rect 674134 885103 674186 885109
rect 674134 885045 674186 885051
rect 674038 876297 674090 876303
rect 674038 876239 674090 876245
rect 674146 867423 674174 885045
rect 674242 876451 674270 887117
rect 676258 887107 676286 887741
rect 674422 887101 674474 887107
rect 674422 887043 674474 887049
rect 676246 887101 676298 887107
rect 676246 887043 676298 887049
rect 674326 884289 674378 884295
rect 674326 884231 674378 884237
rect 674230 876445 674282 876451
rect 674230 876387 674282 876393
rect 674230 876297 674282 876303
rect 674230 876239 674282 876245
rect 674134 867417 674186 867423
rect 674134 867359 674186 867365
rect 674242 865795 674270 876239
rect 674338 869791 674366 884231
rect 674434 876544 674462 887043
rect 679700 886770 679756 886779
rect 679700 886705 679756 886714
rect 676052 885512 676108 885521
rect 676052 885447 676108 885456
rect 676066 885109 676094 885447
rect 676054 885103 676106 885109
rect 676054 885045 676106 885051
rect 676052 884994 676108 885003
rect 676052 884929 676108 884938
rect 676066 884295 676094 884929
rect 676054 884289 676106 884295
rect 676054 884231 676106 884237
rect 676244 884254 676300 884263
rect 674902 884215 674954 884221
rect 676244 884189 676246 884198
rect 674902 884157 674954 884163
rect 676298 884189 676300 884198
rect 676246 884157 676298 884163
rect 674518 883105 674570 883111
rect 674518 883047 674570 883053
rect 674530 876673 674558 883047
rect 674710 881551 674762 881557
rect 674710 881493 674762 881499
rect 674614 881255 674666 881261
rect 674614 881197 674666 881203
rect 674626 876747 674654 881197
rect 674614 876741 674666 876747
rect 674614 876683 674666 876689
rect 674518 876667 674570 876673
rect 674518 876609 674570 876615
rect 674434 876516 674654 876544
rect 674518 876445 674570 876451
rect 674518 876387 674570 876393
rect 674326 869785 674378 869791
rect 674326 869727 674378 869733
rect 674530 869717 674558 876387
rect 674626 870605 674654 876516
rect 674722 872973 674750 881493
rect 674806 881329 674858 881335
rect 674806 881271 674858 881277
rect 674818 873047 674846 881271
rect 674914 873140 674942 884157
rect 676052 884032 676108 884041
rect 676052 883967 676108 883976
rect 675956 883514 676012 883523
rect 675956 883449 676012 883458
rect 675286 883253 675338 883259
rect 675286 883195 675338 883201
rect 674998 882883 675050 882889
rect 674998 882825 675050 882831
rect 675010 877265 675038 882825
rect 675190 880145 675242 880151
rect 675190 880087 675242 880093
rect 675094 877999 675146 878005
rect 675094 877941 675146 877947
rect 674998 877259 675050 877265
rect 674998 877201 675050 877207
rect 675106 873214 675134 877941
rect 675202 873880 675230 880087
rect 675298 877537 675326 883195
rect 675970 881557 675998 883449
rect 675958 881551 676010 881557
rect 675958 881493 676010 881499
rect 675478 881403 675530 881409
rect 675478 881345 675530 881351
rect 675490 878084 675518 881345
rect 676066 881335 676094 883967
rect 679714 882889 679742 886705
rect 679796 886178 679852 886187
rect 679796 886113 679852 886122
rect 679702 882883 679754 882889
rect 679702 882825 679754 882831
rect 679700 882774 679756 882783
rect 679700 882709 679756 882718
rect 679714 882191 679742 882709
rect 679700 882182 679756 882191
rect 679700 882117 679756 882126
rect 679714 881483 679742 882117
rect 679702 881477 679754 881483
rect 679702 881419 679754 881425
rect 676054 881329 676106 881335
rect 676054 881271 676106 881277
rect 679810 880151 679838 886113
rect 679892 885734 679948 885743
rect 679892 885669 679948 885678
rect 679798 880145 679850 880151
rect 679798 880087 679850 880093
rect 679906 878523 679934 885669
rect 680002 883259 680030 888629
rect 680084 888250 680140 888259
rect 680084 888185 680140 888194
rect 679990 883253 680042 883259
rect 679990 883195 680042 883201
rect 680098 881261 680126 888185
rect 680194 883111 680222 890109
rect 680182 883105 680234 883111
rect 680182 883047 680234 883053
rect 685460 882182 685516 882191
rect 685460 882117 685516 882126
rect 685474 881747 685502 882117
rect 685460 881738 685516 881747
rect 685460 881673 685516 881682
rect 680086 881255 680138 881261
rect 680086 881197 680138 881203
rect 679894 878517 679946 878523
rect 679894 878459 679946 878465
rect 675298 877509 675408 877537
rect 675478 877259 675530 877265
rect 675478 877201 675530 877207
rect 675490 876900 675518 877201
rect 675286 876741 675338 876747
rect 675286 876683 675338 876689
rect 675298 874398 675326 876683
rect 675382 876667 675434 876673
rect 675382 876609 675434 876615
rect 675394 876234 675422 876609
rect 675298 874370 675408 874398
rect 675202 873852 675326 873880
rect 675298 873732 675326 873852
rect 675394 873732 675422 873866
rect 675298 873704 675422 873732
rect 675106 873186 675408 873214
rect 674914 873112 675422 873140
rect 674806 873041 674858 873047
rect 674806 872983 674858 872989
rect 675286 873041 675338 873047
rect 675286 872983 675338 872989
rect 674710 872967 674762 872973
rect 674710 872909 674762 872915
rect 675190 872967 675242 872973
rect 675190 872909 675242 872915
rect 675094 872671 675146 872677
rect 675094 872613 675146 872619
rect 674614 870599 674666 870605
rect 674614 870541 674666 870547
rect 674518 869711 674570 869717
rect 674518 869653 674570 869659
rect 674998 869711 675050 869717
rect 674998 869653 675050 869659
rect 674230 865789 674282 865795
rect 674230 865731 674282 865737
rect 675010 863372 675038 869653
rect 675106 867693 675134 872613
rect 675202 868256 675230 872909
rect 675298 869884 675326 872983
rect 675394 872534 675422 873112
rect 675478 870599 675530 870605
rect 675478 870541 675530 870547
rect 675490 870092 675518 870541
rect 675298 869856 675422 869884
rect 675286 869785 675338 869791
rect 675286 869727 675338 869733
rect 675298 868889 675326 869727
rect 675394 869500 675422 869856
rect 675298 868861 675408 868889
rect 675202 868228 675408 868256
rect 675106 867665 675408 867693
rect 675478 867417 675530 867423
rect 675478 867359 675530 867365
rect 675490 867058 675518 867359
rect 675106 865825 675408 865853
rect 675106 864019 675134 865825
rect 675190 865789 675242 865795
rect 675190 865731 675242 865737
rect 675202 865222 675230 865731
rect 675202 865194 675408 865222
rect 675094 864013 675146 864019
rect 675094 863955 675146 863961
rect 675010 863344 675408 863372
rect 675382 792085 675434 792091
rect 675382 792027 675434 792033
rect 675394 788875 675422 792027
rect 675092 788350 675148 788359
rect 675148 788308 675408 788336
rect 675092 788285 675148 788294
rect 675490 787175 675518 787656
rect 675476 787166 675532 787175
rect 675476 787101 675532 787110
rect 675106 787021 675408 787049
rect 675106 786287 675134 787021
rect 675092 786278 675148 786287
rect 675092 786213 675148 786222
rect 675394 784807 675422 785214
rect 675380 784798 675436 784807
rect 675380 784733 675436 784742
rect 675490 784363 675518 784622
rect 675476 784354 675532 784363
rect 675476 784289 675532 784298
rect 675106 783985 675408 784013
rect 675106 783475 675134 783985
rect 675092 783466 675148 783475
rect 675092 783401 675148 783410
rect 675190 783427 675242 783433
rect 675190 783369 675242 783375
rect 675094 780541 675146 780547
rect 675094 780483 675146 780489
rect 674902 778617 674954 778623
rect 674902 778559 674954 778565
rect 674806 777359 674858 777365
rect 674806 777301 674858 777307
rect 674326 774325 674378 774331
rect 674326 774267 674378 774273
rect 674230 732367 674282 732373
rect 674230 732309 674282 732315
rect 673846 722969 673898 722975
rect 673846 722911 673898 722917
rect 673750 692925 673802 692931
rect 673750 692867 673802 692873
rect 673654 660661 673706 660667
rect 673654 660603 673706 660609
rect 673762 615675 673790 692867
rect 674242 662369 674270 732309
rect 674338 711357 674366 774267
rect 674422 767147 674474 767153
rect 674422 767089 674474 767095
rect 674326 711351 674378 711357
rect 674326 711293 674378 711299
rect 674434 710543 674462 767089
rect 674710 742801 674762 742807
rect 674710 742743 674762 742749
rect 674722 734339 674750 742743
rect 674708 734330 674764 734339
rect 674708 734265 674764 734274
rect 674710 730517 674762 730523
rect 674710 730459 674762 730465
rect 674614 728667 674666 728673
rect 674614 728609 674666 728615
rect 674422 710537 674474 710543
rect 674422 710479 674474 710485
rect 674326 686783 674378 686789
rect 674326 686725 674378 686731
rect 674230 662363 674282 662369
rect 674230 662305 674282 662311
rect 673846 648081 673898 648087
rect 673846 648023 673898 648029
rect 673750 615669 673802 615675
rect 673750 615611 673802 615617
rect 673558 614485 673610 614491
rect 673558 614427 673610 614433
rect 673750 603311 673802 603317
rect 673750 603253 673802 603259
rect 673654 602719 673706 602725
rect 673654 602661 673706 602667
rect 673462 599833 673514 599839
rect 673462 599775 673514 599781
rect 673366 569567 673418 569573
rect 673366 569509 673418 569515
rect 673270 569197 673322 569203
rect 673270 569139 673322 569145
rect 673174 567717 673226 567723
rect 673174 567659 673226 567665
rect 672982 526351 673034 526357
rect 672982 526293 673034 526299
rect 673474 524877 673502 599775
rect 673558 599315 673610 599321
rect 673558 599257 673610 599263
rect 673570 525987 673598 599257
rect 673558 525981 673610 525987
rect 673558 525923 673610 525929
rect 673666 525247 673694 602661
rect 673762 526727 673790 603253
rect 673858 568463 673886 648023
rect 674230 639127 674282 639133
rect 674230 639069 674282 639075
rect 674134 629137 674186 629143
rect 674134 629079 674186 629085
rect 674146 573125 674174 629079
rect 674242 576011 674270 639069
rect 674338 618635 674366 686725
rect 674422 683675 674474 683681
rect 674422 683617 674474 683623
rect 674434 618857 674462 683617
rect 674518 682861 674570 682867
rect 674518 682803 674570 682809
rect 674530 622039 674558 682803
rect 674626 665181 674654 728609
rect 674722 668141 674750 730459
rect 674818 708101 674846 777301
rect 674914 708397 674942 778559
rect 675106 776644 675134 780483
rect 675202 778494 675230 783369
rect 675778 783031 675806 783364
rect 675764 783022 675820 783031
rect 675764 782957 675820 782966
rect 675778 780663 675806 780848
rect 675764 780654 675820 780663
rect 675764 780589 675820 780598
rect 675778 780071 675806 780330
rect 675764 780062 675820 780071
rect 675764 779997 675820 780006
rect 675298 779650 675408 779678
rect 675298 778623 675326 779650
rect 675778 778887 675806 779031
rect 675764 778878 675820 778887
rect 675764 778813 675820 778822
rect 675286 778617 675338 778623
rect 675286 778559 675338 778565
rect 675202 778466 675408 778494
rect 675490 777365 675518 777814
rect 675478 777359 675530 777365
rect 675478 777301 675530 777307
rect 675106 776616 675408 776644
rect 675106 775981 675408 776009
rect 675106 774331 675134 775981
rect 675094 774325 675146 774331
rect 675094 774267 675146 774273
rect 675106 774141 675408 774169
rect 675106 767153 675134 774141
rect 675284 771922 675340 771931
rect 675284 771857 675340 771866
rect 675094 767147 675146 767153
rect 675094 767089 675146 767095
rect 675298 751694 675326 771857
rect 675202 751666 675326 751694
rect 674998 737473 675050 737479
rect 674998 737415 675050 737421
rect 675010 732077 675038 737415
rect 675094 737399 675146 737405
rect 675094 737341 675146 737347
rect 675106 733927 675134 737341
rect 675202 735777 675230 751666
rect 675382 748869 675434 748875
rect 675382 748811 675434 748817
rect 675394 743848 675422 748811
rect 675394 742807 675422 743330
rect 675382 742801 675434 742807
rect 675382 742743 675434 742749
rect 675490 742479 675518 742664
rect 675476 742470 675532 742479
rect 675476 742405 675532 742414
rect 675682 741739 675710 742035
rect 675668 741730 675724 741739
rect 675668 741665 675724 741674
rect 675394 740111 675422 740222
rect 675380 740102 675436 740111
rect 675380 740037 675436 740046
rect 675778 739223 675806 739630
rect 675764 739214 675820 739223
rect 675764 739149 675820 739158
rect 675394 738631 675422 738999
rect 675380 738622 675436 738631
rect 675380 738557 675436 738566
rect 675394 737923 675422 738372
rect 675382 737917 675434 737923
rect 675382 737859 675434 737865
rect 675190 735771 675242 735777
rect 675190 735713 675242 735719
rect 675490 735648 675518 735856
rect 675202 735620 675518 735648
rect 675094 733921 675146 733927
rect 675094 733863 675146 733869
rect 675202 733724 675230 735620
rect 675286 735549 675338 735555
rect 675286 735491 675338 735497
rect 675106 733696 675230 733724
rect 674998 732071 675050 732077
rect 674998 732013 675050 732019
rect 675106 731534 675134 733696
rect 675010 731506 675134 731534
rect 674902 708391 674954 708397
rect 674902 708333 674954 708339
rect 674806 708095 674858 708101
rect 674806 708037 674858 708043
rect 674902 690483 674954 690489
rect 674902 690425 674954 690431
rect 674806 689151 674858 689157
rect 674806 689093 674858 689099
rect 674710 668135 674762 668141
rect 674710 668077 674762 668083
rect 674614 665175 674666 665181
rect 674614 665117 674666 665123
rect 674518 622033 674570 622039
rect 674518 621975 674570 621981
rect 674422 618851 674474 618857
rect 674422 618793 674474 618799
rect 674326 618629 674378 618635
rect 674326 618571 674378 618577
rect 674818 616341 674846 689093
rect 674914 619079 674942 690425
rect 675010 665255 675038 731506
rect 675298 708471 675326 735491
rect 675778 735079 675806 735338
rect 675764 735070 675820 735079
rect 675764 735005 675820 735014
rect 675490 734487 675518 734672
rect 675476 734478 675532 734487
rect 675476 734413 675532 734422
rect 675382 733921 675434 733927
rect 675382 733863 675434 733869
rect 675394 733576 675422 733863
rect 675490 733779 675518 734006
rect 675478 733773 675530 733779
rect 675478 733715 675530 733721
rect 675394 733548 675518 733576
rect 675490 733488 675518 733548
rect 675490 732373 675518 732822
rect 675478 732367 675530 732373
rect 675478 732309 675530 732315
rect 675382 732071 675434 732077
rect 675382 732013 675434 732019
rect 675394 731638 675422 732013
rect 675490 730523 675518 730972
rect 675478 730517 675530 730523
rect 675478 730459 675530 730465
rect 675394 728673 675422 729155
rect 675382 728667 675434 728673
rect 675382 728609 675434 728615
rect 679702 722969 679754 722975
rect 679702 722911 679754 722917
rect 676340 715534 676396 715543
rect 676340 715469 676396 715478
rect 676148 714942 676204 714951
rect 676148 714877 676204 714886
rect 676162 714613 676190 714877
rect 676244 714794 676300 714803
rect 676244 714729 676246 714738
rect 676298 714729 676300 714738
rect 676246 714697 676298 714703
rect 676150 714607 676202 714613
rect 676150 714549 676202 714555
rect 676354 714465 676382 715469
rect 676342 714459 676394 714465
rect 676342 714401 676394 714407
rect 679714 713915 679742 722911
rect 679700 713906 679756 713915
rect 679700 713841 679756 713850
rect 679700 713314 679756 713323
rect 679700 713249 679756 713258
rect 676052 713166 676108 713175
rect 676052 713101 676054 713110
rect 676106 713101 676108 713110
rect 676054 713069 676106 713075
rect 676052 712722 676108 712731
rect 676052 712657 676054 712666
rect 676106 712657 676108 712666
rect 676054 712625 676106 712631
rect 676244 711982 676300 711991
rect 676244 711917 676246 711926
rect 676298 711917 676300 711926
rect 676246 711885 676298 711891
rect 676052 711612 676108 711621
rect 676052 711547 676054 711556
rect 676106 711547 676108 711556
rect 676054 711515 676106 711521
rect 676054 711351 676106 711357
rect 676054 711293 676106 711299
rect 676066 710659 676094 711293
rect 676052 710650 676108 710659
rect 676052 710585 676108 710594
rect 676054 710537 676106 710543
rect 676054 710479 676106 710485
rect 676066 708587 676094 710479
rect 676052 708578 676108 708587
rect 676052 708513 676108 708522
rect 675286 708465 675338 708471
rect 675286 708407 675338 708413
rect 676054 708465 676106 708471
rect 676054 708407 676106 708413
rect 676066 708217 676094 708407
rect 676246 708391 676298 708397
rect 676246 708333 676298 708339
rect 676052 708208 676108 708217
rect 676052 708143 676108 708152
rect 676054 708095 676106 708101
rect 676054 708037 676106 708043
rect 676066 706737 676094 708037
rect 676052 706728 676108 706737
rect 676052 706663 676108 706672
rect 676258 706367 676286 708333
rect 676244 706358 676300 706367
rect 676244 706293 676300 706302
rect 675382 702841 675434 702847
rect 675382 702783 675434 702789
rect 675394 698856 675422 702783
rect 679714 699887 679742 713249
rect 679988 704434 680044 704443
rect 679988 704369 680044 704378
rect 680002 703407 680030 704369
rect 679796 703398 679852 703407
rect 679796 703333 679852 703342
rect 679988 703398 680044 703407
rect 679988 703333 680044 703342
rect 679810 702963 679838 703333
rect 679796 702954 679852 702963
rect 679796 702889 679852 702898
rect 680002 702773 680030 703333
rect 679990 702767 680042 702773
rect 679990 702709 680042 702715
rect 679702 699881 679754 699887
rect 679702 699823 679754 699829
rect 675394 697931 675422 698338
rect 675380 697922 675436 697931
rect 675380 697857 675436 697866
rect 675106 697658 675408 697686
rect 675106 697191 675134 697658
rect 675092 697182 675148 697191
rect 675092 697117 675148 697126
rect 675106 697043 675408 697049
rect 675092 697034 675408 697043
rect 675148 697021 675408 697034
rect 675092 696969 675148 696978
rect 675778 694971 675806 695195
rect 675764 694962 675820 694971
rect 675764 694897 675820 694906
rect 675092 694666 675148 694675
rect 675148 694624 675408 694652
rect 675092 694601 675148 694610
rect 675286 694183 675338 694189
rect 675286 694125 675338 694131
rect 675094 691297 675146 691303
rect 675094 691239 675146 691245
rect 675106 686660 675134 691239
rect 675190 689817 675242 689823
rect 675190 689759 675242 689765
rect 675202 686831 675230 689759
rect 675298 688436 675326 694125
rect 675490 693491 675518 693972
rect 675476 693482 675532 693491
rect 675476 693417 675532 693426
rect 675394 692931 675422 693380
rect 675382 692925 675434 692931
rect 675382 692867 675434 692873
rect 675490 690489 675518 690864
rect 675478 690483 675530 690489
rect 675478 690425 675530 690431
rect 675394 689823 675422 690346
rect 675382 689817 675434 689823
rect 675382 689759 675434 689765
rect 675394 689157 675422 689680
rect 675382 689151 675434 689157
rect 675382 689093 675434 689099
rect 675490 688787 675518 689014
rect 675478 688781 675530 688787
rect 675478 688723 675530 688729
rect 675394 688436 675422 688496
rect 675298 688408 675422 688436
rect 675298 687816 675408 687844
rect 675188 686822 675244 686831
rect 675298 686789 675326 687816
rect 675188 686757 675244 686766
rect 675286 686783 675338 686789
rect 675286 686725 675338 686731
rect 675106 686632 675408 686660
rect 675298 686040 675422 686068
rect 675298 685994 675326 686040
rect 675202 685966 675326 685994
rect 675394 685980 675422 686040
rect 675202 682867 675230 685966
rect 675490 683681 675518 684130
rect 675478 683675 675530 683681
rect 675478 683617 675530 683623
rect 675190 682861 675242 682867
rect 675190 682803 675242 682809
rect 676148 670394 676204 670403
rect 676148 670329 676204 670338
rect 676054 669245 676106 669251
rect 676052 669210 676054 669219
rect 676106 669210 676108 669219
rect 676052 669145 676108 669154
rect 676052 668618 676108 668627
rect 676162 668585 676190 670329
rect 676340 669802 676396 669811
rect 676340 669737 676396 669746
rect 676244 669358 676300 669367
rect 676244 669293 676300 669302
rect 676052 668553 676108 668562
rect 676150 668579 676202 668585
rect 676066 668289 676094 668553
rect 676150 668521 676202 668527
rect 676258 668437 676286 669293
rect 676246 668431 676298 668437
rect 676246 668373 676298 668379
rect 675094 668283 675146 668289
rect 675094 668225 675146 668231
rect 676054 668283 676106 668289
rect 676054 668225 676106 668231
rect 674998 665249 675050 665255
rect 674998 665191 675050 665197
rect 675106 659534 675134 668225
rect 676354 668215 676382 669737
rect 676342 668209 676394 668215
rect 676342 668151 676394 668157
rect 676054 668135 676106 668141
rect 675956 668100 676012 668109
rect 676054 668077 676106 668083
rect 675956 668035 675958 668044
rect 676010 668035 676012 668044
rect 675958 668003 676010 668009
rect 675956 667730 676012 667739
rect 675956 667665 675958 667674
rect 676010 667665 676012 667674
rect 675958 667633 676010 667639
rect 676066 665667 676094 668077
rect 676244 666990 676300 666999
rect 676244 666925 676300 666934
rect 676258 666809 676286 666925
rect 676246 666803 676298 666809
rect 676246 666745 676298 666751
rect 676244 666398 676300 666407
rect 676244 666333 676246 666342
rect 676298 666333 676300 666342
rect 676246 666301 676298 666307
rect 676052 665658 676108 665667
rect 676052 665593 676108 665602
rect 676246 665249 676298 665255
rect 676246 665191 676298 665197
rect 676054 665175 676106 665181
rect 676054 665117 676106 665123
rect 676066 663595 676094 665117
rect 676258 664335 676286 665191
rect 676244 664326 676300 664335
rect 676244 664261 676300 664270
rect 676052 663586 676108 663595
rect 676052 663521 676108 663530
rect 676054 662363 676106 662369
rect 676054 662305 676106 662311
rect 676066 661671 676094 662305
rect 676052 661662 676108 661671
rect 676052 661597 676108 661606
rect 676054 660661 676106 660667
rect 676052 660626 676054 660635
rect 676106 660626 676108 660635
rect 676052 660561 676108 660570
rect 676246 659921 676298 659927
rect 676244 659886 676246 659895
rect 676298 659886 676300 659895
rect 676244 659821 676300 659830
rect 675010 659506 675134 659534
rect 675010 635063 675038 659506
rect 679796 659294 679852 659303
rect 679796 659229 679852 659238
rect 679810 658415 679838 659229
rect 679796 658406 679852 658415
rect 679796 658341 679852 658350
rect 685460 658406 685516 658415
rect 685460 658341 685516 658350
rect 675382 656813 675434 656819
rect 675382 656755 675434 656761
rect 675394 653675 675422 656755
rect 679810 656745 679838 658341
rect 685474 657971 685502 658341
rect 685460 657962 685516 657971
rect 685460 657897 685516 657906
rect 679798 656739 679850 656745
rect 679798 656681 679850 656687
rect 675106 653110 675408 653138
rect 675106 651015 675134 653110
rect 675490 652199 675518 652458
rect 675476 652190 675532 652199
rect 675476 652125 675532 652134
rect 675490 651459 675518 651835
rect 675476 651450 675532 651459
rect 675476 651385 675532 651394
rect 675092 651006 675148 651015
rect 675092 650941 675148 650950
rect 675682 649831 675710 650016
rect 675668 649822 675724 649831
rect 675668 649757 675724 649766
rect 675298 649484 675422 649512
rect 675298 649438 675326 649484
rect 675202 649410 675326 649438
rect 675394 649424 675422 649484
rect 675202 648351 675230 649410
rect 675778 648351 675806 648799
rect 675188 648342 675244 648351
rect 675188 648277 675244 648286
rect 675764 648342 675820 648351
rect 675764 648277 675820 648286
rect 675190 648229 675242 648235
rect 675190 648171 675242 648177
rect 675094 645195 675146 645201
rect 675094 645137 675146 645143
rect 675106 641446 675134 645137
rect 675202 643296 675230 648171
rect 675298 648152 675408 648180
rect 675298 648087 675326 648152
rect 675286 648081 675338 648087
rect 675286 648023 675338 648029
rect 675778 645391 675806 645650
rect 675764 645382 675820 645391
rect 675764 645317 675820 645326
rect 675298 645118 675408 645146
rect 675298 644609 675326 645118
rect 675286 644603 675338 644609
rect 675286 644545 675338 644551
rect 675298 644452 675408 644480
rect 675298 643943 675326 644452
rect 675286 643937 675338 643943
rect 675286 643879 675338 643885
rect 675298 643817 675408 643845
rect 675298 643425 675326 643817
rect 675286 643419 675338 643425
rect 675286 643361 675338 643367
rect 675202 643268 675408 643296
rect 675298 642676 675422 642704
rect 675298 642630 675326 642676
rect 675202 642602 675326 642630
rect 675394 642616 675422 642676
rect 675202 642315 675230 642602
rect 675190 642309 675242 642315
rect 675190 642251 675242 642257
rect 675106 641418 675408 641446
rect 675106 640781 675408 640809
rect 675106 639133 675134 640781
rect 675094 639127 675146 639133
rect 675094 639069 675146 639075
rect 675106 638941 675408 638969
rect 674998 635057 675050 635063
rect 674998 634999 675050 635005
rect 675106 629143 675134 638941
rect 679702 635057 679754 635063
rect 679702 634999 679754 635005
rect 675094 629137 675146 629143
rect 675094 629079 675146 629085
rect 676244 625106 676300 625115
rect 676244 625041 676300 625050
rect 676258 624999 676286 625041
rect 676246 624993 676298 624999
rect 676246 624935 676298 624941
rect 676148 624662 676204 624671
rect 676148 624597 676204 624606
rect 676052 623478 676108 623487
rect 676052 623413 676054 623422
rect 676106 623413 676108 623422
rect 676054 623381 676106 623387
rect 676054 623143 676106 623149
rect 676054 623085 676106 623091
rect 676066 622895 676094 623085
rect 676052 622886 676108 622895
rect 676052 622821 676108 622830
rect 676052 622516 676108 622525
rect 676052 622451 676054 622460
rect 676106 622451 676108 622460
rect 676054 622419 676106 622425
rect 676162 622409 676190 624597
rect 679714 624227 679742 634999
rect 676244 624218 676300 624227
rect 676244 624153 676300 624162
rect 679700 624218 679756 624227
rect 679700 624153 679756 624162
rect 676258 622557 676286 624153
rect 676246 622551 676298 622557
rect 676246 622493 676298 622499
rect 676150 622403 676202 622409
rect 676150 622345 676202 622351
rect 676246 622033 676298 622039
rect 676052 621998 676108 622007
rect 676246 621975 676298 621981
rect 676052 621933 676054 621942
rect 676106 621933 676108 621942
rect 676054 621901 676106 621907
rect 676052 621406 676108 621415
rect 676052 621341 676054 621350
rect 676106 621341 676108 621350
rect 676054 621309 676106 621315
rect 676258 620675 676286 621975
rect 676244 620666 676300 620675
rect 676244 620601 676300 620610
rect 674902 619073 674954 619079
rect 674902 619015 674954 619021
rect 676054 619073 676106 619079
rect 676054 619015 676106 619021
rect 676066 618973 676094 619015
rect 676052 618964 676108 618973
rect 676052 618899 676108 618908
rect 676246 618851 676298 618857
rect 676246 618793 676298 618799
rect 676054 618629 676106 618635
rect 676258 618603 676286 618793
rect 676054 618571 676106 618577
rect 676244 618594 676300 618603
rect 676066 616531 676094 618571
rect 676244 618529 676300 618538
rect 676052 616522 676108 616531
rect 676052 616457 676108 616466
rect 674806 616335 674858 616341
rect 674806 616277 674858 616283
rect 676054 616335 676106 616341
rect 676054 616277 676106 616283
rect 676066 615939 676094 616277
rect 676052 615930 676108 615939
rect 676052 615865 676108 615874
rect 676246 615669 676298 615675
rect 676244 615634 676246 615643
rect 676298 615634 676300 615643
rect 676244 615569 676300 615578
rect 676054 614485 676106 614491
rect 676052 614450 676054 614459
rect 676106 614450 676108 614459
rect 676052 614385 676108 614394
rect 679988 613710 680044 613719
rect 679988 613645 680044 613654
rect 675382 613523 675434 613529
rect 675382 613465 675434 613471
rect 675394 608650 675422 613465
rect 680002 613275 680030 613645
rect 679796 613266 679852 613275
rect 679796 613201 679852 613210
rect 679988 613266 680044 613275
rect 679988 613201 680044 613210
rect 679810 612831 679838 613201
rect 679796 612822 679852 612831
rect 679796 612757 679852 612766
rect 680002 610643 680030 613201
rect 679990 610637 680042 610643
rect 679990 610579 680042 610585
rect 675106 608118 675408 608146
rect 675106 607799 675134 608118
rect 675092 607790 675148 607799
rect 675092 607725 675148 607734
rect 675092 607494 675148 607503
rect 675148 607452 675408 607480
rect 675092 607429 675148 607438
rect 675778 606467 675806 606835
rect 675764 606458 675820 606467
rect 675764 606393 675820 606402
rect 675106 604981 675408 605009
rect 675106 604839 675134 604981
rect 675092 604830 675148 604839
rect 675092 604765 675148 604774
rect 675298 604418 675408 604446
rect 674902 602127 674954 602133
rect 674902 602069 674954 602075
rect 674914 596454 674942 602069
rect 674998 602053 675050 602059
rect 675298 602027 675326 604418
rect 675394 603317 675422 603799
rect 675382 603311 675434 603317
rect 675382 603253 675434 603259
rect 675394 602725 675422 603174
rect 675382 602719 675434 602725
rect 675382 602661 675434 602667
rect 674998 601995 675050 602001
rect 675284 602018 675340 602027
rect 675010 599192 675038 601995
rect 675284 601953 675340 601962
rect 675778 600251 675806 600658
rect 675764 600242 675820 600251
rect 675764 600177 675820 600186
rect 675394 599839 675422 600140
rect 675382 599833 675434 599839
rect 675382 599775 675434 599781
rect 675106 599460 675408 599488
rect 675106 599321 675134 599460
rect 675094 599315 675146 599321
rect 675094 599257 675146 599263
rect 675010 599164 675134 599192
rect 675106 598304 675134 599164
rect 675298 598868 675422 598896
rect 675298 598822 675326 598868
rect 675202 598794 675326 598822
rect 675394 598808 675422 598868
rect 675202 598433 675230 598794
rect 675190 598427 675242 598433
rect 675190 598369 675242 598375
rect 675106 598276 675408 598304
rect 675106 597610 675408 597638
rect 675106 596583 675134 597610
rect 675094 596577 675146 596583
rect 675094 596519 675146 596525
rect 674914 596426 675408 596454
rect 675298 595908 675422 595936
rect 675298 595788 675326 595908
rect 674722 595760 675326 595788
rect 675394 595774 675422 595908
rect 674614 586439 674666 586445
rect 674614 586381 674666 586387
rect 674230 576005 674282 576011
rect 674230 575947 674282 575953
rect 674134 573119 674186 573125
rect 674134 573061 674186 573067
rect 673846 568457 673898 568463
rect 673846 568399 673898 568405
rect 674038 559577 674090 559583
rect 674038 559519 674090 559525
rect 673846 553361 673898 553367
rect 673846 553303 673898 553309
rect 673750 526721 673802 526727
rect 673750 526663 673802 526669
rect 673654 525241 673706 525247
rect 673654 525183 673706 525189
rect 673462 524871 673514 524877
rect 673462 524813 673514 524819
rect 672886 524501 672938 524507
rect 672886 524443 672938 524449
rect 673858 480107 673886 553303
rect 674050 486619 674078 559519
rect 674326 555285 674378 555291
rect 674326 555227 674378 555233
rect 674230 551955 674282 551961
rect 674230 551897 674282 551903
rect 674038 486613 674090 486619
rect 674038 486555 674090 486561
rect 674242 482179 674270 551897
rect 674338 485731 674366 555227
rect 674518 548921 674570 548927
rect 674518 548863 674570 548869
rect 674422 543667 674474 543673
rect 674422 543609 674474 543615
rect 674326 485725 674378 485731
rect 674326 485667 674378 485673
rect 674434 483733 674462 543609
rect 674530 486693 674558 548863
rect 674626 529909 674654 586381
rect 674722 532795 674750 595760
rect 675106 593941 675408 593969
rect 675106 586445 675134 593941
rect 679702 590361 679754 590367
rect 679702 590303 679754 590309
rect 675094 586439 675146 586445
rect 675094 586381 675146 586387
rect 676340 578338 676396 578347
rect 676340 578273 676396 578282
rect 676148 577598 676204 577607
rect 676148 577533 676204 577542
rect 676162 576529 676190 577533
rect 676244 577154 676300 577163
rect 676244 577089 676300 577098
rect 676258 576677 676286 577089
rect 676246 576671 676298 576677
rect 676246 576613 676298 576619
rect 676150 576523 676202 576529
rect 676150 576465 676202 576471
rect 676354 576381 676382 578273
rect 679714 577163 679742 590303
rect 679700 577154 679756 577163
rect 679700 577089 679756 577098
rect 676342 576375 676394 576381
rect 676342 576317 676394 576323
rect 676244 576266 676300 576275
rect 676244 576201 676246 576210
rect 676298 576201 676300 576210
rect 676246 576169 676298 576175
rect 676054 576005 676106 576011
rect 675956 575970 676012 575979
rect 676054 575947 676106 575953
rect 675956 575905 675958 575914
rect 676010 575905 676012 575914
rect 675958 575873 676010 575879
rect 675956 575526 676012 575535
rect 675956 575461 675958 575470
rect 676010 575461 676012 575470
rect 675958 575429 676010 575435
rect 675958 574969 676010 574975
rect 675956 574934 675958 574943
rect 676010 574934 676012 574943
rect 675956 574869 676012 574878
rect 676066 573463 676094 575947
rect 676244 574194 676300 574203
rect 676244 574129 676246 574138
rect 676298 574129 676300 574138
rect 676246 574097 676298 574103
rect 676052 573454 676108 573463
rect 676052 573389 676108 573398
rect 676054 573119 676106 573125
rect 676054 573061 676106 573067
rect 676066 571391 676094 573061
rect 676052 571382 676108 571391
rect 676052 571317 676108 571326
rect 676054 569567 676106 569573
rect 676052 569532 676054 569541
rect 676106 569532 676108 569541
rect 676052 569467 676108 569476
rect 676246 569197 676298 569203
rect 676244 569162 676246 569171
rect 676298 569162 676300 569171
rect 676244 569097 676300 569106
rect 676054 568457 676106 568463
rect 676052 568422 676054 568431
rect 676106 568422 676108 568431
rect 676052 568357 676108 568366
rect 676054 568013 676106 568019
rect 676052 567978 676054 567987
rect 676106 567978 676108 567987
rect 676052 567913 676108 567922
rect 676246 567717 676298 567723
rect 676244 567682 676246 567691
rect 676298 567682 676300 567691
rect 676244 567617 676300 567626
rect 675382 567495 675434 567501
rect 675382 567437 675434 567443
rect 675394 563475 675422 567437
rect 679796 567090 679852 567099
rect 679796 567025 679852 567034
rect 679810 566211 679838 567025
rect 679796 566202 679852 566211
rect 679796 566137 679852 566146
rect 685460 566202 685516 566211
rect 685460 566137 685516 566146
rect 679810 564541 679838 566137
rect 685474 565767 685502 566137
rect 685460 565758 685516 565767
rect 685460 565693 685516 565702
rect 679798 564535 679850 564541
rect 679798 564477 679850 564483
rect 675092 562946 675148 562955
rect 675148 562904 675408 562932
rect 675092 562881 675148 562890
rect 675490 561771 675518 562252
rect 675476 561762 675532 561771
rect 675476 561697 675532 561706
rect 675394 561475 675422 561660
rect 675380 561466 675436 561475
rect 675380 561401 675436 561410
rect 675394 559583 675422 559810
rect 675382 559577 675434 559583
rect 675382 559519 675434 559525
rect 675490 558959 675518 559218
rect 675476 558950 675532 558959
rect 675476 558885 675532 558894
rect 675190 558837 675242 558843
rect 675190 558779 675242 558785
rect 674806 558097 674858 558103
rect 674806 558039 674858 558045
rect 674710 532789 674762 532795
rect 674710 532731 674762 532737
rect 674614 529903 674666 529909
rect 674614 529845 674666 529851
rect 674518 486687 674570 486693
rect 674518 486629 674570 486635
rect 674818 483807 674846 558039
rect 675094 555877 675146 555883
rect 675094 555819 675146 555825
rect 674998 553805 675050 553811
rect 674998 553747 675050 553753
rect 674806 483801 674858 483807
rect 674806 483743 674858 483749
rect 674422 483727 674474 483733
rect 674422 483669 674474 483675
rect 675010 483659 675038 553747
rect 675106 551240 675134 555819
rect 675202 553090 675230 558779
rect 675394 558103 675422 558626
rect 675382 558097 675434 558103
rect 675382 558039 675434 558045
rect 675298 557946 675408 557974
rect 675298 553335 675326 557946
rect 675490 555291 675518 555444
rect 675478 555285 675530 555291
rect 675478 555227 675530 555233
rect 675778 554667 675806 554926
rect 675764 554658 675820 554667
rect 675764 554593 675820 554602
rect 675490 553811 675518 554260
rect 675478 553805 675530 553811
rect 675478 553747 675530 553753
rect 675394 553367 675422 553631
rect 675382 553361 675434 553367
rect 675284 553326 675340 553335
rect 675382 553303 675434 553309
rect 675284 553261 675340 553270
rect 675202 553062 675408 553090
rect 675490 551961 675518 552410
rect 675478 551955 675530 551961
rect 675478 551897 675530 551903
rect 675106 551212 675408 551240
rect 675106 550581 675408 550609
rect 675106 548927 675134 550581
rect 675094 548921 675146 548927
rect 675094 548863 675146 548869
rect 675106 548741 675408 548769
rect 675106 543673 675134 548741
rect 679702 547219 679754 547225
rect 679702 547161 679754 547167
rect 675094 543667 675146 543673
rect 675094 543609 675146 543615
rect 676244 534974 676300 534983
rect 676244 534909 676300 534918
rect 676148 534382 676204 534391
rect 676148 534317 676204 534326
rect 676052 534234 676108 534243
rect 676052 534169 676108 534178
rect 676066 533461 676094 534169
rect 676054 533455 676106 533461
rect 676054 533397 676106 533403
rect 676162 533165 676190 534317
rect 676258 533313 676286 534909
rect 679714 533651 679742 547161
rect 679700 533642 679756 533651
rect 679700 533577 679756 533586
rect 676246 533307 676298 533313
rect 676246 533249 676298 533255
rect 676150 533159 676202 533165
rect 676150 533101 676202 533107
rect 676532 533050 676588 533059
rect 676532 532985 676588 532994
rect 676054 532789 676106 532795
rect 675956 532754 676012 532763
rect 676054 532731 676106 532737
rect 675956 532689 675958 532698
rect 676010 532689 676012 532698
rect 675958 532657 676010 532663
rect 676066 530247 676094 532731
rect 676244 531570 676300 531579
rect 676244 531505 676246 531514
rect 676298 531505 676300 531514
rect 676246 531473 676298 531479
rect 676052 530238 676108 530247
rect 676052 530173 676108 530182
rect 676054 529903 676106 529909
rect 676054 529845 676106 529851
rect 676066 528175 676094 529845
rect 676052 528166 676108 528175
rect 676052 528101 676108 528110
rect 676054 526721 676106 526727
rect 676052 526686 676054 526695
rect 676106 526686 676108 526695
rect 676052 526621 676108 526630
rect 676054 526351 676106 526357
rect 676052 526316 676054 526325
rect 676106 526316 676108 526325
rect 676052 526251 676108 526260
rect 676246 525981 676298 525987
rect 676244 525946 676246 525955
rect 676298 525946 676300 525955
rect 676244 525881 676300 525890
rect 676054 525241 676106 525247
rect 676052 525206 676054 525215
rect 676106 525206 676108 525215
rect 676052 525141 676108 525150
rect 676054 524871 676106 524877
rect 676052 524836 676054 524845
rect 676106 524836 676108 524845
rect 676052 524771 676108 524780
rect 676246 524501 676298 524507
rect 676244 524466 676246 524475
rect 676298 524466 676300 524475
rect 676244 524401 676300 524410
rect 676546 498311 676574 532985
rect 676628 532014 676684 532023
rect 676628 531949 676684 531958
rect 676534 498305 676586 498311
rect 676534 498247 676586 498253
rect 676244 490574 676300 490583
rect 676244 490509 676300 490518
rect 676148 490130 676204 490139
rect 676258 490097 676286 490509
rect 676148 490065 676204 490074
rect 676246 490091 676298 490097
rect 676162 489801 676190 490065
rect 676246 490033 676298 490039
rect 676244 489982 676300 489991
rect 676244 489917 676246 489926
rect 676298 489917 676300 489926
rect 676246 489885 676298 489891
rect 676150 489795 676202 489801
rect 676150 489737 676202 489743
rect 676246 488759 676298 488765
rect 676246 488701 676298 488707
rect 676052 488354 676108 488363
rect 676052 488289 676108 488298
rect 676066 488173 676094 488289
rect 676054 488167 676106 488173
rect 676054 488109 676106 488115
rect 675284 487910 675340 487919
rect 675284 487845 675340 487854
rect 674998 483653 675050 483659
rect 674998 483595 675050 483601
rect 674230 482173 674282 482179
rect 674230 482115 674282 482121
rect 673846 480101 673898 480107
rect 673846 480043 673898 480049
rect 675298 440665 675326 487845
rect 676258 487179 676286 488701
rect 676642 488173 676670 531949
rect 676724 530978 676780 530987
rect 676724 530913 676780 530922
rect 676738 488765 676766 530913
rect 679796 523578 679852 523587
rect 679796 523513 679852 523522
rect 679810 522995 679838 523513
rect 679796 522986 679852 522995
rect 679796 522921 679852 522930
rect 685460 522986 685516 522995
rect 685460 522921 685516 522930
rect 679810 521325 679838 522921
rect 685474 522551 685502 522921
rect 685460 522542 685516 522551
rect 685460 522477 685516 522486
rect 679798 521319 679850 521325
rect 679798 521261 679850 521267
rect 679702 498305 679754 498311
rect 679702 498247 679754 498253
rect 679714 489251 679742 498247
rect 679700 489242 679756 489251
rect 679700 489177 679756 489186
rect 676726 488759 676778 488765
rect 676726 488701 676778 488707
rect 676724 488650 676780 488659
rect 676724 488585 676780 488594
rect 676630 488167 676682 488173
rect 676630 488109 676682 488115
rect 676244 487170 676300 487179
rect 676244 487105 676246 487114
rect 676298 487105 676300 487114
rect 676246 487073 676298 487079
rect 676052 486874 676108 486883
rect 676052 486809 676054 486818
rect 676106 486809 676108 486818
rect 676054 486777 676106 486783
rect 676054 486687 676106 486693
rect 676054 486629 676106 486635
rect 676066 485847 676094 486629
rect 676246 486613 676298 486619
rect 676246 486555 676298 486561
rect 676052 485838 676108 485847
rect 676052 485773 676108 485782
rect 676054 485725 676106 485731
rect 676054 485667 676106 485673
rect 676066 484367 676094 485667
rect 676258 485107 676286 486555
rect 676244 485098 676300 485107
rect 676244 485033 676300 485042
rect 676052 484358 676108 484367
rect 676052 484293 676108 484302
rect 676054 483801 676106 483807
rect 675956 483766 676012 483775
rect 676054 483743 676106 483749
rect 675956 483701 675958 483710
rect 676010 483701 676012 483710
rect 675958 483669 676010 483675
rect 676066 482295 676094 483743
rect 676246 483653 676298 483659
rect 676246 483595 676298 483601
rect 676052 482286 676108 482295
rect 676052 482221 676108 482230
rect 676054 482173 676106 482179
rect 676054 482115 676106 482121
rect 676066 481925 676094 482115
rect 676052 481916 676108 481925
rect 676052 481851 676108 481860
rect 676258 481555 676286 483595
rect 676244 481546 676300 481555
rect 676244 481481 676300 481490
rect 676246 480101 676298 480107
rect 676244 480066 676246 480075
rect 676298 480066 676300 480075
rect 676244 480001 676300 480010
rect 673846 440659 673898 440665
rect 673846 440601 673898 440607
rect 675286 440659 675338 440665
rect 675286 440601 675338 440607
rect 673750 400625 673802 400631
rect 673750 400567 673802 400573
rect 673762 356823 673790 400567
rect 673858 400335 673886 440601
rect 676148 402366 676204 402375
rect 676148 402301 676204 402310
rect 676052 401626 676108 401635
rect 676052 401561 676108 401570
rect 675956 400664 676012 400673
rect 675956 400599 675958 400608
rect 676010 400599 676012 400608
rect 675958 400567 676010 400573
rect 676066 400557 676094 401561
rect 676054 400551 676106 400557
rect 676054 400493 676106 400499
rect 676162 400409 676190 402301
rect 676244 401922 676300 401931
rect 676244 401857 676300 401866
rect 676258 400483 676286 401857
rect 676738 401043 676766 488585
rect 679892 479178 679948 479187
rect 679892 479113 679948 479122
rect 679906 478595 679934 479113
rect 679700 478586 679756 478595
rect 679700 478521 679756 478530
rect 679892 478586 679948 478595
rect 679892 478521 679948 478530
rect 679714 478151 679742 478521
rect 679906 478183 679934 478521
rect 679894 478177 679946 478183
rect 679700 478142 679756 478151
rect 679894 478119 679946 478125
rect 679700 478077 679756 478086
rect 676724 401034 676780 401043
rect 676724 400969 676780 400978
rect 676246 400477 676298 400483
rect 676246 400419 676298 400425
rect 676150 400403 676202 400409
rect 676150 400345 676202 400351
rect 673846 400329 673898 400335
rect 676246 400329 676298 400335
rect 673846 400271 673898 400277
rect 676244 400294 676246 400303
rect 676298 400294 676300 400303
rect 676244 400229 676300 400238
rect 676052 399110 676108 399119
rect 676052 399045 676054 399054
rect 676106 399045 676108 399054
rect 676054 399013 676106 399019
rect 675572 397038 675628 397047
rect 675572 396973 675628 396982
rect 675284 395262 675340 395271
rect 675284 395197 675340 395206
rect 675190 392559 675242 392565
rect 675190 392501 675242 392507
rect 674998 391745 675050 391751
rect 674998 391687 675050 391693
rect 675010 388814 675038 391687
rect 674914 388786 675038 388814
rect 674914 381040 674942 388786
rect 675202 387552 675230 392501
rect 675010 387524 675230 387552
rect 675010 381410 675038 387524
rect 675298 387404 675326 395197
rect 675202 387376 675326 387404
rect 675094 385973 675146 385979
rect 675094 385915 675146 385921
rect 675106 381613 675134 385915
rect 675202 385110 675230 387376
rect 675586 387256 675614 396973
rect 676244 393930 676300 393939
rect 676244 393865 676300 393874
rect 676258 392565 676286 393865
rect 676246 392559 676298 392565
rect 676246 392501 676298 392507
rect 676244 392450 676300 392459
rect 676244 392385 676300 392394
rect 676258 391751 676286 392385
rect 676246 391745 676298 391751
rect 676246 391687 676298 391693
rect 679796 390970 679852 390979
rect 679796 390905 679852 390914
rect 679810 390387 679838 390905
rect 679796 390378 679852 390387
rect 679796 390313 679852 390322
rect 685460 390378 685516 390387
rect 685460 390313 685516 390322
rect 679810 388865 679838 390313
rect 685474 389943 685502 390313
rect 685460 389934 685516 389943
rect 685460 389869 685516 389878
rect 679798 388859 679850 388865
rect 679798 388801 679850 388807
rect 675298 387228 675614 387256
rect 675298 385737 675326 387228
rect 675394 385979 675422 386280
rect 675382 385973 675434 385979
rect 675382 385915 675434 385921
rect 675298 385709 675408 385737
rect 675202 385082 675326 385110
rect 675298 385036 675326 385082
rect 675394 385036 675422 385096
rect 675298 385008 675422 385036
rect 675764 384754 675820 384763
rect 675764 384689 675820 384698
rect 675778 384430 675806 384689
rect 675764 382978 675820 382987
rect 675764 382913 675820 382922
rect 675778 382580 675806 382913
rect 675476 382386 675532 382395
rect 675476 382321 675532 382330
rect 675490 382062 675518 382321
rect 675094 381607 675146 381613
rect 675094 381549 675146 381555
rect 675010 381382 675408 381410
rect 674914 381012 675422 381040
rect 675394 380730 675422 381012
rect 675764 378834 675820 378843
rect 675764 378769 675820 378778
rect 675778 378288 675806 378769
rect 675764 378094 675820 378103
rect 675764 378029 675820 378038
rect 675778 377696 675806 378029
rect 675476 377206 675532 377215
rect 675476 377141 675532 377150
rect 675490 377075 675518 377141
rect 675188 376466 675244 376475
rect 675244 376424 675408 376452
rect 675188 376401 675244 376410
rect 675476 375726 675532 375735
rect 675476 375661 675532 375670
rect 675490 375254 675518 375661
rect 675092 374394 675148 374403
rect 675092 374329 675148 374338
rect 675106 373418 675134 374329
rect 675106 373390 675408 373418
rect 675764 372026 675820 372035
rect 675764 371961 675820 371970
rect 675778 371554 675806 371961
rect 676148 358114 676204 358123
rect 676148 358049 676204 358058
rect 676162 357341 676190 358049
rect 676244 357374 676300 357383
rect 676150 357335 676202 357341
rect 676244 357309 676300 357318
rect 676150 357277 676202 357283
rect 676258 357267 676286 357309
rect 676246 357261 676298 357267
rect 676052 357226 676108 357235
rect 676246 357203 676298 357209
rect 676052 357161 676054 357170
rect 676106 357161 676108 357170
rect 676054 357129 676106 357135
rect 673750 356817 673802 356823
rect 676054 356817 676106 356823
rect 673750 356759 673802 356765
rect 676052 356782 676054 356791
rect 676106 356782 676108 356791
rect 676052 356717 676108 356726
rect 676052 353822 676108 353831
rect 676052 353757 676108 353766
rect 675572 352638 675628 352647
rect 675572 352573 675628 352582
rect 674518 352451 674570 352457
rect 674518 352393 674570 352399
rect 674134 348603 674186 348609
rect 674134 348545 674186 348551
rect 674146 336621 674174 348545
rect 674530 339581 674558 352393
rect 674806 351415 674858 351421
rect 674806 351357 674858 351363
rect 674818 339803 674846 351357
rect 675284 350862 675340 350871
rect 675284 350797 675340 350806
rect 675190 348529 675242 348535
rect 675190 348471 675242 348477
rect 674902 345791 674954 345797
rect 674902 345733 674954 345739
rect 674806 339797 674858 339803
rect 674806 339739 674858 339745
rect 674518 339575 674570 339581
rect 674518 339517 674570 339523
rect 674134 336615 674186 336621
rect 674134 336557 674186 336563
rect 674914 331312 674942 345733
rect 674998 345717 675050 345723
rect 674998 345659 675050 345665
rect 675010 332533 675038 345659
rect 675094 345643 675146 345649
rect 675094 345585 675146 345591
rect 675106 335569 675134 345585
rect 675202 336862 675230 348471
rect 675298 339896 675326 350797
rect 675586 348494 675614 352573
rect 676066 352457 676094 353757
rect 676054 352451 676106 352457
rect 676054 352393 676106 352399
rect 676052 352342 676108 352351
rect 676052 352277 676108 352286
rect 676066 351421 676094 352277
rect 676916 351602 676972 351611
rect 676916 351537 676972 351546
rect 676054 351415 676106 351421
rect 676054 351357 676106 351363
rect 676052 350270 676108 350279
rect 676052 350205 676108 350214
rect 676066 348535 676094 350205
rect 676244 349530 676300 349539
rect 676244 349465 676300 349474
rect 676258 348609 676286 349465
rect 676820 349086 676876 349095
rect 676820 349021 676876 349030
rect 676246 348603 676298 348609
rect 676246 348545 676298 348551
rect 676054 348529 676106 348535
rect 675586 348466 675806 348494
rect 676054 348471 676106 348477
rect 675778 341431 675806 348466
rect 676244 348050 676300 348059
rect 676244 347985 676300 347994
rect 676052 347828 676108 347837
rect 676052 347763 676108 347772
rect 675956 347310 676012 347319
rect 675956 347245 676012 347254
rect 675970 345797 675998 347245
rect 675958 345791 676010 345797
rect 675958 345733 676010 345739
rect 676066 345723 676094 347763
rect 676054 345717 676106 345723
rect 676054 345659 676106 345665
rect 676258 345649 676286 347985
rect 676246 345643 676298 345649
rect 676246 345585 676298 345591
rect 676834 343027 676862 349021
rect 676820 343018 676876 343027
rect 676820 342953 676876 342962
rect 676930 342879 676958 351537
rect 679892 346570 679948 346579
rect 679892 346505 679948 346514
rect 679906 346135 679934 346505
rect 679892 346126 679948 346135
rect 679892 346061 679948 346070
rect 679700 345978 679756 345987
rect 679700 345913 679756 345922
rect 679714 345543 679742 345913
rect 679906 345871 679934 346061
rect 679894 345865 679946 345871
rect 679894 345807 679946 345813
rect 679700 345534 679756 345543
rect 679700 345469 679756 345478
rect 676916 342870 676972 342879
rect 676916 342805 676972 342814
rect 675766 341425 675818 341431
rect 675766 341367 675818 341373
rect 675490 340691 675518 341066
rect 675766 340759 675818 340765
rect 675766 340701 675818 340707
rect 675478 340685 675530 340691
rect 675478 340627 675530 340633
rect 675778 340548 675806 340701
rect 675298 339868 675408 339896
rect 675286 339797 675338 339803
rect 675286 339739 675338 339745
rect 675298 337409 675326 339739
rect 675382 339575 675434 339581
rect 675382 339517 675434 339523
rect 675394 339216 675422 339517
rect 675298 337381 675408 337409
rect 675202 336834 675408 336862
rect 675382 336615 675434 336621
rect 675382 336557 675434 336563
rect 675394 336182 675422 336557
rect 675106 335541 675408 335569
rect 675764 333546 675820 333555
rect 675764 333481 675820 333490
rect 675778 333074 675806 333481
rect 675010 332505 675408 332533
rect 675476 332362 675532 332371
rect 675476 332297 675532 332306
rect 675490 331890 675518 332297
rect 674914 331284 675038 331312
rect 675010 331238 675038 331284
rect 675010 331210 675408 331238
rect 675764 330586 675820 330595
rect 675764 330521 675820 330530
rect 675778 330040 675806 330521
rect 675092 328218 675148 328227
rect 675148 328176 675408 328204
rect 675092 328153 675148 328162
rect 675380 326886 675436 326895
rect 675380 326821 675436 326830
rect 675394 326340 675422 326821
rect 676340 312234 676396 312243
rect 676340 312169 676396 312178
rect 676148 311642 676204 311651
rect 676148 311577 676204 311586
rect 676162 311165 676190 311577
rect 676246 311233 676298 311239
rect 676244 311198 676246 311207
rect 676298 311198 676300 311207
rect 676150 311159 676202 311165
rect 676244 311133 676300 311142
rect 676150 311101 676202 311107
rect 676354 311091 676382 312169
rect 676342 311085 676394 311091
rect 676342 311027 676394 311033
rect 676244 306758 676300 306767
rect 676244 306693 676300 306702
rect 676258 305319 676286 306693
rect 674134 305313 674186 305319
rect 674134 305255 674186 305261
rect 676246 305313 676298 305319
rect 676246 305255 676298 305261
rect 673942 302575 673994 302581
rect 673942 302517 673994 302523
rect 673954 291777 673982 302517
rect 674038 302501 674090 302507
rect 674038 302443 674090 302449
rect 674050 294293 674078 302443
rect 674146 295995 674174 305255
rect 676244 304834 676300 304843
rect 676244 304769 676300 304778
rect 676052 304464 676108 304473
rect 676052 304399 676108 304408
rect 675956 303946 676012 303955
rect 675956 303881 676012 303890
rect 675970 302581 675998 303881
rect 675958 302575 676010 302581
rect 675958 302517 676010 302523
rect 676066 302507 676094 304399
rect 676054 302501 676106 302507
rect 676054 302443 676106 302449
rect 676258 302433 676286 304769
rect 674230 302427 674282 302433
rect 674230 302369 674282 302375
rect 676246 302427 676298 302433
rect 676246 302369 676298 302375
rect 674134 295989 674186 295995
rect 674134 295931 674186 295937
rect 674242 295773 674270 302369
rect 679988 300690 680044 300699
rect 679988 300625 680044 300634
rect 680002 300255 680030 300625
rect 679796 300246 679852 300255
rect 679796 300181 679852 300190
rect 679988 300246 680044 300255
rect 679988 300181 680044 300190
rect 679810 299811 679838 300181
rect 679796 299802 679852 299811
rect 679796 299737 679852 299746
rect 680002 299621 680030 300181
rect 679990 299615 680042 299621
rect 679990 299557 680042 299563
rect 675106 296060 675408 296088
rect 674230 295767 674282 295773
rect 674230 295709 674282 295715
rect 674038 294287 674090 294293
rect 674038 294229 674090 294235
rect 673942 291771 673994 291777
rect 673942 291713 673994 291719
rect 675106 290889 675134 296060
rect 675286 295989 675338 295995
rect 675286 295931 675338 295937
rect 675190 295767 675242 295773
rect 675190 295709 675242 295715
rect 675202 294904 675230 295709
rect 675298 295537 675326 295931
rect 675298 295509 675408 295537
rect 675202 294876 675408 294904
rect 675764 294622 675820 294631
rect 675764 294557 675820 294566
rect 675190 294287 675242 294293
rect 675190 294229 675242 294235
rect 675202 291870 675230 294229
rect 675778 294224 675806 294557
rect 675380 292846 675436 292855
rect 675380 292781 675436 292790
rect 675394 292374 675422 292781
rect 675202 291842 675408 291870
rect 675190 291771 675242 291777
rect 675190 291713 675242 291719
rect 675202 291204 675230 291713
rect 675202 291176 675408 291204
rect 675094 290883 675146 290889
rect 675094 290825 675146 290831
rect 675764 290774 675820 290783
rect 675764 290709 675820 290718
rect 675778 290555 675806 290709
rect 675668 288554 675724 288563
rect 675668 288489 675724 288498
rect 675682 288082 675710 288489
rect 675572 287814 675628 287823
rect 675572 287749 675628 287758
rect 675586 287519 675614 287749
rect 675476 287222 675532 287231
rect 675476 287157 675532 287166
rect 675490 286898 675518 287157
rect 675764 286630 675820 286639
rect 675764 286565 675820 286574
rect 675778 286232 675806 286565
rect 675476 285594 675532 285603
rect 675476 285529 675532 285538
rect 675490 285048 675518 285529
rect 675092 283226 675148 283235
rect 675148 283184 675408 283212
rect 675092 283161 675148 283170
rect 675092 282190 675148 282199
rect 675092 282125 675148 282134
rect 675106 281362 675134 282125
rect 675106 281334 675408 281362
rect 675092 278342 675148 278351
rect 675092 278277 675148 278286
rect 672596 278194 672652 278203
rect 672596 278129 672652 278138
rect 675106 278013 675134 278277
rect 675094 278007 675146 278013
rect 675094 277949 675146 277955
rect 679798 278007 679850 278013
rect 679798 277949 679850 277955
rect 672500 273458 672556 273467
rect 672500 273393 672556 273402
rect 679700 270646 679756 270655
rect 679700 270581 679756 270590
rect 676148 266946 676204 266955
rect 676148 266881 676204 266890
rect 672404 266798 672460 266807
rect 672404 266733 672460 266742
rect 669814 264983 669866 264989
rect 669814 264925 669866 264931
rect 669622 264909 669674 264915
rect 669622 264851 669674 264857
rect 665878 250701 665930 250707
rect 665878 250643 665930 250649
rect 665890 247673 665918 250643
rect 665878 247667 665930 247673
rect 665878 247609 665930 247615
rect 672418 174751 672446 266733
rect 672596 266650 672652 266659
rect 672596 266585 672652 266594
rect 672404 174742 672460 174751
rect 672404 174677 672460 174686
rect 672610 173567 672638 266585
rect 673750 266389 673802 266395
rect 673750 266331 673802 266337
rect 673762 265063 673790 266331
rect 676052 266206 676108 266215
rect 676052 266141 676108 266150
rect 676066 265433 676094 266141
rect 676054 265427 676106 265433
rect 676054 265369 676106 265375
rect 676162 265137 676190 266881
rect 676244 266502 676300 266511
rect 676244 266437 676300 266446
rect 676258 265285 676286 266437
rect 676246 265279 676298 265285
rect 676246 265221 676298 265227
rect 676150 265131 676202 265137
rect 676150 265073 676202 265079
rect 673750 265057 673802 265063
rect 673750 264999 673802 265005
rect 676054 265057 676106 265063
rect 676054 264999 676106 265005
rect 673762 247694 673790 264999
rect 676066 264291 676094 264999
rect 679714 264883 679742 270581
rect 679700 264874 679756 264883
rect 679700 264809 679756 264818
rect 676052 264282 676108 264291
rect 676052 264217 676108 264226
rect 679810 264143 679838 277949
rect 679796 264134 679852 264143
rect 679796 264069 679852 264078
rect 676244 262654 676300 262663
rect 676244 262589 676300 262598
rect 676258 262177 676286 262589
rect 674806 262171 674858 262177
rect 674806 262113 674858 262119
rect 676246 262171 676298 262177
rect 676246 262113 676298 262119
rect 674614 259433 674666 259439
rect 674614 259375 674666 259381
rect 674518 256991 674570 256997
rect 674518 256933 674570 256939
rect 673762 247666 673886 247694
rect 673858 219553 673886 247666
rect 674530 247525 674558 256933
rect 674626 249153 674654 259375
rect 674710 256473 674762 256479
rect 674710 256415 674762 256421
rect 674614 249147 674666 249153
rect 674614 249089 674666 249095
rect 674518 247519 674570 247525
rect 674518 247461 674570 247467
rect 674722 242789 674750 256415
rect 674818 250263 674846 262113
rect 676052 261322 676108 261331
rect 676052 261257 676108 261266
rect 675284 259842 675340 259851
rect 675284 259777 675340 259786
rect 675190 259285 675242 259291
rect 675190 259227 675242 259233
rect 674998 256399 675050 256405
rect 674998 256341 675050 256347
rect 674902 253587 674954 253593
rect 674902 253529 674954 253535
rect 674806 250257 674858 250263
rect 674806 250199 674858 250205
rect 674710 242783 674762 242789
rect 674710 242725 674762 242731
rect 674914 241328 674942 253529
rect 675010 245546 675038 256341
rect 675094 247519 675146 247525
rect 675094 247461 675146 247467
rect 675106 246212 675134 247461
rect 675202 246878 675230 259227
rect 675298 250356 675326 259777
rect 676066 259439 676094 261257
rect 676820 259990 676876 259999
rect 676820 259925 676876 259934
rect 676054 259433 676106 259439
rect 676054 259375 676106 259381
rect 676054 259285 676106 259291
rect 676052 259250 676054 259259
rect 676106 259250 676108 259259
rect 676052 259185 676108 259194
rect 676052 258732 676108 258741
rect 676052 258667 676108 258676
rect 676066 256997 676094 258667
rect 676244 257030 676300 257039
rect 676054 256991 676106 256997
rect 676244 256965 676300 256974
rect 676054 256933 676106 256939
rect 676052 256882 676108 256891
rect 676052 256817 676108 256826
rect 676066 256479 676094 256817
rect 676054 256473 676106 256479
rect 676054 256415 676106 256421
rect 676258 256405 676286 256965
rect 676246 256399 676298 256405
rect 676246 256341 676298 256347
rect 676052 256290 676108 256299
rect 676052 256225 676108 256234
rect 676066 253593 676094 256225
rect 676054 253587 676106 253593
rect 676054 253529 676106 253535
rect 676834 253339 676862 259925
rect 679700 255550 679756 255559
rect 679700 255485 679756 255494
rect 679714 254967 679742 255485
rect 679700 254958 679756 254967
rect 679700 254893 679756 254902
rect 685460 254958 685516 254967
rect 685460 254893 685516 254902
rect 679714 253519 679742 254893
rect 685474 254523 685502 254893
rect 685460 254514 685516 254523
rect 685460 254449 685516 254458
rect 679702 253513 679754 253519
rect 679702 253455 679754 253461
rect 676820 253330 676876 253339
rect 676820 253265 676876 253274
rect 675394 250707 675422 251082
rect 675764 250814 675820 250823
rect 675764 250749 675820 250758
rect 675382 250701 675434 250707
rect 675382 250643 675434 250649
rect 675778 250523 675806 250749
rect 675298 250328 675518 250356
rect 675286 250257 675338 250263
rect 675286 250199 675338 250205
rect 675298 249246 675326 250199
rect 675490 249898 675518 250328
rect 675298 249218 675408 249246
rect 675286 249147 675338 249153
rect 675286 249089 675338 249095
rect 675298 247396 675326 249089
rect 675298 247368 675408 247396
rect 675202 246850 675326 246878
rect 675298 246804 675326 246850
rect 675394 246804 675422 246864
rect 675298 246776 675422 246804
rect 675106 246184 675408 246212
rect 675298 245592 675422 245620
rect 675298 245546 675326 245592
rect 675010 245518 675326 245546
rect 675394 245532 675422 245592
rect 675668 243562 675724 243571
rect 675668 243497 675724 243506
rect 675682 243090 675710 243497
rect 675382 242783 675434 242789
rect 675382 242725 675434 242731
rect 675394 242498 675422 242725
rect 675092 241934 675148 241943
rect 675148 241878 675408 241889
rect 675092 241869 675408 241878
rect 675106 241861 675408 241869
rect 674914 241300 675038 241328
rect 675010 241254 675038 241300
rect 675010 241226 675408 241254
rect 675188 241046 675244 241055
rect 675188 240981 675244 240990
rect 675202 240070 675230 240981
rect 675202 240042 675326 240070
rect 675298 239996 675326 240042
rect 675394 239996 675422 240056
rect 675298 239968 675422 239996
rect 675092 238234 675148 238243
rect 675148 238192 675408 238220
rect 675092 238169 675148 238178
rect 675764 236902 675820 236911
rect 675764 236837 675820 236846
rect 675778 236356 675806 236837
rect 676246 221841 676298 221847
rect 676244 221806 676246 221815
rect 676298 221806 676300 221815
rect 676244 221741 676300 221750
rect 676148 221214 676204 221223
rect 676148 221149 676204 221158
rect 673846 219547 673898 219553
rect 676054 219547 676106 219553
rect 673846 219489 673898 219495
rect 676052 219512 676054 219521
rect 676106 219512 676108 219521
rect 676052 219447 676108 219456
rect 676162 219109 676190 221149
rect 676244 220770 676300 220779
rect 676244 220705 676300 220714
rect 676258 219257 676286 220705
rect 676246 219251 676298 219257
rect 676246 219193 676298 219199
rect 676150 219103 676202 219109
rect 676150 219045 676202 219051
rect 676916 216774 676972 216783
rect 676916 216709 676972 216718
rect 675764 216478 675820 216487
rect 675764 216413 675820 216422
rect 675094 216069 675146 216075
rect 675094 216011 675146 216017
rect 674710 213331 674762 213337
rect 674710 213273 674762 213279
rect 674518 212147 674570 212153
rect 674518 212089 674570 212095
rect 674530 197205 674558 212089
rect 674614 210445 674666 210451
rect 674614 210387 674666 210393
rect 674518 197199 674570 197205
rect 674518 197141 674570 197147
rect 674626 196188 674654 210387
rect 674722 201349 674750 213273
rect 674806 213257 674858 213263
rect 674806 213199 674858 213205
rect 674818 202089 674846 213199
rect 674902 210371 674954 210377
rect 674902 210313 674954 210319
rect 674806 202083 674858 202089
rect 674806 202025 674858 202031
rect 674710 201343 674762 201349
rect 674710 201285 674762 201291
rect 674914 197372 674942 210313
rect 674998 210297 675050 210303
rect 674998 210239 675050 210245
rect 675010 200369 675038 210239
rect 675106 205808 675134 216011
rect 675286 213183 675338 213189
rect 675286 213125 675338 213131
rect 675106 205780 675230 205808
rect 675094 205709 675146 205715
rect 675094 205651 675146 205657
rect 675106 201571 675134 205651
rect 675202 202182 675230 205780
rect 675298 204698 675326 213125
rect 675778 206159 675806 216413
rect 676052 216108 676108 216117
rect 676052 216043 676054 216052
rect 676106 216043 676108 216052
rect 676054 216011 676106 216017
rect 676820 214850 676876 214859
rect 676820 214785 676876 214794
rect 676052 214628 676108 214637
rect 676052 214563 676108 214572
rect 675956 214110 676012 214119
rect 675956 214045 676012 214054
rect 675970 213263 675998 214045
rect 675958 213257 676010 213263
rect 675958 213199 676010 213205
rect 676066 213189 676094 214563
rect 676244 213370 676300 213379
rect 676244 213305 676246 213314
rect 676298 213305 676300 213314
rect 676246 213273 676298 213279
rect 676054 213183 676106 213189
rect 676054 213125 676106 213131
rect 676052 212630 676108 212639
rect 676052 212565 676108 212574
rect 676066 212153 676094 212565
rect 676054 212147 676106 212153
rect 676054 212089 676106 212095
rect 676052 212038 676108 212047
rect 676052 211973 676108 211982
rect 675956 211076 676012 211085
rect 675956 211011 676012 211020
rect 675970 210451 675998 211011
rect 675958 210445 676010 210451
rect 675958 210387 676010 210393
rect 676066 210303 676094 211973
rect 676244 211446 676300 211455
rect 676244 211381 676300 211390
rect 676258 210377 676286 211381
rect 676246 210371 676298 210377
rect 676246 210313 676298 210319
rect 676054 210297 676106 210303
rect 676054 210239 676106 210245
rect 676834 207607 676862 214785
rect 676820 207598 676876 207607
rect 676820 207533 676876 207542
rect 676930 207459 676958 216709
rect 679796 210706 679852 210715
rect 679796 210641 679852 210650
rect 679810 209827 679838 210641
rect 679796 209818 679852 209827
rect 679796 209753 679852 209762
rect 685460 209818 685516 209827
rect 685460 209753 685516 209762
rect 676916 207450 676972 207459
rect 679810 207417 679838 209753
rect 685474 209383 685502 209753
rect 685460 209374 685516 209383
rect 685460 209309 685516 209318
rect 676916 207385 676972 207394
rect 679798 207411 679850 207417
rect 679798 207353 679850 207359
rect 675766 206153 675818 206159
rect 675766 206095 675818 206101
rect 675490 205715 675518 205868
rect 675478 205709 675530 205715
rect 675478 205651 675530 205657
rect 675766 205635 675818 205641
rect 675766 205577 675818 205583
rect 675778 205350 675806 205577
rect 675298 204670 675408 204698
rect 675668 204490 675724 204499
rect 675668 204425 675724 204434
rect 675682 204018 675710 204425
rect 675298 202228 675422 202256
rect 675298 202182 675326 202228
rect 675202 202154 675326 202182
rect 675394 202168 675422 202228
rect 675190 202083 675242 202089
rect 675190 202025 675242 202031
rect 675202 201664 675230 202025
rect 675202 201636 675408 201664
rect 675094 201565 675146 201571
rect 675094 201507 675146 201513
rect 675382 201343 675434 201349
rect 675382 201285 675434 201291
rect 675394 200984 675422 201285
rect 675010 200341 675408 200369
rect 675764 198422 675820 198431
rect 675764 198357 675820 198366
rect 675778 197876 675806 198357
rect 674914 197344 675038 197372
rect 675010 197333 675038 197344
rect 675010 197305 675408 197333
rect 675190 197199 675242 197205
rect 675190 197141 675242 197147
rect 675202 196706 675230 197141
rect 675202 196678 675326 196706
rect 675298 196632 675326 196678
rect 675394 196632 675422 196692
rect 675298 196604 675422 196632
rect 674626 196160 675038 196188
rect 675010 196040 675038 196160
rect 675010 196012 675408 196040
rect 675092 194870 675148 194879
rect 675148 194828 675408 194856
rect 675092 194805 675148 194814
rect 675764 193538 675820 193547
rect 675764 193473 675820 193482
rect 675778 192992 675806 193473
rect 675764 191614 675820 191623
rect 675764 191549 675820 191558
rect 675778 191142 675806 191549
rect 676148 177406 676204 177415
rect 676148 177341 676204 177350
rect 676162 176189 676190 177341
rect 676340 176814 676396 176823
rect 676340 176749 676396 176758
rect 676244 176370 676300 176379
rect 676244 176305 676300 176314
rect 676150 176183 676202 176189
rect 676150 176125 676202 176131
rect 676258 176041 676286 176305
rect 676246 176035 676298 176041
rect 676246 175977 676298 175983
rect 676354 175893 676382 176749
rect 676342 175887 676394 175893
rect 676342 175829 676394 175835
rect 672596 173558 672652 173567
rect 672596 173493 672652 173502
rect 675572 172078 675628 172087
rect 675572 172013 675628 172022
rect 675286 169967 675338 169973
rect 675286 169909 675338 169915
rect 674998 167155 675050 167161
rect 674998 167097 675050 167103
rect 670390 160495 670442 160501
rect 670390 160437 670442 160443
rect 670402 155543 670430 160437
rect 675010 156524 675038 167097
rect 675190 167081 675242 167087
rect 675106 167029 675190 167054
rect 675106 167026 675242 167029
rect 675106 156672 675134 167026
rect 675190 167023 675242 167026
rect 675298 159706 675326 169909
rect 675586 167054 675614 172013
rect 676052 170228 676108 170237
rect 676052 170163 676108 170172
rect 676066 169973 676094 170163
rect 676054 169967 676106 169973
rect 676054 169909 676106 169915
rect 676052 169710 676108 169719
rect 676052 169645 676108 169654
rect 676066 167087 676094 169645
rect 676244 168970 676300 168979
rect 676244 168905 676300 168914
rect 676258 167161 676286 168905
rect 676246 167155 676298 167161
rect 676246 167097 676298 167103
rect 676054 167081 676106 167087
rect 675586 167026 675710 167054
rect 675682 161167 675710 167026
rect 676054 167023 676106 167029
rect 676052 166158 676108 166167
rect 676052 166093 676108 166102
rect 676066 164201 676094 166093
rect 676148 165418 676204 165427
rect 676148 165353 676204 165362
rect 676162 164275 676190 165353
rect 676244 164826 676300 164835
rect 676244 164761 676300 164770
rect 676258 164349 676286 164761
rect 676246 164343 676298 164349
rect 676246 164285 676298 164291
rect 676150 164269 676202 164275
rect 676150 164211 676202 164217
rect 676054 164195 676106 164201
rect 676054 164137 676106 164143
rect 675670 161161 675722 161167
rect 675670 161103 675722 161109
rect 675394 160501 675422 160876
rect 675670 160643 675722 160649
rect 675670 160585 675722 160591
rect 675382 160495 675434 160501
rect 675382 160437 675434 160443
rect 675682 160323 675710 160585
rect 675298 159678 675408 159706
rect 675764 159350 675820 159359
rect 675764 159285 675820 159294
rect 675778 159026 675806 159285
rect 675476 157722 675532 157731
rect 675476 157657 675532 157666
rect 675490 157176 675518 157657
rect 675106 156644 675326 156672
rect 675298 156524 675326 156644
rect 675394 156524 675422 156658
rect 675010 156496 675230 156524
rect 675298 156496 675422 156524
rect 675202 156006 675230 156496
rect 675202 155978 675408 156006
rect 670390 155537 670442 155543
rect 670390 155479 670442 155485
rect 675764 155502 675820 155511
rect 675764 155437 675820 155446
rect 675092 155354 675148 155363
rect 675778 155355 675806 155437
rect 675092 155289 675148 155298
rect 675106 152898 675134 155289
rect 675106 152870 675408 152898
rect 675188 152542 675244 152551
rect 675188 152477 675244 152486
rect 675668 152542 675724 152551
rect 675668 152477 675724 152486
rect 675202 151714 675230 152477
rect 675682 152292 675710 152477
rect 675202 151686 675326 151714
rect 675298 151640 675326 151686
rect 675394 151640 675422 151700
rect 675298 151612 675422 151640
rect 675764 151358 675820 151367
rect 675764 151293 675820 151302
rect 675778 151034 675806 151293
rect 675476 150322 675532 150331
rect 675476 150257 675532 150266
rect 675490 149850 675518 150257
rect 675092 149730 675148 149739
rect 675092 149665 675148 149674
rect 675106 148014 675134 149665
rect 675106 147986 675408 148014
rect 675764 146622 675820 146631
rect 675764 146557 675820 146566
rect 675778 146150 675806 146557
rect 676148 131822 676204 131831
rect 676148 131757 676204 131766
rect 676162 130161 676190 131757
rect 676340 131230 676396 131239
rect 676340 131165 676396 131174
rect 676244 130786 676300 130795
rect 676244 130721 676300 130730
rect 676150 130155 676202 130161
rect 676150 130097 676202 130103
rect 676258 130013 676286 130721
rect 676246 130007 676298 130013
rect 676246 129949 676298 129955
rect 676354 129865 676382 131165
rect 676342 129859 676394 129865
rect 676342 129801 676394 129807
rect 676244 129750 676300 129759
rect 676244 129685 676300 129694
rect 676258 129643 676286 129685
rect 676246 129637 676298 129643
rect 676246 129579 676298 129585
rect 676148 128862 676204 128871
rect 676148 128797 676204 128806
rect 676052 127604 676108 127613
rect 676052 127539 676108 127548
rect 676066 126757 676094 127539
rect 676162 126831 676190 128797
rect 676244 127826 676300 127835
rect 676244 127761 676300 127770
rect 676258 126905 676286 127761
rect 676246 126899 676298 126905
rect 676246 126841 676298 126847
rect 676150 126825 676202 126831
rect 676150 126767 676202 126773
rect 676916 126790 676972 126799
rect 674134 126751 674186 126757
rect 674134 126693 674186 126699
rect 676054 126751 676106 126757
rect 676916 126725 676972 126734
rect 676054 126693 676106 126699
rect 674038 124087 674090 124093
rect 674038 124029 674090 124035
rect 665302 115281 665354 115287
rect 665302 115223 665354 115229
rect 663766 115207 663818 115213
rect 663766 115149 663818 115155
rect 665206 115207 665258 115213
rect 665206 115149 665258 115155
rect 646484 113174 646540 113183
rect 646484 113109 646540 113118
rect 186164 107846 186220 107855
rect 186164 107781 186220 107790
rect 184436 107106 184492 107115
rect 184436 107041 184492 107050
rect 182998 106549 183050 106555
rect 182998 106491 183050 106497
rect 184534 106549 184586 106555
rect 184534 106491 184586 106497
rect 184342 106475 184394 106481
rect 184342 106417 184394 106423
rect 179926 106401 179978 106407
rect 179926 106343 179978 106349
rect 184354 105635 184382 106417
rect 184438 106327 184490 106333
rect 184438 106269 184490 106275
rect 184340 105626 184396 105635
rect 184340 105561 184396 105570
rect 184450 104007 184478 106269
rect 184546 104895 184574 106491
rect 185302 106401 185354 106407
rect 185300 106366 185302 106375
rect 185354 106366 185356 106375
rect 185300 106301 185356 106310
rect 646100 106070 646156 106079
rect 646100 106005 646156 106014
rect 184726 105143 184778 105149
rect 184726 105085 184778 105091
rect 184532 104886 184588 104895
rect 184532 104821 184588 104830
rect 184436 103998 184492 104007
rect 184436 103933 184492 103942
rect 184438 103663 184490 103669
rect 184438 103605 184490 103611
rect 184342 103441 184394 103447
rect 184450 103415 184478 103605
rect 184630 103589 184682 103595
rect 184630 103531 184682 103537
rect 184534 103515 184586 103521
rect 184534 103457 184586 103463
rect 184342 103383 184394 103389
rect 184436 103406 184492 103415
rect 184354 102527 184382 103383
rect 184436 103341 184492 103350
rect 184340 102518 184396 102527
rect 184340 102453 184396 102462
rect 184546 101935 184574 103457
rect 184532 101926 184588 101935
rect 184532 101861 184588 101870
rect 184642 101047 184670 103531
rect 184628 101038 184684 101047
rect 184628 100973 184684 100982
rect 184438 100777 184490 100783
rect 184438 100719 184490 100725
rect 184342 100555 184394 100561
rect 184342 100497 184394 100503
rect 184354 100307 184382 100497
rect 184340 100298 184396 100307
rect 184340 100233 184396 100242
rect 184450 99567 184478 100719
rect 184534 100703 184586 100709
rect 184534 100645 184586 100651
rect 184436 99558 184492 99567
rect 184436 99493 184492 99502
rect 184546 98679 184574 100645
rect 184630 100629 184682 100635
rect 184630 100571 184682 100577
rect 184532 98670 184588 98679
rect 184532 98605 184588 98614
rect 184642 98087 184670 100571
rect 184628 98078 184684 98087
rect 184246 98039 184298 98045
rect 184628 98013 184684 98022
rect 184246 97981 184298 97987
rect 179926 95079 179978 95085
rect 179926 95021 179978 95027
rect 177142 91897 177194 91903
rect 177142 91839 177194 91845
rect 171286 83461 171338 83467
rect 171286 83403 171338 83409
rect 165238 80501 165290 80507
rect 165238 80443 165290 80449
rect 179938 80433 179966 95021
rect 184258 81955 184286 97981
rect 184438 97891 184490 97897
rect 184438 97833 184490 97839
rect 184342 97817 184394 97823
rect 184342 97759 184394 97765
rect 184354 97199 184382 97759
rect 184340 97190 184396 97199
rect 184340 97125 184396 97134
rect 184450 96459 184478 97833
rect 184436 96450 184492 96459
rect 184436 96385 184492 96394
rect 184738 95719 184766 105085
rect 646114 103891 646142 106005
rect 646102 103885 646154 103891
rect 646102 103827 646154 103833
rect 643606 103737 643658 103743
rect 643606 103679 643658 103685
rect 186166 97965 186218 97971
rect 186166 97907 186218 97913
rect 184724 95710 184780 95719
rect 184724 95645 184780 95654
rect 184630 95005 184682 95011
rect 184630 94947 184682 94953
rect 184534 94931 184586 94937
rect 184534 94873 184586 94879
rect 184438 94857 184490 94863
rect 184340 94822 184396 94831
rect 184438 94799 184490 94805
rect 184340 94757 184342 94766
rect 184394 94757 184396 94766
rect 184342 94725 184394 94731
rect 184450 94239 184478 94799
rect 184436 94230 184492 94239
rect 184436 94165 184492 94174
rect 184546 93499 184574 94873
rect 184532 93490 184588 93499
rect 184532 93425 184588 93434
rect 184642 92759 184670 94947
rect 184628 92750 184684 92759
rect 184628 92685 184684 92694
rect 184438 92119 184490 92125
rect 184438 92061 184490 92067
rect 184340 92010 184396 92019
rect 184340 91945 184342 91954
rect 184394 91945 184396 91954
rect 184342 91913 184394 91919
rect 184450 90391 184478 92061
rect 184534 92045 184586 92051
rect 184534 91987 184586 91993
rect 184436 90382 184492 90391
rect 184436 90317 184492 90326
rect 184546 89651 184574 91987
rect 184630 91897 184682 91903
rect 184630 91839 184682 91845
rect 184642 91131 184670 91839
rect 184628 91122 184684 91131
rect 184628 91057 184684 91066
rect 184532 89642 184588 89651
rect 184532 89577 184588 89586
rect 184534 89233 184586 89239
rect 184534 89175 184586 89181
rect 184438 89085 184490 89091
rect 184438 89027 184490 89033
rect 184342 89011 184394 89017
rect 184342 88953 184394 88959
rect 184354 88911 184382 88953
rect 184340 88902 184396 88911
rect 184340 88837 184396 88846
rect 184450 88171 184478 89027
rect 184436 88162 184492 88171
rect 184436 88097 184492 88106
rect 184546 87283 184574 89175
rect 184630 89159 184682 89165
rect 184630 89101 184682 89107
rect 184532 87274 184588 87283
rect 184532 87209 184588 87218
rect 184642 86691 184670 89101
rect 184628 86682 184684 86691
rect 184628 86617 184684 86626
rect 184438 86421 184490 86427
rect 184438 86363 184490 86369
rect 184342 86273 184394 86279
rect 184342 86215 184394 86221
rect 184354 85211 184382 86215
rect 184450 85803 184478 86363
rect 184534 86347 184586 86353
rect 184534 86289 184586 86295
rect 184436 85794 184492 85803
rect 184436 85729 184492 85738
rect 184340 85202 184396 85211
rect 184340 85137 184396 85146
rect 184546 84323 184574 86289
rect 184532 84314 184588 84323
rect 184532 84249 184588 84258
rect 184438 83535 184490 83541
rect 184438 83477 184490 83483
rect 184342 83461 184394 83467
rect 184340 83426 184342 83435
rect 184394 83426 184396 83435
rect 184340 83361 184396 83370
rect 184244 81946 184300 81955
rect 184244 81881 184300 81890
rect 184450 81363 184478 83477
rect 186178 82843 186206 97907
rect 643618 85021 643646 103679
rect 645140 102222 645196 102231
rect 645140 102157 645196 102166
rect 645154 102115 645182 102157
rect 645142 102109 645194 102115
rect 645142 102051 645194 102057
rect 645428 96006 645484 96015
rect 645428 95941 645430 95950
rect 645482 95941 645484 95950
rect 645430 95909 645482 95915
rect 646390 92415 646442 92421
rect 646390 92357 646442 92363
rect 645908 88902 645964 88911
rect 645908 88837 645964 88846
rect 645922 87537 645950 88837
rect 645910 87531 645962 87537
rect 645910 87473 645962 87479
rect 640726 85015 640778 85021
rect 640726 84957 640778 84963
rect 643606 85015 643658 85021
rect 643606 84957 643658 84963
rect 186164 82834 186220 82843
rect 186164 82769 186220 82778
rect 184436 81354 184492 81363
rect 184436 81289 184492 81298
rect 184438 80649 184490 80655
rect 184438 80591 184490 80597
rect 184342 80501 184394 80507
rect 184342 80443 184394 80449
rect 179926 80427 179978 80433
rect 179926 80369 179978 80375
rect 184354 78995 184382 80443
rect 184450 79883 184478 80591
rect 184534 80575 184586 80581
rect 184534 80517 184586 80523
rect 184436 79874 184492 79883
rect 184436 79809 184492 79818
rect 184340 78986 184396 78995
rect 184340 78921 184396 78930
rect 184546 78255 184574 80517
rect 184628 80466 184684 80475
rect 184628 80401 184630 80410
rect 184682 80401 184684 80410
rect 184630 80369 184682 80375
rect 184532 78246 184588 78255
rect 184532 78181 184588 78190
rect 184630 77763 184682 77769
rect 184630 77705 184682 77711
rect 184438 77689 184490 77695
rect 184438 77631 184490 77637
rect 159766 77541 159818 77547
rect 159766 77483 159818 77489
rect 184342 77541 184394 77547
rect 184450 77515 184478 77631
rect 184534 77615 184586 77621
rect 184534 77557 184586 77563
rect 184342 77483 184394 77489
rect 184436 77506 184492 77515
rect 184354 76775 184382 77483
rect 184436 77441 184492 77450
rect 184340 76766 184396 76775
rect 184340 76701 184396 76710
rect 184546 75147 184574 77557
rect 184642 76035 184670 77705
rect 184628 76026 184684 76035
rect 184628 75961 184684 75970
rect 184532 75138 184588 75147
rect 184532 75073 184588 75082
rect 184534 74877 184586 74883
rect 184534 74819 184586 74825
rect 184438 74729 184490 74735
rect 184438 74671 184490 74677
rect 154102 74655 154154 74661
rect 154102 74597 154154 74603
rect 184342 74655 184394 74661
rect 184342 74597 184394 74603
rect 184354 74407 184382 74597
rect 184340 74398 184396 74407
rect 184340 74333 184396 74342
rect 149684 73066 149740 73075
rect 149684 73001 149740 73010
rect 149590 71843 149642 71849
rect 149590 71785 149642 71791
rect 149506 70952 149630 70980
rect 149492 70846 149548 70855
rect 149492 70781 149548 70790
rect 149396 69514 149452 69523
rect 149396 69449 149452 69458
rect 149302 68957 149354 68963
rect 149302 68899 149354 68905
rect 149206 68883 149258 68889
rect 149206 68825 149258 68831
rect 149300 68330 149356 68339
rect 149300 68265 149356 68274
rect 149204 67146 149260 67155
rect 149204 67081 149260 67090
rect 149110 66219 149162 66225
rect 149110 66161 149162 66167
rect 149218 63191 149246 67081
rect 149314 63339 149342 68265
rect 149410 66003 149438 69449
rect 149506 66077 149534 70781
rect 149602 69111 149630 70952
rect 149590 69105 149642 69111
rect 149590 69047 149642 69053
rect 149698 66151 149726 73001
rect 184450 72927 184478 74671
rect 184546 73667 184574 74819
rect 184630 74803 184682 74809
rect 184630 74745 184682 74751
rect 184532 73658 184588 73667
rect 184532 73593 184588 73602
rect 184436 72918 184492 72927
rect 184436 72853 184492 72862
rect 184642 72187 184670 74745
rect 184628 72178 184684 72187
rect 184628 72113 184684 72122
rect 184342 71991 184394 71997
rect 184342 71933 184394 71939
rect 184354 71447 184382 71933
rect 184438 71917 184490 71923
rect 184438 71859 184490 71865
rect 184340 71438 184396 71447
rect 184340 71373 184396 71382
rect 184450 70559 184478 71859
rect 184534 71843 184586 71849
rect 184534 71785 184586 71791
rect 184436 70550 184492 70559
rect 184436 70485 184492 70494
rect 184546 69967 184574 71785
rect 184532 69958 184588 69967
rect 184532 69893 184588 69902
rect 184534 69105 184586 69111
rect 184340 69070 184396 69079
rect 184534 69047 184586 69053
rect 184340 69005 184342 69014
rect 184394 69005 184396 69014
rect 184342 68973 184394 68979
rect 184438 68957 184490 68963
rect 184438 68899 184490 68905
rect 184342 68883 184394 68889
rect 184342 68825 184394 68831
rect 184354 68487 184382 68825
rect 184340 68478 184396 68487
rect 184340 68413 184396 68422
rect 184450 66859 184478 68899
rect 184546 67599 184574 69047
rect 184532 67590 184588 67599
rect 184532 67525 184588 67534
rect 184436 66850 184492 66859
rect 184436 66785 184492 66794
rect 184534 66219 184586 66225
rect 184534 66161 184586 66167
rect 149686 66145 149738 66151
rect 184342 66145 184394 66151
rect 149686 66087 149738 66093
rect 184340 66110 184342 66119
rect 184394 66110 184396 66119
rect 149494 66071 149546 66077
rect 184340 66045 184396 66054
rect 184438 66071 184490 66077
rect 149494 66013 149546 66019
rect 184438 66013 184490 66019
rect 149398 65997 149450 66003
rect 149398 65939 149450 65945
rect 184342 65997 184394 66003
rect 184342 65939 184394 65945
rect 149396 65370 149452 65379
rect 149396 65305 149452 65314
rect 149302 63333 149354 63339
rect 149302 63275 149354 63281
rect 149410 63265 149438 65305
rect 149492 64630 149548 64639
rect 149492 64565 149548 64574
rect 149398 63259 149450 63265
rect 149398 63201 149450 63207
rect 149206 63185 149258 63191
rect 149206 63127 149258 63133
rect 149506 63117 149534 64565
rect 184354 63751 184382 65939
rect 184450 64639 184478 66013
rect 184546 65231 184574 66161
rect 184532 65222 184588 65231
rect 184532 65157 184588 65166
rect 184436 64630 184492 64639
rect 184436 64565 184492 64574
rect 184340 63742 184396 63751
rect 184340 63677 184396 63686
rect 149588 63446 149644 63455
rect 149588 63381 149644 63390
rect 149494 63111 149546 63117
rect 149494 63053 149546 63059
rect 149396 62262 149452 62271
rect 149396 62197 149452 62206
rect 149300 60634 149356 60643
rect 149300 60569 149356 60578
rect 149314 60305 149342 60569
rect 149410 60453 149438 62197
rect 149398 60447 149450 60453
rect 149398 60389 149450 60395
rect 149602 60379 149630 63381
rect 184438 63333 184490 63339
rect 184438 63275 184490 63281
rect 184342 63185 184394 63191
rect 184450 63159 184478 63275
rect 184630 63259 184682 63265
rect 184630 63201 184682 63207
rect 184342 63127 184394 63133
rect 184436 63150 184492 63159
rect 184354 62271 184382 63127
rect 184436 63085 184492 63094
rect 184534 63111 184586 63117
rect 184534 63053 184586 63059
rect 184340 62262 184396 62271
rect 184340 62197 184396 62206
rect 184546 60791 184574 63053
rect 184642 61531 184670 63201
rect 184628 61522 184684 61531
rect 184628 61457 184684 61466
rect 184532 60782 184588 60791
rect 184532 60717 184588 60726
rect 184438 60447 184490 60453
rect 184438 60389 184490 60395
rect 149590 60373 149642 60379
rect 149590 60315 149642 60321
rect 184342 60373 184394 60379
rect 184342 60315 184394 60321
rect 149302 60299 149354 60305
rect 149302 60241 149354 60247
rect 184354 60051 184382 60315
rect 184340 60042 184396 60051
rect 184340 59977 184396 59986
rect 149396 59746 149452 59755
rect 149396 59681 149452 59690
rect 149410 59047 149438 59681
rect 184450 59311 184478 60389
rect 184534 60299 184586 60305
rect 184534 60241 184586 60247
rect 184436 59302 184492 59311
rect 184436 59237 184492 59246
rect 149398 59041 149450 59047
rect 149398 58983 149450 58989
rect 184342 59041 184394 59047
rect 184342 58983 184394 58989
rect 149396 58562 149452 58571
rect 149396 58497 149452 58506
rect 149410 57567 149438 58497
rect 184354 57683 184382 58983
rect 184546 58423 184574 60241
rect 184532 58414 184588 58423
rect 184532 58349 184588 58358
rect 184340 57674 184396 57683
rect 184340 57609 184396 57618
rect 149398 57561 149450 57567
rect 149398 57503 149450 57509
rect 184342 57561 184394 57567
rect 184342 57503 184394 57509
rect 149492 57378 149548 57387
rect 149492 57313 149548 57322
rect 149506 56235 149534 57313
rect 184354 56943 184382 57503
rect 184340 56934 184396 56943
rect 184340 56869 184396 56878
rect 149494 56229 149546 56235
rect 149396 56194 149452 56203
rect 184342 56229 184394 56235
rect 149494 56171 149546 56177
rect 184340 56194 184342 56203
rect 184394 56194 184396 56203
rect 149396 56129 149398 56138
rect 149450 56129 149452 56138
rect 184340 56129 184396 56138
rect 184438 56155 184490 56161
rect 149398 56097 149450 56103
rect 184438 56097 184490 56103
rect 184450 55463 184478 56097
rect 184436 55454 184492 55463
rect 184436 55389 184492 55398
rect 149684 54862 149740 54871
rect 149684 54797 149740 54806
rect 149698 54681 149726 54797
rect 184340 54714 184396 54723
rect 149686 54675 149738 54681
rect 184340 54649 184342 54658
rect 149686 54617 149738 54623
rect 184394 54649 184396 54658
rect 184342 54617 184394 54623
rect 184340 53974 184396 53983
rect 184340 53909 184396 53918
rect 149396 53826 149452 53835
rect 149396 53761 149452 53770
rect 149410 53275 149438 53761
rect 184354 53275 184382 53909
rect 149398 53269 149450 53275
rect 149398 53211 149450 53217
rect 184342 53269 184394 53275
rect 184342 53211 184394 53217
rect 145104 49788 145406 49816
rect 145378 47133 145406 49788
rect 199138 47133 199166 53650
rect 145366 47127 145418 47133
rect 145366 47069 145418 47075
rect 199126 47127 199178 47133
rect 199126 47069 199178 47075
rect 142114 46680 142416 46708
rect 142114 40367 142142 46680
rect 216418 46171 216446 53650
rect 233698 47651 233726 53650
rect 233686 47645 233738 47651
rect 233686 47587 233738 47593
rect 250978 47577 251006 53650
rect 268320 53636 268574 53664
rect 285600 53636 285854 53664
rect 268546 47725 268574 53636
rect 285826 47799 285854 53636
rect 302914 47873 302942 53650
rect 311158 48089 311210 48095
rect 311158 48031 311210 48037
rect 311062 48015 311114 48021
rect 311062 47957 311114 47963
rect 302902 47867 302954 47873
rect 302902 47809 302954 47815
rect 285814 47793 285866 47799
rect 285814 47735 285866 47741
rect 268534 47719 268586 47725
rect 268534 47661 268586 47667
rect 250966 47571 251018 47577
rect 250966 47513 251018 47519
rect 207382 46165 207434 46171
rect 207382 46107 207434 46113
rect 216406 46165 216458 46171
rect 216406 46107 216458 46113
rect 145078 41873 145130 41879
rect 145078 41815 145130 41821
rect 142100 40358 142156 40367
rect 142100 40293 142156 40302
rect 145090 40196 145118 41815
rect 187344 41805 187646 41824
rect 194064 41805 194366 41824
rect 187344 41799 187658 41805
rect 187344 41796 187606 41799
rect 194064 41799 194378 41805
rect 194064 41796 194326 41799
rect 187606 41741 187658 41747
rect 194326 41741 194378 41747
rect 207394 41509 207422 46107
rect 311074 42268 311102 47957
rect 310498 42240 311102 42268
rect 302900 42134 302956 42143
rect 302688 42092 302900 42120
rect 310498 42120 310526 42240
rect 311170 42143 311198 48031
rect 320194 47947 320222 53650
rect 320182 47941 320234 47947
rect 320182 47883 320234 47889
rect 337474 46985 337502 53650
rect 354850 48095 354878 53650
rect 371938 53636 372192 53664
rect 389218 53636 389472 53664
rect 354838 48089 354890 48095
rect 354838 48031 354890 48037
rect 371938 48021 371966 53636
rect 371926 48015 371978 48021
rect 371926 47957 371978 47963
rect 334102 46979 334154 46985
rect 334102 46921 334154 46927
rect 337462 46979 337514 46985
rect 337462 46921 337514 46927
rect 310128 42092 310526 42120
rect 311156 42134 311212 42143
rect 302900 42069 302956 42078
rect 311156 42069 311212 42078
rect 307008 41953 307262 41972
rect 307008 41947 307274 41953
rect 307008 41944 307222 41947
rect 307222 41889 307274 41895
rect 311062 41947 311114 41953
rect 311062 41889 311114 41895
rect 207382 41503 207434 41509
rect 207382 41445 207434 41451
rect 145090 40168 145131 40196
rect 145103 39960 145131 40168
rect 311074 37259 311102 41889
rect 334114 37259 334142 46921
rect 365314 42240 365726 42268
rect 365314 42120 365342 42240
rect 364944 42092 365342 42120
rect 357716 41838 357772 41847
rect 357456 41796 357716 41824
rect 362036 41838 362092 41847
rect 361776 41796 362036 41824
rect 357716 41773 357772 41782
rect 365698 41824 365726 42240
rect 389218 41847 389246 53636
rect 405526 48015 405578 48021
rect 405526 47957 405578 47963
rect 403222 46387 403274 46393
rect 403222 46329 403274 46335
rect 394582 41947 394634 41953
rect 394582 41889 394634 41895
rect 389204 41838 389260 41847
rect 365698 41796 365918 41824
rect 362036 41773 362092 41782
rect 365890 37439 365918 41796
rect 389204 41773 389260 41782
rect 394594 37439 394622 41889
rect 403234 40515 403262 46329
rect 405538 42106 405566 47957
rect 406786 46393 406814 53650
rect 406774 46387 406826 46393
rect 406774 46329 406826 46335
rect 420130 42240 420446 42268
rect 412532 42134 412588 42143
rect 412272 42092 412532 42120
rect 420130 42120 420158 42240
rect 419712 42092 420158 42120
rect 412532 42069 412588 42078
rect 416852 41986 416908 41995
rect 416592 41944 416852 41972
rect 416852 41921 416908 41930
rect 420418 41824 420446 42240
rect 424066 41953 424094 53650
rect 441346 48021 441374 53650
rect 441334 48015 441386 48021
rect 441334 47957 441386 47963
rect 424054 41947 424106 41953
rect 424054 41889 424106 41895
rect 449302 41947 449354 41953
rect 449302 41889 449354 41895
rect 420418 41796 420734 41824
rect 403220 40506 403276 40515
rect 403220 40441 403276 40450
rect 420706 37439 420734 41796
rect 449314 37439 449342 41889
rect 458626 40515 458654 53650
rect 475714 53636 475968 53664
rect 492994 53636 493248 53664
rect 510370 53636 510624 53664
rect 460342 48015 460394 48021
rect 460342 47957 460394 47963
rect 460354 42106 460382 47957
rect 475222 47645 475274 47651
rect 475222 47587 475274 47593
rect 474946 42240 475166 42268
rect 474946 42120 474974 42240
rect 474528 42092 474974 42120
rect 467348 41838 467404 41847
rect 467088 41796 467348 41824
rect 471668 41838 471724 41847
rect 471408 41796 471668 41824
rect 467348 41773 467404 41782
rect 475138 41824 475166 42240
rect 475234 41953 475262 47587
rect 475606 47571 475658 47577
rect 475606 47513 475658 47519
rect 475222 41947 475274 41953
rect 475222 41889 475274 41895
rect 475138 41796 475550 41824
rect 471668 41773 471724 41782
rect 458612 40506 458668 40515
rect 458612 40441 458668 40450
rect 365878 37433 365930 37439
rect 365878 37375 365930 37381
rect 394582 37433 394634 37439
rect 394582 37375 394634 37381
rect 420694 37433 420746 37439
rect 420694 37375 420746 37381
rect 449302 37433 449354 37439
rect 449302 37375 449354 37381
rect 475522 37365 475550 41796
rect 475618 37439 475646 47513
rect 475714 40663 475742 53636
rect 492994 47651 493022 53636
rect 510370 48021 510398 53636
rect 510358 48015 510410 48021
rect 510358 47957 510410 47963
rect 521110 47867 521162 47873
rect 521110 47809 521162 47815
rect 515542 47793 515594 47799
rect 515542 47735 515594 47741
rect 503926 47719 503978 47725
rect 503926 47661 503978 47667
rect 492982 47645 493034 47651
rect 492982 47587 493034 47593
rect 503938 43285 503966 47661
rect 515554 44691 515582 47735
rect 521122 44839 521150 47809
rect 521206 47571 521258 47577
rect 521206 47513 521258 47519
rect 521110 44833 521162 44839
rect 521110 44775 521162 44781
rect 515542 44685 515594 44691
rect 515542 44627 515594 44633
rect 521218 43304 521246 47513
rect 527938 46171 527966 53650
rect 529270 47941 529322 47947
rect 529270 47883 529322 47889
rect 522838 46165 522890 46171
rect 522838 46107 522890 46113
rect 527926 46165 527978 46171
rect 527926 46107 527978 46113
rect 503926 43279 503978 43285
rect 521218 43276 521534 43304
rect 503926 43221 503978 43227
rect 520342 43205 520394 43211
rect 520342 43147 520394 43153
rect 520354 42120 520382 43147
rect 521506 42120 521534 43276
rect 520354 42092 520656 42120
rect 521506 42092 521856 42120
rect 506806 42021 506858 42027
rect 506806 41963 506858 41969
rect 475700 40654 475756 40663
rect 475700 40589 475756 40598
rect 475606 37433 475658 37439
rect 475606 37375 475658 37381
rect 506818 37365 506846 41963
rect 514882 41953 515136 41972
rect 514006 41947 514058 41953
rect 514006 41889 514058 41895
rect 514870 41947 515136 41953
rect 514922 41944 515136 41947
rect 514870 41889 514922 41895
rect 514018 37439 514046 41889
rect 522850 41847 522878 46107
rect 525910 44833 525962 44839
rect 525910 44775 525962 44781
rect 524950 44685 525002 44691
rect 524950 44627 525002 44633
rect 524962 42106 524990 44627
rect 525922 42120 525950 44775
rect 525922 42092 526176 42120
rect 529282 42106 529310 47883
rect 545218 43359 545246 53650
rect 541462 43353 541514 43359
rect 541462 43295 541514 43301
rect 545206 43353 545258 43359
rect 545206 43295 545258 43301
rect 522836 41838 522892 41847
rect 522836 41773 522892 41782
rect 541474 40515 541502 43295
rect 562498 41953 562526 53650
rect 579796 53602 579852 54402
rect 597092 53602 597148 54402
rect 614388 53602 614444 54402
rect 631684 53602 631740 54402
rect 636502 46757 636554 46763
rect 636502 46699 636554 46705
rect 562486 41947 562538 41953
rect 562486 41889 562538 41895
rect 636514 41879 636542 46699
rect 636502 41873 636554 41879
rect 636502 41815 636554 41821
rect 640738 41805 640766 84957
rect 645716 84462 645772 84471
rect 645716 84397 645772 84406
rect 645730 84207 645758 84397
rect 645718 84201 645770 84207
rect 645718 84143 645770 84149
rect 646294 75691 646346 75697
rect 646294 75633 646346 75639
rect 646306 75591 646334 75633
rect 646292 75582 646348 75591
rect 646292 75517 646348 75526
rect 646402 74894 646430 92357
rect 646498 77695 646526 113109
rect 665218 112327 665246 115149
rect 665206 112321 665258 112327
rect 665206 112263 665258 112269
rect 647156 111398 647212 111407
rect 647156 111333 647212 111342
rect 646676 109474 646732 109483
rect 646676 109409 646732 109418
rect 646690 92440 646718 109409
rect 646772 107994 646828 108003
rect 646772 107929 646828 107938
rect 646786 92717 646814 107929
rect 647060 98078 647116 98087
rect 647060 98013 647116 98022
rect 646774 92711 646826 92717
rect 646774 92653 646826 92659
rect 646594 92412 646718 92440
rect 646486 77689 646538 77695
rect 646486 77631 646538 77637
rect 646594 77621 646622 92412
rect 646678 92341 646730 92347
rect 646678 92283 646730 92289
rect 646690 79439 646718 92283
rect 646870 92267 646922 92273
rect 646870 92209 646922 92215
rect 646774 83609 646826 83615
rect 646774 83551 646826 83557
rect 646676 79430 646732 79439
rect 646676 79365 646732 79374
rect 646582 77615 646634 77621
rect 646582 77557 646634 77563
rect 646402 74866 646526 74894
rect 646004 66258 646060 66267
rect 646004 66193 646006 66202
rect 646058 66193 646060 66202
rect 646006 66161 646058 66167
rect 646006 59115 646058 59121
rect 646006 59057 646058 59063
rect 646018 59015 646046 59057
rect 646004 59006 646060 59015
rect 646004 58941 646060 58950
rect 646498 54723 646526 74866
rect 646786 57091 646814 83551
rect 646882 68635 646910 92209
rect 646966 92193 647018 92199
rect 646966 92135 647018 92141
rect 646978 71891 647006 92135
rect 647074 77769 647102 98013
rect 647170 87093 647198 111333
rect 665204 105626 665260 105635
rect 665204 105561 665260 105570
rect 665218 104557 665246 105561
rect 665314 105191 665342 115223
rect 674050 111735 674078 124029
rect 674146 114177 674174 126693
rect 676244 126346 676300 126355
rect 676244 126281 676300 126290
rect 676052 126124 676108 126133
rect 676052 126059 676108 126068
rect 676066 124685 676094 126059
rect 674326 124679 674378 124685
rect 674326 124621 674378 124627
rect 676054 124679 676106 124685
rect 676054 124621 676106 124627
rect 674230 121127 674282 121133
rect 674230 121069 674282 121075
rect 674134 114171 674186 114177
rect 674134 114113 674186 114119
rect 674038 111729 674090 111735
rect 674038 111671 674090 111677
rect 674242 110107 674270 121069
rect 674338 112549 674366 124621
rect 676052 124570 676108 124579
rect 676052 124505 676108 124514
rect 675956 124126 676012 124135
rect 675956 124061 675958 124070
rect 676010 124061 676012 124070
rect 675958 124029 676010 124035
rect 676066 124019 676094 124505
rect 674422 124013 674474 124019
rect 674422 123955 674474 123961
rect 676054 124013 676106 124019
rect 676054 123955 676106 123961
rect 674434 114991 674462 123955
rect 676258 123945 676286 126281
rect 676820 124866 676876 124875
rect 676820 124801 676876 124810
rect 675094 123939 675146 123945
rect 675094 123881 675146 123887
rect 676246 123939 676298 123945
rect 676246 123881 676298 123887
rect 674614 122163 674666 122169
rect 674614 122105 674666 122111
rect 674518 121201 674570 121207
rect 674518 121143 674570 121149
rect 674422 114985 674474 114991
rect 674422 114927 674474 114933
rect 674326 112543 674378 112549
rect 674326 112485 674378 112491
rect 674530 112179 674558 121143
rect 674626 114621 674654 122105
rect 674806 121053 674858 121059
rect 674806 120995 674858 121001
rect 674818 115214 674846 120995
rect 675106 115528 675134 123881
rect 676052 123534 676108 123543
rect 676052 123469 676108 123478
rect 676066 122169 676094 123469
rect 676054 122163 676106 122169
rect 676054 122105 676106 122111
rect 676052 122054 676108 122063
rect 676052 121989 676108 121998
rect 676066 121207 676094 121989
rect 676244 121462 676300 121471
rect 676244 121397 676300 121406
rect 676054 121201 676106 121207
rect 676054 121143 676106 121149
rect 676258 121133 676286 121397
rect 676246 121127 676298 121133
rect 676052 121092 676108 121101
rect 676246 121069 676298 121075
rect 676052 121027 676054 121036
rect 676106 121027 676108 121036
rect 676054 120995 676106 121001
rect 676052 120574 676108 120583
rect 676052 120509 676108 120518
rect 676066 118173 676094 120509
rect 676148 119834 676204 119843
rect 676148 119769 676204 119778
rect 676162 118247 676190 119769
rect 676244 119242 676300 119251
rect 676244 119177 676300 119186
rect 676258 118395 676286 119177
rect 676246 118389 676298 118395
rect 676246 118331 676298 118337
rect 676150 118241 676202 118247
rect 676150 118183 676202 118189
rect 676054 118167 676106 118173
rect 676054 118109 676106 118115
rect 676834 118067 676862 124801
rect 676820 118058 676876 118067
rect 676820 117993 676876 118002
rect 676930 117919 676958 126725
rect 676916 117910 676972 117919
rect 676916 117845 676972 117854
rect 675298 115648 675408 115676
rect 675106 115500 675230 115528
rect 675094 115429 675146 115435
rect 675094 115371 675146 115377
rect 674818 115186 675038 115214
rect 674614 114615 674666 114621
rect 674614 114557 674666 114563
rect 674518 112173 674570 112179
rect 674518 112115 674570 112121
rect 674230 110101 674282 110107
rect 674230 110043 674282 110049
rect 675010 105834 675038 115186
rect 675106 112327 675134 115371
rect 675202 115158 675230 115500
rect 675298 115435 675326 115648
rect 675286 115429 675338 115435
rect 675286 115371 675338 115377
rect 675202 115130 675326 115158
rect 675298 115084 675326 115130
rect 675394 115084 675422 115144
rect 675298 115056 675422 115084
rect 675190 114985 675242 114991
rect 675190 114927 675242 114933
rect 675202 114492 675230 114927
rect 675202 114464 675408 114492
rect 675286 114393 675338 114399
rect 675286 114335 675338 114341
rect 675094 112321 675146 112327
rect 675094 112263 675146 112269
rect 675094 112173 675146 112179
rect 675094 112115 675146 112121
rect 675106 110169 675134 112115
rect 675298 111384 675326 114335
rect 675382 114171 675434 114177
rect 675382 114113 675434 114119
rect 675394 113812 675422 114113
rect 675382 112543 675434 112549
rect 675382 112485 675434 112491
rect 675394 111995 675422 112485
rect 675382 111729 675434 111735
rect 675382 111671 675434 111677
rect 675394 111444 675422 111671
rect 675298 111356 675422 111384
rect 675394 110778 675422 111356
rect 675106 110141 675408 110169
rect 675094 110101 675146 110107
rect 675094 110043 675146 110049
rect 675106 107133 675134 110043
rect 675188 107698 675244 107707
rect 675244 107656 675408 107684
rect 675188 107633 675244 107642
rect 675106 107105 675408 107133
rect 675092 106514 675148 106523
rect 675148 106472 675408 106500
rect 675092 106449 675148 106458
rect 675010 105806 675408 105834
rect 675092 105626 675148 105635
rect 675092 105561 675148 105570
rect 665588 105330 665644 105339
rect 665588 105265 665644 105274
rect 665300 105182 665356 105191
rect 665300 105117 665356 105126
rect 654070 104551 654122 104557
rect 654070 104493 654122 104499
rect 665206 104551 665258 104557
rect 665206 104493 665258 104499
rect 647924 104146 647980 104155
rect 647924 104081 647980 104090
rect 647938 103965 647966 104081
rect 647926 103959 647978 103965
rect 647926 103901 647978 103907
rect 652438 102109 652490 102115
rect 652438 102051 652490 102057
rect 647924 99706 647980 99715
rect 647924 99641 647980 99650
rect 647938 97971 647966 99641
rect 647926 97965 647978 97971
rect 647926 97907 647978 97913
rect 647732 94082 647788 94091
rect 647732 94017 647788 94026
rect 647158 87087 647210 87093
rect 647158 87029 647210 87035
rect 647746 81617 647774 94017
rect 647828 92750 647884 92759
rect 647828 92685 647884 92694
rect 647842 81839 647870 92685
rect 650902 87531 650954 87537
rect 650902 87473 650954 87479
rect 647926 87309 647978 87315
rect 647926 87251 647978 87257
rect 647938 87135 647966 87251
rect 647924 87126 647980 87135
rect 647924 87061 647980 87070
rect 650914 86247 650942 87473
rect 650900 86238 650956 86247
rect 650900 86173 650956 86182
rect 652340 85350 652396 85359
rect 652340 85285 652396 85294
rect 652244 83426 652300 83435
rect 652244 83361 652300 83370
rect 647924 82686 647980 82695
rect 647924 82621 647980 82630
rect 647938 81913 647966 82621
rect 647926 81907 647978 81913
rect 647926 81849 647978 81855
rect 647830 81833 647882 81839
rect 647830 81775 647882 81781
rect 647734 81611 647786 81617
rect 647734 81553 647786 81559
rect 647924 81058 647980 81067
rect 647924 80993 647980 81002
rect 647938 80803 647966 80993
rect 647926 80797 647978 80803
rect 647926 80739 647978 80745
rect 647062 77763 647114 77769
rect 647062 77705 647114 77711
rect 647926 77541 647978 77547
rect 647924 77506 647926 77515
rect 647978 77506 647980 77515
rect 647924 77441 647980 77450
rect 647158 74951 647210 74957
rect 647158 74893 647210 74899
rect 646964 71882 647020 71891
rect 646964 71817 647020 71826
rect 646868 68626 646924 68635
rect 646868 68561 646924 68570
rect 647170 60347 647198 74893
rect 647924 73658 647980 73667
rect 647924 73593 647980 73602
rect 647938 72145 647966 73593
rect 647926 72139 647978 72145
rect 647926 72081 647978 72087
rect 647924 69662 647980 69671
rect 647924 69597 647926 69606
rect 647978 69597 647980 69606
rect 647926 69565 647978 69571
rect 647924 64186 647980 64195
rect 647924 64121 647980 64130
rect 647938 63487 647966 64121
rect 647926 63481 647978 63487
rect 647926 63423 647978 63429
rect 647924 62262 647980 62271
rect 647924 62197 647980 62206
rect 647938 61045 647966 62197
rect 647926 61039 647978 61045
rect 647926 60981 647978 60987
rect 647156 60338 647212 60347
rect 647156 60273 647212 60282
rect 652258 59121 652286 83361
rect 652354 66225 652382 85285
rect 652450 82695 652478 102051
rect 653686 95967 653738 95973
rect 653686 95909 653738 95915
rect 653698 86987 653726 95909
rect 653684 86978 653740 86987
rect 653684 86913 653740 86922
rect 653684 84314 653740 84323
rect 653684 84249 653740 84258
rect 653698 83615 653726 84249
rect 653686 83609 653738 83615
rect 653686 83551 653738 83557
rect 652436 82686 652492 82695
rect 652436 82621 652492 82630
rect 652342 66219 652394 66225
rect 652342 66161 652394 66167
rect 652246 59115 652298 59121
rect 652246 59057 652298 59063
rect 646772 57082 646828 57091
rect 646772 57017 646828 57026
rect 646484 54714 646540 54723
rect 646484 54649 646540 54658
rect 654082 51943 654110 104493
rect 661174 103959 661226 103965
rect 661174 103901 661226 103907
rect 657526 103885 657578 103891
rect 657526 103827 657578 103833
rect 657538 88000 657566 103827
rect 660694 92415 660746 92421
rect 660694 92357 660746 92363
rect 659830 92267 659882 92273
rect 659830 92209 659882 92215
rect 658870 92193 658922 92199
rect 658870 92135 658922 92141
rect 657538 87972 657792 88000
rect 658882 87986 658910 92135
rect 659348 90826 659404 90835
rect 659348 90761 659404 90770
rect 659362 88000 659390 90761
rect 659842 88000 659870 92209
rect 659362 87972 659616 88000
rect 659842 87972 660144 88000
rect 660706 87986 660734 92357
rect 661186 88000 661214 103901
rect 665602 103743 665630 105265
rect 675106 104650 675134 105561
rect 675106 104622 675408 104650
rect 665590 103737 665642 103743
rect 665590 103679 665642 103685
rect 675764 103258 675820 103267
rect 675764 103193 675820 103202
rect 675778 102786 675806 103193
rect 675764 101482 675820 101491
rect 675764 101417 675820 101426
rect 675778 100936 675806 101417
rect 662518 97965 662570 97971
rect 662518 97907 662570 97913
rect 661750 92341 661802 92347
rect 661750 92283 661802 92289
rect 661762 88000 661790 92283
rect 661186 87972 661440 88000
rect 661762 87972 662016 88000
rect 662530 87986 662558 97907
rect 663094 92711 663146 92717
rect 663094 92653 663146 92659
rect 663106 87986 663134 92653
rect 658006 87309 658058 87315
rect 658058 87257 658320 87260
rect 658006 87251 658320 87257
rect 658018 87232 658320 87251
rect 663286 87087 663338 87093
rect 663286 87029 663338 87035
rect 663298 86395 663326 87029
rect 663284 86386 663340 86395
rect 663284 86321 663340 86330
rect 663284 84758 663340 84767
rect 663202 84716 663284 84744
rect 657046 84201 657098 84207
rect 657046 84143 657098 84149
rect 657058 81691 657086 84143
rect 657046 81685 657098 81691
rect 657046 81627 657098 81633
rect 658582 81685 658634 81691
rect 662420 81650 662476 81659
rect 658634 81633 658896 81636
rect 658582 81627 658896 81633
rect 658594 81608 658896 81627
rect 662420 81585 662422 81594
rect 662474 81585 662476 81594
rect 662422 81553 662474 81559
rect 656962 81016 657216 81044
rect 657538 81016 657792 81044
rect 656962 77547 656990 81016
rect 656950 77541 657002 77547
rect 656950 77483 657002 77489
rect 657538 75697 657566 81016
rect 658306 77769 658334 81030
rect 659602 80748 659630 81030
rect 659554 80720 659630 80748
rect 658294 77763 658346 77769
rect 658294 77705 658346 77711
rect 659554 77695 659582 80720
rect 659542 77689 659594 77695
rect 659542 77631 659594 77637
rect 657526 75691 657578 75697
rect 657526 75633 657578 75639
rect 660130 74957 660158 81030
rect 660118 74951 660170 74957
rect 660118 74893 660170 74899
rect 660706 72145 660734 81030
rect 661186 81016 661440 81044
rect 661762 81016 662016 81044
rect 660694 72139 660746 72145
rect 660694 72081 660746 72087
rect 661186 69629 661214 81016
rect 661762 77621 661790 81016
rect 662530 80803 662558 81030
rect 662518 80797 662570 80803
rect 662518 80739 662570 80745
rect 661750 77615 661802 77621
rect 661750 77557 661802 77563
rect 661174 69623 661226 69629
rect 661174 69565 661226 69571
rect 663202 63487 663230 84716
rect 663284 84693 663340 84702
rect 663476 84018 663532 84027
rect 663476 83953 663532 83962
rect 663380 82834 663436 82843
rect 663380 82769 663436 82778
rect 663284 82094 663340 82103
rect 663284 82029 663340 82038
rect 663298 81913 663326 82029
rect 663286 81907 663338 81913
rect 663286 81849 663338 81855
rect 663394 81839 663422 82769
rect 663382 81833 663434 81839
rect 663382 81775 663434 81781
rect 663190 63481 663242 63487
rect 663190 63423 663242 63429
rect 663490 61045 663518 83953
rect 663478 61039 663530 61045
rect 663478 60981 663530 60987
rect 643606 51937 643658 51943
rect 643606 51879 643658 51885
rect 654070 51937 654122 51943
rect 654070 51879 654122 51885
rect 643618 46763 643646 51879
rect 643606 46757 643658 46763
rect 643606 46699 643658 46705
rect 640726 41799 640778 41805
rect 640726 41741 640778 41747
rect 541460 40506 541516 40515
rect 541460 40441 541516 40450
rect 514006 37433 514058 37439
rect 514006 37375 514058 37381
rect 475510 37359 475562 37365
rect 475510 37301 475562 37307
rect 506806 37359 506858 37365
rect 506806 37301 506858 37307
rect 311060 37250 311116 37259
rect 311060 37185 311116 37194
rect 334100 37250 334156 37259
rect 334100 37185 334156 37194
<< via2 >>
rect 483668 1005153 483670 1005170
rect 483670 1005153 483722 1005170
rect 483722 1005153 483724 1005170
rect 483668 1005114 483724 1005153
rect 535028 1005153 535030 1005170
rect 535030 1005153 535082 1005170
rect 535082 1005153 535084 1005170
rect 535028 1005114 535084 1005153
rect 636884 1005153 636886 1005170
rect 636886 1005153 636938 1005170
rect 636938 1005153 636940 1005170
rect 636884 1005114 636940 1005153
rect 679700 964118 679756 964174
rect 649460 961602 649516 961658
rect 676148 894114 676204 894170
rect 676052 893374 676108 893430
rect 655220 867622 655276 867678
rect 655124 866438 655180 866494
rect 676244 893522 676300 893578
rect 676052 892429 676108 892468
rect 676052 892412 676054 892429
rect 676054 892412 676106 892429
rect 676106 892412 676108 892429
rect 655412 868806 655468 868862
rect 655316 865254 655372 865310
rect 654164 863922 654220 863978
rect 653780 862886 653836 862942
rect 41780 817933 41782 817950
rect 41782 817933 41834 817950
rect 41834 817933 41836 817950
rect 41780 817894 41836 817933
rect 41780 817319 41836 817358
rect 41780 817302 41782 817319
rect 41782 817302 41834 817319
rect 41834 817302 41836 817319
rect 41588 816579 41644 816618
rect 41588 816562 41590 816579
rect 41590 816562 41642 816579
rect 41642 816562 41644 816579
rect 41780 815839 41836 815878
rect 41780 815822 41782 815839
rect 41782 815822 41834 815839
rect 41834 815822 41836 815839
rect 41780 814877 41836 814916
rect 41780 814860 41782 814877
rect 41782 814860 41834 814877
rect 41834 814860 41836 814877
rect 41588 813619 41644 813658
rect 41588 813602 41590 813619
rect 41590 813602 41642 813619
rect 41642 813602 41644 813619
rect 41588 813158 41644 813214
rect 40244 812418 40300 812474
rect 42260 812862 42316 812918
rect 28820 805610 28876 805666
rect 28820 805166 28876 805222
rect 41492 811678 41548 811734
rect 40244 802258 40300 802314
rect 41780 811308 41836 811364
rect 41876 810790 41932 810846
rect 41780 808866 41836 808922
rect 41588 808126 41644 808182
rect 41588 806663 41644 806702
rect 41588 806646 41590 806663
rect 41590 806646 41642 806663
rect 41642 806646 41644 806663
rect 42164 809754 42220 809810
rect 42068 809310 42124 809366
rect 41972 807830 42028 807886
rect 41588 806054 41644 806110
rect 41588 805183 41644 805222
rect 41588 805166 41590 805183
rect 41590 805166 41642 805183
rect 41642 805166 41644 805183
rect 41492 800430 41548 800486
rect 42164 800430 42220 800486
rect 42068 800282 42124 800338
rect 42836 807386 42892 807442
rect 42740 796730 42796 796786
rect 42260 791846 42316 791902
rect 42356 791698 42412 791754
rect 42644 794362 42700 794418
rect 42644 792882 42700 792938
rect 41780 774695 41836 774734
rect 41780 774678 41782 774695
rect 41782 774678 41834 774695
rect 41834 774678 41836 774695
rect 41588 773955 41644 773994
rect 41588 773938 41590 773955
rect 41590 773938 41642 773955
rect 41642 773938 41644 773955
rect 41780 773511 41836 773550
rect 41780 773494 41782 773511
rect 41782 773494 41834 773511
rect 41834 773494 41836 773511
rect 41588 773385 41590 773402
rect 41590 773385 41642 773402
rect 41642 773385 41644 773402
rect 41588 773346 41644 773385
rect 41780 772623 41836 772662
rect 41780 772606 41782 772623
rect 41782 772606 41834 772623
rect 41834 772606 41836 772623
rect 41588 772310 41644 772366
rect 43124 771866 43180 771922
rect 41588 770830 41644 770886
rect 42452 770090 42508 770146
rect 41972 769646 42028 769702
rect 38804 768906 38860 768962
rect 33044 766982 33100 767038
rect 28820 762394 28876 762450
rect 28820 761950 28876 762006
rect 33044 758842 33100 758898
rect 41588 768462 41644 768518
rect 41780 768166 41836 768222
rect 41780 766629 41836 766668
rect 41780 766612 41782 766629
rect 41782 766612 41834 766629
rect 41834 766612 41836 766629
rect 41876 766094 41932 766150
rect 41588 765502 41644 765558
rect 41780 765132 41836 765188
rect 41780 764614 41836 764670
rect 41588 763447 41644 763486
rect 41588 763430 41590 763447
rect 41590 763430 41642 763447
rect 41642 763430 41644 763447
rect 41588 762838 41644 762894
rect 41588 761967 41644 762006
rect 41588 761950 41590 761967
rect 41590 761950 41642 761967
rect 41642 761950 41644 761967
rect 38804 757510 38860 757566
rect 42356 767574 42412 767630
rect 42068 764170 42124 764226
rect 42356 746262 42412 746318
rect 42548 745966 42604 746022
rect 41780 731479 41836 731518
rect 41780 731462 41782 731479
rect 41782 731462 41834 731479
rect 41834 731462 41836 731479
rect 41588 730739 41644 730778
rect 41588 730722 41590 730739
rect 41590 730722 41642 730739
rect 41642 730722 41644 730739
rect 41780 730369 41836 730408
rect 41780 730352 41782 730369
rect 41782 730352 41834 730369
rect 41834 730352 41836 730369
rect 41588 730169 41590 730186
rect 41590 730169 41642 730186
rect 41642 730169 41644 730186
rect 41588 730130 41644 730169
rect 41780 729407 41836 729446
rect 41780 729390 41782 729407
rect 41782 729390 41834 729407
rect 41834 729390 41836 729407
rect 42260 729242 42316 729298
rect 41780 728815 41836 728854
rect 41780 728798 41782 728815
rect 41782 728798 41834 728815
rect 41834 728798 41836 728815
rect 40436 728689 40438 728706
rect 40438 728689 40490 728706
rect 40490 728689 40492 728706
rect 40436 728650 40492 728689
rect 41780 727927 41836 727966
rect 41780 727910 41782 727927
rect 41782 727910 41834 727927
rect 41834 727910 41836 727927
rect 41780 726948 41836 727004
rect 41780 726447 41836 726486
rect 41780 726430 41782 726447
rect 41782 726430 41834 726447
rect 41834 726430 41836 726447
rect 40244 725690 40300 725746
rect 34484 723766 34540 723822
rect 28820 719178 28876 719234
rect 28820 718734 28876 718790
rect 41684 725246 41740 725302
rect 41588 722286 41644 722342
rect 41588 720806 41644 720862
rect 41972 724950 42028 725006
rect 41780 723470 41836 723526
rect 41780 721916 41836 721972
rect 41876 721398 41932 721454
rect 41780 720436 41836 720492
rect 41588 718751 41644 718790
rect 41588 718734 41590 718751
rect 41590 718734 41642 718751
rect 41642 718734 41644 718751
rect 40244 717308 40300 717364
rect 34484 715774 34540 715830
rect 42260 724358 42316 724414
rect 42452 722878 42508 722934
rect 42452 711630 42508 711686
rect 42356 711038 42412 711094
rect 42836 711332 42892 711388
rect 42356 702898 42412 702954
rect 42548 702750 42604 702806
rect 42932 711186 42988 711242
rect 41780 688263 41836 688302
rect 41780 688246 41782 688263
rect 41782 688246 41834 688263
rect 41834 688246 41836 688263
rect 41588 687523 41644 687562
rect 41588 687506 41590 687523
rect 41590 687506 41642 687523
rect 41642 687506 41644 687523
rect 41780 687227 41836 687266
rect 41780 687210 41782 687227
rect 41782 687210 41834 687227
rect 41834 687210 41836 687227
rect 41588 686953 41590 686970
rect 41590 686953 41642 686970
rect 41642 686953 41644 686970
rect 41588 686914 41644 686953
rect 41588 686043 41644 686082
rect 41588 686026 41590 686043
rect 41590 686026 41642 686043
rect 41642 686026 41644 686043
rect 41780 685325 41782 685342
rect 41782 685325 41834 685342
rect 41834 685325 41836 685342
rect 41780 685286 41836 685325
rect 41780 684141 41782 684158
rect 41782 684141 41834 684158
rect 41834 684141 41836 684158
rect 41780 684102 41836 684141
rect 42068 683806 42124 683862
rect 39860 682474 39916 682530
rect 34484 680550 34540 680606
rect 28820 675962 28876 676018
rect 28820 675518 28876 675574
rect 34484 672860 34540 672916
rect 41780 681734 41836 681790
rect 41780 680254 41836 680310
rect 41780 679701 41782 679718
rect 41782 679701 41834 679718
rect 41834 679701 41836 679718
rect 41780 679662 41836 679701
rect 41588 679070 41644 679126
rect 41780 678774 41836 678830
rect 41972 678182 42028 678238
rect 41780 677738 41836 677794
rect 41780 677220 41836 677276
rect 41780 676702 41836 676758
rect 41780 675757 41836 675796
rect 41780 675740 41782 675757
rect 41782 675740 41834 675757
rect 41834 675740 41836 675757
rect 39860 671078 39916 671134
rect 41972 670634 42028 670690
rect 42548 683214 42604 683270
rect 42164 682178 42220 682234
rect 42356 681142 42412 681198
rect 42452 671226 42508 671282
rect 42548 668414 42604 668470
rect 42452 667674 42508 667730
rect 42548 660866 42604 660922
rect 42356 659386 42412 659442
rect 41588 644899 41644 644938
rect 41588 644882 41590 644899
rect 41590 644882 41642 644899
rect 41642 644882 41644 644899
rect 41492 644734 41548 644790
rect 41588 644307 41644 644346
rect 41588 644290 41590 644307
rect 41590 644290 41642 644307
rect 41642 644290 41644 644307
rect 41780 644011 41836 644050
rect 41780 643994 41782 644011
rect 41782 643994 41834 644011
rect 41834 643994 41836 644011
rect 41588 643737 41590 643754
rect 41590 643737 41642 643754
rect 41642 643737 41644 643754
rect 41588 643698 41644 643737
rect 41588 642827 41644 642866
rect 41588 642810 41590 642827
rect 41590 642810 41642 642827
rect 41642 642810 41644 642827
rect 41588 641347 41644 641386
rect 41588 641330 41590 641347
rect 41590 641330 41642 641347
rect 41642 641330 41644 641347
rect 41492 641182 41548 641238
rect 41780 640607 41836 640646
rect 41780 640590 41782 640607
rect 41782 640590 41834 640607
rect 41834 640590 41836 640607
rect 42164 639998 42220 640054
rect 39860 639258 39916 639314
rect 34484 637334 34540 637390
rect 28820 632746 28876 632802
rect 28820 632302 28876 632358
rect 42068 639110 42124 639166
rect 41780 638518 41836 638574
rect 41876 637926 41932 637982
rect 41588 636298 41644 636354
rect 41780 636093 41836 636132
rect 41780 636076 41782 636093
rect 41782 636076 41834 636093
rect 41834 636076 41836 636093
rect 41588 635262 41644 635318
rect 41684 634818 41740 634874
rect 41588 634374 41644 634430
rect 41780 633486 41836 633542
rect 41780 632541 41836 632580
rect 41780 632524 41782 632541
rect 41782 632524 41834 632541
rect 41834 632524 41836 632541
rect 42164 637038 42220 637094
rect 42356 634078 42412 634134
rect 39860 628010 39916 628066
rect 34484 627862 34540 627918
rect 42836 616466 42892 616522
rect 42740 616318 42796 616374
rect 41684 602110 41740 602166
rect 41588 601683 41644 601722
rect 41588 601666 41590 601683
rect 41590 601666 41642 601683
rect 41642 601666 41644 601683
rect 41780 601387 41836 601426
rect 41780 601370 41782 601387
rect 41782 601370 41834 601387
rect 41834 601370 41836 601387
rect 41780 600795 41836 600834
rect 41780 600778 41782 600795
rect 41782 600778 41834 600795
rect 41834 600778 41836 600795
rect 41780 600373 41782 600390
rect 41782 600373 41834 600390
rect 41834 600373 41836 600390
rect 41780 600334 41836 600373
rect 41780 599833 41836 599872
rect 41780 599816 41782 599833
rect 41782 599816 41834 599833
rect 41834 599816 41836 599833
rect 41780 599315 41836 599354
rect 41780 599298 41782 599315
rect 41782 599298 41834 599315
rect 41834 599298 41836 599315
rect 39860 598706 39916 598762
rect 41780 598353 41836 598392
rect 41780 598336 41782 598353
rect 41782 598336 41834 598353
rect 41834 598336 41836 598353
rect 41780 597857 41782 597874
rect 41782 597857 41834 597874
rect 41834 597857 41836 597874
rect 41780 597818 41836 597857
rect 41876 597374 41932 597430
rect 41588 596651 41644 596690
rect 41588 596634 41590 596651
rect 41590 596634 41642 596651
rect 41642 596634 41644 596651
rect 34388 596042 34444 596098
rect 28820 589530 28876 589586
rect 28820 589086 28876 589142
rect 41780 595894 41836 595950
rect 41588 595154 41644 595210
rect 41780 594784 41836 594840
rect 34484 594118 34540 594174
rect 41588 593691 41644 593730
rect 41588 593674 41590 593691
rect 41590 593674 41642 593691
rect 41642 593674 41644 593691
rect 41684 592211 41740 592250
rect 41684 592194 41686 592211
rect 41686 592194 41738 592211
rect 41738 592194 41740 592211
rect 41588 591158 41644 591214
rect 41588 589086 41644 589142
rect 34484 586216 34540 586272
rect 34388 585920 34444 585976
rect 42068 593304 42124 593360
rect 41972 590879 42028 590918
rect 41972 590862 41974 590879
rect 41974 590862 42026 590879
rect 42026 590862 42028 590879
rect 42260 592934 42316 592990
rect 42356 591750 42412 591806
rect 42932 587458 42988 587514
rect 42836 577246 42892 577302
rect 42260 573990 42316 574046
rect 42548 573842 42604 573898
rect 41780 539802 41836 539858
rect 41780 538026 41836 538082
rect 41780 536250 41836 536306
rect 41780 535066 41836 535122
rect 41780 534178 41836 534234
rect 41780 533882 41836 533938
rect 41876 532994 41932 533050
rect 41780 530774 41836 530830
rect 41780 530034 41836 530090
rect 42164 529294 42220 529350
rect 42164 527222 42220 527278
rect 42260 527074 42316 527130
rect 41488 476049 41548 476109
rect 41511 475531 41571 475591
rect 41098 474949 41158 475009
rect 41469 474569 41529 474629
rect 40340 473794 40396 473850
rect 39764 473202 39820 473258
rect 39668 472314 39724 472370
rect 34484 464322 34540 464378
rect 23060 463730 23116 463786
rect 23060 463286 23116 463342
rect 42260 472166 42316 472222
rect 42260 469946 42316 470002
rect 43212 478086 43268 478142
rect 43124 472166 43180 472222
rect 42452 470538 42508 470594
rect 42356 468614 42412 468670
rect 41780 463599 41836 463638
rect 41780 463582 41782 463599
rect 41782 463582 41834 463599
rect 41834 463582 41836 463599
rect 41588 428495 41644 428534
rect 41588 428478 41590 428495
rect 41590 428478 41642 428495
rect 41642 428478 41644 428495
rect 41780 428125 41836 428164
rect 41780 428108 41782 428125
rect 41782 428108 41834 428125
rect 41834 428108 41836 428125
rect 40340 426850 40396 426906
rect 34292 425814 34348 425870
rect 25844 424926 25900 424982
rect 41780 427607 41836 427646
rect 41780 427590 41782 427607
rect 41782 427590 41834 427607
rect 41834 427590 41836 427607
rect 41780 426571 41836 426610
rect 41780 426554 41782 426571
rect 41782 426554 41834 426571
rect 41834 426554 41836 426571
rect 41588 425370 41644 425426
rect 34484 424778 34540 424834
rect 34388 423446 34444 423502
rect 34292 420782 34348 420838
rect 34484 423298 34540 423354
rect 42260 421522 42316 421578
rect 39956 420338 40012 420394
rect 39860 419894 39916 419950
rect 40148 419450 40204 419506
rect 41588 418858 41644 418914
rect 41780 418562 41836 418618
rect 41588 417970 41644 418026
rect 41780 417082 41836 417138
rect 23060 416342 23116 416398
rect 41780 416137 41836 416176
rect 41780 416120 41782 416137
rect 41782 416120 41834 416137
rect 41834 416120 41836 416137
rect 23060 415898 23116 415954
rect 42548 417674 42604 417730
rect 42068 406010 42124 406066
rect 41780 402014 41836 402070
rect 41780 400090 41836 400146
rect 41780 399498 41836 399554
rect 41780 398758 41836 398814
rect 41780 388084 41836 388140
rect 41780 386030 41836 386086
rect 41588 385921 41590 385938
rect 41590 385921 41642 385938
rect 41642 385921 41644 385938
rect 41588 385882 41644 385921
rect 41588 385307 41644 385346
rect 41588 385290 41590 385307
rect 41590 385290 41642 385307
rect 41642 385290 41644 385307
rect 41588 384737 41590 384754
rect 41590 384737 41642 384754
rect 41642 384737 41644 384754
rect 41588 384698 41644 384737
rect 41588 383827 41644 383866
rect 41588 383810 41590 383827
rect 41590 383810 41642 383827
rect 41642 383810 41644 383827
rect 34484 383218 34540 383274
rect 41876 385011 41932 385050
rect 41876 384994 41878 385011
rect 41878 384994 41930 385011
rect 41930 384994 41932 385011
rect 41876 383218 41932 383274
rect 41780 383070 41836 383126
rect 41588 382347 41644 382386
rect 41588 382330 41590 382347
rect 41590 382330 41642 382347
rect 41642 382330 41644 382347
rect 41876 381960 41932 382016
rect 39956 380850 40012 380906
rect 37364 379222 37420 379278
rect 34484 378778 34540 378834
rect 28820 373746 28876 373802
rect 28820 373302 28876 373358
rect 41780 379535 41836 379574
rect 41780 379518 41782 379535
rect 41782 379518 41834 379535
rect 41834 379518 41836 379535
rect 41588 377315 41644 377354
rect 41588 377298 41590 377315
rect 41590 377298 41642 377315
rect 41642 377298 41644 377315
rect 42452 377002 42508 377058
rect 41492 376262 41548 376318
rect 41780 375966 41836 376022
rect 41684 375374 41740 375430
rect 41588 374782 41644 374838
rect 41588 373319 41644 373358
rect 41588 373302 41590 373319
rect 41590 373302 41642 373319
rect 41642 373302 41644 373319
rect 41780 359242 41836 359298
rect 41780 358798 41836 358854
rect 41780 356874 41836 356930
rect 41780 356430 41836 356486
rect 41780 355542 41836 355598
rect 41684 343110 41740 343166
rect 41588 340611 41644 340650
rect 41588 340594 41590 340611
rect 41590 340594 41642 340611
rect 41642 340594 41644 340611
rect 41780 342831 41836 342870
rect 41780 342814 41782 342831
rect 41782 342814 41834 342831
rect 41834 342814 41836 342831
rect 41780 342313 41836 342352
rect 41780 342296 41782 342313
rect 41782 342296 41834 342313
rect 41834 342296 41836 342313
rect 41780 341795 41836 341834
rect 41780 341778 41782 341795
rect 41782 341778 41834 341795
rect 41834 341778 41836 341795
rect 41780 341373 41782 341390
rect 41782 341373 41834 341390
rect 41834 341373 41836 341390
rect 41780 341334 41836 341373
rect 41780 340315 41836 340354
rect 41780 340298 41782 340315
rect 41782 340298 41834 340315
rect 41834 340298 41836 340315
rect 41684 340002 41740 340058
rect 41588 339131 41644 339170
rect 41588 339114 41590 339131
rect 41590 339114 41642 339131
rect 41642 339114 41644 339131
rect 43124 338818 43180 338874
rect 39764 337634 39820 337690
rect 41588 336154 41644 336210
rect 41780 335710 41836 335766
rect 41492 333046 41548 333102
rect 41396 332602 41452 332658
rect 41684 332158 41740 332214
rect 41588 331566 41644 331622
rect 28820 330530 28876 330586
rect 28820 330086 28876 330142
rect 41876 334230 41932 334286
rect 42452 333786 42508 333842
rect 41876 330399 41932 330438
rect 41876 330382 41878 330399
rect 41878 330382 41930 330399
rect 41930 330382 41932 330399
rect 41780 316174 41836 316230
rect 41780 315434 41836 315490
rect 41780 313658 41836 313714
rect 41780 313214 41836 313270
rect 41780 312326 41836 312382
rect 39668 298710 39724 298766
rect 41780 299615 41836 299654
rect 41780 299598 41782 299615
rect 41782 299598 41834 299615
rect 41834 299598 41836 299615
rect 41780 299171 41836 299210
rect 41780 299154 41782 299171
rect 41782 299154 41834 299171
rect 41834 299154 41836 299171
rect 41780 298157 41782 298174
rect 41782 298157 41834 298174
rect 41834 298157 41836 298174
rect 41780 298118 41836 298157
rect 41780 297617 41836 297656
rect 41780 297600 41782 297617
rect 41782 297600 41834 297617
rect 41834 297600 41836 297617
rect 41780 297099 41836 297138
rect 41780 297082 41782 297099
rect 41782 297082 41834 297099
rect 41834 297082 41836 297099
rect 39764 296490 39820 296546
rect 39956 295898 40012 295954
rect 41588 295915 41644 295954
rect 41588 295898 41590 295915
rect 41590 295898 41642 295915
rect 41642 295898 41644 295915
rect 40244 294418 40300 294474
rect 41588 292938 41644 292994
rect 41780 292568 41836 292624
rect 41588 290905 41590 290922
rect 41590 290905 41642 290922
rect 41642 290905 41644 290922
rect 41588 290866 41644 290905
rect 41492 289386 41548 289442
rect 41588 288942 41644 288998
rect 28820 287314 28876 287370
rect 28820 286870 28876 286926
rect 42356 290718 42412 290774
rect 42260 288646 42316 288702
rect 41876 287183 41932 287222
rect 41876 287166 41878 287183
rect 41878 287166 41930 287183
rect 41930 287166 41932 287183
rect 42548 290126 42604 290182
rect 41780 272958 41836 273014
rect 41780 272366 41836 272422
rect 41780 270590 41836 270646
rect 41780 269998 41836 270054
rect 41780 269110 41836 269166
rect 23156 254162 23212 254218
rect 23060 253274 23116 253330
rect 43316 261886 43372 261942
rect 40244 256234 40300 256290
rect 41588 255642 41644 255698
rect 41780 255385 41782 255402
rect 41782 255385 41834 255402
rect 41834 255385 41836 255402
rect 41780 255346 41836 255385
rect 41780 254941 41782 254958
rect 41782 254941 41834 254958
rect 41834 254941 41836 254958
rect 41780 254902 41836 254941
rect 41780 254475 41836 254514
rect 41780 254458 41782 254475
rect 41782 254458 41834 254475
rect 41834 254458 41836 254475
rect 23348 253274 23404 253330
rect 23252 252682 23308 252738
rect 40244 251202 40300 251258
rect 34484 249722 34540 249778
rect 41780 249426 41836 249482
rect 41492 246614 41548 246670
rect 41684 245726 41740 245782
rect 41588 245151 41644 245190
rect 41588 245134 41590 245151
rect 41590 245134 41642 245151
rect 41642 245134 41644 245151
rect 41588 244690 41644 244746
rect 41588 243654 41644 243710
rect 41876 247889 41932 247928
rect 41876 247872 41878 247889
rect 41878 247872 41930 247889
rect 41930 247872 41932 247889
rect 42260 247502 42316 247558
rect 41876 246318 41932 246374
rect 42548 245430 42604 245486
rect 41780 229742 41836 229798
rect 41780 229150 41836 229206
rect 41780 227374 41836 227430
rect 41780 226782 41836 226838
rect 41780 225894 41836 225950
rect 41780 213279 41782 213296
rect 41782 213279 41834 213296
rect 41834 213279 41836 213296
rect 41780 213240 41836 213279
rect 41588 212909 41590 212926
rect 41590 212909 41642 212926
rect 41642 212909 41644 212926
rect 41588 212870 41644 212909
rect 41780 212169 41782 212186
rect 41782 212169 41834 212186
rect 41834 212169 41836 212186
rect 41780 212130 41836 212169
rect 41780 211725 41782 211742
rect 41782 211725 41834 211742
rect 41834 211725 41836 211742
rect 41780 211686 41836 211725
rect 41588 211429 41590 211446
rect 41590 211429 41642 211446
rect 41642 211429 41644 211446
rect 41588 211390 41644 211429
rect 41780 210689 41782 210706
rect 41782 210689 41834 210706
rect 41834 210689 41836 210706
rect 41780 210650 41836 210689
rect 41780 210223 41836 210262
rect 43508 266890 43564 266946
rect 41780 210206 41782 210223
rect 41782 210206 41834 210223
rect 41834 210206 41836 210223
rect 41588 209949 41590 209966
rect 41590 209949 41642 209966
rect 41642 209949 41644 209966
rect 41588 209910 41644 209949
rect 57716 790810 57772 790866
rect 57620 789626 57676 789682
rect 58196 788442 58252 788498
rect 58388 787258 58444 787314
rect 59636 785482 59692 785538
rect 59156 784890 59212 784946
rect 44756 275326 44812 275382
rect 44660 267038 44716 267094
rect 58676 747594 58732 747650
rect 54740 745983 54796 746022
rect 54740 745966 54742 745983
rect 54742 745966 54794 745983
rect 54794 745966 54796 745983
rect 54644 745818 54700 745874
rect 57620 745226 57676 745282
rect 58580 745374 58636 745430
rect 58100 744042 58156 744098
rect 59636 742858 59692 742914
rect 59732 741674 59788 741730
rect 45140 276214 45196 276270
rect 44948 261642 45004 261698
rect 41588 209357 41590 209374
rect 41590 209357 41642 209374
rect 41642 209357 41644 209374
rect 41588 209318 41644 209357
rect 41780 208208 41836 208264
rect 34100 206506 34156 206562
rect 42260 206210 42316 206266
rect 34196 204434 34252 204490
rect 34292 203990 34348 204046
rect 41588 203546 41644 203602
rect 34484 202954 34540 203010
rect 34388 201918 34444 201974
rect 41876 202806 41932 202862
rect 41972 201661 41974 201678
rect 41974 201661 42026 201678
rect 42026 201661 42028 201678
rect 41972 201622 42028 201661
rect 41588 201513 41590 201530
rect 41590 201513 41642 201530
rect 41642 201513 41644 201530
rect 41588 201474 41644 201513
rect 41588 200921 41590 200938
rect 41590 200921 41642 200938
rect 41642 200921 41644 200938
rect 41588 200882 41644 200921
rect 59636 704378 59692 704434
rect 58772 702641 58774 702658
rect 58774 702641 58826 702658
rect 58826 702641 58828 702658
rect 58772 702602 58828 702641
rect 58868 702010 58924 702066
rect 58676 700826 58732 700882
rect 59252 699642 59308 699698
rect 58868 698458 58924 698514
rect 59636 661162 59692 661218
rect 58772 659403 58828 659442
rect 58772 659386 58774 659403
rect 58774 659386 58826 659403
rect 58826 659386 58828 659403
rect 57716 658794 57772 658850
rect 59156 657610 59212 657666
rect 58196 656426 58252 656482
rect 58388 655242 58444 655298
rect 58964 617946 59020 618002
rect 58196 615578 58252 615634
rect 59636 616209 59638 616226
rect 59638 616209 59690 616226
rect 59690 616209 59692 616226
rect 59636 616170 59692 616209
rect 58964 614394 59020 614450
rect 59636 613210 59692 613266
rect 59540 612026 59596 612082
rect 41780 186674 41836 186730
rect 41780 185786 41836 185842
rect 41780 184158 41836 184214
rect 41780 183566 41836 183622
rect 41780 182826 41836 182882
rect 50612 275178 50668 275234
rect 50420 275030 50476 275086
rect 58964 574730 59020 574786
rect 58196 572362 58252 572418
rect 59636 572993 59638 573010
rect 59638 572993 59690 573010
rect 59690 572993 59692 573010
rect 59636 572954 59692 572993
rect 58964 571178 59020 571234
rect 59348 569994 59404 570050
rect 59540 568810 59596 568866
rect 57716 531662 57772 531718
rect 57620 530478 57676 530534
rect 58196 529294 58252 529350
rect 58964 527074 59020 527130
rect 58580 525890 58636 525946
rect 59348 524706 59404 524762
rect 58484 404086 58540 404142
rect 58772 402902 58828 402958
rect 57620 400534 57676 400590
rect 58772 399942 58828 399998
rect 58196 399350 58252 399406
rect 59732 398166 59788 398222
rect 58484 360870 58540 360926
rect 59156 359686 59212 359742
rect 57620 357466 57676 357522
rect 58196 356134 58252 356190
rect 59636 356726 59692 356782
rect 58580 354950 58636 355006
rect 58484 317654 58540 317710
rect 59156 316470 59212 316526
rect 59156 314102 59212 314158
rect 58868 312918 58924 312974
rect 59636 313845 59638 313862
rect 59638 313845 59690 313862
rect 59690 313845 59692 313862
rect 59636 313806 59692 313845
rect 59636 311734 59692 311790
rect 59348 295158 59404 295214
rect 59252 293974 59308 294030
rect 58196 292642 58252 292698
rect 58868 289238 58924 289294
rect 59156 288071 59212 288110
rect 59156 288054 59158 288071
rect 59158 288054 59210 288071
rect 59210 288054 59212 288071
rect 59060 285686 59116 285742
rect 57620 284502 57676 284558
rect 58868 283318 58924 283374
rect 58964 282282 59020 282338
rect 59252 286870 59308 286926
rect 59252 280950 59308 281006
rect 59444 292790 59500 292846
rect 59636 291458 59692 291514
rect 59540 279766 59596 279822
rect 61652 277842 61708 277898
rect 61940 278286 61996 278342
rect 62132 602110 62188 602166
rect 62132 278434 62188 278490
rect 62036 266742 62092 266798
rect 61844 266594 61900 266650
rect 62324 536990 62380 537046
rect 62324 270590 62380 270646
rect 62516 277990 62572 278046
rect 62708 386030 62764 386086
rect 62900 383218 62956 383274
rect 63092 343110 63148 343166
rect 63092 278138 63148 278194
rect 62900 277694 62956 277750
rect 62708 277546 62764 277602
rect 63284 277398 63340 277454
rect 62612 273402 62668 273458
rect 65876 269258 65932 269314
rect 70580 272070 70636 272126
rect 69428 269554 69484 269610
rect 72980 272218 73036 272274
rect 71732 269406 71788 269462
rect 78836 272366 78892 272422
rect 77588 269702 77644 269758
rect 62420 266446 62476 266502
rect 62228 266298 62284 266354
rect 88340 272514 88396 272570
rect 91892 272662 91948 272718
rect 139124 269850 139180 269906
rect 148532 244542 148588 244598
rect 148340 242026 148396 242082
rect 148244 239658 148300 239714
rect 147860 232258 147916 232314
rect 146900 229890 146956 229946
rect 147188 226355 147244 226394
rect 147188 226338 147190 226355
rect 147190 226338 147242 226355
rect 147242 226338 147244 226355
rect 146900 221471 146956 221510
rect 146900 221454 146902 221471
rect 146902 221454 146954 221471
rect 146954 221454 146956 221471
rect 147668 218938 147724 218994
rect 147092 214071 147148 214110
rect 147092 214054 147094 214071
rect 147094 214054 147146 214071
rect 147146 214054 147148 214071
rect 146900 212887 146956 212926
rect 146900 212870 146902 212887
rect 146902 212870 146954 212887
rect 146954 212870 146956 212887
rect 147380 211686 147436 211742
rect 147476 210371 147532 210410
rect 147476 210354 147478 210371
rect 147478 210354 147530 210371
rect 147530 210354 147532 210371
rect 146900 209170 146956 209226
rect 147188 207986 147244 208042
rect 147284 206358 147340 206414
rect 147476 199550 147532 199606
rect 147380 190966 147436 191022
rect 147764 176462 147820 176518
rect 148436 234774 148492 234830
rect 148724 243358 148780 243414
rect 148628 238474 148684 238530
rect 149012 240842 149068 240898
rect 148916 236698 148972 236754
rect 148820 233590 148876 233646
rect 148916 173946 148972 174002
rect 149108 235958 149164 236014
rect 148916 168026 148972 168082
rect 148532 166250 148588 166306
rect 148340 165510 148396 165566
rect 148244 161810 148300 161866
rect 147092 159442 147148 159498
rect 146900 156926 146956 156982
rect 147668 146122 147724 146178
rect 147668 144494 147724 144550
rect 147284 143606 147340 143662
rect 147476 142422 147532 142478
rect 147476 139906 147532 139962
rect 147668 138722 147724 138778
rect 147476 130286 147532 130342
rect 147668 127918 147724 127974
rect 148436 163142 148492 163198
rect 148724 164326 148780 164382
rect 148628 160626 148684 160682
rect 148820 157666 148876 157722
rect 149396 231074 149452 231130
rect 149396 228114 149452 228170
rect 149396 227374 149452 227430
rect 149396 225154 149452 225210
rect 149492 223822 149548 223878
rect 149396 222638 149452 222694
rect 149396 219678 149452 219734
rect 149396 217754 149452 217810
rect 149492 216570 149548 216626
rect 149396 214794 149452 214850
rect 149396 205618 149452 205674
rect 149300 204434 149356 204490
rect 149492 203250 149548 203306
rect 149396 201918 149452 201974
rect 149396 200734 149452 200790
rect 149492 198366 149548 198422
rect 149396 197034 149452 197090
rect 149396 195867 149452 195906
rect 149396 195850 149398 195867
rect 149398 195850 149450 195867
rect 149450 195850 149452 195867
rect 149492 194666 149548 194722
rect 149396 193334 149452 193390
rect 149396 192150 149452 192206
rect 149396 189782 149452 189838
rect 149300 187414 149356 187470
rect 149204 186230 149260 186286
rect 149492 188006 149548 188062
rect 149396 183714 149452 183770
rect 149588 184454 149644 184510
rect 149492 182530 149548 182586
rect 149300 181346 149356 181402
rect 149492 179570 149548 179626
rect 149396 178830 149452 178886
rect 149396 177646 149452 177702
rect 149396 175130 149452 175186
rect 149300 172762 149356 172818
rect 149204 170246 149260 170302
rect 148916 133838 148972 133894
rect 148820 132654 148876 132710
rect 147476 120518 147532 120574
rect 148436 111934 148492 111990
rect 147188 108399 147244 108438
rect 147188 108382 147190 108399
rect 147190 108382 147242 108399
rect 147242 108382 147244 108399
rect 148340 107198 148396 107254
rect 148244 104682 148300 104738
rect 148628 109583 148684 109622
rect 148628 109566 148630 109583
rect 148630 109566 148682 109583
rect 148682 109566 148684 109583
rect 148628 106014 148684 106070
rect 148532 102314 148588 102370
rect 149588 170986 149644 171042
rect 149492 169062 149548 169118
rect 149300 154558 149356 154614
rect 149300 149822 149356 149878
rect 149300 148490 149356 148546
rect 149108 129102 149164 129158
rect 148916 121702 148972 121758
rect 148724 103498 148780 103554
rect 148628 86495 148684 86534
rect 148628 86478 148630 86495
rect 148630 86478 148682 86495
rect 148682 86478 148684 86495
rect 149492 153078 149548 153134
rect 149492 150858 149548 150914
rect 149492 147306 149548 147362
rect 149684 155742 149740 155798
rect 149684 152042 149740 152098
rect 149684 141255 149740 141294
rect 149684 141238 149686 141255
rect 149686 141238 149738 141255
rect 149738 141238 149740 141255
rect 149588 137538 149644 137594
rect 149684 135910 149740 135966
rect 149684 135022 149740 135078
rect 149684 130878 149740 130934
rect 149300 126586 149356 126642
rect 149204 122442 149260 122498
rect 149108 115190 149164 115246
rect 149588 125402 149644 125458
rect 149396 124218 149452 124274
rect 149492 119334 149548 119390
rect 149396 118189 149398 118206
rect 149398 118189 149450 118206
rect 149450 118189 149452 118206
rect 149396 118150 149452 118189
rect 149492 116818 149548 116874
rect 149396 115634 149452 115690
rect 149396 115190 149452 115246
rect 149492 114450 149548 114506
rect 149396 113118 149452 113174
rect 149396 110898 149452 110954
rect 149396 100851 149452 100890
rect 149396 100834 149398 100851
rect 149398 100834 149450 100851
rect 149450 100834 149452 100851
rect 149492 99798 149548 99854
rect 149396 98614 149452 98670
rect 149492 97430 149548 97486
rect 149396 95654 149452 95710
rect 149300 94914 149356 94970
rect 148436 85294 148492 85350
rect 146996 84110 147052 84166
rect 148340 81594 148396 81650
rect 149204 82334 149260 82390
rect 148820 77894 148876 77950
rect 149492 93730 149548 93786
rect 149396 92546 149452 92602
rect 149684 91362 149740 91418
rect 149396 90178 149452 90234
rect 149396 88994 149452 89050
rect 149300 80410 149356 80466
rect 149108 71974 149164 72030
rect 149492 87218 149548 87274
rect 149588 79226 149644 79282
rect 149396 76710 149452 76766
rect 149492 75526 149548 75582
rect 149300 73750 149356 73806
rect 184340 219530 184396 219586
rect 184340 218829 184342 218846
rect 184342 218829 184394 218846
rect 184394 218829 184396 218846
rect 184340 218790 184396 218829
rect 194420 272218 194476 272274
rect 193748 272070 193804 272126
rect 192404 269258 192460 269314
rect 193076 269554 193132 269610
rect 194228 269406 194284 269462
rect 196628 272366 196684 272422
rect 196148 269702 196204 269758
rect 199220 272514 199276 272570
rect 200180 272662 200236 272718
rect 209588 268074 209644 268130
rect 213332 269850 213388 269906
rect 214292 268074 214348 268130
rect 284276 270294 284332 270350
rect 284660 270311 284716 270350
rect 284660 270294 284662 270311
rect 284662 270294 284714 270311
rect 284714 270294 284716 270311
rect 341684 274438 341740 274494
rect 347636 274586 347692 274642
rect 350228 274734 350284 274790
rect 353396 274882 353452 274938
rect 370100 271774 370156 271830
rect 369620 271626 369676 271682
rect 368372 269110 368428 269166
rect 367892 268962 367948 269018
rect 374324 270442 374380 270498
rect 375572 271922 375628 271978
rect 377012 270294 377068 270350
rect 379028 276066 379084 276122
rect 378644 273254 378700 273310
rect 383444 275918 383500 275974
rect 382964 273106 383020 273162
rect 385556 268814 385612 268870
rect 388436 270146 388492 270202
rect 390356 275770 390412 275826
rect 390164 272958 390220 273014
rect 391508 269998 391564 270054
rect 392756 272810 392812 272866
rect 395156 276510 395212 276566
rect 397076 269850 397132 269906
rect 398900 275622 398956 275678
rect 398708 272662 398764 272718
rect 402548 276658 402604 276714
rect 403028 269702 403084 269758
rect 404180 272514 404236 272570
rect 405428 276806 405484 276862
rect 405620 269554 405676 269610
rect 407828 275474 407884 275530
rect 407252 272366 407308 272422
rect 410900 272218 410956 272274
rect 410420 269406 410476 269462
rect 411764 272070 411820 272126
rect 411572 269258 411628 269314
rect 474836 274438 474892 274494
rect 489044 274586 489100 274642
rect 496052 274734 496108 274790
rect 503156 274882 503212 274938
rect 521300 276806 521356 276862
rect 523028 268814 523084 268870
rect 529844 276658 529900 276714
rect 540980 269110 541036 269166
rect 539828 268962 539884 269018
rect 544532 271774 544588 271830
rect 543380 271626 543436 271682
rect 558740 271922 558796 271978
rect 555188 270442 555244 270498
rect 566996 276066 567052 276122
rect 565844 273254 565900 273310
rect 562292 270294 562348 270350
rect 577652 275918 577708 275974
rect 576500 273106 576556 273162
rect 595412 275770 595468 275826
rect 594164 272958 594220 273014
rect 590612 270146 590668 270202
rect 601268 272810 601324 272866
rect 597716 269998 597772 270054
rect 607220 276510 607276 276566
rect 611924 269850 611980 269906
rect 616628 275622 616684 275678
rect 615476 272662 615532 272718
rect 626132 269702 626188 269758
rect 629684 272514 629740 272570
rect 633236 269554 633292 269610
rect 637940 275474 637996 275530
rect 636788 272366 636844 272422
rect 646484 275326 646540 275382
rect 646196 272218 646252 272274
rect 645044 269406 645100 269462
rect 420404 262171 420460 262210
rect 420404 262154 420406 262171
rect 420406 262154 420458 262171
rect 420458 262154 420460 262171
rect 185588 220270 185644 220326
rect 185492 198218 185548 198274
rect 184244 197626 184300 197682
rect 184340 195258 184396 195314
rect 184436 194370 184492 194426
rect 184532 193778 184588 193834
rect 184436 192890 184492 192946
rect 184340 192298 184396 192354
rect 184532 191410 184588 191466
rect 184628 190670 184684 190726
rect 184340 189969 184342 189986
rect 184342 189969 184394 189986
rect 184394 189969 184396 189986
rect 184340 189930 184396 189969
rect 184340 188450 184396 188506
rect 184532 189190 184588 189246
rect 184436 187562 184492 187618
rect 184340 186822 184396 186878
rect 184436 186082 184492 186138
rect 184628 185342 184684 185398
rect 184532 184602 184588 184658
rect 184340 183862 184396 183918
rect 184436 181494 184492 181550
rect 184340 180754 184396 180810
rect 184436 180014 184492 180070
rect 184628 179274 184684 179330
rect 184532 178534 184588 178590
rect 184436 177646 184492 177702
rect 184340 177054 184396 177110
rect 184532 176166 184588 176222
rect 184340 175591 184396 175630
rect 184340 175574 184342 175591
rect 184342 175574 184394 175591
rect 184394 175574 184396 175591
rect 184436 173946 184492 174002
rect 184340 172466 184396 172522
rect 184436 171726 184492 171782
rect 184628 170838 184684 170894
rect 184532 170246 184588 170302
rect 184436 169358 184492 169414
rect 184340 168618 184396 168674
rect 184628 167878 184684 167934
rect 184532 167138 184588 167194
rect 184340 166398 184396 166454
rect 184436 165658 184492 165714
rect 186068 211982 186124 212038
rect 185972 204286 186028 204342
rect 186260 214942 186316 214998
rect 186452 213462 186508 213518
rect 186356 207246 186412 207302
rect 186644 210502 186700 210558
rect 186932 221010 186988 221066
rect 186836 218050 186892 218106
rect 187124 243358 187180 243414
rect 187028 216422 187084 216478
rect 186740 209022 186796 209078
rect 186548 205914 186604 205970
rect 186164 202806 186220 202862
rect 185972 199698 186028 199754
rect 420404 259786 420460 259842
rect 191540 259342 191596 259398
rect 190196 251646 190252 251702
rect 420404 256974 420460 257030
rect 420404 255198 420460 255254
rect 420404 252830 420460 252886
rect 420308 250462 420364 250518
rect 420404 248094 420460 248150
rect 420404 245282 420460 245338
rect 420404 243506 420460 243562
rect 420404 241138 420460 241194
rect 412148 240102 412204 240158
rect 412052 239971 412108 240010
rect 412052 239954 412054 239971
rect 412054 239954 412106 239971
rect 412106 239954 412108 239971
rect 292148 229002 292204 229058
rect 293108 228854 293164 228910
rect 296564 229150 296620 229206
rect 299444 234922 299500 234978
rect 299348 234626 299404 234682
rect 307604 231074 307660 231130
rect 316724 231222 316780 231278
rect 318932 225302 318988 225358
rect 319508 231370 319564 231426
rect 322484 231518 322540 231574
rect 327284 225450 327340 225506
rect 328052 225598 328108 225654
rect 330260 231666 330316 231722
rect 330836 225746 330892 225802
rect 332564 234034 332620 234090
rect 333812 231814 333868 231870
rect 333044 228114 333100 228170
rect 336884 227374 336940 227430
rect 339380 228262 339436 228318
rect 340148 225894 340204 225950
rect 341588 234182 341644 234238
rect 342548 235662 342604 235718
rect 342164 228410 342220 228466
rect 343124 227226 343180 227282
rect 343988 233146 344044 233202
rect 345428 228558 345484 228614
rect 344756 227078 344812 227134
rect 347636 234774 347692 234830
rect 354068 224562 354124 224618
rect 355892 234922 355948 234978
rect 356852 236106 356908 236162
rect 356756 234922 356812 234978
rect 355604 222638 355660 222694
rect 357236 224414 357292 224470
rect 358964 230038 359020 230094
rect 358580 222934 358636 222990
rect 359828 229002 359884 229058
rect 359732 223970 359788 224026
rect 359444 222786 359500 222842
rect 360788 228706 360844 228762
rect 360308 224266 360364 224322
rect 361460 224118 361516 224174
rect 363572 230186 363628 230242
rect 362804 229150 362860 229206
rect 364052 233738 364108 233794
rect 365684 233294 365740 233350
rect 363764 223822 363820 223878
rect 366644 229890 366700 229946
rect 365684 228854 365740 228910
rect 367220 235514 367276 235570
rect 368948 236402 369004 236458
rect 368660 231814 368716 231870
rect 367604 223674 367660 223730
rect 370388 236698 370444 236754
rect 368660 225154 368716 225210
rect 372212 236994 372268 237050
rect 371156 232998 371212 233054
rect 370772 232850 370828 232906
rect 373460 236846 373516 236902
rect 374036 232702 374092 232758
rect 373076 229742 373132 229798
rect 374900 236254 374956 236310
rect 375380 232554 375436 232610
rect 376724 223378 376780 223434
rect 379508 236550 379564 236606
rect 379124 234478 379180 234534
rect 380084 233294 380140 233350
rect 379892 229594 379948 229650
rect 377588 223526 377644 223582
rect 382388 236550 382444 236606
rect 382580 236550 382636 236606
rect 382100 234330 382156 234386
rect 381716 232406 381772 232462
rect 382676 232110 382732 232166
rect 381332 229446 381388 229502
rect 381236 223230 381292 223286
rect 383540 229298 383596 229354
rect 384980 232258 385036 232314
rect 385268 231962 385324 232018
rect 384404 229150 384460 229206
rect 385844 235958 385900 236014
rect 384308 223082 384364 223138
rect 386996 236994 387052 237050
rect 387092 236550 387148 236606
rect 387188 236402 387244 236458
rect 387476 236994 387532 237050
rect 387572 236698 387628 236754
rect 387476 236402 387532 236458
rect 387476 236293 387478 236310
rect 387478 236293 387530 236310
rect 387530 236293 387532 236310
rect 387476 236254 387532 236293
rect 387860 236994 387916 237050
rect 389876 235810 389932 235866
rect 390740 235662 390796 235718
rect 391604 226930 391660 226986
rect 391220 226782 391276 226838
rect 393044 235662 393100 235718
rect 394100 226634 394156 226690
rect 394484 226486 394540 226542
rect 397076 236254 397132 236310
rect 397460 236698 397516 236754
rect 397364 236254 397420 236310
rect 397460 235514 397516 235570
rect 397748 236994 397804 237050
rect 397844 236863 397900 236902
rect 397844 236846 397846 236863
rect 397846 236846 397898 236863
rect 397898 236846 397900 236863
rect 398036 236846 398092 236902
rect 399860 235514 399916 235570
rect 400244 233886 400300 233942
rect 400244 229002 400300 229058
rect 399476 228854 399532 228910
rect 401396 235366 401452 235422
rect 402740 235218 402796 235274
rect 403124 234922 403180 234978
rect 403988 234922 404044 234978
rect 404372 226338 404428 226394
rect 405428 235070 405484 235126
rect 405332 234774 405388 234830
rect 405524 234774 405580 234830
rect 405716 234626 405772 234682
rect 406484 236106 406540 236162
rect 405908 233738 405964 233794
rect 406004 231814 406060 231870
rect 405812 226190 405868 226246
rect 407444 236698 407500 236754
rect 407444 236254 407500 236310
rect 406484 222490 406540 222546
rect 409940 236106 409996 236162
rect 408500 234626 408556 234682
rect 409844 234478 409900 234534
rect 408116 230334 408172 230390
rect 407636 226042 407692 226098
rect 410036 234330 410092 234386
rect 411380 234478 411436 234534
rect 410804 234330 410860 234386
rect 569012 239954 569068 240010
rect 413396 238918 413452 238974
rect 414068 238770 414124 238826
rect 413684 238622 413740 238678
rect 413972 238326 414028 238382
rect 415220 238178 415276 238234
rect 414452 238030 414508 238086
rect 413684 236254 413740 236310
rect 415220 236254 415276 236310
rect 415412 236254 415468 236310
rect 413876 236106 413932 236162
rect 424724 231074 424780 231130
rect 442868 231222 442924 231278
rect 445172 225302 445228 225358
rect 448916 231370 448972 231426
rect 455156 231518 455212 231574
rect 457268 225450 457324 225506
rect 463316 225598 463372 225654
rect 470132 231666 470188 231722
rect 469364 225746 469420 225802
rect 472340 234034 472396 234090
rect 476180 228114 476236 228170
rect 475316 225154 475372 225210
rect 480884 233886 480940 233942
rect 481460 227374 481516 227430
rect 488276 228262 488332 228318
rect 487508 225894 487564 225950
rect 490484 234182 490540 234238
rect 495092 233146 495148 233202
rect 494228 228410 494284 228466
rect 493460 227226 493516 227282
rect 497972 228558 498028 228614
rect 498836 227078 498892 227134
rect 518420 224562 518476 224618
rect 519860 222638 519916 222694
rect 522932 222490 522988 222546
rect 524468 224414 524524 224470
rect 527540 230038 527596 230094
rect 526004 222934 526060 222990
rect 526676 222786 526732 222842
rect 528308 228706 528364 228762
rect 528980 223970 529036 224026
rect 530516 224266 530572 224322
rect 532052 224118 532108 224174
rect 538004 238030 538060 238086
rect 534260 230186 534316 230242
rect 536564 223822 536620 223878
rect 540308 229890 540364 229946
rect 544340 238326 544396 238382
rect 544052 223674 544108 223730
rect 550196 238622 550252 238678
rect 549428 232998 549484 233054
rect 555380 238918 555436 238974
rect 551636 232850 551692 232906
rect 553940 229742 553996 229798
rect 559892 238178 559948 238234
rect 559220 236550 559276 236606
rect 558452 236402 558508 236458
rect 557684 232702 557740 232758
rect 567476 236846 567532 236902
rect 565268 236698 565324 236754
rect 560756 232554 560812 232610
rect 562964 223526 563020 223582
rect 562196 223378 562252 223434
rect 581780 238770 581836 238826
rect 573140 236994 573196 237050
rect 570452 232406 570508 232462
rect 569780 229594 569836 229650
rect 571316 223230 571372 223286
rect 572756 229446 572812 229502
rect 573524 229298 573580 229354
rect 580340 235958 580396 236014
rect 576596 232258 576652 232314
rect 575828 232110 575884 232166
rect 575060 230334 575116 230390
rect 578036 231962 578092 232018
rect 577268 223082 577324 223138
rect 578900 229150 578956 229206
rect 590420 236106 590476 236162
rect 587924 235810 587980 235866
rect 587444 234330 587500 234386
rect 591476 235662 591532 235718
rect 590900 234478 590956 234534
rect 591668 226930 591724 226986
rect 590900 226782 590956 226838
rect 599924 229002 599980 229058
rect 596180 226634 596236 226690
rect 596948 226486 597004 226542
rect 604532 231814 604588 231870
rect 627188 240102 627244 240158
rect 621140 236254 621196 236310
rect 608276 235514 608332 235570
rect 607508 228854 607564 228910
rect 611252 235366 611308 235422
rect 614324 235218 614380 235274
rect 618836 235070 618892 235126
rect 616628 234922 616684 234978
rect 617300 226338 617356 226394
rect 619604 234774 619660 234830
rect 620372 226190 620428 226246
rect 623348 226042 623404 226098
rect 625556 234626 625612 234682
rect 640148 212278 640204 212334
rect 640148 211538 640204 211594
rect 190292 201326 190348 201382
rect 640148 200882 640204 200938
rect 190292 200512 190348 200568
rect 640148 200142 640204 200198
rect 187220 199106 187276 199162
rect 185972 196738 186028 196794
rect 186068 195998 186124 196054
rect 185780 182382 185836 182438
rect 185588 173206 185644 173262
rect 184532 164770 184588 164826
rect 184340 164047 184396 164086
rect 184340 164030 184342 164047
rect 184342 164030 184394 164047
rect 184394 164030 184396 164047
rect 184340 162550 184396 162606
rect 184532 163290 184588 163346
rect 184436 161810 184492 161866
rect 184436 160922 184492 160978
rect 184532 160330 184588 160386
rect 184340 159442 184396 159498
rect 184628 158850 184684 158906
rect 184340 157962 184396 158018
rect 184436 157370 184492 157426
rect 184532 156482 184588 156538
rect 184628 155594 184684 155650
rect 184340 155002 184396 155058
rect 184436 154114 184492 154170
rect 184532 153522 184588 153578
rect 184628 152634 184684 152690
rect 184340 151894 184396 151950
rect 184436 151154 184492 151210
rect 184532 150414 184588 150470
rect 184340 149674 184396 149730
rect 184436 148934 184492 148990
rect 184532 147306 184588 147362
rect 184340 145826 184396 145882
rect 184436 145086 184492 145142
rect 184628 146605 184630 146622
rect 184630 146605 184682 146622
rect 184682 146605 184684 146622
rect 184628 146566 184684 146605
rect 184532 144346 184588 144402
rect 184340 143606 184396 143662
rect 184436 142718 184492 142774
rect 184628 142126 184684 142182
rect 184532 141238 184588 141294
rect 184340 140498 184396 140554
rect 184436 139758 184492 139814
rect 184532 138870 184588 138926
rect 184340 134430 184396 134486
rect 186068 138278 186124 138334
rect 185972 137390 186028 137446
rect 640244 185638 640300 185694
rect 640244 184898 640300 184954
rect 186740 183122 186796 183178
rect 645140 182974 645196 183030
rect 186260 174686 186316 174742
rect 186164 136798 186220 136854
rect 185780 135170 185836 135226
rect 184436 132950 184492 133006
rect 184340 132227 184396 132266
rect 184340 132210 184342 132227
rect 184342 132210 184394 132227
rect 184394 132210 184396 132227
rect 184436 131470 184492 131526
rect 184532 130582 184588 130638
rect 184628 129842 184684 129898
rect 184340 128362 184396 128418
rect 184436 127622 184492 127678
rect 184532 126882 184588 126938
rect 184436 125994 184492 126050
rect 184340 125402 184396 125458
rect 184532 124514 184588 124570
rect 184340 123791 184396 123830
rect 184340 123774 184342 123791
rect 184342 123774 184394 123791
rect 184394 123774 184396 123791
rect 184436 123034 184492 123090
rect 184340 122146 184396 122202
rect 184532 121554 184588 121610
rect 184340 120666 184396 120722
rect 184436 120074 184492 120130
rect 184532 119186 184588 119242
rect 645140 179274 645196 179330
rect 645140 174873 645142 174890
rect 645142 174873 645194 174890
rect 645194 174873 645196 174890
rect 645140 174834 645196 174873
rect 645140 171025 645142 171042
rect 645142 171025 645194 171042
rect 645194 171025 645196 171042
rect 645140 170986 645196 171025
rect 645140 167730 645196 167786
rect 645140 163329 645142 163346
rect 645142 163329 645194 163346
rect 645194 163329 645196 163346
rect 645140 163290 645196 163329
rect 645140 159442 645196 159498
rect 645140 155446 645196 155502
rect 645140 152525 645142 152542
rect 645142 152525 645194 152542
rect 645194 152525 645196 152542
rect 645140 152486 645196 152525
rect 186740 148046 186796 148102
rect 645140 148046 645196 148102
rect 186452 135910 186508 135966
rect 186260 133690 186316 133746
rect 184724 118594 184780 118650
rect 184340 117706 184396 117762
rect 184436 116966 184492 117022
rect 184532 116226 184588 116282
rect 184628 115338 184684 115394
rect 184340 114746 184396 114802
rect 184436 113858 184492 113914
rect 184532 113118 184588 113174
rect 184628 112378 184684 112434
rect 184340 111638 184396 111694
rect 184436 110898 184492 110954
rect 184532 110158 184588 110214
rect 184340 109309 184342 109326
rect 184342 109309 184394 109326
rect 184394 109309 184396 109326
rect 184340 109270 184396 109309
rect 186740 129102 186796 129158
rect 645716 128954 645772 129010
rect 648596 272070 648652 272126
rect 647348 269258 647404 269314
rect 646580 267038 646636 267094
rect 185684 108678 185740 108734
rect 646676 144198 646732 144254
rect 655412 778230 655468 778286
rect 655220 777638 655276 777694
rect 655124 775862 655180 775918
rect 654356 773494 654412 773550
rect 655124 734422 655180 734478
rect 654164 730130 654220 730186
rect 654068 728502 654124 728558
rect 654740 686914 654796 686970
rect 654164 685286 654220 685342
rect 654068 684546 654124 684602
rect 655316 731610 655372 731666
rect 655220 689430 655276 689486
rect 649748 263486 649804 263542
rect 646772 140942 646828 140998
rect 655124 642366 655180 642422
rect 654164 640590 654220 640646
rect 653972 594118 654028 594174
rect 655604 776010 655660 776066
rect 655508 732646 655564 732702
rect 655412 687062 655468 687118
rect 655316 642958 655372 643014
rect 655220 597818 655276 597874
rect 655124 553270 655180 553326
rect 654164 548534 654220 548590
rect 656564 774678 656620 774734
rect 655700 731314 655756 731370
rect 655604 688394 655660 688450
rect 655508 640738 655564 640794
rect 655412 596634 655468 596690
rect 655316 550902 655372 550958
rect 655796 639110 655852 639166
rect 655988 638222 656044 638278
rect 655604 595450 655660 595506
rect 655508 552086 655564 552142
rect 655796 595302 655852 595358
rect 656564 592934 656620 592990
rect 655700 550754 655756 550810
rect 656564 549718 656620 549774
rect 655316 374338 655372 374394
rect 655124 373302 655180 373358
rect 655508 372118 655564 372174
rect 656564 370934 656620 370990
rect 655220 329790 655276 329846
rect 655316 328014 655372 328070
rect 655124 327422 655180 327478
rect 654164 326238 654220 326294
rect 654164 303298 654220 303354
rect 654068 302114 654124 302170
rect 654260 300930 654316 300986
rect 656564 298710 656620 298766
rect 656276 297526 656332 297582
rect 656084 296786 656140 296842
rect 655892 293974 655948 294030
rect 655796 292790 655852 292846
rect 655604 289238 655660 289294
rect 655412 288054 655468 288110
rect 653780 284502 653836 284558
rect 655124 283318 655180 283374
rect 654164 279766 654220 279822
rect 652244 266890 652300 266946
rect 647060 134726 647116 134782
rect 647828 130878 647884 130934
rect 646964 127622 647020 127678
rect 646868 125698 646924 125754
rect 646580 123774 646636 123830
rect 646484 121998 646540 122054
rect 655316 282282 655372 282338
rect 655220 280950 655276 281006
rect 655508 285686 655564 285742
rect 655700 286870 655756 286926
rect 655988 290866 656044 290922
rect 656180 291606 656236 291662
rect 656372 295158 656428 295214
rect 647924 119482 647980 119538
rect 645236 117558 645292 117614
rect 647924 115634 647980 115690
rect 669524 275430 669580 275486
rect 669716 275578 669772 275634
rect 670004 354654 670060 354710
rect 669908 277842 669964 277898
rect 670196 355986 670252 356042
rect 670100 277398 670156 277454
rect 670388 308922 670444 308978
rect 670292 277546 670348 277602
rect 670196 277162 670252 277218
rect 672404 278582 672460 278638
rect 670676 277990 670732 278046
rect 670484 277694 670540 277750
rect 670388 277014 670444 277070
rect 670004 273550 670060 273606
rect 676052 891467 676108 891506
rect 676052 891450 676054 891467
rect 676054 891450 676106 891467
rect 676106 891450 676108 891467
rect 676052 890431 676108 890470
rect 676052 890414 676054 890431
rect 676054 890414 676106 890431
rect 676106 890414 676108 890431
rect 680180 890118 680236 890174
rect 676244 889230 676300 889286
rect 679988 888638 680044 888694
rect 676244 887750 676300 887806
rect 676052 887380 676108 887436
rect 679700 886714 679756 886770
rect 676052 885456 676108 885512
rect 676052 884938 676108 884994
rect 676244 884215 676300 884254
rect 676244 884198 676246 884215
rect 676246 884198 676298 884215
rect 676298 884198 676300 884215
rect 676052 883976 676108 884032
rect 675956 883458 676012 883514
rect 679796 886122 679852 886178
rect 679700 882718 679756 882774
rect 679700 882126 679756 882182
rect 679892 885678 679948 885734
rect 680084 888194 680140 888250
rect 685460 882126 685516 882182
rect 685460 881682 685516 881738
rect 675092 788294 675148 788350
rect 675476 787110 675532 787166
rect 675092 786222 675148 786278
rect 675380 784742 675436 784798
rect 675476 784298 675532 784354
rect 675092 783410 675148 783466
rect 674708 734274 674764 734330
rect 675764 782966 675820 783022
rect 675764 780598 675820 780654
rect 675764 780006 675820 780062
rect 675764 778822 675820 778878
rect 675284 771866 675340 771922
rect 675476 742414 675532 742470
rect 675668 741674 675724 741730
rect 675380 740046 675436 740102
rect 675764 739158 675820 739214
rect 675380 738566 675436 738622
rect 675764 735014 675820 735070
rect 675476 734422 675532 734478
rect 676340 715478 676396 715534
rect 676148 714886 676204 714942
rect 676244 714755 676300 714794
rect 676244 714738 676246 714755
rect 676298 714738 676300 714755
rect 679700 713850 679756 713906
rect 679700 713258 679756 713314
rect 676052 713127 676108 713166
rect 676052 713110 676054 713127
rect 676106 713110 676108 713127
rect 676052 712683 676108 712722
rect 676052 712666 676054 712683
rect 676106 712666 676108 712683
rect 676244 711943 676300 711982
rect 676244 711926 676246 711943
rect 676298 711926 676300 711943
rect 676052 711573 676108 711612
rect 676052 711556 676054 711573
rect 676106 711556 676108 711573
rect 676052 710594 676108 710650
rect 676052 708522 676108 708578
rect 676052 708152 676108 708208
rect 676052 706672 676108 706728
rect 676244 706302 676300 706358
rect 679988 704378 680044 704434
rect 679796 703342 679852 703398
rect 679988 703342 680044 703398
rect 679796 702898 679852 702954
rect 675380 697866 675436 697922
rect 675092 697126 675148 697182
rect 675092 696978 675148 697034
rect 675764 694906 675820 694962
rect 675092 694610 675148 694666
rect 675476 693426 675532 693482
rect 675188 686766 675244 686822
rect 676148 670338 676204 670394
rect 676052 669193 676054 669210
rect 676106 669193 676108 669210
rect 676052 669154 676108 669193
rect 676052 668562 676108 668618
rect 676340 669746 676396 669802
rect 676244 669302 676300 669358
rect 675956 668061 676012 668100
rect 675956 668044 675958 668061
rect 676010 668044 676012 668061
rect 675956 667691 676012 667730
rect 675956 667674 675958 667691
rect 676010 667674 676012 667691
rect 676244 666934 676300 666990
rect 676244 666359 676300 666398
rect 676244 666342 676246 666359
rect 676298 666342 676300 666359
rect 676052 665602 676108 665658
rect 676244 664270 676300 664326
rect 676052 663530 676108 663586
rect 676052 661606 676108 661662
rect 676052 660609 676054 660626
rect 676106 660609 676108 660626
rect 676052 660570 676108 660609
rect 676244 659869 676246 659886
rect 676298 659869 676300 659886
rect 676244 659830 676300 659869
rect 679796 659238 679852 659294
rect 679796 658350 679852 658406
rect 685460 658350 685516 658406
rect 685460 657906 685516 657962
rect 675476 652134 675532 652190
rect 675476 651394 675532 651450
rect 675092 650950 675148 651006
rect 675668 649766 675724 649822
rect 675188 648286 675244 648342
rect 675764 648286 675820 648342
rect 675764 645326 675820 645382
rect 676244 625050 676300 625106
rect 676148 624606 676204 624662
rect 676052 623439 676108 623478
rect 676052 623422 676054 623439
rect 676106 623422 676108 623439
rect 676052 622830 676108 622886
rect 676052 622477 676108 622516
rect 676052 622460 676054 622477
rect 676106 622460 676108 622477
rect 676244 624162 676300 624218
rect 679700 624162 679756 624218
rect 676052 621959 676108 621998
rect 676052 621942 676054 621959
rect 676106 621942 676108 621959
rect 676052 621367 676108 621406
rect 676052 621350 676054 621367
rect 676106 621350 676108 621367
rect 676244 620610 676300 620666
rect 676052 618908 676108 618964
rect 676244 618538 676300 618594
rect 676052 616466 676108 616522
rect 676052 615874 676108 615930
rect 676244 615617 676246 615634
rect 676298 615617 676300 615634
rect 676244 615578 676300 615617
rect 676052 614433 676054 614450
rect 676106 614433 676108 614450
rect 676052 614394 676108 614433
rect 679988 613654 680044 613710
rect 679796 613210 679852 613266
rect 679988 613210 680044 613266
rect 679796 612766 679852 612822
rect 675092 607734 675148 607790
rect 675092 607438 675148 607494
rect 675764 606402 675820 606458
rect 675092 604774 675148 604830
rect 675284 601962 675340 602018
rect 675764 600186 675820 600242
rect 676340 578282 676396 578338
rect 676148 577542 676204 577598
rect 676244 577098 676300 577154
rect 679700 577098 679756 577154
rect 676244 576227 676300 576266
rect 676244 576210 676246 576227
rect 676298 576210 676300 576227
rect 675956 575931 676012 575970
rect 675956 575914 675958 575931
rect 676010 575914 676012 575931
rect 675956 575487 676012 575526
rect 675956 575470 675958 575487
rect 676010 575470 676012 575487
rect 675956 574917 675958 574934
rect 676010 574917 676012 574934
rect 675956 574878 676012 574917
rect 676244 574155 676300 574194
rect 676244 574138 676246 574155
rect 676298 574138 676300 574155
rect 676052 573398 676108 573454
rect 676052 571326 676108 571382
rect 676052 569515 676054 569532
rect 676106 569515 676108 569532
rect 676052 569476 676108 569515
rect 676244 569145 676246 569162
rect 676298 569145 676300 569162
rect 676244 569106 676300 569145
rect 676052 568405 676054 568422
rect 676106 568405 676108 568422
rect 676052 568366 676108 568405
rect 676052 567961 676054 567978
rect 676106 567961 676108 567978
rect 676052 567922 676108 567961
rect 676244 567665 676246 567682
rect 676298 567665 676300 567682
rect 676244 567626 676300 567665
rect 679796 567034 679852 567090
rect 679796 566146 679852 566202
rect 685460 566146 685516 566202
rect 685460 565702 685516 565758
rect 675092 562890 675148 562946
rect 675476 561706 675532 561762
rect 675380 561410 675436 561466
rect 675476 558894 675532 558950
rect 675764 554602 675820 554658
rect 675284 553270 675340 553326
rect 676244 534918 676300 534974
rect 676148 534326 676204 534382
rect 676052 534178 676108 534234
rect 679700 533586 679756 533642
rect 676532 532994 676588 533050
rect 675956 532715 676012 532754
rect 675956 532698 675958 532715
rect 676010 532698 676012 532715
rect 676244 531531 676300 531570
rect 676244 531514 676246 531531
rect 676298 531514 676300 531531
rect 676052 530182 676108 530238
rect 676052 528110 676108 528166
rect 676052 526669 676054 526686
rect 676106 526669 676108 526686
rect 676052 526630 676108 526669
rect 676052 526299 676054 526316
rect 676106 526299 676108 526316
rect 676052 526260 676108 526299
rect 676244 525929 676246 525946
rect 676298 525929 676300 525946
rect 676244 525890 676300 525929
rect 676052 525189 676054 525206
rect 676106 525189 676108 525206
rect 676052 525150 676108 525189
rect 676052 524819 676054 524836
rect 676106 524819 676108 524836
rect 676052 524780 676108 524819
rect 676244 524449 676246 524466
rect 676298 524449 676300 524466
rect 676244 524410 676300 524449
rect 676628 531958 676684 532014
rect 676244 490518 676300 490574
rect 676148 490074 676204 490130
rect 676244 489943 676300 489982
rect 676244 489926 676246 489943
rect 676298 489926 676300 489943
rect 676052 488298 676108 488354
rect 675284 487854 675340 487910
rect 676724 530922 676780 530978
rect 679796 523522 679852 523578
rect 679796 522930 679852 522986
rect 685460 522930 685516 522986
rect 685460 522486 685516 522542
rect 679700 489186 679756 489242
rect 676724 488594 676780 488650
rect 676244 487131 676300 487170
rect 676244 487114 676246 487131
rect 676298 487114 676300 487131
rect 676052 486835 676108 486874
rect 676052 486818 676054 486835
rect 676106 486818 676108 486835
rect 676052 485782 676108 485838
rect 676244 485042 676300 485098
rect 676052 484302 676108 484358
rect 675956 483727 676012 483766
rect 675956 483710 675958 483727
rect 676010 483710 676012 483727
rect 676052 482230 676108 482286
rect 676052 481860 676108 481916
rect 676244 481490 676300 481546
rect 676244 480049 676246 480066
rect 676298 480049 676300 480066
rect 676244 480010 676300 480049
rect 676148 402310 676204 402366
rect 676052 401570 676108 401626
rect 675956 400625 676012 400664
rect 675956 400608 675958 400625
rect 676010 400608 676012 400625
rect 676244 401866 676300 401922
rect 679892 479122 679948 479178
rect 679700 478530 679756 478586
rect 679892 478530 679948 478586
rect 679700 478086 679756 478142
rect 676724 400978 676780 401034
rect 676244 400277 676246 400294
rect 676298 400277 676300 400294
rect 676244 400238 676300 400277
rect 676052 399071 676108 399110
rect 676052 399054 676054 399071
rect 676106 399054 676108 399071
rect 675572 396982 675628 397038
rect 675284 395206 675340 395262
rect 676244 393874 676300 393930
rect 676244 392394 676300 392450
rect 679796 390914 679852 390970
rect 679796 390322 679852 390378
rect 685460 390322 685516 390378
rect 685460 389878 685516 389934
rect 675764 384698 675820 384754
rect 675764 382922 675820 382978
rect 675476 382330 675532 382386
rect 675764 378778 675820 378834
rect 675764 378038 675820 378094
rect 675476 377150 675532 377206
rect 675188 376410 675244 376466
rect 675476 375670 675532 375726
rect 675092 374338 675148 374394
rect 675764 371970 675820 372026
rect 676148 358058 676204 358114
rect 676244 357318 676300 357374
rect 676052 357187 676108 357226
rect 676052 357170 676054 357187
rect 676106 357170 676108 357187
rect 676052 356765 676054 356782
rect 676106 356765 676108 356782
rect 676052 356726 676108 356765
rect 676052 353766 676108 353822
rect 675572 352582 675628 352638
rect 675284 350806 675340 350862
rect 676052 352286 676108 352342
rect 676916 351546 676972 351602
rect 676052 350214 676108 350270
rect 676244 349474 676300 349530
rect 676820 349030 676876 349086
rect 676244 347994 676300 348050
rect 676052 347772 676108 347828
rect 675956 347254 676012 347310
rect 676820 342962 676876 343018
rect 679892 346514 679948 346570
rect 679892 346070 679948 346126
rect 679700 345922 679756 345978
rect 679700 345478 679756 345534
rect 676916 342814 676972 342870
rect 675764 333490 675820 333546
rect 675476 332306 675532 332362
rect 675764 330530 675820 330586
rect 675092 328162 675148 328218
rect 675380 326830 675436 326886
rect 676340 312178 676396 312234
rect 676148 311586 676204 311642
rect 676244 311181 676246 311198
rect 676298 311181 676300 311198
rect 676244 311142 676300 311181
rect 676244 306702 676300 306758
rect 676244 304778 676300 304834
rect 676052 304408 676108 304464
rect 675956 303890 676012 303946
rect 679988 300634 680044 300690
rect 679796 300190 679852 300246
rect 679988 300190 680044 300246
rect 679796 299746 679852 299802
rect 675764 294566 675820 294622
rect 675380 292790 675436 292846
rect 675764 290718 675820 290774
rect 675668 288498 675724 288554
rect 675572 287758 675628 287814
rect 675476 287166 675532 287222
rect 675764 286574 675820 286630
rect 675476 285538 675532 285594
rect 675092 283170 675148 283226
rect 675092 282134 675148 282190
rect 675092 278286 675148 278342
rect 672596 278138 672652 278194
rect 672500 273402 672556 273458
rect 679700 270590 679756 270646
rect 676148 266890 676204 266946
rect 672404 266742 672460 266798
rect 672596 266594 672652 266650
rect 672404 174686 672460 174742
rect 676052 266150 676108 266206
rect 676244 266446 676300 266502
rect 679700 264818 679756 264874
rect 676052 264226 676108 264282
rect 679796 264078 679852 264134
rect 676244 262598 676300 262654
rect 676052 261266 676108 261322
rect 675284 259786 675340 259842
rect 676820 259934 676876 259990
rect 676052 259233 676054 259250
rect 676106 259233 676108 259250
rect 676052 259194 676108 259233
rect 676052 258676 676108 258732
rect 676244 256974 676300 257030
rect 676052 256826 676108 256882
rect 676052 256234 676108 256290
rect 679700 255494 679756 255550
rect 679700 254902 679756 254958
rect 685460 254902 685516 254958
rect 685460 254458 685516 254514
rect 676820 253274 676876 253330
rect 675764 250758 675820 250814
rect 675668 243506 675724 243562
rect 675092 241878 675148 241934
rect 675188 240990 675244 241046
rect 675092 238178 675148 238234
rect 675764 236846 675820 236902
rect 676244 221789 676246 221806
rect 676298 221789 676300 221806
rect 676244 221750 676300 221789
rect 676148 221158 676204 221214
rect 676052 219495 676054 219512
rect 676106 219495 676108 219512
rect 676052 219456 676108 219495
rect 676244 220714 676300 220770
rect 676916 216718 676972 216774
rect 675764 216422 675820 216478
rect 676052 216069 676108 216108
rect 676052 216052 676054 216069
rect 676106 216052 676108 216069
rect 676820 214794 676876 214850
rect 676052 214572 676108 214628
rect 675956 214054 676012 214110
rect 676244 213331 676300 213370
rect 676244 213314 676246 213331
rect 676298 213314 676300 213331
rect 676052 212574 676108 212630
rect 676052 211982 676108 212038
rect 675956 211020 676012 211076
rect 676244 211390 676300 211446
rect 676820 207542 676876 207598
rect 679796 210650 679852 210706
rect 679796 209762 679852 209818
rect 685460 209762 685516 209818
rect 676916 207394 676972 207450
rect 685460 209318 685516 209374
rect 675668 204434 675724 204490
rect 675764 198366 675820 198422
rect 675092 194814 675148 194870
rect 675764 193482 675820 193538
rect 675764 191558 675820 191614
rect 676148 177350 676204 177406
rect 676340 176758 676396 176814
rect 676244 176314 676300 176370
rect 672596 173502 672652 173558
rect 675572 172022 675628 172078
rect 676052 170172 676108 170228
rect 676052 169654 676108 169710
rect 676244 168914 676300 168970
rect 676052 166102 676108 166158
rect 676148 165362 676204 165418
rect 676244 164770 676300 164826
rect 675764 159294 675820 159350
rect 675476 157666 675532 157722
rect 675764 155446 675820 155502
rect 675092 155298 675148 155354
rect 675188 152486 675244 152542
rect 675668 152486 675724 152542
rect 675764 151302 675820 151358
rect 675476 150266 675532 150322
rect 675092 149674 675148 149730
rect 675764 146566 675820 146622
rect 676148 131766 676204 131822
rect 676340 131174 676396 131230
rect 676244 130730 676300 130786
rect 676244 129694 676300 129750
rect 676148 128806 676204 128862
rect 676052 127548 676108 127604
rect 676244 127770 676300 127826
rect 676916 126734 676972 126790
rect 646484 113118 646540 113174
rect 186164 107790 186220 107846
rect 184436 107050 184492 107106
rect 184340 105570 184396 105626
rect 185300 106349 185302 106366
rect 185302 106349 185354 106366
rect 185354 106349 185356 106366
rect 185300 106310 185356 106349
rect 646100 106014 646156 106070
rect 184532 104830 184588 104886
rect 184436 103942 184492 103998
rect 184436 103350 184492 103406
rect 184340 102462 184396 102518
rect 184532 101870 184588 101926
rect 184628 100982 184684 101038
rect 184340 100242 184396 100298
rect 184436 99502 184492 99558
rect 184532 98614 184588 98670
rect 184628 98022 184684 98078
rect 184340 97134 184396 97190
rect 184436 96394 184492 96450
rect 184724 95654 184780 95710
rect 184340 94783 184396 94822
rect 184340 94766 184342 94783
rect 184342 94766 184394 94783
rect 184394 94766 184396 94783
rect 184436 94174 184492 94230
rect 184532 93434 184588 93490
rect 184628 92694 184684 92750
rect 184340 91971 184396 92010
rect 184340 91954 184342 91971
rect 184342 91954 184394 91971
rect 184394 91954 184396 91971
rect 184436 90326 184492 90382
rect 184628 91066 184684 91122
rect 184532 89586 184588 89642
rect 184340 88846 184396 88902
rect 184436 88106 184492 88162
rect 184532 87218 184588 87274
rect 184628 86626 184684 86682
rect 184436 85738 184492 85794
rect 184340 85146 184396 85202
rect 184532 84258 184588 84314
rect 184340 83409 184342 83426
rect 184342 83409 184394 83426
rect 184394 83409 184396 83426
rect 184340 83370 184396 83409
rect 184244 81890 184300 81946
rect 645140 102166 645196 102222
rect 645428 95967 645484 96006
rect 645428 95950 645430 95967
rect 645430 95950 645482 95967
rect 645482 95950 645484 95967
rect 645908 88846 645964 88902
rect 186164 82778 186220 82834
rect 184436 81298 184492 81354
rect 184436 79818 184492 79874
rect 184340 78930 184396 78986
rect 184628 80427 184684 80466
rect 184628 80410 184630 80427
rect 184630 80410 184682 80427
rect 184682 80410 184684 80427
rect 184532 78190 184588 78246
rect 184436 77450 184492 77506
rect 184340 76710 184396 76766
rect 184628 75970 184684 76026
rect 184532 75082 184588 75138
rect 184340 74342 184396 74398
rect 149684 73010 149740 73066
rect 149492 70790 149548 70846
rect 149396 69458 149452 69514
rect 149300 68274 149356 68330
rect 149204 67090 149260 67146
rect 184532 73602 184588 73658
rect 184436 72862 184492 72918
rect 184628 72122 184684 72178
rect 184340 71382 184396 71438
rect 184436 70494 184492 70550
rect 184532 69902 184588 69958
rect 184340 69031 184396 69070
rect 184340 69014 184342 69031
rect 184342 69014 184394 69031
rect 184394 69014 184396 69031
rect 184340 68422 184396 68478
rect 184532 67534 184588 67590
rect 184436 66794 184492 66850
rect 184340 66093 184342 66110
rect 184342 66093 184394 66110
rect 184394 66093 184396 66110
rect 184340 66054 184396 66093
rect 149396 65314 149452 65370
rect 149492 64574 149548 64630
rect 184532 65166 184588 65222
rect 184436 64574 184492 64630
rect 184340 63686 184396 63742
rect 149588 63390 149644 63446
rect 149396 62206 149452 62262
rect 149300 60578 149356 60634
rect 184436 63094 184492 63150
rect 184340 62206 184396 62262
rect 184628 61466 184684 61522
rect 184532 60726 184588 60782
rect 184340 59986 184396 60042
rect 149396 59690 149452 59746
rect 184436 59246 184492 59302
rect 149396 58506 149452 58562
rect 184532 58358 184588 58414
rect 184340 57618 184396 57674
rect 149492 57322 149548 57378
rect 184340 56878 184396 56934
rect 149396 56155 149452 56194
rect 184340 56177 184342 56194
rect 184342 56177 184394 56194
rect 184394 56177 184396 56194
rect 149396 56138 149398 56155
rect 149398 56138 149450 56155
rect 149450 56138 149452 56155
rect 184340 56138 184396 56177
rect 184436 55398 184492 55454
rect 149684 54806 149740 54862
rect 184340 54675 184396 54714
rect 184340 54658 184342 54675
rect 184342 54658 184394 54675
rect 184394 54658 184396 54675
rect 184340 53918 184396 53974
rect 149396 53770 149452 53826
rect 142100 40302 142156 40358
rect 302900 42078 302956 42134
rect 311156 42078 311212 42134
rect 357716 41782 357772 41838
rect 362036 41782 362092 41838
rect 389204 41782 389260 41838
rect 412532 42078 412588 42134
rect 416852 41930 416908 41986
rect 403220 40450 403276 40506
rect 467348 41782 467404 41838
rect 471668 41782 471724 41838
rect 458612 40450 458668 40506
rect 475700 40598 475756 40654
rect 522836 41782 522892 41838
rect 645716 84406 645772 84462
rect 646292 75526 646348 75582
rect 647156 111342 647212 111398
rect 646676 109418 646732 109474
rect 646772 107938 646828 107994
rect 647060 98022 647116 98078
rect 646676 79374 646732 79430
rect 646004 66219 646060 66258
rect 646004 66202 646006 66219
rect 646006 66202 646058 66219
rect 646058 66202 646060 66219
rect 646004 58950 646060 59006
rect 665204 105570 665260 105626
rect 676244 126290 676300 126346
rect 676052 126068 676108 126124
rect 676052 124514 676108 124570
rect 675956 124087 676012 124126
rect 675956 124070 675958 124087
rect 676010 124070 676012 124087
rect 676820 124810 676876 124866
rect 676052 123478 676108 123534
rect 676052 121998 676108 122054
rect 676244 121406 676300 121462
rect 676052 121053 676108 121092
rect 676052 121036 676054 121053
rect 676106 121036 676108 121053
rect 676052 120518 676108 120574
rect 676148 119778 676204 119834
rect 676244 119186 676300 119242
rect 676820 118002 676876 118058
rect 676916 117854 676972 117910
rect 675188 107642 675244 107698
rect 675092 106458 675148 106514
rect 675092 105570 675148 105626
rect 665588 105274 665644 105330
rect 665300 105126 665356 105182
rect 647924 104090 647980 104146
rect 647924 99650 647980 99706
rect 647732 94026 647788 94082
rect 647828 92694 647884 92750
rect 647924 87070 647980 87126
rect 650900 86182 650956 86238
rect 652340 85294 652396 85350
rect 652244 83370 652300 83426
rect 647924 82630 647980 82686
rect 647924 81002 647980 81058
rect 647924 77489 647926 77506
rect 647926 77489 647978 77506
rect 647978 77489 647980 77506
rect 647924 77450 647980 77489
rect 646964 71826 647020 71882
rect 646868 68570 646924 68626
rect 647924 73602 647980 73658
rect 647924 69623 647980 69662
rect 647924 69606 647926 69623
rect 647926 69606 647978 69623
rect 647978 69606 647980 69623
rect 647924 64130 647980 64186
rect 647924 62206 647980 62262
rect 647156 60282 647212 60338
rect 653684 86922 653740 86978
rect 653684 84258 653740 84314
rect 652436 82630 652492 82686
rect 646772 57026 646828 57082
rect 646484 54658 646540 54714
rect 659348 90770 659404 90826
rect 675764 103202 675820 103258
rect 675764 101426 675820 101482
rect 663284 86330 663340 86386
rect 662420 81611 662476 81650
rect 662420 81594 662422 81611
rect 662422 81594 662474 81611
rect 662474 81594 662476 81611
rect 663284 84702 663340 84758
rect 663476 83962 663532 84018
rect 663380 82778 663436 82834
rect 663284 82038 663340 82094
rect 541460 40450 541516 40506
rect 311060 37194 311116 37250
rect 334100 37194 334156 37250
<< metal3 >>
rect 483663 1005172 483729 1005175
rect 535023 1005172 535089 1005175
rect 636879 1005172 636945 1005175
rect 483663 1005170 483744 1005172
rect 483663 1005114 483668 1005170
rect 483724 1005114 483744 1005170
rect 483663 1005112 483744 1005114
rect 535008 1005170 535089 1005172
rect 535008 1005114 535028 1005170
rect 535084 1005114 535089 1005170
rect 535008 1005112 535089 1005114
rect 636768 1005170 636945 1005172
rect 636768 1005114 636884 1005170
rect 636940 1005114 636945 1005170
rect 636768 1005112 636945 1005114
rect 483663 1005109 483729 1005112
rect 535023 1005109 535089 1005112
rect 636879 1005109 636945 1005112
rect 241218 997740 241278 997742
rect 679695 964176 679761 964179
rect 679695 964174 679806 964176
rect 679695 964118 679700 964174
rect 679756 964118 679806 964174
rect 679695 964113 679806 964118
rect 679746 963554 679806 964113
rect 649455 961660 649521 961663
rect 649248 961658 649521 961660
rect 649248 961602 649460 961658
rect 649516 961602 649521 961658
rect 649248 961600 649521 961602
rect 649455 961597 649521 961600
rect 676143 894172 676209 894175
rect 676290 894172 676350 894438
rect 676143 894170 676350 894172
rect 676143 894114 676148 894170
rect 676204 894114 676350 894170
rect 676143 894112 676350 894114
rect 676143 894109 676209 894112
rect 676290 893583 676350 893920
rect 676239 893578 676350 893583
rect 676239 893522 676244 893578
rect 676300 893522 676350 893578
rect 676239 893520 676350 893522
rect 676239 893517 676305 893520
rect 676047 893432 676113 893435
rect 676047 893430 676320 893432
rect 676047 893374 676052 893430
rect 676108 893374 676320 893430
rect 676047 893372 676320 893374
rect 676047 893369 676113 893372
rect 676047 892470 676113 892473
rect 676047 892468 676320 892470
rect 676047 892412 676052 892468
rect 676108 892412 676320 892468
rect 676047 892410 676320 892412
rect 676047 892407 676113 892410
rect 676047 891508 676113 891511
rect 676047 891506 676320 891508
rect 676047 891450 676052 891506
rect 676108 891450 676320 891506
rect 676047 891448 676320 891450
rect 676047 891445 676113 891448
rect 676047 890472 676113 890475
rect 676047 890470 676320 890472
rect 676047 890414 676052 890470
rect 676108 890414 676320 890470
rect 676047 890412 676320 890414
rect 676047 890409 676113 890412
rect 680175 890176 680241 890179
rect 680130 890174 680241 890176
rect 680130 890118 680180 890174
rect 680236 890118 680241 890174
rect 680130 890113 680241 890118
rect 680130 889998 680190 890113
rect 676290 889291 676350 889406
rect 676239 889286 676350 889291
rect 676239 889230 676244 889286
rect 676300 889230 676350 889286
rect 676239 889228 676350 889230
rect 676239 889225 676305 889228
rect 679938 888699 679998 888888
rect 679938 888694 680049 888699
rect 679938 888638 679988 888694
rect 680044 888638 680049 888694
rect 679938 888636 680049 888638
rect 679983 888633 680049 888636
rect 680130 888255 680190 888518
rect 680079 888250 680190 888255
rect 680079 888194 680084 888250
rect 680140 888194 680190 888250
rect 680079 888192 680190 888194
rect 680079 888189 680145 888192
rect 676290 887811 676350 887926
rect 676239 887806 676350 887811
rect 676239 887750 676244 887806
rect 676300 887750 676350 887806
rect 676239 887748 676350 887750
rect 676239 887745 676305 887748
rect 676047 887438 676113 887441
rect 676047 887436 676320 887438
rect 676047 887380 676052 887436
rect 676108 887380 676320 887436
rect 676047 887378 676320 887380
rect 676047 887375 676113 887378
rect 679746 886775 679806 887038
rect 679695 886770 679806 886775
rect 679695 886714 679700 886770
rect 679756 886714 679806 886770
rect 679695 886712 679806 886714
rect 679695 886709 679761 886712
rect 679746 886183 679806 886446
rect 679746 886178 679857 886183
rect 679746 886122 679796 886178
rect 679852 886122 679857 886178
rect 679746 886120 679857 886122
rect 679791 886117 679857 886120
rect 679938 885739 679998 885854
rect 679887 885734 679998 885739
rect 679887 885678 679892 885734
rect 679948 885678 679998 885734
rect 679887 885676 679998 885678
rect 679887 885673 679953 885676
rect 676047 885514 676113 885517
rect 676047 885512 676320 885514
rect 676047 885456 676052 885512
rect 676108 885456 676320 885512
rect 676047 885454 676320 885456
rect 676047 885451 676113 885454
rect 676047 884996 676113 884999
rect 676047 884994 676320 884996
rect 676047 884938 676052 884994
rect 676108 884938 676320 884994
rect 676047 884936 676320 884938
rect 676047 884933 676113 884936
rect 676290 884259 676350 884374
rect 676239 884254 676350 884259
rect 676239 884198 676244 884254
rect 676300 884198 676350 884254
rect 676239 884196 676350 884198
rect 676239 884193 676305 884196
rect 676047 884034 676113 884037
rect 676047 884032 676320 884034
rect 676047 883976 676052 884032
rect 676108 883976 676320 884032
rect 676047 883974 676320 883976
rect 676047 883971 676113 883974
rect 675951 883516 676017 883519
rect 675951 883514 676320 883516
rect 675951 883458 675956 883514
rect 676012 883458 676320 883514
rect 675951 883456 676320 883458
rect 675951 883453 676017 883456
rect 679746 882779 679806 882894
rect 679695 882774 679806 882779
rect 679695 882718 679700 882774
rect 679756 882718 679806 882774
rect 679695 882716 679806 882718
rect 679695 882713 679761 882716
rect 685506 882187 685566 882450
rect 679695 882184 679761 882187
rect 679695 882182 679806 882184
rect 679695 882126 679700 882182
rect 679756 882126 679806 882182
rect 679695 882121 679806 882126
rect 685455 882182 685566 882187
rect 685455 882126 685460 882182
rect 685516 882126 685566 882182
rect 685455 882124 685566 882126
rect 685455 882121 685521 882124
rect 679746 882006 679806 882121
rect 685455 881740 685521 881743
rect 685455 881738 685566 881740
rect 685455 881682 685460 881738
rect 685516 881682 685566 881738
rect 685455 881677 685566 881682
rect 685506 881414 685566 881677
rect 655407 868864 655473 868867
rect 649986 868862 655473 868864
rect 649986 868806 655412 868862
rect 655468 868806 655473 868862
rect 649986 868804 655473 868806
rect 649986 868246 650046 868804
rect 655407 868801 655473 868804
rect 655215 867680 655281 867683
rect 649986 867678 655281 867680
rect 649986 867622 655220 867678
rect 655276 867622 655281 867678
rect 649986 867620 655281 867622
rect 649986 867064 650046 867620
rect 655215 867617 655281 867620
rect 655119 866496 655185 866499
rect 649986 866494 655185 866496
rect 649986 866438 655124 866494
rect 655180 866438 655185 866494
rect 649986 866436 655185 866438
rect 649986 865882 650046 866436
rect 655119 866433 655185 866436
rect 655311 865312 655377 865315
rect 649986 865310 655377 865312
rect 649986 865254 655316 865310
rect 655372 865254 655377 865310
rect 649986 865252 655377 865254
rect 649986 864700 650046 865252
rect 655311 865249 655377 865252
rect 654159 863980 654225 863983
rect 649986 863978 654225 863980
rect 649986 863922 654164 863978
rect 654220 863922 654225 863978
rect 649986 863920 654225 863922
rect 649986 863518 650046 863920
rect 654159 863917 654225 863920
rect 653775 862944 653841 862947
rect 649986 862942 653841 862944
rect 649986 862886 653780 862942
rect 653836 862886 653841 862942
rect 649986 862884 653841 862886
rect 649986 862336 650046 862884
rect 653775 862881 653841 862884
rect 41775 817952 41841 817955
rect 41568 817950 41841 817952
rect 41568 817894 41780 817950
rect 41836 817894 41841 817950
rect 41568 817892 41841 817894
rect 41775 817889 41841 817892
rect 41775 817360 41841 817363
rect 41568 817358 41841 817360
rect 41568 817302 41780 817358
rect 41836 817302 41841 817358
rect 41568 817300 41841 817302
rect 41775 817297 41841 817300
rect 41538 816623 41598 816738
rect 41538 816618 41649 816623
rect 41538 816562 41588 816618
rect 41644 816562 41649 816618
rect 41538 816560 41649 816562
rect 41583 816557 41649 816560
rect 41775 815880 41841 815883
rect 41568 815878 41841 815880
rect 41568 815822 41780 815878
rect 41836 815822 41841 815878
rect 41568 815820 41841 815822
rect 41775 815817 41841 815820
rect 40386 815142 40446 815258
rect 40378 815078 40384 815142
rect 40448 815078 40454 815142
rect 41775 814918 41841 814921
rect 41568 814916 41841 814918
rect 41568 814860 41780 814916
rect 41836 814860 41841 814916
rect 41568 814858 41841 814860
rect 41775 814855 41841 814858
rect 40578 814106 40638 814370
rect 40570 814042 40576 814106
rect 40640 814042 40646 814106
rect 41538 813663 41598 813778
rect 41538 813658 41649 813663
rect 41538 813602 41588 813658
rect 41644 813602 41649 813658
rect 41538 813600 41649 813602
rect 41583 813597 41649 813600
rect 41538 813219 41598 813334
rect 41538 813214 41649 813219
rect 41538 813158 41588 813214
rect 41644 813158 41649 813214
rect 41538 813156 41649 813158
rect 41583 813153 41649 813156
rect 42255 812920 42321 812923
rect 41568 812918 42321 812920
rect 41568 812862 42260 812918
rect 42316 812862 42321 812918
rect 41568 812860 42321 812862
rect 42255 812857 42321 812860
rect 40239 812476 40305 812479
rect 40194 812474 40305 812476
rect 40194 812418 40244 812474
rect 40300 812418 40305 812474
rect 40194 812413 40305 812418
rect 40194 812298 40254 812413
rect 41538 811739 41598 811854
rect 41487 811734 41598 811739
rect 41487 811678 41492 811734
rect 41548 811678 41598 811734
rect 41487 811676 41598 811678
rect 41487 811673 41553 811676
rect 41775 811366 41841 811369
rect 41568 811364 41841 811366
rect 41568 811308 41780 811364
rect 41836 811308 41841 811364
rect 41568 811306 41841 811308
rect 41775 811303 41841 811306
rect 41871 810848 41937 810851
rect 41568 810846 41937 810848
rect 41568 810790 41876 810846
rect 41932 810790 41937 810846
rect 41568 810788 41937 810790
rect 41871 810785 41937 810788
rect 41346 810258 41406 810374
rect 41338 810194 41344 810258
rect 41408 810194 41414 810258
rect 41538 809812 41598 809856
rect 42159 809812 42225 809815
rect 41538 809810 42225 809812
rect 41538 809754 42164 809810
rect 42220 809754 42225 809810
rect 41538 809752 42225 809754
rect 42159 809749 42225 809752
rect 42063 809368 42129 809371
rect 41568 809366 42129 809368
rect 41568 809310 42068 809366
rect 42124 809310 42129 809366
rect 41568 809308 42129 809310
rect 42063 809305 42129 809308
rect 41775 808924 41841 808927
rect 41568 808922 41841 808924
rect 41568 808866 41780 808922
rect 41836 808866 41841 808922
rect 41568 808864 41841 808866
rect 41775 808861 41841 808864
rect 41538 808187 41598 808302
rect 41538 808182 41649 808187
rect 41538 808126 41588 808182
rect 41644 808126 41649 808182
rect 41538 808124 41649 808126
rect 41583 808121 41649 808124
rect 41967 807888 42033 807891
rect 41568 807886 42033 807888
rect 41568 807830 41972 807886
rect 42028 807830 42033 807886
rect 41568 807828 42033 807830
rect 41967 807825 42033 807828
rect 42831 807444 42897 807447
rect 41568 807442 42897 807444
rect 41568 807386 42836 807442
rect 42892 807386 42897 807442
rect 41568 807384 42897 807386
rect 42831 807381 42897 807384
rect 41538 806707 41598 806822
rect 41538 806702 41649 806707
rect 41538 806646 41588 806702
rect 41644 806646 41649 806702
rect 41538 806644 41649 806646
rect 41583 806641 41649 806644
rect 41538 806115 41598 806304
rect 41538 806110 41649 806115
rect 41538 806054 41588 806110
rect 41644 806054 41649 806110
rect 41538 806052 41649 806054
rect 41583 806049 41649 806052
rect 28866 805671 28926 805934
rect 28815 805666 28926 805671
rect 28815 805610 28820 805666
rect 28876 805610 28926 805666
rect 28815 805608 28926 805610
rect 28815 805605 28881 805608
rect 41538 805227 41598 805342
rect 28815 805224 28881 805227
rect 28815 805222 28926 805224
rect 28815 805166 28820 805222
rect 28876 805166 28926 805222
rect 28815 805161 28926 805166
rect 41538 805222 41649 805227
rect 41538 805166 41588 805222
rect 41644 805166 41649 805222
rect 41538 805164 41649 805166
rect 41583 805161 41649 805164
rect 28866 804824 28926 805161
rect 40239 802316 40305 802319
rect 41530 802316 41536 802318
rect 40239 802314 41536 802316
rect 40239 802258 40244 802314
rect 40300 802258 41536 802314
rect 40239 802256 41536 802258
rect 40239 802253 40305 802256
rect 41530 802254 41536 802256
rect 41600 802254 41606 802318
rect 41487 800488 41553 800491
rect 41722 800488 41728 800490
rect 41487 800486 41728 800488
rect 41487 800430 41492 800486
rect 41548 800430 41728 800486
rect 41487 800428 41728 800430
rect 41487 800425 41553 800428
rect 41722 800426 41728 800428
rect 41792 800426 41798 800490
rect 42159 800488 42225 800491
rect 42490 800488 42496 800490
rect 42159 800486 42496 800488
rect 42159 800430 42164 800486
rect 42220 800430 42496 800486
rect 42159 800428 42496 800430
rect 42159 800425 42225 800428
rect 42490 800426 42496 800428
rect 42560 800426 42566 800490
rect 42063 800340 42129 800343
rect 42298 800340 42304 800342
rect 42063 800338 42304 800340
rect 42063 800282 42068 800338
rect 42124 800282 42304 800338
rect 42063 800280 42304 800282
rect 42063 800277 42129 800280
rect 42298 800278 42304 800280
rect 42368 800278 42374 800342
rect 42298 796726 42304 796790
rect 42368 796788 42374 796790
rect 42735 796788 42801 796791
rect 42368 796786 42801 796788
rect 42368 796730 42740 796786
rect 42796 796730 42801 796786
rect 42368 796728 42801 796730
rect 42368 796726 42374 796728
rect 42735 796725 42801 796728
rect 42490 794358 42496 794422
rect 42560 794420 42566 794422
rect 42639 794420 42705 794423
rect 42560 794418 42705 794420
rect 42560 794362 42644 794418
rect 42700 794362 42705 794418
rect 42560 794360 42705 794362
rect 42560 794358 42566 794360
rect 42639 794357 42705 794360
rect 41722 792878 41728 792942
rect 41792 792940 41798 792942
rect 42639 792940 42705 792943
rect 41792 792938 42705 792940
rect 41792 792882 42644 792938
rect 42700 792882 42705 792938
rect 41792 792880 42705 792882
rect 41792 792878 41798 792880
rect 42639 792877 42705 792880
rect 41530 791842 41536 791906
rect 41600 791904 41606 791906
rect 42255 791904 42321 791907
rect 41600 791902 42321 791904
rect 41600 791846 42260 791902
rect 42316 791846 42321 791902
rect 41600 791844 42321 791846
rect 41600 791842 41606 791844
rect 42255 791841 42321 791844
rect 41338 791694 41344 791758
rect 41408 791756 41414 791758
rect 42351 791756 42417 791759
rect 41408 791754 42417 791756
rect 41408 791698 42356 791754
rect 42412 791698 42417 791754
rect 41408 791696 42417 791698
rect 41408 791694 41414 791696
rect 42351 791693 42417 791696
rect 57711 790868 57777 790871
rect 57711 790866 64638 790868
rect 57711 790810 57716 790866
rect 57772 790810 64638 790866
rect 57711 790808 64638 790810
rect 57711 790805 57777 790808
rect 64578 790304 64638 790808
rect 57615 789684 57681 789687
rect 57615 789682 64638 789684
rect 57615 789626 57620 789682
rect 57676 789626 64638 789682
rect 57615 789624 64638 789626
rect 57615 789621 57681 789624
rect 64578 789122 64638 789624
rect 58191 788500 58257 788503
rect 58191 788498 64638 788500
rect 58191 788442 58196 788498
rect 58252 788442 64638 788498
rect 58191 788440 64638 788442
rect 58191 788437 58257 788440
rect 64578 787940 64638 788440
rect 674938 788290 674944 788354
rect 675008 788352 675014 788354
rect 675087 788352 675153 788355
rect 675008 788350 675153 788352
rect 675008 788294 675092 788350
rect 675148 788294 675153 788350
rect 675008 788292 675153 788294
rect 675008 788290 675014 788292
rect 675087 788289 675153 788292
rect 58383 787316 58449 787319
rect 58383 787314 64638 787316
rect 58383 787258 58388 787314
rect 58444 787258 64638 787314
rect 58383 787256 64638 787258
rect 58383 787253 58449 787256
rect 64578 786758 64638 787256
rect 675471 787170 675537 787171
rect 675471 787166 675520 787170
rect 675584 787168 675590 787170
rect 675471 787110 675476 787166
rect 675471 787106 675520 787110
rect 675584 787108 675628 787168
rect 675584 787106 675590 787108
rect 675471 787105 675537 787106
rect 674746 786218 674752 786282
rect 674816 786280 674822 786282
rect 675087 786280 675153 786283
rect 674816 786278 675153 786280
rect 674816 786222 675092 786278
rect 675148 786222 675153 786278
rect 674816 786220 675153 786222
rect 674816 786218 674822 786220
rect 675087 786217 675153 786220
rect 59631 785540 59697 785543
rect 64578 785540 64638 785576
rect 59631 785538 64638 785540
rect 59631 785482 59636 785538
rect 59692 785482 64638 785538
rect 59631 785480 64638 785482
rect 59631 785477 59697 785480
rect 59151 784948 59217 784951
rect 59151 784946 64638 784948
rect 59151 784890 59156 784946
rect 59212 784890 64638 784946
rect 59151 784888 64638 784890
rect 59151 784885 59217 784888
rect 64578 784394 64638 784888
rect 675375 784802 675441 784803
rect 675322 784800 675328 784802
rect 675284 784740 675328 784800
rect 675392 784798 675441 784802
rect 675436 784742 675441 784798
rect 675322 784738 675328 784740
rect 675392 784738 675441 784742
rect 675375 784737 675441 784738
rect 674170 784294 674176 784358
rect 674240 784356 674246 784358
rect 675471 784356 675537 784359
rect 674240 784354 675537 784356
rect 674240 784298 675476 784354
rect 675532 784298 675537 784354
rect 674240 784296 675537 784298
rect 674240 784294 674246 784296
rect 675471 784293 675537 784296
rect 673978 783406 673984 783470
rect 674048 783468 674054 783470
rect 675087 783468 675153 783471
rect 674048 783466 675153 783468
rect 674048 783410 675092 783466
rect 675148 783410 675153 783466
rect 674048 783408 675153 783410
rect 674048 783406 674054 783408
rect 675087 783405 675153 783408
rect 675759 783024 675825 783027
rect 676666 783024 676672 783026
rect 675759 783022 676672 783024
rect 675759 782966 675764 783022
rect 675820 782966 676672 783022
rect 675759 782964 676672 782966
rect 675759 782961 675825 782964
rect 676666 782962 676672 782964
rect 676736 782962 676742 783026
rect 675759 780656 675825 780659
rect 676090 780656 676096 780658
rect 675759 780654 676096 780656
rect 675759 780598 675764 780654
rect 675820 780598 676096 780654
rect 675759 780596 676096 780598
rect 675759 780593 675825 780596
rect 676090 780594 676096 780596
rect 676160 780594 676166 780658
rect 675759 780064 675825 780067
rect 676474 780064 676480 780066
rect 675759 780062 676480 780064
rect 675759 780006 675764 780062
rect 675820 780006 676480 780062
rect 675759 780004 676480 780006
rect 675759 780001 675825 780004
rect 676474 780002 676480 780004
rect 676544 780002 676550 780066
rect 675759 778880 675825 778883
rect 676282 778880 676288 778882
rect 675759 778878 676288 778880
rect 649986 778288 650046 778824
rect 675759 778822 675764 778878
rect 675820 778822 676288 778878
rect 675759 778820 676288 778822
rect 675759 778817 675825 778820
rect 676282 778818 676288 778820
rect 676352 778818 676358 778882
rect 655407 778288 655473 778291
rect 649986 778286 655473 778288
rect 649986 778230 655412 778286
rect 655468 778230 655473 778286
rect 649986 778228 655473 778230
rect 655407 778225 655473 778228
rect 655215 777696 655281 777699
rect 649986 777694 655281 777696
rect 649986 777638 655220 777694
rect 655276 777638 655281 777694
rect 649986 777636 655281 777638
rect 655215 777633 655281 777636
rect 649986 776068 650046 776460
rect 655599 776068 655665 776071
rect 649986 776066 655665 776068
rect 649986 776010 655604 776066
rect 655660 776010 655665 776066
rect 649986 776008 655665 776010
rect 655599 776005 655665 776008
rect 655119 775920 655185 775923
rect 649986 775918 655185 775920
rect 649986 775862 655124 775918
rect 655180 775862 655185 775918
rect 649986 775860 655185 775862
rect 649986 775278 650046 775860
rect 655119 775857 655185 775860
rect 41775 774736 41841 774739
rect 656559 774736 656625 774739
rect 41568 774734 41841 774736
rect 41568 774678 41780 774734
rect 41836 774678 41841 774734
rect 41568 774676 41841 774678
rect 41775 774673 41841 774676
rect 649986 774734 656625 774736
rect 649986 774678 656564 774734
rect 656620 774678 656625 774734
rect 649986 774676 656625 774678
rect 41538 773999 41598 774114
rect 649986 774096 650046 774676
rect 656559 774673 656625 774676
rect 41538 773994 41649 773999
rect 41538 773938 41588 773994
rect 41644 773938 41649 773994
rect 41538 773936 41649 773938
rect 41583 773933 41649 773936
rect 41775 773552 41841 773555
rect 654351 773552 654417 773555
rect 41568 773550 41841 773552
rect 41568 773494 41780 773550
rect 41836 773494 41841 773550
rect 41568 773492 41841 773494
rect 41775 773489 41841 773492
rect 649986 773550 654417 773552
rect 649986 773494 654356 773550
rect 654412 773494 654417 773550
rect 649986 773492 654417 773494
rect 41583 773404 41649 773407
rect 41538 773402 41649 773404
rect 41538 773346 41588 773402
rect 41644 773346 41649 773402
rect 41538 773341 41649 773346
rect 41538 773226 41598 773341
rect 649986 772914 650046 773492
rect 654351 773489 654417 773492
rect 41775 772664 41841 772667
rect 41568 772662 41841 772664
rect 41568 772606 41780 772662
rect 41836 772606 41841 772662
rect 41568 772604 41841 772606
rect 41775 772601 41841 772604
rect 40570 772306 40576 772370
rect 40640 772368 40646 772370
rect 41583 772368 41649 772371
rect 40640 772366 41649 772368
rect 40640 772310 41588 772366
rect 41644 772310 41649 772366
rect 40640 772308 41649 772310
rect 40640 772306 40646 772308
rect 41583 772305 41649 772308
rect 40194 771926 40254 772042
rect 40186 771862 40192 771926
rect 40256 771862 40262 771926
rect 40378 771862 40384 771926
rect 40448 771924 40454 771926
rect 43119 771924 43185 771927
rect 40448 771922 43185 771924
rect 40448 771866 43124 771922
rect 43180 771866 43185 771922
rect 40448 771864 43185 771866
rect 40448 771862 40454 771864
rect 41538 771672 41598 771864
rect 43119 771861 43185 771864
rect 675279 771924 675345 771927
rect 675514 771924 675520 771926
rect 675279 771922 675520 771924
rect 675279 771866 675284 771922
rect 675340 771866 675520 771922
rect 675279 771864 675520 771866
rect 675279 771861 675345 771864
rect 675514 771862 675520 771864
rect 675584 771862 675590 771926
rect 40578 770890 40638 771154
rect 40570 770826 40576 770890
rect 40640 770826 40646 770890
rect 41583 770888 41649 770891
rect 41538 770886 41649 770888
rect 41538 770830 41588 770886
rect 41644 770830 41649 770886
rect 41538 770825 41649 770830
rect 41538 770562 41598 770825
rect 41538 770148 41598 770192
rect 42447 770148 42513 770151
rect 41538 770146 42513 770148
rect 41538 770090 42452 770146
rect 42508 770090 42513 770146
rect 41538 770088 42513 770090
rect 42447 770085 42513 770088
rect 41967 769704 42033 769707
rect 41568 769702 42033 769704
rect 41568 769646 41972 769702
rect 42028 769646 42033 769702
rect 41568 769644 42033 769646
rect 41967 769641 42033 769644
rect 38850 768967 38910 769082
rect 38799 768962 38910 768967
rect 38799 768906 38804 768962
rect 38860 768906 38910 768962
rect 38799 768904 38910 768906
rect 38799 768901 38865 768904
rect 41538 768523 41598 768638
rect 41538 768518 41649 768523
rect 41538 768462 41588 768518
rect 41644 768462 41649 768518
rect 41538 768460 41649 768462
rect 41583 768457 41649 768460
rect 41775 768224 41841 768227
rect 41568 768222 41841 768224
rect 41568 768166 41780 768222
rect 41836 768166 41841 768222
rect 41568 768164 41841 768166
rect 41775 768161 41841 768164
rect 42351 767632 42417 767635
rect 41568 767630 42417 767632
rect 41568 767574 42356 767630
rect 42412 767574 42417 767630
rect 41568 767572 42417 767574
rect 42351 767569 42417 767572
rect 33090 767043 33150 767158
rect 33039 767038 33150 767043
rect 33039 766982 33044 767038
rect 33100 766982 33150 767038
rect 33039 766980 33150 766982
rect 33039 766977 33105 766980
rect 41775 766670 41841 766673
rect 41568 766668 41841 766670
rect 41568 766612 41780 766668
rect 41836 766612 41841 766668
rect 41568 766610 41841 766612
rect 41775 766607 41841 766610
rect 41871 766152 41937 766155
rect 41568 766150 41937 766152
rect 41568 766094 41876 766150
rect 41932 766094 41937 766150
rect 41568 766092 41937 766094
rect 41871 766089 41937 766092
rect 41538 765563 41598 765678
rect 41538 765558 41649 765563
rect 41538 765502 41588 765558
rect 41644 765502 41649 765558
rect 41538 765500 41649 765502
rect 41583 765497 41649 765500
rect 41775 765190 41841 765193
rect 41568 765188 41841 765190
rect 41568 765132 41780 765188
rect 41836 765132 41841 765188
rect 41568 765130 41841 765132
rect 41775 765127 41841 765130
rect 41775 764672 41841 764675
rect 41568 764670 41841 764672
rect 41568 764614 41780 764670
rect 41836 764614 41841 764670
rect 41568 764612 41841 764614
rect 41775 764609 41841 764612
rect 42063 764228 42129 764231
rect 41568 764226 42129 764228
rect 41568 764170 42068 764226
rect 42124 764170 42129 764226
rect 41568 764168 42129 764170
rect 42063 764165 42129 764168
rect 41538 763491 41598 763606
rect 41538 763486 41649 763491
rect 41538 763430 41588 763486
rect 41644 763430 41649 763486
rect 41538 763428 41649 763430
rect 41583 763425 41649 763428
rect 41538 762899 41598 763162
rect 41538 762894 41649 762899
rect 41538 762838 41588 762894
rect 41644 762838 41649 762894
rect 41538 762836 41649 762838
rect 41583 762833 41649 762836
rect 28866 762455 28926 762718
rect 28815 762450 28926 762455
rect 28815 762394 28820 762450
rect 28876 762394 28926 762450
rect 28815 762392 28926 762394
rect 28815 762389 28881 762392
rect 41538 762011 41598 762126
rect 28815 762008 28881 762011
rect 28815 762006 28926 762008
rect 28815 761950 28820 762006
rect 28876 761950 28926 762006
rect 28815 761945 28926 761950
rect 41538 762006 41649 762011
rect 41538 761950 41588 762006
rect 41644 761950 41649 762006
rect 41538 761948 41649 761950
rect 41583 761945 41649 761948
rect 28866 761608 28926 761945
rect 33039 758900 33105 758903
rect 40762 758900 40768 758902
rect 33039 758898 40768 758900
rect 33039 758842 33044 758898
rect 33100 758842 40768 758898
rect 33039 758840 40768 758842
rect 33039 758837 33105 758840
rect 40762 758838 40768 758840
rect 40832 758838 40838 758902
rect 38799 757568 38865 757571
rect 40954 757568 40960 757570
rect 38799 757566 40960 757568
rect 38799 757510 38804 757566
rect 38860 757510 40960 757566
rect 38799 757508 40960 757510
rect 38799 757505 38865 757508
rect 40954 757506 40960 757508
rect 41024 757506 41030 757570
rect 58671 747652 58737 747655
rect 58671 747650 64638 747652
rect 58671 747594 58676 747650
rect 58732 747594 64638 747650
rect 58671 747592 64638 747594
rect 58671 747589 58737 747592
rect 64578 747082 64638 747592
rect 40762 746258 40768 746322
rect 40832 746320 40838 746322
rect 42351 746320 42417 746323
rect 40832 746318 42417 746320
rect 40832 746262 42356 746318
rect 42412 746262 42417 746318
rect 40832 746260 42417 746262
rect 40832 746258 40838 746260
rect 42351 746257 42417 746260
rect 40954 745962 40960 746026
rect 41024 746024 41030 746026
rect 42543 746024 42609 746027
rect 54735 746024 54801 746027
rect 41024 746022 42609 746024
rect 41024 745966 42548 746022
rect 42604 745966 42609 746022
rect 41024 745964 42609 745966
rect 41024 745962 41030 745964
rect 42543 745961 42609 745964
rect 54690 746022 54801 746024
rect 54690 745966 54740 746022
rect 54796 745966 54801 746022
rect 54690 745961 54801 745966
rect 54690 745879 54750 745961
rect 54639 745874 54750 745879
rect 54639 745818 54644 745874
rect 54700 745818 54750 745874
rect 54639 745816 54750 745818
rect 54639 745813 54705 745816
rect 58575 745432 58641 745435
rect 64578 745432 64638 745900
rect 58575 745430 64638 745432
rect 58575 745374 58580 745430
rect 58636 745374 64638 745430
rect 58575 745372 64638 745374
rect 58575 745369 58641 745372
rect 676282 745370 676288 745434
rect 676352 745432 676358 745434
rect 676858 745432 676864 745434
rect 676352 745372 676864 745432
rect 676352 745370 676358 745372
rect 676858 745370 676864 745372
rect 676928 745370 676934 745434
rect 57615 745284 57681 745287
rect 57615 745282 64638 745284
rect 57615 745226 57620 745282
rect 57676 745226 64638 745282
rect 57615 745224 64638 745226
rect 57615 745221 57681 745224
rect 64578 744718 64638 745224
rect 58095 744100 58161 744103
rect 58095 744098 64638 744100
rect 58095 744042 58100 744098
rect 58156 744042 64638 744098
rect 58095 744040 64638 744042
rect 58095 744037 58161 744040
rect 64578 743536 64638 744040
rect 59631 742916 59697 742919
rect 59631 742914 64638 742916
rect 59631 742858 59636 742914
rect 59692 742858 64638 742914
rect 59631 742856 64638 742858
rect 59631 742853 59697 742856
rect 64578 742354 64638 742856
rect 674362 742410 674368 742474
rect 674432 742472 674438 742474
rect 675471 742472 675537 742475
rect 674432 742470 675537 742472
rect 674432 742414 675476 742470
rect 675532 742414 675537 742470
rect 674432 742412 675537 742414
rect 674432 742410 674438 742412
rect 675471 742409 675537 742412
rect 59727 741732 59793 741735
rect 675663 741734 675729 741735
rect 59727 741730 64638 741732
rect 59727 741674 59732 741730
rect 59788 741674 64638 741730
rect 59727 741672 64638 741674
rect 59727 741669 59793 741672
rect 64578 741172 64638 741672
rect 675663 741730 675712 741734
rect 675776 741732 675782 741734
rect 675663 741674 675668 741730
rect 675663 741670 675712 741674
rect 675776 741672 675820 741732
rect 675776 741670 675782 741672
rect 675663 741669 675729 741670
rect 676474 741522 676480 741586
rect 676544 741584 676550 741586
rect 677050 741584 677056 741586
rect 676544 741524 677056 741584
rect 676544 741522 676550 741524
rect 677050 741522 677056 741524
rect 677120 741522 677126 741586
rect 675130 740042 675136 740106
rect 675200 740104 675206 740106
rect 675375 740104 675441 740107
rect 675200 740102 675441 740104
rect 675200 740046 675380 740102
rect 675436 740046 675441 740102
rect 675200 740044 675441 740046
rect 675200 740042 675206 740044
rect 675375 740041 675441 740044
rect 675759 739216 675825 739219
rect 675898 739216 675904 739218
rect 675759 739214 675904 739216
rect 675759 739158 675764 739214
rect 675820 739158 675904 739214
rect 675759 739156 675904 739158
rect 675759 739153 675825 739156
rect 675898 739154 675904 739156
rect 675968 739154 675974 739218
rect 674554 738562 674560 738626
rect 674624 738624 674630 738626
rect 675375 738624 675441 738627
rect 674624 738622 675441 738624
rect 674624 738566 675380 738622
rect 675436 738566 675441 738622
rect 674624 738564 675441 738566
rect 674624 738562 674630 738564
rect 675375 738561 675441 738564
rect 675759 735072 675825 735075
rect 676474 735072 676480 735074
rect 675759 735070 676480 735072
rect 675759 735014 675764 735070
rect 675820 735014 676480 735070
rect 675759 735012 676480 735014
rect 675759 735009 675825 735012
rect 676474 735010 676480 735012
rect 676544 735010 676550 735074
rect 655119 734480 655185 734483
rect 649986 734478 655185 734480
rect 649986 734422 655124 734478
rect 655180 734422 655185 734478
rect 649986 734420 655185 734422
rect 649986 734402 650046 734420
rect 655119 734417 655185 734420
rect 675471 734482 675537 734483
rect 675471 734478 675520 734482
rect 675584 734480 675590 734482
rect 675471 734422 675476 734478
rect 675471 734418 675520 734422
rect 675584 734420 675628 734480
rect 675584 734418 675590 734420
rect 675471 734417 675537 734418
rect 674703 734332 674769 734335
rect 676282 734332 676288 734334
rect 674703 734330 676288 734332
rect 674703 734274 674708 734330
rect 674764 734274 676288 734330
rect 674703 734272 676288 734274
rect 674703 734269 674769 734272
rect 676282 734270 676288 734272
rect 676352 734270 676358 734334
rect 649986 732704 650046 733220
rect 655503 732704 655569 732707
rect 649986 732702 655569 732704
rect 649986 732646 655508 732702
rect 655564 732646 655569 732702
rect 649986 732644 655569 732646
rect 655503 732641 655569 732644
rect 649986 731668 650046 732038
rect 655311 731668 655377 731671
rect 649986 731666 655377 731668
rect 649986 731610 655316 731666
rect 655372 731610 655377 731666
rect 649986 731608 655377 731610
rect 655311 731605 655377 731608
rect 41775 731520 41841 731523
rect 41568 731518 41841 731520
rect 41568 731462 41780 731518
rect 41836 731462 41841 731518
rect 41568 731460 41841 731462
rect 41775 731457 41841 731460
rect 655695 731372 655761 731375
rect 649986 731370 655761 731372
rect 649986 731314 655700 731370
rect 655756 731314 655761 731370
rect 649986 731312 655761 731314
rect 41538 730783 41598 730898
rect 649986 730856 650046 731312
rect 655695 731309 655761 731312
rect 41538 730778 41649 730783
rect 41538 730722 41588 730778
rect 41644 730722 41649 730778
rect 41538 730720 41649 730722
rect 41583 730717 41649 730720
rect 41775 730410 41841 730413
rect 41568 730408 41841 730410
rect 41568 730352 41780 730408
rect 41836 730352 41841 730408
rect 41568 730350 41841 730352
rect 41775 730347 41841 730350
rect 41583 730188 41649 730191
rect 654159 730188 654225 730191
rect 41538 730186 41649 730188
rect 41538 730130 41588 730186
rect 41644 730130 41649 730186
rect 41538 730125 41649 730130
rect 649986 730186 654225 730188
rect 649986 730130 654164 730186
rect 654220 730130 654225 730186
rect 649986 730128 654225 730130
rect 41538 730010 41598 730125
rect 649986 729674 650046 730128
rect 654159 730125 654225 730128
rect 41775 729448 41841 729451
rect 41568 729446 41841 729448
rect 41568 729390 41780 729446
rect 41836 729390 41841 729446
rect 41568 729388 41841 729390
rect 41775 729385 41841 729388
rect 40570 729238 40576 729302
rect 40640 729300 40646 729302
rect 42255 729300 42321 729303
rect 40640 729298 42321 729300
rect 40640 729242 42260 729298
rect 42316 729242 42321 729298
rect 40640 729240 42321 729242
rect 40640 729238 40646 729240
rect 42255 729237 42321 729240
rect 41775 728856 41841 728859
rect 41568 728854 41841 728856
rect 41568 728798 41780 728854
rect 41836 728798 41841 728854
rect 41568 728796 41841 728798
rect 41775 728793 41841 728796
rect 40431 728710 40497 728711
rect 40378 728646 40384 728710
rect 40448 728708 40497 728710
rect 40448 728706 40576 728708
rect 40492 728650 40576 728706
rect 40448 728648 40576 728650
rect 40448 728646 40497 728648
rect 40386 728645 40497 728646
rect 40386 728530 40446 728645
rect 654063 728560 654129 728563
rect 649986 728558 654129 728560
rect 649986 728502 654068 728558
rect 654124 728502 654129 728558
rect 649986 728500 654129 728502
rect 649986 728492 650046 728500
rect 654063 728497 654129 728500
rect 676858 728054 676864 728118
rect 676928 728116 676934 728118
rect 677434 728116 677440 728118
rect 676928 728056 677440 728116
rect 676928 728054 676934 728056
rect 677434 728054 677440 728056
rect 677504 728054 677510 728118
rect 41775 727968 41841 727971
rect 41568 727966 41841 727968
rect 41568 727910 41780 727966
rect 41836 727910 41841 727966
rect 41568 727908 41841 727910
rect 41775 727905 41841 727908
rect 40570 727610 40576 727674
rect 40640 727610 40646 727674
rect 40578 727346 40638 727610
rect 41775 727006 41841 727009
rect 41568 727004 41841 727006
rect 41568 726948 41780 727004
rect 41836 726948 41841 727004
rect 41568 726946 41841 726948
rect 41775 726943 41841 726946
rect 41775 726488 41841 726491
rect 41568 726486 41841 726488
rect 41568 726430 41780 726486
rect 41836 726430 41841 726486
rect 41568 726428 41841 726430
rect 41775 726425 41841 726428
rect 40194 725751 40254 725866
rect 40194 725746 40305 725751
rect 40194 725690 40244 725746
rect 40300 725690 40305 725746
rect 40194 725688 40305 725690
rect 40239 725685 40305 725688
rect 41538 725304 41598 725496
rect 41679 725304 41745 725307
rect 41538 725302 41745 725304
rect 41538 725246 41684 725302
rect 41740 725246 41745 725302
rect 41538 725244 41745 725246
rect 41679 725241 41745 725244
rect 41967 725008 42033 725011
rect 41568 725006 42033 725008
rect 41568 724950 41972 725006
rect 42028 724950 42033 725006
rect 41568 724948 42033 724950
rect 41967 724945 42033 724948
rect 42255 724416 42321 724419
rect 41568 724414 42321 724416
rect 41568 724358 42260 724414
rect 42316 724358 42321 724414
rect 41568 724356 42321 724358
rect 42255 724353 42321 724356
rect 34434 723827 34494 723942
rect 34434 723822 34545 723827
rect 34434 723766 34484 723822
rect 34540 723766 34545 723822
rect 34434 723764 34545 723766
rect 34479 723761 34545 723764
rect 41775 723528 41841 723531
rect 41568 723526 41841 723528
rect 41568 723470 41780 723526
rect 41836 723470 41841 723526
rect 41568 723468 41841 723470
rect 41775 723465 41841 723468
rect 42447 722936 42513 722939
rect 41568 722934 42513 722936
rect 41568 722878 42452 722934
rect 42508 722878 42513 722934
rect 41568 722876 42513 722878
rect 42447 722873 42513 722876
rect 41538 722347 41598 722462
rect 41538 722342 41649 722347
rect 41538 722286 41588 722342
rect 41644 722286 41649 722342
rect 41538 722284 41649 722286
rect 41583 722281 41649 722284
rect 41775 721974 41841 721977
rect 41568 721972 41841 721974
rect 41568 721916 41780 721972
rect 41836 721916 41841 721972
rect 41568 721914 41841 721916
rect 41775 721911 41841 721914
rect 41871 721456 41937 721459
rect 41568 721454 41937 721456
rect 41568 721398 41876 721454
rect 41932 721398 41937 721454
rect 41568 721396 41937 721398
rect 41871 721393 41937 721396
rect 41538 720867 41598 720982
rect 41538 720862 41649 720867
rect 41538 720806 41588 720862
rect 41644 720806 41649 720862
rect 41538 720804 41649 720806
rect 41583 720801 41649 720804
rect 41775 720494 41841 720497
rect 41568 720492 41841 720494
rect 41568 720436 41780 720492
rect 41836 720436 41841 720492
rect 41568 720434 41841 720436
rect 41775 720431 41841 720434
rect 41538 719680 41598 719946
rect 41538 719620 41790 719680
rect 28866 719239 28926 719502
rect 28815 719234 28926 719239
rect 41730 719236 41790 719620
rect 28815 719178 28820 719234
rect 28876 719178 28926 719234
rect 28815 719176 28926 719178
rect 41538 719176 41790 719236
rect 28815 719173 28881 719176
rect 41538 718795 41598 719176
rect 28815 718792 28881 718795
rect 28815 718790 28926 718792
rect 28815 718734 28820 718790
rect 28876 718734 28926 718790
rect 28815 718729 28926 718734
rect 41538 718790 41649 718795
rect 41538 718734 41588 718790
rect 41644 718734 41649 718790
rect 41538 718732 41649 718734
rect 41583 718729 41649 718732
rect 28866 718466 28926 718729
rect 40239 717366 40305 717369
rect 40570 717366 40576 717368
rect 40239 717364 40576 717366
rect 40239 717308 40244 717364
rect 40300 717308 40576 717364
rect 40239 717306 40576 717308
rect 40239 717303 40305 717306
rect 40570 717304 40576 717306
rect 40640 717304 40646 717368
rect 34479 715832 34545 715835
rect 40378 715832 40384 715834
rect 34479 715830 40384 715832
rect 34479 715774 34484 715830
rect 34540 715774 40384 715830
rect 34479 715772 40384 715774
rect 34479 715769 34545 715772
rect 40378 715770 40384 715772
rect 40448 715770 40454 715834
rect 676290 715539 676350 715654
rect 676290 715534 676401 715539
rect 676290 715478 676340 715534
rect 676396 715478 676401 715534
rect 676290 715476 676401 715478
rect 676335 715473 676401 715476
rect 676143 714944 676209 714947
rect 676290 714944 676350 715136
rect 676143 714942 676350 714944
rect 676143 714886 676148 714942
rect 676204 714886 676350 714942
rect 676143 714884 676350 714886
rect 676143 714881 676209 714884
rect 676239 714796 676305 714799
rect 676239 714794 676350 714796
rect 676239 714738 676244 714794
rect 676300 714738 676350 714794
rect 676239 714733 676350 714738
rect 676290 714618 676350 714733
rect 679746 713911 679806 714174
rect 679695 713906 679806 713911
rect 679695 713850 679700 713906
rect 679756 713850 679806 713906
rect 679695 713848 679806 713850
rect 679695 713845 679761 713848
rect 679746 713319 679806 713582
rect 679695 713314 679806 713319
rect 679695 713258 679700 713314
rect 679756 713258 679806 713314
rect 679695 713256 679806 713258
rect 679695 713253 679761 713256
rect 676047 713168 676113 713171
rect 676047 713166 676320 713168
rect 676047 713110 676052 713166
rect 676108 713110 676320 713166
rect 676047 713108 676320 713110
rect 676047 713105 676113 713108
rect 676047 712724 676113 712727
rect 676047 712722 676320 712724
rect 676047 712666 676052 712722
rect 676108 712666 676320 712722
rect 676047 712664 676320 712666
rect 676047 712661 676113 712664
rect 676290 711987 676350 712102
rect 676239 711982 676350 711987
rect 676239 711926 676244 711982
rect 676300 711926 676350 711982
rect 676239 711924 676350 711926
rect 676239 711921 676305 711924
rect 42447 711688 42513 711691
rect 42682 711688 42688 711690
rect 42447 711686 42688 711688
rect 42447 711630 42452 711686
rect 42508 711630 42688 711686
rect 42447 711628 42688 711630
rect 42447 711625 42513 711628
rect 42682 711626 42688 711628
rect 42752 711626 42758 711690
rect 676047 711614 676113 711617
rect 676047 711612 676320 711614
rect 676047 711556 676052 711612
rect 676108 711556 676320 711612
rect 676047 711554 676320 711556
rect 676047 711551 676113 711554
rect 42831 711390 42897 711393
rect 42498 711388 42897 711390
rect 42498 711332 42836 711388
rect 42892 711332 42897 711388
rect 42498 711330 42897 711332
rect 42351 711096 42417 711099
rect 42498 711096 42558 711330
rect 42831 711327 42897 711330
rect 42682 711182 42688 711246
rect 42752 711244 42758 711246
rect 42927 711244 42993 711247
rect 42752 711242 42993 711244
rect 42752 711186 42932 711242
rect 42988 711186 42993 711242
rect 42752 711184 42993 711186
rect 42752 711182 42758 711184
rect 42927 711181 42993 711184
rect 674746 711182 674752 711246
rect 674816 711244 674822 711246
rect 674816 711184 676320 711244
rect 674816 711182 674822 711184
rect 42351 711094 42558 711096
rect 42351 711038 42356 711094
rect 42412 711038 42558 711094
rect 42351 711036 42558 711038
rect 42351 711033 42417 711036
rect 676047 710652 676113 710655
rect 676047 710650 676320 710652
rect 676047 710594 676052 710650
rect 676108 710594 676320 710650
rect 676047 710592 676320 710594
rect 676047 710589 676113 710592
rect 674938 710442 674944 710506
rect 675008 710504 675014 710506
rect 675008 710444 676350 710504
rect 675008 710442 675014 710444
rect 676290 710104 676350 710444
rect 675322 709702 675328 709766
rect 675392 709764 675398 709766
rect 675392 709704 676320 709764
rect 675392 709702 675398 709704
rect 676090 709406 676096 709470
rect 676160 709468 676166 709470
rect 676160 709408 676350 709468
rect 676160 709406 676166 709408
rect 676290 709142 676350 709408
rect 676047 708580 676113 708583
rect 676047 708578 676320 708580
rect 676047 708522 676052 708578
rect 676108 708522 676320 708578
rect 676047 708520 676320 708522
rect 676047 708517 676113 708520
rect 676047 708210 676113 708213
rect 676047 708208 676320 708210
rect 676047 708152 676052 708208
rect 676108 708152 676320 708208
rect 676047 708150 676320 708152
rect 676047 708147 676113 708150
rect 674170 707630 674176 707694
rect 674240 707692 674246 707694
rect 674240 707632 676320 707692
rect 674240 707630 674246 707632
rect 673978 707038 673984 707102
rect 674048 707100 674054 707102
rect 674048 707040 676320 707100
rect 674048 707038 674054 707040
rect 676047 706730 676113 706733
rect 676047 706728 676320 706730
rect 676047 706672 676052 706728
rect 676108 706672 676320 706728
rect 676047 706670 676320 706672
rect 676047 706667 676113 706670
rect 676239 706360 676305 706363
rect 676239 706358 676350 706360
rect 676239 706302 676244 706358
rect 676300 706302 676350 706358
rect 676239 706297 676350 706302
rect 676290 706182 676350 706297
rect 677434 705854 677440 705918
rect 677504 705854 677510 705918
rect 677442 705590 677502 705854
rect 677242 705410 677248 705474
rect 677312 705410 677318 705474
rect 677250 705146 677310 705410
rect 677050 704966 677056 705030
rect 677120 704966 677126 705030
rect 677058 704702 677118 704966
rect 59631 704436 59697 704439
rect 679983 704436 680049 704439
rect 59631 704434 64638 704436
rect 59631 704378 59636 704434
rect 59692 704378 64638 704434
rect 59631 704376 64638 704378
rect 59631 704373 59697 704376
rect 64578 703860 64638 704376
rect 679938 704434 680049 704436
rect 679938 704378 679988 704434
rect 680044 704378 680049 704434
rect 679938 704373 680049 704378
rect 679938 704110 679998 704373
rect 679746 703403 679806 703666
rect 679746 703398 679857 703403
rect 679983 703400 680049 703403
rect 679746 703342 679796 703398
rect 679852 703342 679857 703398
rect 679746 703340 679857 703342
rect 679791 703337 679857 703340
rect 679938 703398 680049 703400
rect 679938 703342 679988 703398
rect 680044 703342 680049 703398
rect 679938 703337 680049 703342
rect 679938 703148 679998 703337
rect 40570 702894 40576 702958
rect 40640 702956 40646 702958
rect 42351 702956 42417 702959
rect 679791 702956 679857 702959
rect 40640 702954 42417 702956
rect 40640 702898 42356 702954
rect 42412 702898 42417 702954
rect 40640 702896 42417 702898
rect 40640 702894 40646 702896
rect 42351 702893 42417 702896
rect 679746 702954 679857 702956
rect 679746 702898 679796 702954
rect 679852 702898 679857 702954
rect 679746 702893 679857 702898
rect 40378 702746 40384 702810
rect 40448 702808 40454 702810
rect 42543 702808 42609 702811
rect 40448 702806 42609 702808
rect 40448 702750 42548 702806
rect 42604 702750 42609 702806
rect 40448 702748 42609 702750
rect 40448 702746 40454 702748
rect 42543 702745 42609 702748
rect 58767 702660 58833 702663
rect 64578 702660 64638 702678
rect 58767 702658 64638 702660
rect 58767 702602 58772 702658
rect 58828 702602 64638 702658
rect 679746 702630 679806 702893
rect 58767 702600 64638 702602
rect 58767 702597 58833 702600
rect 58863 702068 58929 702071
rect 58863 702066 64638 702068
rect 58863 702010 58868 702066
rect 58924 702010 64638 702066
rect 58863 702008 64638 702010
rect 58863 702005 58929 702008
rect 64578 701496 64638 702008
rect 58671 700884 58737 700887
rect 58671 700882 64638 700884
rect 58671 700826 58676 700882
rect 58732 700826 64638 700882
rect 58671 700824 64638 700826
rect 58671 700821 58737 700824
rect 64578 700314 64638 700824
rect 59247 699700 59313 699703
rect 59247 699698 64638 699700
rect 59247 699642 59252 699698
rect 59308 699642 64638 699698
rect 59247 699640 64638 699642
rect 59247 699637 59313 699640
rect 64578 699132 64638 699640
rect 58863 698516 58929 698519
rect 58863 698514 64638 698516
rect 58863 698458 58868 698514
rect 58924 698458 64638 698514
rect 58863 698456 64638 698458
rect 58863 698453 58929 698456
rect 64578 697950 64638 698456
rect 675375 697926 675441 697927
rect 675322 697924 675328 697926
rect 675284 697864 675328 697924
rect 675392 697922 675441 697926
rect 675436 697866 675441 697922
rect 675322 697862 675328 697864
rect 675392 697862 675441 697866
rect 675375 697861 675441 697862
rect 674170 697122 674176 697186
rect 674240 697184 674246 697186
rect 675087 697184 675153 697187
rect 674240 697182 675153 697184
rect 674240 697126 675092 697182
rect 675148 697126 675153 697182
rect 674240 697124 675153 697126
rect 674240 697122 674246 697124
rect 675087 697121 675153 697124
rect 674746 696974 674752 697038
rect 674816 697036 674822 697038
rect 675087 697036 675153 697039
rect 674816 697034 675153 697036
rect 674816 696978 675092 697034
rect 675148 696978 675153 697034
rect 674816 696976 675153 696978
rect 674816 696974 674822 696976
rect 675087 696973 675153 696976
rect 675759 694964 675825 694967
rect 676282 694964 676288 694966
rect 675759 694962 676288 694964
rect 675759 694906 675764 694962
rect 675820 694906 676288 694962
rect 675759 694904 676288 694906
rect 675759 694901 675825 694904
rect 676282 694902 676288 694904
rect 676352 694902 676358 694966
rect 674938 694606 674944 694670
rect 675008 694668 675014 694670
rect 675087 694668 675153 694671
rect 675008 694666 675153 694668
rect 675008 694610 675092 694666
rect 675148 694610 675153 694666
rect 675008 694608 675153 694610
rect 675008 694606 675014 694608
rect 675087 694605 675153 694608
rect 673978 693422 673984 693486
rect 674048 693484 674054 693486
rect 675471 693484 675537 693487
rect 674048 693482 675537 693484
rect 674048 693426 675476 693482
rect 675532 693426 675537 693482
rect 674048 693424 675537 693426
rect 674048 693422 674054 693424
rect 675471 693421 675537 693424
rect 649986 689488 650046 689980
rect 655215 689488 655281 689491
rect 649986 689486 655281 689488
rect 649986 689430 655220 689486
rect 655276 689430 655281 689486
rect 649986 689428 655281 689430
rect 655215 689425 655281 689428
rect 649986 688452 650046 688798
rect 655599 688452 655665 688455
rect 649986 688450 655665 688452
rect 649986 688394 655604 688450
rect 655660 688394 655665 688450
rect 649986 688392 655665 688394
rect 655599 688389 655665 688392
rect 41775 688304 41841 688307
rect 41568 688302 41841 688304
rect 41568 688246 41780 688302
rect 41836 688246 41841 688302
rect 41568 688244 41841 688246
rect 41775 688241 41841 688244
rect 41538 687567 41598 687682
rect 41538 687562 41649 687567
rect 41538 687506 41588 687562
rect 41644 687506 41649 687562
rect 41538 687504 41649 687506
rect 41583 687501 41649 687504
rect 41775 687268 41841 687271
rect 41568 687266 41841 687268
rect 41568 687210 41780 687266
rect 41836 687210 41841 687266
rect 41568 687208 41841 687210
rect 41775 687205 41841 687208
rect 649986 687120 650046 687616
rect 655407 687120 655473 687123
rect 649986 687118 655473 687120
rect 649986 687062 655412 687118
rect 655468 687062 655473 687118
rect 649986 687060 655473 687062
rect 655407 687057 655473 687060
rect 41583 686972 41649 686975
rect 654735 686972 654801 686975
rect 41538 686970 41649 686972
rect 41538 686914 41588 686970
rect 41644 686914 41649 686970
rect 41538 686909 41649 686914
rect 649986 686970 654801 686972
rect 649986 686914 654740 686970
rect 654796 686914 654801 686970
rect 649986 686912 654801 686914
rect 41538 686794 41598 686909
rect 649986 686434 650046 686912
rect 654735 686909 654801 686912
rect 675183 686824 675249 686827
rect 677050 686824 677056 686826
rect 675183 686822 677056 686824
rect 675183 686766 675188 686822
rect 675244 686766 677056 686822
rect 675183 686764 677056 686766
rect 675183 686761 675249 686764
rect 677050 686762 677056 686764
rect 677120 686762 677126 686826
rect 41538 686087 41598 686202
rect 41538 686082 41649 686087
rect 41538 686026 41588 686082
rect 41644 686026 41649 686082
rect 41538 686024 41649 686026
rect 41583 686021 41649 686024
rect 40386 685494 40446 685684
rect 40378 685430 40384 685494
rect 40448 685430 40454 685494
rect 41775 685344 41841 685347
rect 654159 685344 654225 685347
rect 41568 685342 41841 685344
rect 41568 685286 41780 685342
rect 41836 685286 41841 685342
rect 41568 685284 41841 685286
rect 41775 685281 41841 685284
rect 649986 685342 654225 685344
rect 649986 685286 654164 685342
rect 654220 685286 654225 685342
rect 649986 685284 654225 685286
rect 649986 685252 650046 685284
rect 654159 685281 654225 685284
rect 40578 684458 40638 684722
rect 654063 684604 654129 684607
rect 649986 684602 654129 684604
rect 649986 684546 654068 684602
rect 654124 684546 654129 684602
rect 649986 684544 654129 684546
rect 40570 684394 40576 684458
rect 40640 684394 40646 684458
rect 41775 684160 41841 684163
rect 41568 684158 41841 684160
rect 41568 684102 41780 684158
rect 41836 684102 41841 684158
rect 41568 684100 41841 684102
rect 41775 684097 41841 684100
rect 649986 684070 650046 684544
rect 654063 684541 654129 684544
rect 42063 683864 42129 683867
rect 41568 683862 42129 683864
rect 41568 683806 42068 683862
rect 42124 683806 42129 683862
rect 41568 683804 42129 683806
rect 42063 683801 42129 683804
rect 42543 683272 42609 683275
rect 41568 683270 42609 683272
rect 41568 683214 42548 683270
rect 42604 683214 42609 683270
rect 41568 683212 42609 683214
rect 42543 683209 42609 683212
rect 39810 682535 39870 682650
rect 39810 682530 39921 682535
rect 39810 682474 39860 682530
rect 39916 682474 39921 682530
rect 39810 682472 39921 682474
rect 39855 682469 39921 682472
rect 41538 682236 41598 682280
rect 42159 682236 42225 682239
rect 41538 682234 42225 682236
rect 41538 682178 42164 682234
rect 42220 682178 42225 682234
rect 41538 682176 42225 682178
rect 42159 682173 42225 682176
rect 41775 681792 41841 681795
rect 41568 681790 41841 681792
rect 41568 681734 41780 681790
rect 41836 681734 41841 681790
rect 41568 681732 41841 681734
rect 41775 681729 41841 681732
rect 42351 681200 42417 681203
rect 41568 681198 42417 681200
rect 41568 681142 42356 681198
rect 42412 681142 42417 681198
rect 41568 681140 42417 681142
rect 42351 681137 42417 681140
rect 34434 680611 34494 680800
rect 34434 680606 34545 680611
rect 34434 680550 34484 680606
rect 34540 680550 34545 680606
rect 34434 680548 34545 680550
rect 34479 680545 34545 680548
rect 41775 680312 41841 680315
rect 41568 680310 41841 680312
rect 41568 680254 41780 680310
rect 41836 680254 41841 680310
rect 41568 680252 41841 680254
rect 41775 680249 41841 680252
rect 41775 679720 41841 679723
rect 41568 679718 41841 679720
rect 41568 679662 41780 679718
rect 41836 679662 41841 679718
rect 41568 679660 41841 679662
rect 41775 679657 41841 679660
rect 41538 679131 41598 679246
rect 41538 679126 41649 679131
rect 41538 679070 41588 679126
rect 41644 679070 41649 679126
rect 41538 679068 41649 679070
rect 41583 679065 41649 679068
rect 41775 678832 41841 678835
rect 41568 678830 41841 678832
rect 41568 678774 41780 678830
rect 41836 678774 41841 678830
rect 41568 678772 41841 678774
rect 41775 678769 41841 678772
rect 41967 678240 42033 678243
rect 41568 678238 42033 678240
rect 41568 678182 41972 678238
rect 42028 678182 42033 678238
rect 41568 678180 42033 678182
rect 41967 678177 42033 678180
rect 41775 677796 41841 677799
rect 41568 677794 41841 677796
rect 41568 677738 41780 677794
rect 41836 677738 41841 677794
rect 41568 677736 41841 677738
rect 41775 677733 41841 677736
rect 41775 677278 41841 677281
rect 41568 677276 41841 677278
rect 41568 677220 41780 677276
rect 41836 677220 41841 677276
rect 41568 677218 41841 677220
rect 41775 677215 41841 677218
rect 41775 676760 41841 676763
rect 41568 676758 41841 676760
rect 41568 676702 41780 676758
rect 41836 676702 41841 676758
rect 41568 676700 41841 676702
rect 41775 676697 41841 676700
rect 28866 676023 28926 676286
rect 28815 676018 28926 676023
rect 28815 675962 28820 676018
rect 28876 675962 28926 676018
rect 28815 675960 28926 675962
rect 28815 675957 28881 675960
rect 41775 675798 41841 675801
rect 41568 675796 41841 675798
rect 41568 675740 41780 675796
rect 41836 675740 41841 675796
rect 41568 675738 41841 675740
rect 41775 675735 41841 675738
rect 28815 675576 28881 675579
rect 28815 675574 28926 675576
rect 28815 675518 28820 675574
rect 28876 675518 28926 675574
rect 28815 675513 28926 675518
rect 28866 675250 28926 675513
rect 34479 672918 34545 672921
rect 40762 672918 40768 672920
rect 34479 672916 40768 672918
rect 34479 672860 34484 672916
rect 34540 672860 40768 672916
rect 34479 672858 40768 672860
rect 34479 672855 34545 672858
rect 40762 672856 40768 672858
rect 40832 672856 40838 672920
rect 42447 671286 42513 671287
rect 42447 671282 42496 671286
rect 42560 671284 42566 671286
rect 42447 671226 42452 671282
rect 42447 671222 42496 671226
rect 42560 671224 42604 671284
rect 42560 671222 42566 671224
rect 42447 671221 42513 671222
rect 39855 671136 39921 671139
rect 42298 671136 42304 671138
rect 39855 671134 42304 671136
rect 39855 671078 39860 671134
rect 39916 671078 42304 671134
rect 39855 671076 42304 671078
rect 39855 671073 39921 671076
rect 42298 671074 42304 671076
rect 42368 671074 42374 671138
rect 41967 670692 42033 670695
rect 42106 670692 42112 670694
rect 41967 670690 42112 670692
rect 41967 670634 41972 670690
rect 42028 670634 42112 670690
rect 41967 670632 42112 670634
rect 41967 670629 42033 670632
rect 42106 670630 42112 670632
rect 42176 670630 42182 670694
rect 676143 670396 676209 670399
rect 676290 670396 676350 670662
rect 676143 670394 676350 670396
rect 676143 670338 676148 670394
rect 676204 670338 676350 670394
rect 676143 670336 676350 670338
rect 676143 670333 676209 670336
rect 676290 669807 676350 670070
rect 676290 669802 676401 669807
rect 676290 669746 676340 669802
rect 676396 669746 676401 669802
rect 676290 669744 676401 669746
rect 676335 669741 676401 669744
rect 676290 669363 676350 669626
rect 676239 669358 676350 669363
rect 676239 669302 676244 669358
rect 676300 669302 676350 669358
rect 676239 669300 676350 669302
rect 676239 669297 676305 669300
rect 676047 669212 676113 669215
rect 676047 669210 676320 669212
rect 676047 669154 676052 669210
rect 676108 669154 676320 669210
rect 676047 669152 676320 669154
rect 676047 669149 676113 669152
rect 676047 668620 676113 668623
rect 676047 668618 676320 668620
rect 676047 668562 676052 668618
rect 676108 668562 676320 668618
rect 676047 668560 676320 668562
rect 676047 668557 676113 668560
rect 42106 668410 42112 668474
rect 42176 668472 42182 668474
rect 42543 668472 42609 668475
rect 42176 668470 42609 668472
rect 42176 668414 42548 668470
rect 42604 668414 42609 668470
rect 42176 668412 42609 668414
rect 42176 668410 42182 668412
rect 42543 668409 42609 668412
rect 675951 668102 676017 668105
rect 675951 668100 676320 668102
rect 675951 668044 675956 668100
rect 676012 668044 676320 668100
rect 675951 668042 676320 668044
rect 675951 668039 676017 668042
rect 42447 667734 42513 667735
rect 42447 667732 42496 667734
rect 42404 667730 42496 667732
rect 42404 667674 42452 667730
rect 42404 667672 42496 667674
rect 42447 667670 42496 667672
rect 42560 667670 42566 667734
rect 675951 667732 676017 667735
rect 675951 667730 676320 667732
rect 675951 667674 675956 667730
rect 676012 667674 676320 667730
rect 675951 667672 676320 667674
rect 42447 667669 42513 667670
rect 675951 667669 676017 667672
rect 676290 666995 676350 667110
rect 676239 666990 676350 666995
rect 676239 666934 676244 666990
rect 676300 666934 676350 666990
rect 676239 666932 676350 666934
rect 676239 666929 676305 666932
rect 676290 666403 676350 666592
rect 676239 666398 676350 666403
rect 676239 666342 676244 666398
rect 676300 666342 676350 666398
rect 676239 666340 676350 666342
rect 676239 666337 676305 666340
rect 675706 666190 675712 666254
rect 675776 666252 675782 666254
rect 675776 666192 676320 666252
rect 675776 666190 675782 666192
rect 676047 665660 676113 665663
rect 676047 665658 676320 665660
rect 676047 665602 676052 665658
rect 676108 665602 676320 665658
rect 676047 665600 676320 665602
rect 676047 665597 676113 665600
rect 676474 665302 676480 665366
rect 676544 665302 676550 665366
rect 676482 665038 676542 665302
rect 675130 664710 675136 664774
rect 675200 664772 675206 664774
rect 675200 664712 676320 664772
rect 675200 664710 675206 664712
rect 676239 664328 676305 664331
rect 676239 664326 676350 664328
rect 676239 664270 676244 664326
rect 676300 664270 676350 664326
rect 676239 664265 676350 664270
rect 676290 664150 676350 664265
rect 676047 663588 676113 663591
rect 676047 663586 676320 663588
rect 676047 663530 676052 663586
rect 676108 663530 676320 663586
rect 676047 663528 676320 663530
rect 676047 663525 676113 663528
rect 674362 663378 674368 663442
rect 674432 663440 674438 663442
rect 674432 663380 676350 663440
rect 674432 663378 674438 663380
rect 676290 663188 676350 663380
rect 675898 662638 675904 662702
rect 675968 662700 675974 662702
rect 675968 662640 676320 662700
rect 675968 662638 675974 662640
rect 674554 662046 674560 662110
rect 674624 662108 674630 662110
rect 674624 662048 676320 662108
rect 674624 662046 674630 662048
rect 676047 661664 676113 661667
rect 676047 661662 676320 661664
rect 676047 661606 676052 661662
rect 676108 661606 676320 661662
rect 676047 661604 676320 661606
rect 676047 661601 676113 661604
rect 59631 661220 59697 661223
rect 59631 661218 64638 661220
rect 59631 661162 59636 661218
rect 59692 661162 64638 661218
rect 59631 661160 64638 661162
rect 59631 661157 59697 661160
rect 40762 660862 40768 660926
rect 40832 660924 40838 660926
rect 42543 660924 42609 660927
rect 40832 660922 42609 660924
rect 40832 660866 42548 660922
rect 42604 660866 42609 660922
rect 40832 660864 42609 660866
rect 40832 660862 40838 660864
rect 42543 660861 42609 660864
rect 64578 660638 64638 661160
rect 675514 661158 675520 661222
rect 675584 661220 675590 661222
rect 675584 661160 676320 661220
rect 675584 661158 675590 661160
rect 676047 660628 676113 660631
rect 676047 660626 676320 660628
rect 676047 660570 676052 660626
rect 676108 660570 676320 660626
rect 676047 660568 676320 660570
rect 676047 660565 676113 660568
rect 676858 660418 676864 660482
rect 676928 660418 676934 660482
rect 676866 660154 676926 660418
rect 676239 659888 676305 659891
rect 676239 659886 676350 659888
rect 676239 659830 676244 659886
rect 676300 659830 676350 659886
rect 676239 659825 676350 659830
rect 676290 659710 676350 659825
rect 42298 659530 42304 659594
rect 42368 659530 42374 659594
rect 42306 659447 42366 659530
rect 42306 659442 42417 659447
rect 42306 659386 42356 659442
rect 42412 659386 42417 659442
rect 42306 659384 42417 659386
rect 42351 659381 42417 659384
rect 58767 659444 58833 659447
rect 64578 659444 64638 659456
rect 58767 659442 64638 659444
rect 58767 659386 58772 659442
rect 58828 659386 64638 659442
rect 58767 659384 64638 659386
rect 58767 659381 58833 659384
rect 679791 659296 679857 659299
rect 679746 659294 679857 659296
rect 679746 659238 679796 659294
rect 679852 659238 679857 659294
rect 679746 659233 679857 659238
rect 679746 659118 679806 659233
rect 57711 658852 57777 658855
rect 57711 658850 64638 658852
rect 57711 658794 57716 658850
rect 57772 658794 64638 658850
rect 57711 658792 64638 658794
rect 57711 658789 57777 658792
rect 64578 658274 64638 658792
rect 685506 658411 685566 658674
rect 679791 658408 679857 658411
rect 679746 658406 679857 658408
rect 679746 658350 679796 658406
rect 679852 658350 679857 658406
rect 679746 658345 679857 658350
rect 685455 658406 685566 658411
rect 685455 658350 685460 658406
rect 685516 658350 685566 658406
rect 685455 658348 685566 658350
rect 685455 658345 685521 658348
rect 679746 658156 679806 658345
rect 685455 657964 685521 657967
rect 685455 657962 685566 657964
rect 685455 657906 685460 657962
rect 685516 657906 685566 657962
rect 685455 657901 685566 657906
rect 59151 657668 59217 657671
rect 59151 657666 64638 657668
rect 59151 657610 59156 657666
rect 59212 657610 64638 657666
rect 685506 657638 685566 657901
rect 59151 657608 64638 657610
rect 59151 657605 59217 657608
rect 64578 657092 64638 657608
rect 58191 656484 58257 656487
rect 58191 656482 64638 656484
rect 58191 656426 58196 656482
rect 58252 656426 64638 656482
rect 58191 656424 64638 656426
rect 58191 656421 58257 656424
rect 64578 655910 64638 656424
rect 58383 655300 58449 655303
rect 58383 655298 64638 655300
rect 58383 655242 58388 655298
rect 58444 655242 64638 655298
rect 58383 655240 64638 655242
rect 58383 655237 58449 655240
rect 64578 654728 64638 655240
rect 674362 652130 674368 652194
rect 674432 652192 674438 652194
rect 675471 652192 675537 652195
rect 674432 652190 675537 652192
rect 674432 652134 675476 652190
rect 675532 652134 675537 652190
rect 674432 652132 675537 652134
rect 674432 652130 674438 652132
rect 675471 652129 675537 652132
rect 675471 651454 675537 651455
rect 675471 651450 675520 651454
rect 675584 651452 675590 651454
rect 675471 651394 675476 651450
rect 675471 651390 675520 651394
rect 675584 651392 675628 651452
rect 675584 651390 675590 651392
rect 675471 651389 675537 651390
rect 674554 650946 674560 651010
rect 674624 651008 674630 651010
rect 675087 651008 675153 651011
rect 674624 651006 675153 651008
rect 674624 650950 675092 651006
rect 675148 650950 675153 651006
rect 674624 650948 675153 650950
rect 674624 650946 674630 650948
rect 675087 650945 675153 650948
rect 675663 649826 675729 649827
rect 675663 649822 675712 649826
rect 675776 649824 675782 649826
rect 675663 649766 675668 649822
rect 675663 649762 675712 649766
rect 675776 649764 675820 649824
rect 675776 649762 675782 649764
rect 675663 649761 675729 649762
rect 675183 648346 675249 648347
rect 675130 648344 675136 648346
rect 675092 648284 675136 648344
rect 675200 648342 675249 648346
rect 675244 648286 675249 648342
rect 675130 648282 675136 648284
rect 675200 648282 675249 648286
rect 675183 648281 675249 648282
rect 675759 648344 675825 648347
rect 676474 648344 676480 648346
rect 675759 648342 676480 648344
rect 675759 648286 675764 648342
rect 675820 648286 676480 648342
rect 675759 648284 676480 648286
rect 675759 648281 675825 648284
rect 676474 648282 676480 648284
rect 676544 648282 676550 648346
rect 675759 645384 675825 645387
rect 676090 645384 676096 645386
rect 675759 645382 676096 645384
rect 675759 645326 675764 645382
rect 675820 645326 676096 645382
rect 675759 645324 676096 645326
rect 675759 645321 675825 645324
rect 676090 645322 676096 645324
rect 676160 645322 676166 645386
rect 41538 644943 41598 645058
rect 41538 644938 41649 644943
rect 41538 644882 41588 644938
rect 41644 644882 41649 644938
rect 41538 644880 41649 644882
rect 41583 644877 41649 644880
rect 40570 644730 40576 644794
rect 40640 644792 40646 644794
rect 41487 644792 41553 644795
rect 40640 644790 41553 644792
rect 40640 644734 41492 644790
rect 41548 644734 41553 644790
rect 40640 644732 41553 644734
rect 40640 644730 40646 644732
rect 41487 644729 41553 644732
rect 41538 644351 41598 644466
rect 41538 644346 41649 644351
rect 41538 644290 41588 644346
rect 41644 644290 41649 644346
rect 41538 644288 41649 644290
rect 41583 644285 41649 644288
rect 41775 644052 41841 644055
rect 41568 644050 41841 644052
rect 41568 643994 41780 644050
rect 41836 643994 41841 644050
rect 41568 643992 41841 643994
rect 41775 643989 41841 643992
rect 41583 643756 41649 643759
rect 41538 643754 41649 643756
rect 41538 643698 41588 643754
rect 41644 643698 41649 643754
rect 41538 643693 41649 643698
rect 41538 643578 41598 643693
rect 649986 643016 650046 643558
rect 655311 643016 655377 643019
rect 649986 643014 655377 643016
rect 41538 642871 41598 642986
rect 649986 642958 655316 643014
rect 655372 642958 655377 643014
rect 649986 642956 655377 642958
rect 655311 642953 655377 642956
rect 41538 642866 41649 642871
rect 41538 642810 41588 642866
rect 41644 642810 41649 642866
rect 41538 642808 41649 642810
rect 41583 642805 41649 642808
rect 41722 642572 41728 642574
rect 41568 642512 41728 642572
rect 41722 642510 41728 642512
rect 41792 642510 41798 642574
rect 655119 642424 655185 642427
rect 649986 642422 655185 642424
rect 649986 642366 655124 642422
rect 655180 642366 655185 642422
rect 649986 642364 655185 642366
rect 655119 642361 655185 642364
rect 40378 642214 40384 642278
rect 40448 642276 40454 642278
rect 43066 642276 43072 642278
rect 40448 642216 43072 642276
rect 40448 642214 40454 642216
rect 43066 642214 43072 642216
rect 43136 642214 43142 642278
rect 40386 642098 40446 642214
rect 41538 641391 41598 641506
rect 41538 641386 41649 641391
rect 41538 641330 41588 641386
rect 41644 641330 41649 641386
rect 41538 641328 41649 641330
rect 41583 641325 41649 641328
rect 41487 641240 41553 641243
rect 41487 641238 41598 641240
rect 41487 641182 41492 641238
rect 41548 641182 41598 641238
rect 41487 641177 41598 641182
rect 41538 640988 41598 641177
rect 649986 640796 650046 641194
rect 655503 640796 655569 640799
rect 649986 640794 655569 640796
rect 649986 640738 655508 640794
rect 655564 640738 655569 640794
rect 649986 640736 655569 640738
rect 655503 640733 655569 640736
rect 41775 640648 41841 640651
rect 654159 640648 654225 640651
rect 41568 640646 41841 640648
rect 41568 640590 41780 640646
rect 41836 640590 41841 640646
rect 41568 640588 41841 640590
rect 41775 640585 41841 640588
rect 649986 640646 654225 640648
rect 649986 640590 654164 640646
rect 654220 640590 654225 640646
rect 649986 640588 654225 640590
rect 42159 640056 42225 640059
rect 41568 640054 42225 640056
rect 41568 639998 42164 640054
rect 42220 639998 42225 640054
rect 649986 640012 650046 640588
rect 654159 640585 654225 640588
rect 41568 639996 42225 639998
rect 42159 639993 42225 639996
rect 39810 639319 39870 639434
rect 39810 639314 39921 639319
rect 39810 639258 39860 639314
rect 39916 639258 39921 639314
rect 39810 639256 39921 639258
rect 39855 639253 39921 639256
rect 42063 639168 42129 639171
rect 655791 639168 655857 639171
rect 41568 639166 42129 639168
rect 41568 639110 42068 639166
rect 42124 639110 42129 639166
rect 41568 639108 42129 639110
rect 42063 639105 42129 639108
rect 649986 639166 655857 639168
rect 649986 639110 655796 639166
rect 655852 639110 655857 639166
rect 649986 639108 655857 639110
rect 649986 638830 650046 639108
rect 655791 639105 655857 639108
rect 41775 638576 41841 638579
rect 41568 638574 41841 638576
rect 41568 638518 41780 638574
rect 41836 638518 41841 638574
rect 41568 638516 41841 638518
rect 41775 638513 41841 638516
rect 655983 638280 656049 638283
rect 649986 638278 656049 638280
rect 649986 638222 655988 638278
rect 656044 638222 656049 638278
rect 649986 638220 656049 638222
rect 41871 637984 41937 637987
rect 41568 637982 41937 637984
rect 41568 637926 41876 637982
rect 41932 637926 41937 637982
rect 41568 637924 41937 637926
rect 41871 637921 41937 637924
rect 649986 637648 650046 638220
rect 655983 638217 656049 638220
rect 34434 637395 34494 637584
rect 34434 637390 34545 637395
rect 34434 637334 34484 637390
rect 34540 637334 34545 637390
rect 34434 637332 34545 637334
rect 34479 637329 34545 637332
rect 42159 637096 42225 637099
rect 41568 637094 42225 637096
rect 41568 637038 42164 637094
rect 42220 637038 42225 637094
rect 41568 637036 42225 637038
rect 42159 637033 42225 637036
rect 41538 636359 41598 636474
rect 41538 636354 41649 636359
rect 41538 636298 41588 636354
rect 41644 636298 41649 636354
rect 41538 636296 41649 636298
rect 41583 636293 41649 636296
rect 41775 636134 41841 636137
rect 41568 636132 41841 636134
rect 41568 636076 41780 636132
rect 41836 636076 41841 636132
rect 41568 636074 41841 636076
rect 41775 636071 41841 636074
rect 41538 635323 41598 635586
rect 41538 635318 41649 635323
rect 41538 635262 41588 635318
rect 41644 635262 41649 635318
rect 41538 635260 41649 635262
rect 41583 635257 41649 635260
rect 41538 634876 41598 634994
rect 41679 634876 41745 634879
rect 41538 634874 41745 634876
rect 41538 634818 41684 634874
rect 41740 634818 41745 634874
rect 41538 634816 41745 634818
rect 41679 634813 41745 634816
rect 41538 634435 41598 634550
rect 41538 634430 41649 634435
rect 41538 634374 41588 634430
rect 41644 634374 41649 634430
rect 41538 634372 41649 634374
rect 41583 634369 41649 634372
rect 42351 634136 42417 634139
rect 41568 634134 42417 634136
rect 41568 634078 42356 634134
rect 42412 634078 42417 634134
rect 41568 634076 42417 634078
rect 42351 634073 42417 634076
rect 41775 633544 41841 633547
rect 41568 633542 41841 633544
rect 41568 633486 41780 633542
rect 41836 633486 41841 633542
rect 41568 633484 41841 633486
rect 41775 633481 41841 633484
rect 28866 632807 28926 633070
rect 28815 632802 28926 632807
rect 28815 632746 28820 632802
rect 28876 632746 28926 632802
rect 28815 632744 28926 632746
rect 28815 632741 28881 632744
rect 41775 632582 41841 632585
rect 41568 632580 41841 632582
rect 41568 632524 41780 632580
rect 41836 632524 41841 632580
rect 41568 632522 41841 632524
rect 41775 632519 41841 632522
rect 28815 632360 28881 632363
rect 28815 632358 28926 632360
rect 28815 632302 28820 632358
rect 28876 632302 28926 632358
rect 28815 632297 28926 632302
rect 28866 632034 28926 632297
rect 39855 628068 39921 628071
rect 40570 628068 40576 628070
rect 39855 628066 40576 628068
rect 39855 628010 39860 628066
rect 39916 628010 40576 628066
rect 39855 628008 40576 628010
rect 39855 628005 39921 628008
rect 40570 628006 40576 628008
rect 40640 628006 40646 628070
rect 34479 627920 34545 627923
rect 40378 627920 40384 627922
rect 34479 627918 40384 627920
rect 34479 627862 34484 627918
rect 34540 627862 40384 627918
rect 34479 627860 40384 627862
rect 34479 627857 34545 627860
rect 40378 627858 40384 627860
rect 40448 627858 40454 627922
rect 676290 625111 676350 625522
rect 676239 625106 676350 625111
rect 676239 625050 676244 625106
rect 676300 625050 676350 625106
rect 676239 625048 676350 625050
rect 676239 625045 676305 625048
rect 676143 624664 676209 624667
rect 676290 624664 676350 624930
rect 676143 624662 676350 624664
rect 676143 624606 676148 624662
rect 676204 624606 676350 624662
rect 676143 624604 676350 624606
rect 676143 624601 676209 624604
rect 676290 624223 676350 624338
rect 676239 624218 676350 624223
rect 676239 624162 676244 624218
rect 676300 624162 676350 624218
rect 676239 624160 676350 624162
rect 679695 624220 679761 624223
rect 679695 624218 679806 624220
rect 679695 624162 679700 624218
rect 679756 624162 679806 624218
rect 676239 624157 676305 624160
rect 679695 624157 679806 624162
rect 679746 623968 679806 624157
rect 676047 623480 676113 623483
rect 676047 623478 676320 623480
rect 676047 623422 676052 623478
rect 676108 623422 676320 623478
rect 676047 623420 676320 623422
rect 676047 623417 676113 623420
rect 676047 622888 676113 622891
rect 676047 622886 676320 622888
rect 676047 622830 676052 622886
rect 676108 622830 676320 622886
rect 676047 622828 676320 622830
rect 676047 622825 676113 622828
rect 676047 622518 676113 622521
rect 676047 622516 676320 622518
rect 676047 622460 676052 622516
rect 676108 622460 676320 622516
rect 676047 622458 676320 622460
rect 676047 622455 676113 622458
rect 676047 622000 676113 622003
rect 676047 621998 676320 622000
rect 676047 621942 676052 621998
rect 676108 621942 676320 621998
rect 676047 621940 676320 621942
rect 676047 621937 676113 621940
rect 676047 621408 676113 621411
rect 676047 621406 676320 621408
rect 676047 621350 676052 621406
rect 676108 621350 676320 621406
rect 676047 621348 676320 621350
rect 676047 621345 676113 621348
rect 674746 620902 674752 620966
rect 674816 620964 674822 620966
rect 674816 620904 676320 620964
rect 674816 620902 674822 620904
rect 676239 620668 676305 620671
rect 676239 620666 676350 620668
rect 676239 620610 676244 620666
rect 676300 620610 676350 620666
rect 676239 620605 676350 620610
rect 676290 620490 676350 620605
rect 675322 619866 675328 619930
rect 675392 619928 675398 619930
rect 675392 619868 676320 619928
rect 675392 619866 675398 619868
rect 676290 619338 676350 619454
rect 676282 619274 676288 619338
rect 676352 619274 676358 619338
rect 676047 618966 676113 618969
rect 676047 618964 676320 618966
rect 676047 618908 676052 618964
rect 676108 618908 676320 618964
rect 676047 618906 676320 618908
rect 676047 618903 676113 618906
rect 676239 618596 676305 618599
rect 676239 618594 676350 618596
rect 676239 618538 676244 618594
rect 676300 618538 676350 618594
rect 676239 618533 676350 618538
rect 676290 618418 676350 618533
rect 58959 618004 59025 618007
rect 58959 618002 64638 618004
rect 58959 617946 58964 618002
rect 59020 617946 64638 618002
rect 58959 617944 64638 617946
rect 58959 617941 59025 617944
rect 64578 617416 64638 617944
rect 674170 617942 674176 618006
rect 674240 618004 674246 618006
rect 674240 617944 676320 618004
rect 674240 617942 674246 617944
rect 674938 617794 674944 617858
rect 675008 617856 675014 617858
rect 675008 617796 676350 617856
rect 675008 617794 675014 617796
rect 676290 617456 676350 617796
rect 673978 616906 673984 616970
rect 674048 616968 674054 616970
rect 674048 616908 676320 616968
rect 674048 616906 674054 616908
rect 40570 616462 40576 616526
rect 40640 616524 40646 616526
rect 42831 616524 42897 616527
rect 40640 616522 42897 616524
rect 40640 616466 42836 616522
rect 42892 616466 42897 616522
rect 40640 616464 42897 616466
rect 40640 616462 40646 616464
rect 42831 616461 42897 616464
rect 676047 616524 676113 616527
rect 676047 616522 676320 616524
rect 676047 616466 676052 616522
rect 676108 616466 676320 616522
rect 676047 616464 676320 616466
rect 676047 616461 676113 616464
rect 40378 616314 40384 616378
rect 40448 616376 40454 616378
rect 42735 616376 42801 616379
rect 40448 616374 42801 616376
rect 40448 616318 42740 616374
rect 42796 616318 42801 616374
rect 40448 616316 42801 616318
rect 40448 616314 40454 616316
rect 42735 616313 42801 616316
rect 59631 616228 59697 616231
rect 64578 616228 64638 616234
rect 59631 616226 64638 616228
rect 59631 616170 59636 616226
rect 59692 616170 64638 616226
rect 59631 616168 64638 616170
rect 59631 616165 59697 616168
rect 676047 615932 676113 615935
rect 676047 615930 676320 615932
rect 676047 615874 676052 615930
rect 676108 615874 676320 615930
rect 676047 615872 676320 615874
rect 676047 615869 676113 615872
rect 58191 615636 58257 615639
rect 676239 615636 676305 615639
rect 58191 615634 64638 615636
rect 58191 615578 58196 615634
rect 58252 615578 64638 615634
rect 58191 615576 64638 615578
rect 58191 615573 58257 615576
rect 64578 615052 64638 615576
rect 676239 615634 676350 615636
rect 676239 615578 676244 615634
rect 676300 615578 676350 615634
rect 676239 615573 676350 615578
rect 676290 615458 676350 615573
rect 677050 615130 677056 615194
rect 677120 615130 677126 615194
rect 677058 615014 677118 615130
rect 58959 614452 59025 614455
rect 676047 614452 676113 614455
rect 58959 614450 64638 614452
rect 58959 614394 58964 614450
rect 59020 614394 64638 614450
rect 58959 614392 64638 614394
rect 58959 614389 59025 614392
rect 64578 613870 64638 614392
rect 676047 614450 676320 614452
rect 676047 614394 676052 614450
rect 676108 614394 676320 614450
rect 676047 614392 676320 614394
rect 676047 614389 676113 614392
rect 679938 613715 679998 613904
rect 679938 613710 680049 613715
rect 679938 613654 679988 613710
rect 680044 613654 680049 613710
rect 679938 613652 680049 613654
rect 679983 613649 680049 613652
rect 679746 613271 679806 613534
rect 59631 613268 59697 613271
rect 59631 613266 64638 613268
rect 59631 613210 59636 613266
rect 59692 613210 64638 613266
rect 59631 613208 64638 613210
rect 679746 613266 679857 613271
rect 679983 613268 680049 613271
rect 679746 613210 679796 613266
rect 679852 613210 679857 613266
rect 679746 613208 679857 613210
rect 59631 613205 59697 613208
rect 64578 612688 64638 613208
rect 679791 613205 679857 613208
rect 679938 613266 680049 613268
rect 679938 613210 679988 613266
rect 680044 613210 680049 613266
rect 679938 613205 680049 613210
rect 679938 612942 679998 613205
rect 679791 612824 679857 612827
rect 679746 612822 679857 612824
rect 679746 612766 679796 612822
rect 679852 612766 679857 612822
rect 679746 612761 679857 612766
rect 679746 612424 679806 612761
rect 59535 612084 59601 612087
rect 59535 612082 64638 612084
rect 59535 612026 59540 612082
rect 59596 612026 64638 612082
rect 59535 612024 64638 612026
rect 59535 612021 59601 612024
rect 64578 611506 64638 612024
rect 674170 607730 674176 607794
rect 674240 607792 674246 607794
rect 675087 607792 675153 607795
rect 674240 607790 675153 607792
rect 674240 607734 675092 607790
rect 675148 607734 675153 607790
rect 674240 607732 675153 607734
rect 674240 607730 674246 607732
rect 675087 607729 675153 607732
rect 674938 607434 674944 607498
rect 675008 607496 675014 607498
rect 675087 607496 675153 607499
rect 675008 607494 675153 607496
rect 675008 607438 675092 607494
rect 675148 607438 675153 607494
rect 675008 607436 675153 607438
rect 675008 607434 675014 607436
rect 675087 607433 675153 607436
rect 675759 606460 675825 606463
rect 675898 606460 675904 606462
rect 675759 606458 675904 606460
rect 675759 606402 675764 606458
rect 675820 606402 675904 606458
rect 675759 606400 675904 606402
rect 675759 606397 675825 606400
rect 675898 606398 675904 606400
rect 675968 606398 675974 606462
rect 674746 604770 674752 604834
rect 674816 604832 674822 604834
rect 675087 604832 675153 604835
rect 674816 604830 675153 604832
rect 674816 604774 675092 604830
rect 675148 604774 675153 604830
rect 674816 604772 675153 604774
rect 674816 604770 674822 604772
rect 675087 604769 675153 604772
rect 41679 602170 41745 602171
rect 41679 602168 41728 602170
rect 41636 602166 41728 602168
rect 41792 602168 41798 602170
rect 62127 602168 62193 602171
rect 41792 602166 62193 602168
rect 41636 602110 41684 602166
rect 41792 602110 62132 602166
rect 62188 602110 62193 602166
rect 41636 602108 41728 602110
rect 41679 602106 41728 602108
rect 41792 602108 62193 602110
rect 41792 602106 41798 602108
rect 41679 602105 41745 602106
rect 62127 602105 62193 602108
rect 675279 602022 675345 602023
rect 675279 602018 675328 602022
rect 675392 602020 675398 602022
rect 675279 601962 675284 602018
rect 675279 601958 675328 601962
rect 675392 601960 675436 602020
rect 675392 601958 675398 601960
rect 675279 601957 675345 601958
rect 41538 601727 41598 601842
rect 41538 601722 41649 601727
rect 41538 601666 41588 601722
rect 41644 601666 41649 601722
rect 41538 601664 41649 601666
rect 41583 601661 41649 601664
rect 41775 601428 41841 601431
rect 41568 601426 41841 601428
rect 41568 601370 41780 601426
rect 41836 601370 41841 601426
rect 41568 601368 41841 601370
rect 41775 601365 41841 601368
rect 41775 600836 41841 600839
rect 41568 600834 41841 600836
rect 41568 600778 41780 600834
rect 41836 600778 41841 600834
rect 41568 600776 41841 600778
rect 41775 600773 41841 600776
rect 41775 600392 41841 600395
rect 41568 600390 41841 600392
rect 41568 600334 41780 600390
rect 41836 600334 41841 600390
rect 41568 600332 41841 600334
rect 41775 600329 41841 600332
rect 675759 600244 675825 600247
rect 676282 600244 676288 600246
rect 675759 600242 676288 600244
rect 675759 600186 675764 600242
rect 675820 600186 676288 600242
rect 675759 600184 676288 600186
rect 675759 600181 675825 600184
rect 676282 600182 676288 600184
rect 676352 600182 676358 600246
rect 41775 599874 41841 599877
rect 41568 599872 41841 599874
rect 41568 599816 41780 599872
rect 41836 599816 41841 599872
rect 41568 599814 41841 599816
rect 41775 599811 41841 599814
rect 41775 599356 41841 599359
rect 41568 599354 41841 599356
rect 41568 599298 41780 599354
rect 41836 599298 41841 599354
rect 41568 599296 41841 599298
rect 41775 599293 41841 599296
rect 39810 598767 39870 598882
rect 39810 598762 39921 598767
rect 39810 598706 39860 598762
rect 39916 598706 39921 598762
rect 39810 598704 39921 598706
rect 39855 598701 39921 598704
rect 41775 598394 41841 598397
rect 41568 598392 41841 598394
rect 41568 598336 41780 598392
rect 41836 598336 41841 598392
rect 41568 598334 41841 598336
rect 41775 598331 41841 598334
rect 41775 597876 41841 597879
rect 41568 597874 41841 597876
rect 41568 597818 41780 597874
rect 41836 597818 41841 597874
rect 41568 597816 41841 597818
rect 649986 597876 650046 598336
rect 655215 597876 655281 597879
rect 649986 597874 655281 597876
rect 649986 597818 655220 597874
rect 655276 597818 655281 597874
rect 649986 597816 655281 597818
rect 41775 597813 41841 597816
rect 655215 597813 655281 597816
rect 41871 597432 41937 597435
rect 41568 597430 41937 597432
rect 41568 597374 41876 597430
rect 41932 597374 41937 597430
rect 41568 597372 41937 597374
rect 41871 597369 41937 597372
rect 41538 596695 41598 596810
rect 41538 596690 41649 596695
rect 41538 596634 41588 596690
rect 41644 596634 41649 596690
rect 41538 596632 41649 596634
rect 649986 596692 650046 597154
rect 655407 596692 655473 596695
rect 649986 596690 655473 596692
rect 649986 596634 655412 596690
rect 655468 596634 655473 596690
rect 649986 596632 655473 596634
rect 41583 596629 41649 596632
rect 655407 596629 655473 596632
rect 34434 596103 34494 596366
rect 34383 596098 34494 596103
rect 34383 596042 34388 596098
rect 34444 596042 34494 596098
rect 34383 596040 34494 596042
rect 34383 596037 34449 596040
rect 41775 595952 41841 595955
rect 41568 595950 41841 595952
rect 41568 595894 41780 595950
rect 41836 595894 41841 595950
rect 41568 595892 41841 595894
rect 41775 595889 41841 595892
rect 649986 595508 650046 595972
rect 655599 595508 655665 595511
rect 649986 595506 655665 595508
rect 649986 595450 655604 595506
rect 655660 595450 655665 595506
rect 649986 595448 655665 595450
rect 655599 595445 655665 595448
rect 655791 595360 655857 595363
rect 649986 595358 655857 595360
rect 41538 595215 41598 595330
rect 649986 595302 655796 595358
rect 655852 595302 655857 595358
rect 649986 595300 655857 595302
rect 41538 595210 41649 595215
rect 41538 595154 41588 595210
rect 41644 595154 41649 595210
rect 41538 595152 41649 595154
rect 41583 595149 41649 595152
rect 41775 594842 41841 594845
rect 41568 594840 41841 594842
rect 41568 594784 41780 594840
rect 41836 594784 41841 594840
rect 649986 594790 650046 595300
rect 655791 595297 655857 595300
rect 41568 594782 41841 594784
rect 41775 594779 41841 594782
rect 34434 594179 34494 594442
rect 34434 594174 34545 594179
rect 653967 594176 654033 594179
rect 34434 594118 34484 594174
rect 34540 594118 34545 594174
rect 34434 594116 34545 594118
rect 34479 594113 34545 594116
rect 649986 594174 654033 594176
rect 649986 594118 653972 594174
rect 654028 594118 654033 594174
rect 649986 594116 654033 594118
rect 41538 593735 41598 593850
rect 41538 593730 41649 593735
rect 41538 593674 41588 593730
rect 41644 593674 41649 593730
rect 41538 593672 41649 593674
rect 41583 593669 41649 593672
rect 649986 593608 650046 594116
rect 653967 594113 654033 594116
rect 42063 593362 42129 593365
rect 41568 593360 42129 593362
rect 41568 593304 42068 593360
rect 42124 593304 42129 593360
rect 41568 593302 42129 593304
rect 42063 593299 42129 593302
rect 42255 592992 42321 592995
rect 656559 592992 656625 592995
rect 41568 592990 42321 592992
rect 41568 592934 42260 592990
rect 42316 592934 42321 592990
rect 41568 592932 42321 592934
rect 42255 592929 42321 592932
rect 649986 592990 656625 592992
rect 649986 592934 656564 592990
rect 656620 592934 656625 592990
rect 649986 592932 656625 592934
rect 649986 592426 650046 592932
rect 656559 592929 656625 592932
rect 41538 592252 41598 592370
rect 41679 592252 41745 592255
rect 41538 592250 41745 592252
rect 41538 592194 41684 592250
rect 41740 592194 41745 592250
rect 41538 592192 41745 592194
rect 41679 592189 41745 592192
rect 42351 591808 42417 591811
rect 41568 591806 42417 591808
rect 41568 591750 42356 591806
rect 42412 591750 42417 591806
rect 41568 591748 42417 591750
rect 42351 591745 42417 591748
rect 41538 591219 41598 591408
rect 41538 591214 41649 591219
rect 41538 591158 41588 591214
rect 41644 591158 41649 591214
rect 41538 591156 41649 591158
rect 41583 591153 41649 591156
rect 41967 590920 42033 590923
rect 41568 590918 42033 590920
rect 41568 590862 41972 590918
rect 42028 590862 42033 590918
rect 41568 590860 42033 590862
rect 41967 590857 42033 590860
rect 41538 590180 41598 590298
rect 41538 590120 41790 590180
rect 28866 589591 28926 589928
rect 41730 589736 41790 590120
rect 28815 589586 28926 589591
rect 28815 589530 28820 589586
rect 28876 589530 28926 589586
rect 28815 589528 28926 589530
rect 41538 589676 41790 589736
rect 28815 589525 28881 589528
rect 41538 589147 41598 589676
rect 28815 589144 28881 589147
rect 28815 589142 28926 589144
rect 28815 589086 28820 589142
rect 28876 589086 28926 589142
rect 28815 589081 28926 589086
rect 41538 589142 41649 589147
rect 41538 589086 41588 589142
rect 41644 589086 41649 589142
rect 41538 589084 41649 589086
rect 41583 589081 41649 589084
rect 28866 588818 28926 589081
rect 42927 587518 42993 587519
rect 42874 587516 42880 587518
rect 42836 587456 42880 587516
rect 42944 587514 42993 587518
rect 42988 587458 42993 587514
rect 42874 587454 42880 587456
rect 42944 587454 42993 587458
rect 42927 587453 42993 587454
rect 34479 586274 34545 586277
rect 40378 586274 40384 586276
rect 34479 586272 40384 586274
rect 34479 586216 34484 586272
rect 34540 586216 40384 586272
rect 34479 586214 40384 586216
rect 34479 586211 34545 586214
rect 40378 586212 40384 586214
rect 40448 586212 40454 586276
rect 34383 585978 34449 585981
rect 40570 585978 40576 585980
rect 34383 585976 40576 585978
rect 34383 585920 34388 585976
rect 34444 585920 40576 585976
rect 34383 585918 40576 585920
rect 34383 585915 34449 585918
rect 40570 585916 40576 585918
rect 40640 585916 40646 585980
rect 676290 578343 676350 578458
rect 676290 578338 676401 578343
rect 676290 578282 676340 578338
rect 676396 578282 676401 578338
rect 676290 578280 676401 578282
rect 676335 578277 676401 578280
rect 676143 577600 676209 577603
rect 676290 577600 676350 577866
rect 676143 577598 676350 577600
rect 676143 577542 676148 577598
rect 676204 577542 676350 577598
rect 676143 577540 676350 577542
rect 676143 577537 676209 577540
rect 42831 577306 42897 577307
rect 42831 577304 42880 577306
rect 42788 577302 42880 577304
rect 42788 577246 42836 577302
rect 42788 577244 42880 577246
rect 42831 577242 42880 577244
rect 42944 577242 42950 577306
rect 42831 577241 42897 577242
rect 676290 577159 676350 577422
rect 676239 577154 676350 577159
rect 676239 577098 676244 577154
rect 676300 577098 676350 577154
rect 676239 577096 676350 577098
rect 679695 577156 679761 577159
rect 679695 577154 679806 577156
rect 679695 577098 679700 577154
rect 679756 577098 679806 577154
rect 676239 577093 676305 577096
rect 679695 577093 679806 577098
rect 679746 576978 679806 577093
rect 676290 576271 676350 576386
rect 676239 576266 676350 576271
rect 676239 576210 676244 576266
rect 676300 576210 676350 576266
rect 676239 576208 676350 576210
rect 676239 576205 676305 576208
rect 675951 575972 676017 575975
rect 675951 575970 676320 575972
rect 675951 575914 675956 575970
rect 676012 575914 676320 575970
rect 675951 575912 676320 575914
rect 675951 575909 676017 575912
rect 675951 575528 676017 575531
rect 675951 575526 676320 575528
rect 675951 575470 675956 575526
rect 676012 575470 676320 575526
rect 675951 575468 676320 575470
rect 675951 575465 676017 575468
rect 675951 574936 676017 574939
rect 675951 574934 676320 574936
rect 675951 574878 675956 574934
rect 676012 574878 676320 574934
rect 675951 574876 676320 574878
rect 675951 574873 676017 574876
rect 58959 574788 59025 574791
rect 58959 574786 64638 574788
rect 58959 574730 58964 574786
rect 59020 574730 64638 574786
rect 58959 574728 64638 574730
rect 58959 574725 59025 574728
rect 64578 574194 64638 574728
rect 676290 574199 676350 574388
rect 676239 574194 676350 574199
rect 676239 574138 676244 574194
rect 676300 574138 676350 574194
rect 676239 574136 676350 574138
rect 676239 574133 676305 574136
rect 40378 573986 40384 574050
rect 40448 574048 40454 574050
rect 42255 574048 42321 574051
rect 40448 574046 42321 574048
rect 40448 573990 42260 574046
rect 42316 573990 42321 574046
rect 40448 573988 42321 573990
rect 40448 573986 40454 573988
rect 42255 573985 42321 573988
rect 675514 573986 675520 574050
rect 675584 574048 675590 574050
rect 675584 573988 676320 574048
rect 675584 573986 675590 573988
rect 40570 573838 40576 573902
rect 40640 573900 40646 573902
rect 42543 573900 42609 573903
rect 40640 573898 42609 573900
rect 40640 573842 42548 573898
rect 42604 573842 42609 573898
rect 40640 573840 42609 573842
rect 40640 573838 40646 573840
rect 42543 573837 42609 573840
rect 676047 573456 676113 573459
rect 676047 573454 676320 573456
rect 676047 573398 676052 573454
rect 676108 573398 676320 573454
rect 676047 573396 676320 573398
rect 676047 573393 676113 573396
rect 59631 573012 59697 573015
rect 59631 573010 64638 573012
rect 59631 572954 59636 573010
rect 59692 572954 64638 573010
rect 59631 572952 64638 572954
rect 59631 572949 59697 572952
rect 674554 572802 674560 572866
rect 674624 572864 674630 572866
rect 674624 572804 676320 572864
rect 674624 572802 674630 572804
rect 675706 572506 675712 572570
rect 675776 572568 675782 572570
rect 675776 572508 676320 572568
rect 675776 572506 675782 572508
rect 58191 572420 58257 572423
rect 58191 572418 64638 572420
rect 58191 572362 58196 572418
rect 58252 572362 64638 572418
rect 58191 572360 64638 572362
rect 58191 572357 58257 572360
rect 64578 571830 64638 572360
rect 676090 572210 676096 572274
rect 676160 572272 676166 572274
rect 676160 572212 676350 572272
rect 676160 572210 676166 572212
rect 676290 571946 676350 572212
rect 676047 571384 676113 571387
rect 676047 571382 676320 571384
rect 676047 571326 676052 571382
rect 676108 571326 676320 571382
rect 676047 571324 676320 571326
rect 676047 571321 676113 571324
rect 58959 571236 59025 571239
rect 58959 571234 64638 571236
rect 58959 571178 58964 571234
rect 59020 571178 64638 571234
rect 58959 571176 64638 571178
rect 58959 571173 59025 571176
rect 64578 570648 64638 571176
rect 674362 571174 674368 571238
rect 674432 571236 674438 571238
rect 674432 571176 676350 571236
rect 674432 571174 674438 571176
rect 676290 570984 676350 571176
rect 675130 570434 675136 570498
rect 675200 570496 675206 570498
rect 675200 570436 676320 570496
rect 675200 570434 675206 570436
rect 676474 570138 676480 570202
rect 676544 570138 676550 570202
rect 59343 570052 59409 570055
rect 59343 570050 64638 570052
rect 59343 569994 59348 570050
rect 59404 569994 64638 570050
rect 59343 569992 64638 569994
rect 59343 569989 59409 569992
rect 64578 569466 64638 569992
rect 676482 569874 676542 570138
rect 676047 569534 676113 569537
rect 676047 569532 676320 569534
rect 676047 569476 676052 569532
rect 676108 569476 676320 569532
rect 676047 569474 676320 569476
rect 676047 569471 676113 569474
rect 676239 569164 676305 569167
rect 676239 569162 676350 569164
rect 676239 569106 676244 569162
rect 676300 569106 676350 569162
rect 676239 569101 676350 569106
rect 676290 568986 676350 569101
rect 59535 568868 59601 568871
rect 59535 568866 64638 568868
rect 59535 568810 59540 568866
rect 59596 568810 64638 568866
rect 59535 568808 64638 568810
rect 59535 568805 59601 568808
rect 64578 568284 64638 568808
rect 676047 568424 676113 568427
rect 676047 568422 676320 568424
rect 676047 568366 676052 568422
rect 676108 568366 676320 568422
rect 676047 568364 676320 568366
rect 676047 568361 676113 568364
rect 676047 567980 676113 567983
rect 676047 567978 676320 567980
rect 676047 567922 676052 567978
rect 676108 567922 676320 567978
rect 676047 567920 676320 567922
rect 676047 567917 676113 567920
rect 676239 567684 676305 567687
rect 676239 567682 676350 567684
rect 676239 567626 676244 567682
rect 676300 567626 676350 567682
rect 676239 567621 676350 567626
rect 676290 567506 676350 567621
rect 679791 567092 679857 567095
rect 679746 567090 679857 567092
rect 679746 567034 679796 567090
rect 679852 567034 679857 567090
rect 679746 567029 679857 567034
rect 679746 566914 679806 567029
rect 685506 566207 685566 566470
rect 679791 566204 679857 566207
rect 679746 566202 679857 566204
rect 679746 566146 679796 566202
rect 679852 566146 679857 566202
rect 679746 566141 679857 566146
rect 685455 566202 685566 566207
rect 685455 566146 685460 566202
rect 685516 566146 685566 566202
rect 685455 566144 685566 566146
rect 685455 566141 685521 566144
rect 679746 565952 679806 566141
rect 685455 565760 685521 565763
rect 685455 565758 685566 565760
rect 685455 565702 685460 565758
rect 685516 565702 685566 565758
rect 685455 565697 685566 565702
rect 685506 565434 685566 565697
rect 674362 562886 674368 562950
rect 674432 562948 674438 562950
rect 675087 562948 675153 562951
rect 674432 562946 675153 562948
rect 674432 562890 675092 562946
rect 675148 562890 675153 562946
rect 674432 562888 675153 562890
rect 674432 562886 674438 562888
rect 675087 562885 675153 562888
rect 675471 561766 675537 561767
rect 675471 561762 675520 561766
rect 675584 561764 675590 561766
rect 675471 561706 675476 561762
rect 675471 561702 675520 561706
rect 675584 561704 675628 561764
rect 675584 561702 675590 561704
rect 675471 561701 675537 561702
rect 675130 561406 675136 561470
rect 675200 561468 675206 561470
rect 675375 561468 675441 561471
rect 675200 561466 675441 561468
rect 675200 561410 675380 561466
rect 675436 561410 675441 561466
rect 675200 561408 675441 561410
rect 675200 561406 675206 561408
rect 675375 561405 675441 561408
rect 674554 558890 674560 558954
rect 674624 558952 674630 558954
rect 675471 558952 675537 558955
rect 674624 558950 675537 558952
rect 674624 558894 675476 558950
rect 675532 558894 675537 558950
rect 674624 558892 675537 558894
rect 674624 558890 674630 558892
rect 675471 558889 675537 558892
rect 675759 554660 675825 554663
rect 677050 554660 677056 554662
rect 675759 554658 677056 554660
rect 675759 554602 675764 554658
rect 675820 554602 677056 554658
rect 675759 554600 677056 554602
rect 675759 554597 675825 554600
rect 677050 554598 677056 554600
rect 677120 554598 677126 554662
rect 649986 553328 650046 553914
rect 655119 553328 655185 553331
rect 649986 553326 655185 553328
rect 649986 553270 655124 553326
rect 655180 553270 655185 553326
rect 649986 553268 655185 553270
rect 655119 553265 655185 553268
rect 675279 553328 675345 553331
rect 676858 553328 676864 553330
rect 675279 553326 676864 553328
rect 675279 553270 675284 553326
rect 675340 553270 676864 553326
rect 675279 553268 676864 553270
rect 675279 553265 675345 553268
rect 676858 553266 676864 553268
rect 676928 553266 676934 553330
rect 649986 552144 650046 552732
rect 655503 552144 655569 552147
rect 649986 552142 655569 552144
rect 649986 552086 655508 552142
rect 655564 552086 655569 552142
rect 649986 552084 655569 552086
rect 655503 552081 655569 552084
rect 649986 550960 650046 551550
rect 655311 550960 655377 550963
rect 649986 550958 655377 550960
rect 649986 550902 655316 550958
rect 655372 550902 655377 550958
rect 649986 550900 655377 550902
rect 655311 550897 655377 550900
rect 655695 550812 655761 550815
rect 649986 550810 655761 550812
rect 649986 550754 655700 550810
rect 655756 550754 655761 550810
rect 649986 550752 655761 550754
rect 649986 550368 650046 550752
rect 655695 550749 655761 550752
rect 656559 549776 656625 549779
rect 649986 549774 656625 549776
rect 649986 549718 656564 549774
rect 656620 549718 656625 549774
rect 649986 549716 656625 549718
rect 649986 549186 650046 549716
rect 656559 549713 656625 549716
rect 654159 548592 654225 548595
rect 649986 548590 654225 548592
rect 649986 548534 654164 548590
rect 654220 548534 654225 548590
rect 649986 548532 654225 548534
rect 649986 548004 650046 548532
rect 654159 548529 654225 548532
rect 40378 539798 40384 539862
rect 40448 539860 40454 539862
rect 41775 539860 41841 539863
rect 40448 539858 41841 539860
rect 40448 539802 41780 539858
rect 41836 539802 41841 539858
rect 40448 539800 41841 539802
rect 40448 539798 40454 539800
rect 41775 539797 41841 539800
rect 41530 538022 41536 538086
rect 41600 538084 41606 538086
rect 41775 538084 41841 538087
rect 41600 538082 41841 538084
rect 41600 538026 41780 538082
rect 41836 538026 41841 538082
rect 41600 538024 41841 538026
rect 41600 538022 41606 538024
rect 41775 538021 41841 538024
rect 43066 536986 43072 537050
rect 43136 537048 43142 537050
rect 62319 537048 62385 537051
rect 43136 537046 62385 537048
rect 43136 536990 62324 537046
rect 62380 536990 62385 537046
rect 43136 536988 62385 536990
rect 43136 536986 43142 536988
rect 62319 536985 62385 536988
rect 40954 536246 40960 536310
rect 41024 536308 41030 536310
rect 41775 536308 41841 536311
rect 41024 536306 41841 536308
rect 41024 536250 41780 536306
rect 41836 536250 41841 536306
rect 41024 536248 41841 536250
rect 41024 536246 41030 536248
rect 41775 536245 41841 536248
rect 40762 535062 40768 535126
rect 40832 535124 40838 535126
rect 41775 535124 41841 535127
rect 40832 535122 41841 535124
rect 40832 535066 41780 535122
rect 41836 535066 41841 535122
rect 40832 535064 41841 535066
rect 40832 535062 40838 535064
rect 41775 535061 41841 535064
rect 676290 534979 676350 535242
rect 676239 534974 676350 534979
rect 676239 534918 676244 534974
rect 676300 534918 676350 534974
rect 676239 534916 676350 534918
rect 676239 534913 676305 534916
rect 676143 534384 676209 534387
rect 676290 534384 676350 534724
rect 676143 534382 676350 534384
rect 676143 534326 676148 534382
rect 676204 534326 676350 534382
rect 676143 534324 676350 534326
rect 676143 534321 676209 534324
rect 41338 534174 41344 534238
rect 41408 534236 41414 534238
rect 41775 534236 41841 534239
rect 41408 534234 41841 534236
rect 41408 534178 41780 534234
rect 41836 534178 41841 534234
rect 41408 534176 41841 534178
rect 41408 534174 41414 534176
rect 41775 534173 41841 534176
rect 676047 534236 676113 534239
rect 676047 534234 676320 534236
rect 676047 534178 676052 534234
rect 676108 534178 676320 534234
rect 676047 534176 676320 534178
rect 676047 534173 676113 534176
rect 40570 533878 40576 533942
rect 40640 533940 40646 533942
rect 41775 533940 41841 533943
rect 40640 533938 41841 533940
rect 40640 533882 41780 533938
rect 41836 533882 41841 533938
rect 40640 533880 41841 533882
rect 40640 533878 40646 533880
rect 41775 533877 41841 533880
rect 679746 533647 679806 533762
rect 679695 533642 679806 533647
rect 679695 533586 679700 533642
rect 679756 533586 679806 533642
rect 679695 533584 679806 533586
rect 679695 533581 679761 533584
rect 676482 533055 676542 533170
rect 41871 533054 41937 533055
rect 41871 533050 41920 533054
rect 41984 533052 41990 533054
rect 41871 532994 41876 533050
rect 41871 532990 41920 532994
rect 41984 532992 42028 533052
rect 676482 533050 676593 533055
rect 676482 532994 676532 533050
rect 676588 532994 676593 533050
rect 676482 532992 676593 532994
rect 41984 532990 41990 532992
rect 41871 532989 41937 532990
rect 676527 532989 676593 532992
rect 675951 532756 676017 532759
rect 675951 532754 676320 532756
rect 675951 532698 675956 532754
rect 676012 532698 676320 532754
rect 675951 532696 676320 532698
rect 675951 532693 676017 532696
rect 676674 532019 676734 532282
rect 676623 532014 676734 532019
rect 676623 531958 676628 532014
rect 676684 531958 676734 532014
rect 676623 531956 676734 531958
rect 676623 531953 676689 531956
rect 57711 531720 57777 531723
rect 57711 531718 64638 531720
rect 57711 531662 57716 531718
rect 57772 531662 64638 531718
rect 57711 531660 64638 531662
rect 57711 531657 57777 531660
rect 64578 531172 64638 531660
rect 676290 531575 676350 531690
rect 676239 531570 676350 531575
rect 676239 531514 676244 531570
rect 676300 531514 676350 531570
rect 676239 531512 676350 531514
rect 676239 531509 676305 531512
rect 676674 530983 676734 531246
rect 676674 530978 676785 530983
rect 676674 530922 676724 530978
rect 676780 530922 676785 530978
rect 676674 530920 676785 530922
rect 676719 530917 676785 530920
rect 41146 530770 41152 530834
rect 41216 530832 41222 530834
rect 41775 530832 41841 530835
rect 41216 530830 41841 530832
rect 41216 530774 41780 530830
rect 41836 530774 41841 530830
rect 41216 530772 41841 530774
rect 41216 530770 41222 530772
rect 41775 530769 41841 530772
rect 675898 530770 675904 530834
rect 675968 530832 675974 530834
rect 675968 530772 676320 530832
rect 675968 530770 675974 530772
rect 57615 530536 57681 530539
rect 57615 530534 64638 530536
rect 57615 530478 57620 530534
rect 57676 530478 64638 530534
rect 57615 530476 64638 530478
rect 57615 530473 57681 530476
rect 41775 530094 41841 530095
rect 41722 530092 41728 530094
rect 41684 530032 41728 530092
rect 41792 530090 41841 530094
rect 41836 530034 41841 530090
rect 41722 530030 41728 530032
rect 41792 530030 41841 530034
rect 41775 530029 41841 530030
rect 64578 529990 64638 530476
rect 676047 530240 676113 530243
rect 676047 530238 676320 530240
rect 676047 530182 676052 530238
rect 676108 530182 676320 530238
rect 676047 530180 676320 530182
rect 676047 530177 676113 530180
rect 674170 529882 674176 529946
rect 674240 529944 674246 529946
rect 674240 529884 676350 529944
rect 674240 529882 674246 529884
rect 676290 529692 676350 529884
rect 42159 529354 42225 529355
rect 42106 529352 42112 529354
rect 42068 529292 42112 529352
rect 42176 529350 42225 529354
rect 42220 529294 42225 529350
rect 42106 529290 42112 529292
rect 42176 529290 42225 529294
rect 42159 529289 42225 529290
rect 58191 529352 58257 529355
rect 58191 529350 64638 529352
rect 58191 529294 58196 529350
rect 58252 529294 64638 529350
rect 58191 529292 64638 529294
rect 58191 529289 58257 529292
rect 64578 528808 64638 529292
rect 674746 529290 674752 529354
rect 674816 529352 674822 529354
rect 674816 529292 676320 529352
rect 674816 529290 674822 529292
rect 676282 528994 676288 529058
rect 676352 528994 676358 529058
rect 676290 528730 676350 528994
rect 676047 528168 676113 528171
rect 676047 528166 676320 528168
rect 676047 528110 676052 528166
rect 676108 528110 676320 528166
rect 676047 528108 676320 528110
rect 676047 528105 676113 528108
rect 674938 527810 674944 527874
rect 675008 527872 675014 527874
rect 675008 527812 676320 527872
rect 675008 527810 675014 527812
rect 42159 527280 42225 527283
rect 42490 527280 42496 527282
rect 42159 527278 42496 527280
rect 42159 527222 42164 527278
rect 42220 527222 42496 527278
rect 42159 527220 42496 527222
rect 42159 527217 42225 527220
rect 42490 527218 42496 527220
rect 42560 527218 42566 527282
rect 42255 527134 42321 527135
rect 42255 527130 42304 527134
rect 42368 527132 42374 527134
rect 58959 527132 59025 527135
rect 64578 527132 64638 527626
rect 675322 527218 675328 527282
rect 675392 527280 675398 527282
rect 675392 527220 676320 527280
rect 675392 527218 675398 527220
rect 42255 527074 42260 527130
rect 42255 527070 42304 527074
rect 42368 527072 42412 527132
rect 58959 527130 64638 527132
rect 58959 527074 58964 527130
rect 59020 527074 64638 527130
rect 58959 527072 64638 527074
rect 42368 527070 42374 527072
rect 42255 527069 42321 527070
rect 58959 527069 59025 527072
rect 676047 526688 676113 526691
rect 676047 526686 676320 526688
rect 676047 526630 676052 526686
rect 676108 526630 676320 526686
rect 676047 526628 676320 526630
rect 676047 526625 676113 526628
rect 58575 525948 58641 525951
rect 64578 525948 64638 526444
rect 676047 526318 676113 526321
rect 676047 526316 676320 526318
rect 676047 526260 676052 526316
rect 676108 526260 676320 526316
rect 676047 526258 676320 526260
rect 676047 526255 676113 526258
rect 58575 525946 64638 525948
rect 58575 525890 58580 525946
rect 58636 525890 64638 525946
rect 58575 525888 64638 525890
rect 676239 525948 676305 525951
rect 676239 525946 676350 525948
rect 676239 525890 676244 525946
rect 676300 525890 676350 525946
rect 58575 525885 58641 525888
rect 676239 525885 676350 525890
rect 676290 525770 676350 525885
rect 59343 524764 59409 524767
rect 64578 524764 64638 525262
rect 676047 525208 676113 525211
rect 676047 525206 676320 525208
rect 676047 525150 676052 525206
rect 676108 525150 676320 525206
rect 676047 525148 676320 525150
rect 676047 525145 676113 525148
rect 676047 524838 676113 524841
rect 676047 524836 676320 524838
rect 676047 524780 676052 524836
rect 676108 524780 676320 524836
rect 676047 524778 676320 524780
rect 676047 524775 676113 524778
rect 59343 524762 64638 524764
rect 59343 524706 59348 524762
rect 59404 524706 64638 524762
rect 59343 524704 64638 524706
rect 59343 524701 59409 524704
rect 676239 524468 676305 524471
rect 676239 524466 676350 524468
rect 676239 524410 676244 524466
rect 676300 524410 676350 524466
rect 676239 524405 676350 524410
rect 676290 524290 676350 524405
rect 679746 523583 679806 523698
rect 679746 523578 679857 523583
rect 679746 523522 679796 523578
rect 679852 523522 679857 523578
rect 679746 523520 679857 523522
rect 679791 523517 679857 523520
rect 685506 522991 685566 523254
rect 679791 522988 679857 522991
rect 679746 522986 679857 522988
rect 679746 522930 679796 522986
rect 679852 522930 679857 522986
rect 679746 522925 679857 522930
rect 685455 522986 685566 522991
rect 685455 522930 685460 522986
rect 685516 522930 685566 522986
rect 685455 522928 685566 522930
rect 685455 522925 685521 522928
rect 679746 522810 679806 522925
rect 685455 522544 685521 522547
rect 685455 522542 685566 522544
rect 685455 522486 685460 522542
rect 685516 522486 685566 522542
rect 685455 522481 685566 522486
rect 685506 522218 685566 522481
rect 676290 490579 676350 490842
rect 676239 490574 676350 490579
rect 676239 490518 676244 490574
rect 676300 490518 676350 490574
rect 676239 490516 676350 490518
rect 676239 490513 676305 490516
rect 676143 490132 676209 490135
rect 676290 490132 676350 490324
rect 676143 490130 676350 490132
rect 676143 490074 676148 490130
rect 676204 490074 676350 490130
rect 676143 490072 676350 490074
rect 676143 490069 676209 490072
rect 676239 489984 676305 489987
rect 676239 489982 676350 489984
rect 676239 489926 676244 489982
rect 676300 489926 676350 489982
rect 676239 489921 676350 489926
rect 676290 489806 676350 489921
rect 679746 489247 679806 489362
rect 679695 489242 679806 489247
rect 679695 489186 679700 489242
rect 679756 489186 679806 489242
rect 679695 489184 679806 489186
rect 679695 489181 679761 489184
rect 676674 488655 676734 488770
rect 676674 488650 676785 488655
rect 676674 488594 676724 488650
rect 676780 488594 676785 488650
rect 676674 488592 676785 488594
rect 676719 488589 676785 488592
rect 676047 488356 676113 488359
rect 676047 488354 676320 488356
rect 676047 488298 676052 488354
rect 676108 488298 676320 488354
rect 676047 488296 676320 488298
rect 676047 488293 676113 488296
rect 675279 487912 675345 487915
rect 675279 487910 676320 487912
rect 675279 487854 675284 487910
rect 675340 487854 676320 487910
rect 675279 487852 676320 487854
rect 675279 487849 675345 487852
rect 676290 487175 676350 487290
rect 676239 487170 676350 487175
rect 676239 487114 676244 487170
rect 676300 487114 676350 487170
rect 676239 487112 676350 487114
rect 676239 487109 676305 487112
rect 676047 486876 676113 486879
rect 676047 486874 676320 486876
rect 676047 486818 676052 486874
rect 676108 486818 676320 486874
rect 676047 486816 676320 486818
rect 676047 486813 676113 486816
rect 675130 486370 675136 486434
rect 675200 486432 675206 486434
rect 675200 486372 676320 486432
rect 675200 486370 675206 486372
rect 676047 485840 676113 485843
rect 676047 485838 676320 485840
rect 676047 485782 676052 485838
rect 676108 485782 676320 485838
rect 676047 485780 676320 485782
rect 676047 485777 676113 485780
rect 674362 485630 674368 485694
rect 674432 485692 674438 485694
rect 674432 485632 676350 485692
rect 674432 485630 674438 485632
rect 676290 485292 676350 485632
rect 676239 485100 676305 485103
rect 676239 485098 676350 485100
rect 676239 485042 676244 485098
rect 676300 485042 676350 485098
rect 676239 485037 676350 485042
rect 676290 484922 676350 485037
rect 676047 484360 676113 484363
rect 676047 484358 676320 484360
rect 676047 484302 676052 484358
rect 676108 484302 676320 484358
rect 676047 484300 676320 484302
rect 676047 484297 676113 484300
rect 675951 483768 676017 483771
rect 675951 483766 676320 483768
rect 675951 483710 675956 483766
rect 676012 483710 676320 483766
rect 675951 483708 676320 483710
rect 675951 483705 676017 483708
rect 675514 483410 675520 483474
rect 675584 483472 675590 483474
rect 675584 483412 676320 483472
rect 675584 483410 675590 483412
rect 674554 482818 674560 482882
rect 674624 482880 674630 482882
rect 674624 482820 676320 482880
rect 674624 482818 674630 482820
rect 676047 482288 676113 482291
rect 676047 482286 676320 482288
rect 676047 482230 676052 482286
rect 676108 482230 676320 482286
rect 676047 482228 676320 482230
rect 676047 482225 676113 482228
rect 676047 481918 676113 481921
rect 676047 481916 676320 481918
rect 676047 481860 676052 481916
rect 676108 481860 676320 481916
rect 676047 481858 676320 481860
rect 676047 481855 676113 481858
rect 676239 481548 676305 481551
rect 676239 481546 676350 481548
rect 676239 481490 676244 481546
rect 676300 481490 676350 481546
rect 676239 481485 676350 481490
rect 676290 481370 676350 481485
rect 676858 481042 676864 481106
rect 676928 481042 676934 481106
rect 40762 480746 40768 480810
rect 40832 480808 40838 480810
rect 42682 480808 42688 480810
rect 40832 480748 42688 480808
rect 40832 480746 40838 480748
rect 42682 480746 42688 480748
rect 42752 480746 42758 480810
rect 676866 480778 676926 481042
rect 677050 480598 677056 480662
rect 677120 480598 677126 480662
rect 677058 480408 677118 480598
rect 676239 480068 676305 480071
rect 676239 480066 676350 480068
rect 676239 480010 676244 480066
rect 676300 480010 676350 480066
rect 676239 480005 676350 480010
rect 676290 479890 676350 480005
rect 679938 479183 679998 479298
rect 679887 479178 679998 479183
rect 679887 479122 679892 479178
rect 679948 479122 679998 479178
rect 679887 479120 679998 479122
rect 679887 479117 679953 479120
rect 679746 478591 679806 478854
rect 679695 478586 679806 478591
rect 679695 478530 679700 478586
rect 679756 478530 679806 478586
rect 679695 478528 679806 478530
rect 679887 478588 679953 478591
rect 679887 478586 679998 478588
rect 679887 478530 679892 478586
rect 679948 478530 679998 478586
rect 679695 478525 679761 478528
rect 679887 478525 679998 478530
rect 679938 478410 679998 478525
rect 40570 478082 40576 478146
rect 40640 478144 40646 478146
rect 43207 478144 43273 478147
rect 40640 478142 43273 478144
rect 40640 478086 43212 478142
rect 43268 478086 43273 478142
rect 40640 478084 43273 478086
rect 40640 478082 40646 478084
rect 43207 478081 43273 478084
rect 679695 478144 679761 478147
rect 679695 478142 679806 478144
rect 679695 478086 679700 478142
rect 679756 478086 679806 478142
rect 679695 478081 679806 478086
rect 679746 477818 679806 478081
rect 41483 476109 41553 476114
rect 41483 476049 41488 476109
rect 41548 476049 41553 476109
rect 41483 476044 41553 476049
rect 41506 475591 41576 475596
rect 41506 475531 41511 475591
rect 41571 475531 41576 475591
rect 41506 475526 41576 475531
rect 41093 475009 41163 475014
rect 41093 474949 41098 475009
rect 41158 474949 41163 475009
rect 41093 474944 41163 474949
rect 41464 474629 41534 474634
rect 41464 474569 41469 474629
rect 41529 474569 41534 474629
rect 41464 474564 41534 474569
rect 40386 473855 40446 473970
rect 40335 473850 40446 473855
rect 40335 473794 40340 473850
rect 40396 473794 40446 473850
rect 40335 473792 40446 473794
rect 40335 473789 40401 473792
rect 39810 473263 39870 473526
rect 39759 473258 39870 473263
rect 39759 473202 39764 473258
rect 39820 473202 39870 473258
rect 39759 473200 39870 473202
rect 39759 473197 39825 473200
rect 40570 473198 40576 473262
rect 40640 473198 40646 473262
rect 40578 473112 40638 473198
rect 43066 473112 43072 473114
rect 40578 473082 43072 473112
rect 40608 473052 43072 473082
rect 43066 473050 43072 473052
rect 43136 473050 43142 473114
rect 39618 472375 39678 472490
rect 39618 472370 39729 472375
rect 39618 472314 39668 472370
rect 39724 472314 39729 472370
rect 39618 472312 39729 472314
rect 39663 472309 39729 472312
rect 42255 472224 42321 472227
rect 43119 472224 43185 472227
rect 41538 472222 43185 472224
rect 41538 472166 42260 472222
rect 42316 472166 43124 472222
rect 43180 472166 43185 472222
rect 41538 472164 43185 472166
rect 41538 472046 41598 472164
rect 42255 472161 42321 472164
rect 43119 472161 43185 472164
rect 42490 471632 42496 471634
rect 41568 471572 42496 471632
rect 42490 471570 42496 471572
rect 42560 471570 42566 471634
rect 41530 471274 41536 471338
rect 41600 471274 41606 471338
rect 41538 471010 41598 471274
rect 42447 470596 42513 470599
rect 41538 470594 42513 470596
rect 41538 470538 42452 470594
rect 42508 470538 42513 470594
rect 41538 470536 42513 470538
rect 41538 470492 41598 470536
rect 42447 470533 42513 470536
rect 42298 470152 42304 470154
rect 41568 470092 42304 470152
rect 42298 470090 42304 470092
rect 42368 470090 42374 470154
rect 42255 470006 42321 470007
rect 42255 470002 42304 470006
rect 42368 470004 42374 470006
rect 42255 469946 42260 470002
rect 42255 469942 42304 469946
rect 42368 469944 42412 470004
rect 42368 469942 42374 469944
rect 42255 469941 42321 469942
rect 41914 469560 41920 469562
rect 41568 469500 41920 469560
rect 41914 469498 41920 469500
rect 41984 469498 41990 469562
rect 40570 469350 40576 469414
rect 40640 469350 40646 469414
rect 40578 468938 40638 469350
rect 42351 468672 42417 468675
rect 41568 468670 42417 468672
rect 41568 468614 42356 468670
rect 42412 468614 42417 468670
rect 41568 468612 42417 468614
rect 42351 468609 42417 468612
rect 42106 468080 42112 468082
rect 41568 468020 42112 468080
rect 42106 468018 42112 468020
rect 42176 468018 42182 468082
rect 41722 467488 41728 467490
rect 41568 467428 41728 467488
rect 41722 467426 41728 467428
rect 41792 467426 41798 467490
rect 40954 467278 40960 467342
rect 41024 467278 41030 467342
rect 40962 467088 41022 467278
rect 41338 466834 41344 466898
rect 41408 466834 41414 466898
rect 41346 466570 41406 466834
rect 41146 466242 41152 466306
rect 41216 466242 41222 466306
rect 41154 465978 41214 466242
rect 40762 465798 40768 465862
rect 40832 465798 40838 465862
rect 40770 465608 40830 465798
rect 42682 465120 42688 465122
rect 41568 465060 42688 465120
rect 42682 465058 42688 465060
rect 42752 465058 42758 465122
rect 34434 464383 34494 464498
rect 34434 464378 34545 464383
rect 34434 464322 34484 464378
rect 34540 464322 34545 464378
rect 34434 464320 34545 464322
rect 34479 464317 34545 464320
rect 23106 463791 23166 464054
rect 23055 463786 23166 463791
rect 23055 463730 23060 463786
rect 23116 463730 23166 463786
rect 23055 463728 23166 463730
rect 23055 463725 23121 463728
rect 41775 463640 41841 463643
rect 41568 463638 41841 463640
rect 41568 463582 41780 463638
rect 41836 463582 41841 463638
rect 41568 463580 41841 463582
rect 41775 463577 41841 463580
rect 23055 463344 23121 463347
rect 23055 463342 23166 463344
rect 23055 463286 23060 463342
rect 23116 463286 23166 463342
rect 23055 463281 23166 463286
rect 23106 463018 23166 463281
rect 41538 428539 41598 428654
rect 41538 428534 41649 428539
rect 41538 428478 41588 428534
rect 41644 428478 41649 428534
rect 41538 428476 41649 428478
rect 41583 428473 41649 428476
rect 41775 428166 41841 428169
rect 41568 428164 41841 428166
rect 41568 428108 41780 428164
rect 41836 428108 41841 428164
rect 41568 428106 41841 428108
rect 41775 428103 41841 428106
rect 41775 427648 41841 427651
rect 41568 427646 41841 427648
rect 41568 427590 41780 427646
rect 41836 427590 41841 427646
rect 41568 427588 41841 427590
rect 41775 427585 41841 427588
rect 40386 426911 40446 427174
rect 40335 426906 40446 426911
rect 40335 426850 40340 426906
rect 40396 426850 40446 426906
rect 40335 426848 40446 426850
rect 40335 426845 40401 426848
rect 41775 426612 41841 426615
rect 41568 426610 41841 426612
rect 41568 426554 41780 426610
rect 41836 426554 41841 426610
rect 41568 426552 41841 426554
rect 41775 426549 41841 426552
rect 34242 425875 34302 426138
rect 34242 425870 34353 425875
rect 34242 425814 34292 425870
rect 34348 425814 34353 425870
rect 34242 425812 34353 425814
rect 34287 425809 34353 425812
rect 41538 425431 41598 425694
rect 41538 425426 41649 425431
rect 41538 425370 41588 425426
rect 41644 425370 41649 425426
rect 41538 425368 41649 425370
rect 41583 425365 41649 425368
rect 25839 424984 25905 424987
rect 25794 424982 25905 424984
rect 25794 424926 25844 424982
rect 25900 424926 25905 424982
rect 25794 424921 25905 424926
rect 25794 424584 25854 424921
rect 34434 424839 34494 425102
rect 34434 424834 34545 424839
rect 34434 424778 34484 424834
rect 34540 424778 34545 424834
rect 34434 424776 34545 424778
rect 34479 424773 34545 424776
rect 40578 423950 40638 424214
rect 40570 423886 40576 423950
rect 40640 423886 40646 423950
rect 34242 423504 34302 423622
rect 34383 423504 34449 423507
rect 41722 423504 41728 423506
rect 34242 423502 34449 423504
rect 34242 423446 34388 423502
rect 34444 423446 34449 423502
rect 34242 423444 34449 423446
rect 34383 423441 34449 423444
rect 34530 423444 41728 423504
rect 34530 423359 34590 423444
rect 41722 423442 41728 423444
rect 41792 423442 41798 423506
rect 34479 423354 34590 423359
rect 34479 423298 34484 423354
rect 34540 423298 34590 423354
rect 34479 423296 34590 423298
rect 34479 423293 34545 423296
rect 40770 422914 40830 423104
rect 40762 422850 40768 422914
rect 40832 422850 40838 422914
rect 40962 422470 41022 422734
rect 40954 422406 40960 422470
rect 41024 422406 41030 422470
rect 42106 422172 42112 422174
rect 41568 422112 42112 422172
rect 42106 422110 42112 422112
rect 42176 422110 42182 422174
rect 42255 421580 42321 421583
rect 41568 421578 42321 421580
rect 41568 421522 42260 421578
rect 42316 421522 42321 421578
rect 41568 421520 42321 421522
rect 42255 421517 42321 421520
rect 41154 420990 41214 421180
rect 41146 420926 41152 420990
rect 41216 420926 41222 420990
rect 34287 420840 34353 420843
rect 41914 420840 41920 420842
rect 34287 420838 41920 420840
rect 34287 420782 34292 420838
rect 34348 420782 41920 420838
rect 34287 420780 41920 420782
rect 34287 420777 34353 420780
rect 41914 420778 41920 420780
rect 41984 420778 41990 420842
rect 40002 420399 40062 420662
rect 39951 420394 40062 420399
rect 39951 420338 39956 420394
rect 40012 420338 40062 420394
rect 39951 420336 40062 420338
rect 39951 420333 40017 420336
rect 39810 419955 39870 420070
rect 39810 419950 39921 419955
rect 39810 419894 39860 419950
rect 39916 419894 39921 419950
rect 39810 419892 39921 419894
rect 39855 419889 39921 419892
rect 40194 419511 40254 419700
rect 40143 419506 40254 419511
rect 40143 419450 40148 419506
rect 40204 419450 40254 419506
rect 40143 419448 40254 419450
rect 40143 419445 40209 419448
rect 41538 418919 41598 419182
rect 41538 418914 41649 418919
rect 41538 418858 41588 418914
rect 41644 418858 41649 418914
rect 41538 418856 41649 418858
rect 41583 418853 41649 418856
rect 41775 418620 41841 418623
rect 41568 418618 41841 418620
rect 41568 418562 41780 418618
rect 41836 418562 41841 418618
rect 41568 418560 41841 418562
rect 41775 418557 41841 418560
rect 41538 418031 41598 418146
rect 41538 418026 41649 418031
rect 41538 417970 41588 418026
rect 41644 417970 41649 418026
rect 41538 417968 41649 417970
rect 41583 417965 41649 417968
rect 42543 417732 42609 417735
rect 41568 417730 42609 417732
rect 41568 417674 42548 417730
rect 42604 417674 42609 417730
rect 41568 417672 42609 417674
rect 42543 417669 42609 417672
rect 41775 417140 41841 417143
rect 41568 417138 41841 417140
rect 41568 417082 41780 417138
rect 41836 417082 41841 417138
rect 41568 417080 41841 417082
rect 41775 417077 41841 417080
rect 23106 416403 23166 416666
rect 23055 416398 23166 416403
rect 23055 416342 23060 416398
rect 23116 416342 23166 416398
rect 23055 416340 23166 416342
rect 23055 416337 23121 416340
rect 41775 416178 41841 416181
rect 41568 416176 41841 416178
rect 41568 416120 41780 416176
rect 41836 416120 41841 416176
rect 41568 416118 41841 416120
rect 41775 416115 41841 416118
rect 23055 415956 23121 415959
rect 23055 415954 23166 415956
rect 23055 415898 23060 415954
rect 23116 415898 23166 415954
rect 23055 415893 23166 415898
rect 23106 415630 23166 415893
rect 42063 406070 42129 406071
rect 42063 406066 42112 406070
rect 42176 406068 42182 406070
rect 42063 406010 42068 406066
rect 42063 406006 42112 406010
rect 42176 406008 42220 406068
rect 42176 406006 42182 406008
rect 42063 406005 42129 406006
rect 58479 404144 58545 404147
rect 58479 404142 64638 404144
rect 58479 404086 58484 404142
rect 58540 404086 64638 404142
rect 58479 404084 64638 404086
rect 58479 404081 58545 404084
rect 64578 403550 64638 404084
rect 58767 402960 58833 402963
rect 58767 402958 64638 402960
rect 58767 402902 58772 402958
rect 58828 402902 64638 402958
rect 58767 402900 64638 402902
rect 58767 402897 58833 402900
rect 64578 402368 64638 402900
rect 676143 402368 676209 402371
rect 676290 402368 676350 402634
rect 676143 402366 676350 402368
rect 676143 402310 676148 402366
rect 676204 402310 676350 402366
rect 676143 402308 676350 402310
rect 676143 402305 676209 402308
rect 40954 402010 40960 402074
rect 41024 402072 41030 402074
rect 41775 402072 41841 402075
rect 41024 402070 41841 402072
rect 41024 402014 41780 402070
rect 41836 402014 41841 402070
rect 41024 402012 41841 402014
rect 41024 402010 41030 402012
rect 41775 402009 41841 402012
rect 676290 401927 676350 402116
rect 676239 401922 676350 401927
rect 676239 401866 676244 401922
rect 676300 401866 676350 401922
rect 676239 401864 676350 401866
rect 676239 401861 676305 401864
rect 676047 401628 676113 401631
rect 676047 401626 676320 401628
rect 676047 401570 676052 401626
rect 676108 401570 676320 401626
rect 676047 401568 676320 401570
rect 676047 401565 676113 401568
rect 57615 400592 57681 400595
rect 64578 400592 64638 401186
rect 676674 401039 676734 401154
rect 676674 401034 676785 401039
rect 676674 400978 676724 401034
rect 676780 400978 676785 401034
rect 676674 400976 676785 400978
rect 676719 400973 676785 400976
rect 675951 400666 676017 400669
rect 675951 400664 676320 400666
rect 675951 400608 675956 400664
rect 676012 400608 676320 400664
rect 675951 400606 676320 400608
rect 675951 400603 676017 400606
rect 57615 400590 64638 400592
rect 57615 400534 57620 400590
rect 57676 400534 64638 400590
rect 57615 400532 64638 400534
rect 57615 400529 57681 400532
rect 676239 400296 676305 400299
rect 676239 400294 676350 400296
rect 676239 400238 676244 400294
rect 676300 400238 676350 400294
rect 676239 400233 676350 400238
rect 40570 400086 40576 400150
rect 40640 400148 40646 400150
rect 41775 400148 41841 400151
rect 40640 400146 41841 400148
rect 40640 400090 41780 400146
rect 41836 400090 41841 400146
rect 676290 400118 676350 400233
rect 40640 400088 41841 400090
rect 40640 400086 40646 400088
rect 41775 400085 41841 400088
rect 58767 400000 58833 400003
rect 64578 400000 64638 400004
rect 58767 399998 64638 400000
rect 58767 399942 58772 399998
rect 58828 399942 64638 399998
rect 58767 399940 64638 399942
rect 58767 399937 58833 399940
rect 673978 399642 673984 399706
rect 674048 399704 674054 399706
rect 674048 399644 676320 399704
rect 674048 399642 674054 399644
rect 41146 399494 41152 399558
rect 41216 399556 41222 399558
rect 41775 399556 41841 399559
rect 41216 399554 41841 399556
rect 41216 399498 41780 399554
rect 41836 399498 41841 399554
rect 41216 399496 41841 399498
rect 41216 399494 41222 399496
rect 41775 399493 41841 399496
rect 58191 399408 58257 399411
rect 58191 399406 64638 399408
rect 58191 399350 58196 399406
rect 58252 399350 64638 399406
rect 58191 399348 64638 399350
rect 58191 399345 58257 399348
rect 64578 398822 64638 399348
rect 676047 399112 676113 399115
rect 676047 399110 676320 399112
rect 676047 399054 676052 399110
rect 676108 399054 676320 399110
rect 676047 399052 676320 399054
rect 676047 399049 676113 399052
rect 40762 398754 40768 398818
rect 40832 398816 40838 398818
rect 41775 398816 41841 398819
rect 40832 398814 41841 398816
rect 40832 398758 41780 398814
rect 41836 398758 41841 398814
rect 40832 398756 41841 398758
rect 40832 398754 40838 398756
rect 41775 398753 41841 398756
rect 675706 398606 675712 398670
rect 675776 398668 675782 398670
rect 675776 398608 676320 398668
rect 675776 398606 675782 398608
rect 59727 398224 59793 398227
rect 59727 398222 64638 398224
rect 59727 398166 59732 398222
rect 59788 398166 64638 398222
rect 59727 398164 64638 398166
rect 59727 398161 59793 398164
rect 64578 397640 64638 398164
rect 676290 397930 676350 398194
rect 676282 397866 676288 397930
rect 676352 397866 676358 397930
rect 674362 397570 674368 397634
rect 674432 397632 674438 397634
rect 674432 397572 676320 397632
rect 674432 397570 674438 397572
rect 675567 397040 675633 397043
rect 676290 397040 676350 397084
rect 675567 397038 676350 397040
rect 675567 396982 675572 397038
rect 675628 396982 676350 397038
rect 675567 396980 676350 396982
rect 675567 396977 675633 396980
rect 676290 396450 676350 396714
rect 676282 396386 676288 396450
rect 676352 396386 676358 396450
rect 676674 395858 676734 396122
rect 676666 395794 676672 395858
rect 676736 395794 676742 395858
rect 676090 395350 676096 395414
rect 676160 395412 676166 395414
rect 676290 395412 676350 395604
rect 676160 395352 676350 395412
rect 676160 395350 676166 395352
rect 675279 395264 675345 395267
rect 675279 395262 676320 395264
rect 675279 395206 675284 395262
rect 675340 395206 676320 395262
rect 675279 395204 676320 395206
rect 675279 395201 675345 395204
rect 675322 394610 675328 394674
rect 675392 394672 675398 394674
rect 675392 394612 676320 394672
rect 675392 394610 675398 394612
rect 676290 393935 676350 394050
rect 676239 393930 676350 393935
rect 676239 393874 676244 393930
rect 676300 393874 676350 393930
rect 676239 393872 676350 393874
rect 676239 393869 676305 393872
rect 674746 393278 674752 393342
rect 674816 393340 674822 393342
rect 676290 393340 676350 393680
rect 674816 393280 676350 393340
rect 674816 393278 674822 393280
rect 675514 393130 675520 393194
rect 675584 393192 675590 393194
rect 675584 393132 676320 393192
rect 675584 393130 675590 393132
rect 676290 392455 676350 392570
rect 676239 392450 676350 392455
rect 676239 392394 676244 392450
rect 676300 392394 676350 392450
rect 676239 392392 676350 392394
rect 676239 392389 676305 392392
rect 675898 392168 675904 392232
rect 675968 392230 675974 392232
rect 675968 392170 676320 392230
rect 675968 392168 675974 392170
rect 675130 391650 675136 391714
rect 675200 391712 675206 391714
rect 675200 391652 676320 391712
rect 675200 391650 675206 391652
rect 679746 390975 679806 391090
rect 679746 390970 679857 390975
rect 679746 390914 679796 390970
rect 679852 390914 679857 390970
rect 679746 390912 679857 390914
rect 679791 390909 679857 390912
rect 685506 390383 685566 390646
rect 679791 390380 679857 390383
rect 679746 390378 679857 390380
rect 679746 390322 679796 390378
rect 679852 390322 679857 390378
rect 679746 390317 679857 390322
rect 685455 390378 685566 390383
rect 685455 390322 685460 390378
rect 685516 390322 685566 390378
rect 685455 390320 685566 390322
rect 685455 390317 685521 390320
rect 679746 390202 679806 390317
rect 685455 389936 685521 389939
rect 685455 389934 685566 389936
rect 685455 389878 685460 389934
rect 685516 389878 685566 389934
rect 685455 389873 685566 389878
rect 685506 389610 685566 389873
rect 41775 388142 41841 388145
rect 41914 388142 41920 388144
rect 41775 388140 41920 388142
rect 41775 388084 41780 388140
rect 41836 388084 41920 388140
rect 41775 388082 41920 388084
rect 41775 388079 41841 388082
rect 41914 388080 41920 388082
rect 41984 388080 41990 388144
rect 41775 386088 41841 386091
rect 62703 386088 62769 386091
rect 41775 386086 62769 386088
rect 41538 385943 41598 386058
rect 41775 386030 41780 386086
rect 41836 386030 62708 386086
rect 62764 386030 62769 386086
rect 41775 386028 62769 386030
rect 41775 386025 41841 386028
rect 62703 386025 62769 386028
rect 41538 385938 41649 385943
rect 41538 385882 41588 385938
rect 41644 385882 41649 385938
rect 41538 385880 41649 385882
rect 41583 385877 41649 385880
rect 41538 385351 41598 385466
rect 41538 385346 41649 385351
rect 41538 385290 41588 385346
rect 41644 385290 41649 385346
rect 41538 385288 41649 385290
rect 41583 385285 41649 385288
rect 41871 385052 41937 385055
rect 41568 385050 41937 385052
rect 41568 384994 41876 385050
rect 41932 384994 41937 385050
rect 41568 384992 41937 384994
rect 41871 384989 41937 384992
rect 41583 384756 41649 384759
rect 41538 384754 41649 384756
rect 41538 384698 41588 384754
rect 41644 384698 41649 384754
rect 41538 384693 41649 384698
rect 675759 384756 675825 384759
rect 676474 384756 676480 384758
rect 675759 384754 676480 384756
rect 675759 384698 675764 384754
rect 675820 384698 676480 384754
rect 675759 384696 676480 384698
rect 675759 384693 675825 384696
rect 676474 384694 676480 384696
rect 676544 384694 676550 384758
rect 41538 384578 41598 384693
rect 41538 383871 41598 383986
rect 41538 383866 41649 383871
rect 41538 383810 41588 383866
rect 41644 383810 41649 383866
rect 41538 383808 41649 383810
rect 41583 383805 41649 383808
rect 34434 383279 34494 383542
rect 34434 383274 34545 383279
rect 34434 383218 34484 383274
rect 34540 383218 34545 383274
rect 34434 383216 34545 383218
rect 34479 383213 34545 383216
rect 41722 383214 41728 383278
rect 41792 383276 41798 383278
rect 41871 383276 41937 383279
rect 62895 383276 62961 383279
rect 41792 383274 62961 383276
rect 41792 383218 41876 383274
rect 41932 383218 62900 383274
rect 62956 383218 62961 383274
rect 41792 383216 62961 383218
rect 41792 383214 41798 383216
rect 41871 383213 41937 383216
rect 62895 383213 62961 383216
rect 41775 383128 41841 383131
rect 41568 383126 41841 383128
rect 41568 383070 41780 383126
rect 41836 383070 41841 383126
rect 41568 383068 41841 383070
rect 41775 383065 41841 383068
rect 675759 382980 675825 382983
rect 676282 382980 676288 382982
rect 675759 382978 676288 382980
rect 675759 382922 675764 382978
rect 675820 382922 676288 382978
rect 675759 382920 676288 382922
rect 675759 382917 675825 382920
rect 676282 382918 676288 382920
rect 676352 382918 676358 382982
rect 41538 382391 41598 382506
rect 41538 382386 41649 382391
rect 41538 382330 41588 382386
rect 41644 382330 41649 382386
rect 41538 382328 41649 382330
rect 41583 382325 41649 382328
rect 675322 382326 675328 382390
rect 675392 382388 675398 382390
rect 675471 382388 675537 382391
rect 675392 382386 675537 382388
rect 675392 382330 675476 382386
rect 675532 382330 675537 382386
rect 675392 382328 675537 382330
rect 675392 382326 675398 382328
rect 675471 382325 675537 382328
rect 41871 382018 41937 382021
rect 41568 382016 41937 382018
rect 41568 381960 41876 382016
rect 41932 381960 41937 382016
rect 41568 381958 41937 381960
rect 41871 381955 41937 381958
rect 40578 381354 40638 381618
rect 40570 381290 40576 381354
rect 40640 381290 40646 381354
rect 40002 380911 40062 381026
rect 39951 380906 40062 380911
rect 39951 380850 39956 380906
rect 40012 380850 40062 380906
rect 39951 380848 40062 380850
rect 39951 380845 40017 380848
rect 40770 380318 40830 380434
rect 40762 380254 40768 380318
rect 40832 380254 40838 380318
rect 41346 379726 41406 380138
rect 41338 379662 41344 379726
rect 41408 379662 41414 379726
rect 41775 379576 41841 379579
rect 41568 379574 41841 379576
rect 41568 379518 41780 379574
rect 41836 379518 41841 379574
rect 41568 379516 41841 379518
rect 41775 379513 41841 379516
rect 37359 379280 37425 379283
rect 37314 379278 37425 379280
rect 37314 379222 37364 379278
rect 37420 379222 37425 379278
rect 37314 379217 37425 379222
rect 37314 378954 37374 379217
rect 34479 378836 34545 378839
rect 41722 378836 41728 378838
rect 34479 378834 41728 378836
rect 34479 378778 34484 378834
rect 34540 378778 41728 378834
rect 34479 378776 41728 378778
rect 34479 378773 34545 378776
rect 41722 378774 41728 378776
rect 41792 378774 41798 378838
rect 675759 378836 675825 378839
rect 676666 378836 676672 378838
rect 675759 378834 676672 378836
rect 675759 378778 675764 378834
rect 675820 378778 676672 378834
rect 675759 378776 676672 378778
rect 675759 378773 675825 378776
rect 676666 378774 676672 378776
rect 676736 378774 676742 378838
rect 40962 378246 41022 378584
rect 40954 378182 40960 378246
rect 41024 378182 41030 378246
rect 675759 378096 675825 378099
rect 675898 378096 675904 378098
rect 675759 378094 675904 378096
rect 41154 377802 41214 378066
rect 675759 378038 675764 378094
rect 675820 378038 675904 378094
rect 675759 378036 675904 378038
rect 675759 378033 675825 378036
rect 675898 378034 675904 378036
rect 675968 378034 675974 378098
rect 41146 377738 41152 377802
rect 41216 377738 41222 377802
rect 41538 377359 41598 377474
rect 41538 377354 41649 377359
rect 41538 377298 41588 377354
rect 41644 377298 41649 377354
rect 41538 377296 41649 377298
rect 41583 377293 41649 377296
rect 675471 377210 675537 377211
rect 675471 377206 675520 377210
rect 675584 377208 675590 377210
rect 675471 377150 675476 377206
rect 675471 377146 675520 377150
rect 675584 377148 675628 377208
rect 675584 377146 675590 377148
rect 675471 377145 675537 377146
rect 41538 377060 41598 377104
rect 42447 377060 42513 377063
rect 41538 377058 42513 377060
rect 41538 377002 42452 377058
rect 42508 377002 42513 377058
rect 41538 377000 42513 377002
rect 42447 376997 42513 377000
rect 41538 376323 41598 376586
rect 675183 376470 675249 376471
rect 675130 376468 675136 376470
rect 675092 376408 675136 376468
rect 675200 376466 675249 376470
rect 675244 376410 675249 376466
rect 675130 376406 675136 376408
rect 675200 376406 675249 376410
rect 675183 376405 675249 376406
rect 41487 376318 41598 376323
rect 41487 376262 41492 376318
rect 41548 376262 41598 376318
rect 41487 376260 41598 376262
rect 41487 376257 41553 376260
rect 41775 376024 41841 376027
rect 41568 376022 41841 376024
rect 41568 375966 41780 376022
rect 41836 375966 41841 376022
rect 41568 375964 41841 375966
rect 41775 375961 41841 375964
rect 674746 375666 674752 375730
rect 674816 375728 674822 375730
rect 675471 375728 675537 375731
rect 674816 375726 675537 375728
rect 674816 375670 675476 375726
rect 675532 375670 675537 375726
rect 674816 375668 675537 375670
rect 674816 375666 674822 375668
rect 675471 375665 675537 375668
rect 41538 375432 41598 375550
rect 41679 375432 41745 375435
rect 41538 375430 41745 375432
rect 41538 375374 41684 375430
rect 41740 375374 41745 375430
rect 41538 375372 41745 375374
rect 41679 375369 41745 375372
rect 41538 374843 41598 375106
rect 41538 374838 41649 374843
rect 41538 374782 41588 374838
rect 41644 374782 41649 374838
rect 41538 374780 41649 374782
rect 41583 374777 41649 374780
rect 41568 374484 41790 374544
rect 28866 373807 28926 374070
rect 41730 373952 41790 374484
rect 655311 374396 655377 374399
rect 28815 373802 28926 373807
rect 28815 373746 28820 373802
rect 28876 373746 28926 373802
rect 28815 373744 28926 373746
rect 41538 373892 41790 373952
rect 649986 374394 655377 374396
rect 649986 374338 655316 374394
rect 655372 374338 655377 374394
rect 649986 374336 655377 374338
rect 649986 373892 650046 374336
rect 655311 374333 655377 374336
rect 674362 374334 674368 374398
rect 674432 374396 674438 374398
rect 675087 374396 675153 374399
rect 674432 374394 675153 374396
rect 674432 374338 675092 374394
rect 675148 374338 675153 374394
rect 674432 374336 675153 374338
rect 674432 374334 674438 374336
rect 675087 374333 675153 374336
rect 28815 373741 28881 373744
rect 41538 373363 41598 373892
rect 28815 373360 28881 373363
rect 28815 373358 28926 373360
rect 28815 373302 28820 373358
rect 28876 373302 28926 373358
rect 28815 373297 28926 373302
rect 41538 373358 41649 373363
rect 655119 373360 655185 373363
rect 41538 373302 41588 373358
rect 41644 373302 41649 373358
rect 41538 373300 41649 373302
rect 41583 373297 41649 373300
rect 649986 373358 655185 373360
rect 649986 373302 655124 373358
rect 655180 373302 655185 373358
rect 649986 373300 655185 373302
rect 28866 373034 28926 373297
rect 649986 372710 650046 373300
rect 655119 373297 655185 373300
rect 655503 372176 655569 372179
rect 649986 372174 655569 372176
rect 649986 372118 655508 372174
rect 655564 372118 655569 372174
rect 649986 372116 655569 372118
rect 649986 371528 650046 372116
rect 655503 372113 655569 372116
rect 675759 372028 675825 372031
rect 676090 372028 676096 372030
rect 675759 372026 676096 372028
rect 675759 371970 675764 372026
rect 675820 371970 676096 372026
rect 675759 371968 676096 371970
rect 675759 371965 675825 371968
rect 676090 371966 676096 371968
rect 676160 371966 676166 372030
rect 656559 370992 656625 370995
rect 649986 370990 656625 370992
rect 649986 370934 656564 370990
rect 656620 370934 656625 370990
rect 649986 370932 656625 370934
rect 649986 370346 650046 370932
rect 656559 370929 656625 370932
rect 58479 360928 58545 360931
rect 58479 360926 64638 360928
rect 58479 360870 58484 360926
rect 58540 360870 64638 360926
rect 58479 360868 64638 360870
rect 58479 360865 58545 360868
rect 64578 360328 64638 360868
rect 59151 359744 59217 359747
rect 59151 359742 64638 359744
rect 59151 359686 59156 359742
rect 59212 359686 64638 359742
rect 59151 359684 64638 359686
rect 59151 359681 59217 359684
rect 41146 359238 41152 359302
rect 41216 359300 41222 359302
rect 41775 359300 41841 359303
rect 41216 359298 41841 359300
rect 41216 359242 41780 359298
rect 41836 359242 41841 359298
rect 41216 359240 41841 359242
rect 41216 359238 41222 359240
rect 41775 359237 41841 359240
rect 64578 359146 64638 359684
rect 41338 358794 41344 358858
rect 41408 358856 41414 358858
rect 41775 358856 41841 358859
rect 41408 358854 41841 358856
rect 41408 358798 41780 358854
rect 41836 358798 41841 358854
rect 41408 358796 41841 358798
rect 41408 358794 41414 358796
rect 41775 358793 41841 358796
rect 676143 358116 676209 358119
rect 676290 358116 676350 358234
rect 676143 358114 676350 358116
rect 676143 358058 676148 358114
rect 676204 358058 676350 358114
rect 676143 358056 676350 358058
rect 676143 358053 676209 358056
rect 57615 357524 57681 357527
rect 64578 357524 64638 357964
rect 57615 357522 64638 357524
rect 57615 357466 57620 357522
rect 57676 357466 64638 357522
rect 57615 357464 64638 357466
rect 57615 357461 57681 357464
rect 676290 357379 676350 357716
rect 676239 357374 676350 357379
rect 676239 357318 676244 357374
rect 676300 357318 676350 357374
rect 676239 357316 676350 357318
rect 676239 357313 676305 357316
rect 676047 357228 676113 357231
rect 676047 357226 676320 357228
rect 676047 357170 676052 357226
rect 676108 357170 676320 357226
rect 676047 357168 676320 357170
rect 676047 357165 676113 357168
rect 40570 356870 40576 356934
rect 40640 356932 40646 356934
rect 41775 356932 41841 356935
rect 40640 356930 41841 356932
rect 40640 356874 41780 356930
rect 41836 356874 41841 356930
rect 40640 356872 41841 356874
rect 40640 356870 40646 356872
rect 41775 356869 41841 356872
rect 59631 356784 59697 356787
rect 676047 356784 676113 356787
rect 59631 356782 64638 356784
rect 59631 356726 59636 356782
rect 59692 356726 64638 356782
rect 59631 356724 64638 356726
rect 676047 356782 676320 356784
rect 676047 356726 676052 356782
rect 676108 356726 676320 356782
rect 676047 356724 676320 356726
rect 59631 356721 59697 356724
rect 676047 356721 676113 356724
rect 40954 356426 40960 356490
rect 41024 356488 41030 356490
rect 41775 356488 41841 356491
rect 41024 356486 41841 356488
rect 41024 356430 41780 356486
rect 41836 356430 41841 356486
rect 41024 356428 41841 356430
rect 41024 356426 41030 356428
rect 41775 356425 41841 356428
rect 58191 356192 58257 356195
rect 58191 356190 64638 356192
rect 58191 356134 58196 356190
rect 58252 356134 64638 356190
rect 58191 356132 64638 356134
rect 58191 356129 58257 356132
rect 40762 355538 40768 355602
rect 40832 355600 40838 355602
rect 41775 355600 41841 355603
rect 64578 355600 64638 356132
rect 670191 356044 670257 356047
rect 673978 356044 673984 356046
rect 670191 356042 673984 356044
rect 670191 355986 670196 356042
rect 670252 355986 673984 356042
rect 670191 355984 673984 355986
rect 670191 355981 670257 355984
rect 673794 355748 673854 355984
rect 673978 355982 673984 355984
rect 674048 355982 674054 356046
rect 673978 355834 673984 355898
rect 674048 355896 674054 355898
rect 676290 355896 676350 356236
rect 674048 355836 676350 355896
rect 674048 355834 674054 355836
rect 673794 355688 676320 355748
rect 40832 355598 41841 355600
rect 40832 355542 41780 355598
rect 41836 355542 41841 355598
rect 40832 355540 41841 355542
rect 40832 355538 40838 355540
rect 41775 355537 41841 355540
rect 674170 355242 674176 355306
rect 674240 355304 674246 355306
rect 674240 355244 676320 355304
rect 674240 355242 674246 355244
rect 58575 355008 58641 355011
rect 58575 355006 64638 355008
rect 58575 354950 58580 355006
rect 58636 354950 64638 355006
rect 58575 354948 64638 354950
rect 58575 354945 58641 354948
rect 64578 354418 64638 354948
rect 669999 354712 670065 354715
rect 675706 354712 675712 354714
rect 669999 354710 675712 354712
rect 669999 354654 670004 354710
rect 670060 354654 675712 354710
rect 669999 354652 675712 354654
rect 669999 354649 670065 354652
rect 675706 354650 675712 354652
rect 675776 354712 675782 354714
rect 675776 354652 676320 354712
rect 675776 354650 675782 354652
rect 674362 354206 674368 354270
rect 674432 354268 674438 354270
rect 674432 354208 676320 354268
rect 674432 354206 674438 354208
rect 676047 353824 676113 353827
rect 676047 353822 676320 353824
rect 676047 353766 676052 353822
rect 676108 353766 676320 353822
rect 676047 353764 676320 353766
rect 676047 353761 676113 353764
rect 674554 353170 674560 353234
rect 674624 353232 674630 353234
rect 674624 353172 676320 353232
rect 674624 353170 674630 353172
rect 675567 352640 675633 352643
rect 676290 352640 676350 352684
rect 675567 352638 676350 352640
rect 675567 352582 675572 352638
rect 675628 352582 676350 352638
rect 675567 352580 676350 352582
rect 675567 352577 675633 352580
rect 676047 352344 676113 352347
rect 676047 352342 676320 352344
rect 676047 352286 676052 352342
rect 676108 352286 676320 352342
rect 676047 352284 676320 352286
rect 676047 352281 676113 352284
rect 676866 351607 676926 351722
rect 676866 351602 676977 351607
rect 676866 351546 676916 351602
rect 676972 351546 676977 351602
rect 676866 351544 676977 351546
rect 676911 351541 676977 351544
rect 674746 350950 674752 351014
rect 674816 351012 674822 351014
rect 676290 351012 676350 351204
rect 674816 350952 676350 351012
rect 674816 350950 674822 350952
rect 675279 350864 675345 350867
rect 675279 350862 676320 350864
rect 675279 350806 675284 350862
rect 675340 350806 676320 350862
rect 675279 350804 676320 350806
rect 675279 350801 675345 350804
rect 676047 350272 676113 350275
rect 676047 350270 676320 350272
rect 676047 350214 676052 350270
rect 676108 350214 676320 350270
rect 676047 350212 676320 350214
rect 676047 350209 676113 350212
rect 676290 349535 676350 349650
rect 676239 349530 676350 349535
rect 676239 349474 676244 349530
rect 676300 349474 676350 349530
rect 676239 349472 676350 349474
rect 676239 349469 676305 349472
rect 676866 349091 676926 349280
rect 676815 349086 676926 349091
rect 676815 349030 676820 349086
rect 676876 349030 676926 349086
rect 676815 349028 676926 349030
rect 676815 349025 676881 349028
rect 674938 348730 674944 348794
rect 675008 348792 675014 348794
rect 675008 348732 676320 348792
rect 675008 348730 675014 348732
rect 676290 348055 676350 348170
rect 676239 348050 676350 348055
rect 676239 347994 676244 348050
rect 676300 347994 676350 348050
rect 676239 347992 676350 347994
rect 676239 347989 676305 347992
rect 676047 347830 676113 347833
rect 676047 347828 676320 347830
rect 676047 347772 676052 347828
rect 676108 347772 676320 347828
rect 676047 347770 676320 347772
rect 676047 347767 676113 347770
rect 675951 347312 676017 347315
rect 675951 347310 676320 347312
rect 675951 347254 675956 347310
rect 676012 347254 676320 347310
rect 675951 347252 676320 347254
rect 675951 347249 676017 347252
rect 679938 346575 679998 346690
rect 679887 346570 679998 346575
rect 679887 346514 679892 346570
rect 679948 346514 679998 346570
rect 679887 346512 679998 346514
rect 679887 346509 679953 346512
rect 679746 345983 679806 346246
rect 679887 346128 679953 346131
rect 679887 346126 679998 346128
rect 679887 346070 679892 346126
rect 679948 346070 679998 346126
rect 679887 346065 679998 346070
rect 679695 345978 679806 345983
rect 679695 345922 679700 345978
rect 679756 345922 679806 345978
rect 679695 345920 679806 345922
rect 679695 345917 679761 345920
rect 679938 345802 679998 346065
rect 679695 345536 679761 345539
rect 679695 345534 679806 345536
rect 679695 345478 679700 345534
rect 679756 345478 679806 345534
rect 679695 345473 679806 345478
rect 679746 345210 679806 345473
rect 41679 343170 41745 343171
rect 41679 343168 41728 343170
rect 41600 343166 41728 343168
rect 41792 343168 41798 343170
rect 63087 343168 63153 343171
rect 41792 343166 63153 343168
rect 41600 343110 41684 343166
rect 41792 343110 63092 343166
rect 63148 343110 63153 343166
rect 41600 343108 41728 343110
rect 41679 343106 41728 343108
rect 41792 343108 63153 343110
rect 41792 343106 41798 343108
rect 41679 343105 41745 343106
rect 63087 343105 63153 343108
rect 675898 342958 675904 343022
rect 675968 343020 675974 343022
rect 676815 343020 676881 343023
rect 675968 343018 676881 343020
rect 675968 342962 676820 343018
rect 676876 342962 676881 343018
rect 675968 342960 676881 342962
rect 675968 342958 675974 342960
rect 676815 342957 676881 342960
rect 41775 342872 41841 342875
rect 41568 342870 41841 342872
rect 41568 342814 41780 342870
rect 41836 342814 41841 342870
rect 41568 342812 41841 342814
rect 41775 342809 41841 342812
rect 675706 342810 675712 342874
rect 675776 342872 675782 342874
rect 676911 342872 676977 342875
rect 675776 342870 676977 342872
rect 675776 342814 676916 342870
rect 676972 342814 676977 342870
rect 675776 342812 676977 342814
rect 675776 342810 675782 342812
rect 676911 342809 676977 342812
rect 41775 342354 41841 342357
rect 41568 342352 41841 342354
rect 41568 342296 41780 342352
rect 41836 342296 41841 342352
rect 41568 342294 41841 342296
rect 41775 342291 41841 342294
rect 41775 341836 41841 341839
rect 41568 341834 41841 341836
rect 41568 341778 41780 341834
rect 41836 341778 41841 341834
rect 41568 341776 41841 341778
rect 41775 341773 41841 341776
rect 41775 341392 41841 341395
rect 41568 341390 41841 341392
rect 41568 341334 41780 341390
rect 41836 341334 41841 341390
rect 41568 341332 41841 341334
rect 41775 341329 41841 341332
rect 41538 340655 41598 340770
rect 41538 340650 41649 340655
rect 41538 340594 41588 340650
rect 41644 340594 41649 340650
rect 41538 340592 41649 340594
rect 41583 340589 41649 340592
rect 41775 340356 41841 340359
rect 41568 340354 41841 340356
rect 41568 340298 41780 340354
rect 41836 340298 41841 340354
rect 41568 340296 41841 340298
rect 41775 340293 41841 340296
rect 41679 340060 41745 340063
rect 41538 340058 41745 340060
rect 41538 340002 41684 340058
rect 41740 340002 41745 340058
rect 41538 340000 41745 340002
rect 41538 339882 41598 340000
rect 41679 339997 41745 340000
rect 41538 339175 41598 339290
rect 41538 339170 41649 339175
rect 41538 339114 41588 339170
rect 41644 339114 41649 339170
rect 41538 339112 41649 339114
rect 41583 339109 41649 339112
rect 43119 338876 43185 338879
rect 40608 338874 43185 338876
rect 40608 338846 43124 338874
rect 40578 338818 43124 338846
rect 43180 338818 43185 338874
rect 40578 338816 43185 338818
rect 40578 338582 40638 338816
rect 43119 338813 43185 338816
rect 40570 338518 40576 338582
rect 40640 338518 40646 338582
rect 40770 338138 40830 338402
rect 40762 338074 40768 338138
rect 40832 338074 40838 338138
rect 39810 337695 39870 337810
rect 39759 337690 39870 337695
rect 39759 337634 39764 337690
rect 39820 337634 39870 337690
rect 39759 337632 39870 337634
rect 39759 337629 39825 337632
rect 40962 337102 41022 337292
rect 40954 337038 40960 337102
rect 41024 337038 41030 337102
rect 41346 336658 41406 336922
rect 41338 336594 41344 336658
rect 41408 336594 41414 336658
rect 41538 336215 41598 336330
rect 41538 336210 41649 336215
rect 41538 336154 41588 336210
rect 41644 336154 41649 336210
rect 41538 336152 41649 336154
rect 41583 336149 41649 336152
rect 41775 335768 41841 335771
rect 41568 335766 41841 335768
rect 41568 335710 41780 335766
rect 41836 335710 41841 335766
rect 41568 335708 41841 335710
rect 41775 335705 41841 335708
rect 41154 335030 41214 335442
rect 41146 334966 41152 335030
rect 41216 334966 41222 335030
rect 41538 334586 41598 334850
rect 41530 334522 41536 334586
rect 41600 334522 41606 334586
rect 41871 334288 41937 334291
rect 41568 334286 41937 334288
rect 41568 334230 41876 334286
rect 41932 334230 41937 334286
rect 41568 334228 41937 334230
rect 41871 334225 41937 334228
rect 41538 333844 41598 333888
rect 42447 333844 42513 333847
rect 41538 333842 42513 333844
rect 41538 333786 42452 333842
rect 42508 333786 42513 333842
rect 41538 333784 42513 333786
rect 42447 333781 42513 333784
rect 675759 333550 675825 333551
rect 675706 333486 675712 333550
rect 675776 333548 675825 333550
rect 675776 333546 675868 333548
rect 675820 333490 675868 333546
rect 675776 333488 675868 333490
rect 675776 333486 675825 333488
rect 675759 333485 675825 333486
rect 41538 333107 41598 333370
rect 41487 333102 41598 333107
rect 41487 333046 41492 333102
rect 41548 333046 41598 333102
rect 41487 333044 41598 333046
rect 41487 333041 41553 333044
rect 41346 332663 41406 332778
rect 41346 332658 41457 332663
rect 41346 332602 41396 332658
rect 41452 332602 41457 332658
rect 41346 332600 41457 332602
rect 41391 332597 41457 332600
rect 41538 332216 41598 332408
rect 674938 332302 674944 332366
rect 675008 332364 675014 332366
rect 675471 332364 675537 332367
rect 675008 332362 675537 332364
rect 675008 332306 675476 332362
rect 675532 332306 675537 332362
rect 675008 332304 675537 332306
rect 675008 332302 675014 332304
rect 675471 332301 675537 332304
rect 41679 332216 41745 332219
rect 41538 332214 41745 332216
rect 41538 332158 41684 332214
rect 41740 332158 41745 332214
rect 41538 332156 41745 332158
rect 41679 332153 41745 332156
rect 41538 331627 41598 331890
rect 41538 331622 41649 331627
rect 41538 331566 41588 331622
rect 41644 331566 41649 331622
rect 41538 331564 41649 331566
rect 41583 331561 41649 331564
rect 41538 331180 41598 331298
rect 41538 331120 41790 331180
rect 28866 330591 28926 330854
rect 41730 330736 41790 331120
rect 28815 330586 28926 330591
rect 28815 330530 28820 330586
rect 28876 330530 28926 330586
rect 28815 330528 28926 330530
rect 41538 330676 41790 330736
rect 28815 330525 28881 330528
rect 41538 330440 41598 330676
rect 675759 330588 675825 330591
rect 675898 330588 675904 330590
rect 675759 330586 675904 330588
rect 675759 330530 675764 330586
rect 675820 330530 675904 330586
rect 675759 330528 675904 330530
rect 675759 330525 675825 330528
rect 675898 330526 675904 330528
rect 675968 330526 675974 330590
rect 41871 330440 41937 330443
rect 41538 330438 41937 330440
rect 41538 330410 41876 330438
rect 41568 330382 41876 330410
rect 41932 330382 41937 330438
rect 41568 330380 41937 330382
rect 41871 330377 41937 330380
rect 28815 330144 28881 330147
rect 28815 330142 28926 330144
rect 28815 330086 28820 330142
rect 28876 330086 28926 330142
rect 28815 330081 28926 330086
rect 28866 329818 28926 330081
rect 655215 329848 655281 329851
rect 649986 329846 655281 329848
rect 649986 329790 655220 329846
rect 655276 329790 655281 329846
rect 649986 329788 655281 329790
rect 649986 329234 650046 329788
rect 655215 329785 655281 329788
rect 674554 328158 674560 328222
rect 674624 328220 674630 328222
rect 675087 328220 675153 328223
rect 674624 328218 675153 328220
rect 674624 328162 675092 328218
rect 675148 328162 675153 328218
rect 674624 328160 675153 328162
rect 674624 328158 674630 328160
rect 675087 328157 675153 328160
rect 655311 328072 655377 328075
rect 649986 328070 655377 328072
rect 649986 328014 655316 328070
rect 655372 328014 655377 328070
rect 649986 328012 655377 328014
rect 655311 328009 655377 328012
rect 655119 327480 655185 327483
rect 649986 327478 655185 327480
rect 649986 327422 655124 327478
rect 655180 327422 655185 327478
rect 649986 327420 655185 327422
rect 649986 326870 650046 327420
rect 655119 327417 655185 327420
rect 674746 326826 674752 326890
rect 674816 326888 674822 326890
rect 675375 326888 675441 326891
rect 674816 326886 675441 326888
rect 674816 326830 675380 326886
rect 675436 326830 675441 326886
rect 674816 326828 675441 326830
rect 674816 326826 674822 326828
rect 675375 326825 675441 326828
rect 654159 326296 654225 326299
rect 649986 326294 654225 326296
rect 649986 326238 654164 326294
rect 654220 326238 654225 326294
rect 649986 326236 654225 326238
rect 649986 325688 650046 326236
rect 654159 326233 654225 326236
rect 58479 317712 58545 317715
rect 58479 317710 64638 317712
rect 58479 317654 58484 317710
rect 58540 317654 64638 317710
rect 58479 317652 64638 317654
rect 58479 317649 58545 317652
rect 64578 317106 64638 317652
rect 59151 316528 59217 316531
rect 59151 316526 64638 316528
rect 59151 316470 59156 316526
rect 59212 316470 64638 316526
rect 59151 316468 64638 316470
rect 59151 316465 59217 316468
rect 41530 316170 41536 316234
rect 41600 316232 41606 316234
rect 41775 316232 41841 316235
rect 41600 316230 41841 316232
rect 41600 316174 41780 316230
rect 41836 316174 41841 316230
rect 41600 316172 41841 316174
rect 41600 316170 41606 316172
rect 41775 316169 41841 316172
rect 64578 315924 64638 316468
rect 41338 315430 41344 315494
rect 41408 315492 41414 315494
rect 41775 315492 41841 315495
rect 41408 315490 41841 315492
rect 41408 315434 41780 315490
rect 41836 315434 41841 315490
rect 41408 315432 41841 315434
rect 41408 315430 41414 315432
rect 41775 315429 41841 315432
rect 59151 314160 59217 314163
rect 64578 314160 64638 314742
rect 59151 314158 64638 314160
rect 59151 314102 59156 314158
rect 59212 314102 64638 314158
rect 59151 314100 64638 314102
rect 59151 314097 59217 314100
rect 59631 313864 59697 313867
rect 59631 313862 64638 313864
rect 59631 313806 59636 313862
rect 59692 313806 64638 313862
rect 59631 313804 64638 313806
rect 59631 313801 59697 313804
rect 40762 313654 40768 313718
rect 40832 313716 40838 313718
rect 41775 313716 41841 313719
rect 40832 313714 41841 313716
rect 40832 313658 41780 313714
rect 41836 313658 41841 313714
rect 40832 313656 41841 313658
rect 40832 313654 40838 313656
rect 41775 313653 41841 313656
rect 64578 313560 64638 313804
rect 41146 313210 41152 313274
rect 41216 313272 41222 313274
rect 41775 313272 41841 313275
rect 41216 313270 41841 313272
rect 41216 313214 41780 313270
rect 41836 313214 41841 313270
rect 41216 313212 41841 313214
rect 41216 313210 41222 313212
rect 41775 313209 41841 313212
rect 58863 312976 58929 312979
rect 58863 312974 64638 312976
rect 58863 312918 58868 312974
rect 58924 312918 64638 312974
rect 58863 312916 64638 312918
rect 58863 312913 58929 312916
rect 40954 312322 40960 312386
rect 41024 312384 41030 312386
rect 41775 312384 41841 312387
rect 41024 312382 41841 312384
rect 41024 312326 41780 312382
rect 41836 312326 41841 312382
rect 64578 312378 64638 312916
rect 41024 312324 41841 312326
rect 41024 312322 41030 312324
rect 41775 312321 41841 312324
rect 676290 312239 676350 312502
rect 676290 312234 676401 312239
rect 676290 312178 676340 312234
rect 676396 312178 676401 312234
rect 676290 312176 676401 312178
rect 676335 312173 676401 312176
rect 59631 311792 59697 311795
rect 59631 311790 64638 311792
rect 59631 311734 59636 311790
rect 59692 311734 64638 311790
rect 59631 311732 64638 311734
rect 59631 311729 59697 311732
rect 64578 311196 64638 311732
rect 676143 311644 676209 311647
rect 676290 311644 676350 311910
rect 676143 311642 676350 311644
rect 676143 311586 676148 311642
rect 676204 311586 676350 311642
rect 676143 311584 676350 311586
rect 676143 311581 676209 311584
rect 676290 311203 676350 311392
rect 676239 311198 676350 311203
rect 676239 311142 676244 311198
rect 676300 311142 676350 311198
rect 676239 311140 676350 311142
rect 676239 311137 676305 311140
rect 673978 310990 673984 311054
rect 674048 311052 674054 311054
rect 674048 310992 676320 311052
rect 674048 310990 674054 310992
rect 673978 310398 673984 310462
rect 674048 310460 674054 310462
rect 674048 310400 676320 310460
rect 674048 310398 674054 310400
rect 674170 309806 674176 309870
rect 674240 309868 674246 309870
rect 674240 309838 676896 309868
rect 674240 309808 676926 309838
rect 674240 309806 674246 309808
rect 676866 309722 676926 309808
rect 676858 309658 676864 309722
rect 676928 309658 676934 309722
rect 674554 309066 674560 309130
rect 674624 309128 674630 309130
rect 676290 309128 676350 309468
rect 674624 309068 676350 309128
rect 674624 309066 674630 309068
rect 670383 308980 670449 308983
rect 674362 308980 674368 308982
rect 670383 308978 674368 308980
rect 670383 308922 670388 308978
rect 670444 308922 674368 308978
rect 670383 308920 674368 308922
rect 670383 308917 670449 308920
rect 674362 308918 674368 308920
rect 674432 308980 674438 308982
rect 674432 308920 676320 308980
rect 674432 308918 674438 308920
rect 675898 308326 675904 308390
rect 675968 308388 675974 308390
rect 675968 308328 676320 308388
rect 675968 308326 675974 308328
rect 676290 307650 676350 307988
rect 676282 307586 676288 307650
rect 676352 307586 676358 307650
rect 674746 307438 674752 307502
rect 674816 307500 674822 307502
rect 674816 307440 676320 307500
rect 674816 307438 674822 307440
rect 676290 306763 676350 306878
rect 676239 306758 676350 306763
rect 676239 306702 676244 306758
rect 676300 306702 676350 306758
rect 676239 306700 676350 306702
rect 676239 306697 676305 306700
rect 675322 306402 675328 306466
rect 675392 306464 675398 306466
rect 675392 306404 676320 306464
rect 675392 306402 675398 306404
rect 675706 305958 675712 306022
rect 675776 306020 675782 306022
rect 675776 305960 676320 306020
rect 675776 305958 675782 305960
rect 674170 305366 674176 305430
rect 674240 305428 674246 305430
rect 674240 305368 676320 305428
rect 674240 305366 674246 305368
rect 676290 304839 676350 304954
rect 676239 304834 676350 304839
rect 676239 304778 676244 304834
rect 676300 304778 676350 304834
rect 676239 304776 676350 304778
rect 676239 304773 676305 304776
rect 676047 304466 676113 304469
rect 676047 304464 676320 304466
rect 676047 304408 676052 304464
rect 676108 304408 676320 304464
rect 676047 304406 676320 304408
rect 676047 304403 676113 304406
rect 675951 303948 676017 303951
rect 675951 303946 676320 303948
rect 675951 303890 675956 303946
rect 676012 303890 676320 303946
rect 675951 303888 676320 303890
rect 675951 303885 676017 303888
rect 674938 303442 674944 303506
rect 675008 303504 675014 303506
rect 675008 303444 676320 303504
rect 675008 303442 675014 303444
rect 654159 303356 654225 303359
rect 649986 303354 654225 303356
rect 649986 303298 654164 303354
rect 654220 303298 654225 303354
rect 649986 303296 654225 303298
rect 649986 302776 650046 303296
rect 654159 303293 654225 303296
rect 675130 302702 675136 302766
rect 675200 302764 675206 302766
rect 676290 302764 676350 302956
rect 675200 302704 676350 302764
rect 675200 302702 675206 302704
rect 676090 302554 676096 302618
rect 676160 302616 676166 302618
rect 676160 302556 676350 302616
rect 676160 302554 676166 302556
rect 676290 302438 676350 302556
rect 654063 302172 654129 302175
rect 649986 302170 654129 302172
rect 649986 302114 654068 302170
rect 654124 302114 654129 302170
rect 649986 302112 654129 302114
rect 649986 301594 650046 302112
rect 654063 302109 654129 302112
rect 675514 301962 675520 302026
rect 675584 302024 675590 302026
rect 675584 301964 676320 302024
rect 675584 301962 675590 301964
rect 676482 301138 676542 301402
rect 676474 301074 676480 301138
rect 676544 301074 676550 301138
rect 654255 300988 654321 300991
rect 649986 300986 654321 300988
rect 649986 300930 654260 300986
rect 654316 300930 654321 300986
rect 649986 300928 654321 300930
rect 649986 300412 650046 300928
rect 654255 300925 654321 300928
rect 679938 300695 679998 300958
rect 679938 300690 680049 300695
rect 679938 300634 679988 300690
rect 680044 300634 680049 300690
rect 679938 300632 680049 300634
rect 679983 300629 680049 300632
rect 679746 300251 679806 300514
rect 679746 300246 679857 300251
rect 679983 300248 680049 300251
rect 679746 300190 679796 300246
rect 679852 300190 679857 300246
rect 679746 300188 679857 300190
rect 679791 300185 679857 300188
rect 679938 300246 680049 300248
rect 679938 300190 679988 300246
rect 680044 300190 680049 300246
rect 679938 300185 680049 300190
rect 679938 299922 679998 300185
rect 679791 299804 679857 299807
rect 679746 299802 679857 299804
rect 679746 299746 679796 299802
rect 679852 299746 679857 299802
rect 679746 299741 679857 299746
rect 41775 299656 41841 299659
rect 41568 299654 41841 299656
rect 41568 299598 41780 299654
rect 41836 299598 41841 299654
rect 41568 299596 41841 299598
rect 41775 299593 41841 299596
rect 679746 299404 679806 299741
rect 41775 299212 41841 299215
rect 41568 299210 41841 299212
rect 41568 299154 41780 299210
rect 41836 299154 41841 299210
rect 41568 299152 41841 299154
rect 41775 299149 41841 299152
rect 39663 298768 39729 298771
rect 39618 298766 39729 298768
rect 39618 298710 39668 298766
rect 39724 298710 39729 298766
rect 39618 298705 39729 298710
rect 649986 298768 650046 299230
rect 656559 298768 656625 298771
rect 649986 298766 656625 298768
rect 649986 298710 656564 298766
rect 656620 298710 656625 298766
rect 649986 298708 656625 298710
rect 656559 298705 656625 298708
rect 39618 298590 39678 298705
rect 41775 298176 41841 298179
rect 41568 298174 41841 298176
rect 41568 298118 41780 298174
rect 41836 298118 41841 298174
rect 41568 298116 41841 298118
rect 41775 298113 41841 298116
rect 41775 297658 41841 297661
rect 41568 297656 41841 297658
rect 41568 297600 41780 297656
rect 41836 297600 41841 297656
rect 41568 297598 41841 297600
rect 41775 297595 41841 297598
rect 649986 297584 650046 298048
rect 656271 297584 656337 297587
rect 649986 297582 656337 297584
rect 649986 297526 656276 297582
rect 656332 297526 656337 297582
rect 649986 297524 656337 297526
rect 656271 297521 656337 297524
rect 41775 297140 41841 297143
rect 41568 297138 41841 297140
rect 41568 297082 41780 297138
rect 41836 297082 41841 297138
rect 41568 297080 41841 297082
rect 41775 297077 41841 297080
rect 649986 296844 650046 296866
rect 656079 296844 656145 296847
rect 649986 296842 656145 296844
rect 649986 296786 656084 296842
rect 656140 296786 656145 296842
rect 649986 296784 656145 296786
rect 656079 296781 656145 296784
rect 39810 296551 39870 296670
rect 39759 296546 39870 296551
rect 39759 296490 39764 296546
rect 39820 296490 39870 296546
rect 39759 296488 39870 296490
rect 39759 296485 39825 296488
rect 41538 295959 41598 296074
rect 39951 295956 40017 295959
rect 39951 295954 40062 295956
rect 39951 295898 39956 295954
rect 40012 295898 40062 295954
rect 39951 295893 40062 295898
rect 41538 295954 41649 295959
rect 41538 295898 41588 295954
rect 41644 295898 41649 295954
rect 41538 295896 41649 295898
rect 41583 295893 41649 295896
rect 40002 295630 40062 295893
rect 59343 295216 59409 295219
rect 64578 295216 64638 295684
rect 59343 295214 64638 295216
rect 40962 294922 41022 295186
rect 59343 295158 59348 295214
rect 59404 295158 64638 295214
rect 59343 295156 64638 295158
rect 649986 295216 650046 295684
rect 656367 295216 656433 295219
rect 649986 295214 656433 295216
rect 649986 295158 656372 295214
rect 656428 295158 656433 295214
rect 649986 295156 656433 295158
rect 59343 295153 59409 295156
rect 656367 295153 656433 295156
rect 40954 294858 40960 294922
rect 41024 294858 41030 294922
rect 675759 294624 675825 294627
rect 676282 294624 676288 294626
rect 675759 294622 676288 294624
rect 40194 294479 40254 294594
rect 675759 294566 675764 294622
rect 675820 294566 676288 294622
rect 675759 294564 676288 294566
rect 675759 294561 675825 294564
rect 676282 294562 676288 294564
rect 676352 294562 676358 294626
rect 40194 294474 40305 294479
rect 40194 294418 40244 294474
rect 40300 294418 40305 294474
rect 40194 294416 40305 294418
rect 40239 294413 40305 294416
rect 40770 293886 40830 294150
rect 59247 294032 59313 294035
rect 64578 294032 64638 294502
rect 59247 294030 64638 294032
rect 59247 293974 59252 294030
rect 59308 293974 64638 294030
rect 59247 293972 64638 293974
rect 649986 294032 650046 294502
rect 655887 294032 655953 294035
rect 649986 294030 655953 294032
rect 649986 293974 655892 294030
rect 655948 293974 655953 294030
rect 649986 293972 655953 293974
rect 59247 293969 59313 293972
rect 655887 293969 655953 293972
rect 40762 293822 40768 293886
rect 40832 293822 40838 293886
rect 41538 293442 41598 293706
rect 41530 293378 41536 293442
rect 41600 293378 41606 293442
rect 41538 292999 41598 293114
rect 41538 292994 41649 292999
rect 41538 292938 41588 292994
rect 41644 292938 41649 292994
rect 41538 292936 41649 292938
rect 41583 292933 41649 292936
rect 59439 292848 59505 292851
rect 64578 292848 64638 293320
rect 59439 292846 64638 292848
rect 59439 292790 59444 292846
rect 59500 292790 64638 292846
rect 59439 292788 64638 292790
rect 649986 292848 650046 293320
rect 655791 292848 655857 292851
rect 675375 292850 675441 292851
rect 675322 292848 675328 292850
rect 649986 292846 655857 292848
rect 649986 292790 655796 292846
rect 655852 292790 655857 292846
rect 649986 292788 655857 292790
rect 675284 292788 675328 292848
rect 675392 292846 675441 292850
rect 675436 292790 675441 292846
rect 59439 292785 59505 292788
rect 655791 292785 655857 292788
rect 675322 292786 675328 292788
rect 675392 292786 675441 292790
rect 675375 292785 675441 292786
rect 58191 292700 58257 292703
rect 58191 292698 64638 292700
rect 58191 292642 58196 292698
rect 58252 292642 64638 292698
rect 58191 292640 64638 292642
rect 58191 292637 58257 292640
rect 41775 292626 41841 292629
rect 41568 292624 41841 292626
rect 41568 292568 41780 292624
rect 41836 292568 41841 292624
rect 41568 292566 41841 292568
rect 41775 292563 41841 292566
rect 41154 291962 41214 292226
rect 64578 292138 64638 292640
rect 41146 291898 41152 291962
rect 41216 291898 41222 291962
rect 649986 291664 650046 292138
rect 656175 291664 656241 291667
rect 649986 291662 656241 291664
rect 41346 291370 41406 291634
rect 649986 291606 656180 291662
rect 656236 291606 656241 291662
rect 649986 291604 656241 291606
rect 656175 291601 656241 291604
rect 59631 291516 59697 291519
rect 59631 291514 64638 291516
rect 59631 291458 59636 291514
rect 59692 291458 64638 291514
rect 59631 291456 64638 291458
rect 59631 291453 59697 291456
rect 41338 291306 41344 291370
rect 41408 291306 41414 291370
rect 41538 290927 41598 291042
rect 64578 290956 64638 291456
rect 41538 290922 41649 290927
rect 41538 290866 41588 290922
rect 41644 290866 41649 290922
rect 41538 290864 41649 290866
rect 649986 290924 650046 290956
rect 655983 290924 656049 290927
rect 649986 290922 656049 290924
rect 649986 290866 655988 290922
rect 656044 290866 656049 290922
rect 649986 290864 656049 290866
rect 41583 290861 41649 290864
rect 655983 290861 656049 290864
rect 42351 290776 42417 290779
rect 41568 290774 42417 290776
rect 41568 290718 42356 290774
rect 42412 290718 42417 290774
rect 41568 290716 42417 290718
rect 42351 290713 42417 290716
rect 675759 290776 675825 290779
rect 676090 290776 676096 290778
rect 675759 290774 676096 290776
rect 675759 290718 675764 290774
rect 675820 290718 676096 290774
rect 675759 290716 676096 290718
rect 675759 290713 675825 290716
rect 676090 290714 676096 290716
rect 676160 290714 676166 290778
rect 42543 290184 42609 290187
rect 41568 290182 42609 290184
rect 41568 290126 42548 290182
rect 42604 290126 42609 290182
rect 41568 290124 42609 290126
rect 42543 290121 42609 290124
rect 41538 289447 41598 289562
rect 41487 289442 41598 289447
rect 41487 289386 41492 289442
rect 41548 289386 41598 289442
rect 41487 289384 41598 289386
rect 41487 289381 41553 289384
rect 58863 289296 58929 289299
rect 64578 289296 64638 289774
rect 58863 289294 64638 289296
rect 58863 289238 58868 289294
rect 58924 289238 64638 289294
rect 58863 289236 64638 289238
rect 649986 289296 650046 289774
rect 655599 289296 655665 289299
rect 649986 289294 655665 289296
rect 649986 289238 655604 289294
rect 655660 289238 655665 289294
rect 649986 289236 655665 289238
rect 58863 289233 58929 289236
rect 655599 289233 655665 289236
rect 41538 289003 41598 289192
rect 41538 288998 41649 289003
rect 41538 288942 41588 288998
rect 41644 288942 41649 288998
rect 41538 288940 41649 288942
rect 41583 288937 41649 288940
rect 42255 288704 42321 288707
rect 41568 288702 42321 288704
rect 41568 288646 42260 288702
rect 42316 288646 42321 288702
rect 41568 288644 42321 288646
rect 42255 288641 42321 288644
rect 59151 288112 59217 288115
rect 64578 288112 64638 288592
rect 59151 288110 64638 288112
rect 41538 287964 41598 288082
rect 59151 288054 59156 288110
rect 59212 288054 64638 288110
rect 59151 288052 64638 288054
rect 649986 288112 650046 288592
rect 675663 288558 675729 288559
rect 675663 288554 675712 288558
rect 675776 288556 675782 288558
rect 675663 288498 675668 288554
rect 675663 288494 675712 288498
rect 675776 288496 675820 288556
rect 675776 288494 675782 288496
rect 675663 288493 675729 288494
rect 655407 288112 655473 288115
rect 649986 288110 655473 288112
rect 649986 288054 655412 288110
rect 655468 288054 655473 288110
rect 649986 288052 655473 288054
rect 59151 288049 59217 288052
rect 655407 288049 655473 288052
rect 41538 287904 41790 287964
rect 28866 287375 28926 287712
rect 41730 287520 41790 287904
rect 675567 287818 675633 287819
rect 675514 287816 675520 287818
rect 675476 287756 675520 287816
rect 675584 287814 675633 287818
rect 675628 287758 675633 287814
rect 675514 287754 675520 287756
rect 675584 287754 675633 287758
rect 675567 287753 675633 287754
rect 28815 287370 28926 287375
rect 28815 287314 28820 287370
rect 28876 287314 28926 287370
rect 28815 287312 28926 287314
rect 41538 287460 41790 287520
rect 28815 287309 28881 287312
rect 41538 287224 41598 287460
rect 41871 287224 41937 287227
rect 41538 287222 41937 287224
rect 41538 287194 41876 287222
rect 41568 287166 41876 287194
rect 41932 287166 41937 287222
rect 41568 287164 41937 287166
rect 41871 287161 41937 287164
rect 28815 286928 28881 286931
rect 59247 286928 59313 286931
rect 64578 286928 64638 287410
rect 28815 286926 28926 286928
rect 28815 286870 28820 286926
rect 28876 286870 28926 286926
rect 28815 286865 28926 286870
rect 59247 286926 64638 286928
rect 59247 286870 59252 286926
rect 59308 286870 64638 286926
rect 59247 286868 64638 286870
rect 649986 286928 650046 287410
rect 675130 287162 675136 287226
rect 675200 287224 675206 287226
rect 675471 287224 675537 287227
rect 675200 287222 675537 287224
rect 675200 287166 675476 287222
rect 675532 287166 675537 287222
rect 675200 287164 675537 287166
rect 675200 287162 675206 287164
rect 675471 287161 675537 287164
rect 655695 286928 655761 286931
rect 649986 286926 655761 286928
rect 649986 286870 655700 286926
rect 655756 286870 655761 286926
rect 649986 286868 655761 286870
rect 59247 286865 59313 286868
rect 655695 286865 655761 286868
rect 28866 286602 28926 286865
rect 675759 286632 675825 286635
rect 676474 286632 676480 286634
rect 675759 286630 676480 286632
rect 675759 286574 675764 286630
rect 675820 286574 676480 286630
rect 675759 286572 676480 286574
rect 675759 286569 675825 286572
rect 676474 286570 676480 286572
rect 676544 286570 676550 286634
rect 59055 285744 59121 285747
rect 64578 285744 64638 286228
rect 59055 285742 64638 285744
rect 59055 285686 59060 285742
rect 59116 285686 64638 285742
rect 59055 285684 64638 285686
rect 649986 285744 650046 286228
rect 655503 285744 655569 285747
rect 649986 285742 655569 285744
rect 649986 285686 655508 285742
rect 655564 285686 655569 285742
rect 649986 285684 655569 285686
rect 59055 285681 59121 285684
rect 655503 285681 655569 285684
rect 674938 285534 674944 285598
rect 675008 285596 675014 285598
rect 675471 285596 675537 285599
rect 675008 285594 675537 285596
rect 675008 285538 675476 285594
rect 675532 285538 675537 285594
rect 675008 285536 675537 285538
rect 675008 285534 675014 285536
rect 675471 285533 675537 285536
rect 57615 284560 57681 284563
rect 64578 284560 64638 285046
rect 57615 284558 64638 284560
rect 57615 284502 57620 284558
rect 57676 284502 64638 284558
rect 57615 284500 64638 284502
rect 649986 284560 650046 285046
rect 653775 284560 653841 284563
rect 649986 284558 653841 284560
rect 649986 284502 653780 284558
rect 653836 284502 653841 284558
rect 649986 284500 653841 284502
rect 57615 284497 57681 284500
rect 653775 284497 653841 284500
rect 58863 283376 58929 283379
rect 64578 283376 64638 283864
rect 58863 283374 64638 283376
rect 58863 283318 58868 283374
rect 58924 283318 64638 283374
rect 58863 283316 64638 283318
rect 649986 283376 650046 283864
rect 655119 283376 655185 283379
rect 649986 283374 655185 283376
rect 649986 283318 655124 283374
rect 655180 283318 655185 283374
rect 649986 283316 655185 283318
rect 58863 283313 58929 283316
rect 655119 283313 655185 283316
rect 674746 283166 674752 283230
rect 674816 283228 674822 283230
rect 675087 283228 675153 283231
rect 674816 283226 675153 283228
rect 674816 283170 675092 283226
rect 675148 283170 675153 283226
rect 674816 283168 675153 283170
rect 674816 283166 674822 283168
rect 675087 283165 675153 283168
rect 58959 282340 59025 282343
rect 64578 282340 64638 282682
rect 58959 282338 64638 282340
rect 58959 282282 58964 282338
rect 59020 282282 64638 282338
rect 58959 282280 64638 282282
rect 649986 282340 650046 282682
rect 655311 282340 655377 282343
rect 649986 282338 655377 282340
rect 649986 282282 655316 282338
rect 655372 282282 655377 282338
rect 649986 282280 655377 282282
rect 58959 282277 59025 282280
rect 655311 282277 655377 282280
rect 674170 282130 674176 282194
rect 674240 282192 674246 282194
rect 675087 282192 675153 282195
rect 674240 282190 675153 282192
rect 674240 282134 675092 282190
rect 675148 282134 675153 282190
rect 674240 282132 675153 282134
rect 674240 282130 674246 282132
rect 675087 282129 675153 282132
rect 59247 281008 59313 281011
rect 64578 281008 64638 281500
rect 59247 281006 64638 281008
rect 59247 280950 59252 281006
rect 59308 280950 64638 281006
rect 59247 280948 64638 280950
rect 649986 281008 650046 281500
rect 655215 281008 655281 281011
rect 649986 281006 655281 281008
rect 649986 280950 655220 281006
rect 655276 280950 655281 281006
rect 649986 280948 655281 280950
rect 59247 280945 59313 280948
rect 655215 280945 655281 280948
rect 59535 279824 59601 279827
rect 64578 279824 64638 280318
rect 59535 279822 64638 279824
rect 59535 279766 59540 279822
rect 59596 279766 64638 279822
rect 59535 279764 64638 279766
rect 649986 279824 650046 280318
rect 654159 279824 654225 279827
rect 649986 279822 654225 279824
rect 649986 279766 654164 279822
rect 654220 279766 654225 279822
rect 649986 279764 654225 279766
rect 59535 279761 59601 279764
rect 654159 279761 654225 279764
rect 40570 278578 40576 278642
rect 40640 278640 40646 278642
rect 672399 278640 672465 278643
rect 40640 278638 672465 278640
rect 40640 278582 672404 278638
rect 672460 278582 672465 278638
rect 40640 278580 672465 278582
rect 40640 278578 40646 278580
rect 672399 278577 672465 278580
rect 62127 278492 62193 278495
rect 676858 278492 676864 278494
rect 62127 278490 676864 278492
rect 62127 278434 62132 278490
rect 62188 278434 676864 278490
rect 62127 278432 676864 278434
rect 62127 278429 62193 278432
rect 676858 278430 676864 278432
rect 676928 278430 676934 278494
rect 61935 278344 62001 278347
rect 675087 278344 675153 278347
rect 675898 278344 675904 278346
rect 61935 278342 675904 278344
rect 61935 278286 61940 278342
rect 61996 278286 675092 278342
rect 675148 278286 675904 278342
rect 61935 278284 675904 278286
rect 61935 278281 62001 278284
rect 675087 278281 675153 278284
rect 675898 278282 675904 278284
rect 675968 278282 675974 278346
rect 63087 278196 63153 278199
rect 672591 278196 672657 278199
rect 63087 278194 672657 278196
rect 63087 278138 63092 278194
rect 63148 278138 672596 278194
rect 672652 278138 672657 278194
rect 63087 278136 672657 278138
rect 63087 278133 63153 278136
rect 672591 278133 672657 278136
rect 62511 278048 62577 278051
rect 670671 278048 670737 278051
rect 62511 278046 670737 278048
rect 62511 277990 62516 278046
rect 62572 277990 670676 278046
rect 670732 277990 670737 278046
rect 62511 277988 670737 277990
rect 62511 277985 62577 277988
rect 670671 277985 670737 277988
rect 61647 277900 61713 277903
rect 669903 277900 669969 277903
rect 61647 277898 669969 277900
rect 61647 277842 61652 277898
rect 61708 277842 669908 277898
rect 669964 277842 669969 277898
rect 61647 277840 669969 277842
rect 61647 277837 61713 277840
rect 669903 277837 669969 277840
rect 62895 277752 62961 277755
rect 670479 277752 670545 277755
rect 62895 277750 670545 277752
rect 62895 277694 62900 277750
rect 62956 277694 670484 277750
rect 670540 277694 670545 277750
rect 62895 277692 670545 277694
rect 62895 277689 62961 277692
rect 670479 277689 670545 277692
rect 62703 277604 62769 277607
rect 670287 277604 670353 277607
rect 62703 277602 670353 277604
rect 62703 277546 62708 277602
rect 62764 277546 670292 277602
rect 670348 277546 670353 277602
rect 62703 277544 670353 277546
rect 62703 277541 62769 277544
rect 670287 277541 670353 277544
rect 63279 277456 63345 277459
rect 670095 277456 670161 277459
rect 63279 277454 670161 277456
rect 63279 277398 63284 277454
rect 63340 277398 670100 277454
rect 670156 277398 670161 277454
rect 63279 277396 670161 277398
rect 63279 277393 63345 277396
rect 670095 277393 670161 277396
rect 670191 277220 670257 277223
rect 658227 277219 670257 277220
rect 658217 277218 670257 277219
rect 658217 277162 670196 277218
rect 670252 277162 670257 277218
rect 658217 277160 670257 277162
rect 405423 276864 405489 276867
rect 521295 276864 521361 276867
rect 405423 276862 521361 276864
rect 405423 276806 405428 276862
rect 405484 276806 521300 276862
rect 521356 276806 521361 276862
rect 405423 276804 521361 276806
rect 405423 276801 405489 276804
rect 521295 276801 521361 276804
rect 402543 276716 402609 276719
rect 529839 276716 529905 276719
rect 402543 276714 529905 276716
rect 402543 276658 402548 276714
rect 402604 276658 529844 276714
rect 529900 276658 529905 276714
rect 402543 276656 529905 276658
rect 402543 276653 402609 276656
rect 529839 276653 529905 276656
rect 395151 276568 395217 276571
rect 607215 276568 607281 276571
rect 395151 276566 607281 276568
rect 395151 276510 395156 276566
rect 395212 276510 607220 276566
rect 607276 276510 607281 276566
rect 395151 276508 607281 276510
rect 395151 276505 395217 276508
rect 607215 276505 607281 276508
rect 43066 276358 43072 276422
rect 43136 276420 43142 276422
rect 658217 276420 658277 277160
rect 670191 277157 670257 277160
rect 670383 277072 670449 277075
rect 43136 276360 658277 276420
rect 658550 277070 670449 277072
rect 658550 277014 670388 277070
rect 670444 277014 670449 277070
rect 658550 277012 670449 277014
rect 43136 276358 43142 276360
rect 45135 276272 45201 276275
rect 658550 276272 658610 277012
rect 670383 277009 670449 277012
rect 45135 276270 658611 276272
rect 45135 276214 45140 276270
rect 45196 276214 658611 276270
rect 45135 276212 658611 276214
rect 45135 276209 45201 276212
rect 379023 276124 379089 276127
rect 566991 276124 567057 276127
rect 379023 276122 567057 276124
rect 379023 276066 379028 276122
rect 379084 276066 566996 276122
rect 567052 276066 567057 276122
rect 379023 276064 567057 276066
rect 379023 276061 379089 276064
rect 566991 276061 567057 276064
rect 383439 275976 383505 275979
rect 577647 275976 577713 275979
rect 383439 275974 577713 275976
rect 383439 275918 383444 275974
rect 383500 275918 577652 275974
rect 577708 275918 577713 275974
rect 383439 275916 577713 275918
rect 383439 275913 383505 275916
rect 577647 275913 577713 275916
rect 390351 275828 390417 275831
rect 595407 275828 595473 275831
rect 390351 275826 595473 275828
rect 390351 275770 390356 275826
rect 390412 275770 595412 275826
rect 595468 275770 595473 275826
rect 390351 275768 595473 275770
rect 390351 275765 390417 275768
rect 595407 275765 595473 275768
rect 398895 275680 398961 275683
rect 616623 275680 616689 275683
rect 398895 275678 616689 275680
rect 398895 275622 398900 275678
rect 398956 275622 616628 275678
rect 616684 275622 616689 275678
rect 398895 275620 616689 275622
rect 398895 275617 398961 275620
rect 616623 275617 616689 275620
rect 658346 275636 658406 275637
rect 669711 275636 669777 275639
rect 658346 275634 669777 275636
rect 658346 275578 669716 275634
rect 669772 275578 669777 275634
rect 658346 275576 669777 275578
rect 407823 275532 407889 275535
rect 637935 275532 638001 275535
rect 407823 275530 638001 275532
rect 407823 275474 407828 275530
rect 407884 275474 637940 275530
rect 637996 275474 638001 275530
rect 407823 275472 638001 275474
rect 407823 275469 407889 275472
rect 637935 275469 638001 275472
rect 44751 275384 44817 275387
rect 646479 275384 646545 275387
rect 44751 275382 646545 275384
rect 44751 275326 44756 275382
rect 44812 275326 646484 275382
rect 646540 275326 646545 275382
rect 44751 275324 646545 275326
rect 44751 275321 44817 275324
rect 646479 275321 646545 275324
rect 50607 275236 50673 275239
rect 658346 275236 658406 275576
rect 669711 275573 669777 275576
rect 669519 275488 669585 275491
rect 50607 275234 658406 275236
rect 50607 275178 50612 275234
rect 50668 275178 658406 275234
rect 50607 275176 658406 275178
rect 658660 275486 669585 275488
rect 658660 275430 669524 275486
rect 669580 275430 669585 275486
rect 658660 275428 669585 275430
rect 50607 275173 50673 275176
rect 50415 275088 50481 275091
rect 658660 275088 658720 275428
rect 669519 275425 669585 275428
rect 50415 275086 658720 275088
rect 50415 275030 50420 275086
rect 50476 275030 658720 275086
rect 50415 275028 658720 275030
rect 50415 275025 50481 275028
rect 353391 274940 353457 274943
rect 503151 274940 503217 274943
rect 353391 274938 503217 274940
rect 353391 274882 353396 274938
rect 353452 274882 503156 274938
rect 503212 274882 503217 274938
rect 353391 274880 503217 274882
rect 353391 274877 353457 274880
rect 503151 274877 503217 274880
rect 350223 274792 350289 274795
rect 496047 274792 496113 274795
rect 350223 274790 496113 274792
rect 350223 274734 350228 274790
rect 350284 274734 496052 274790
rect 496108 274734 496113 274790
rect 350223 274732 496113 274734
rect 350223 274729 350289 274732
rect 496047 274729 496113 274732
rect 347631 274644 347697 274647
rect 489039 274644 489105 274647
rect 347631 274642 489105 274644
rect 347631 274586 347636 274642
rect 347692 274586 489044 274642
rect 489100 274586 489105 274642
rect 347631 274584 489105 274586
rect 347631 274581 347697 274584
rect 489039 274581 489105 274584
rect 341679 274496 341745 274499
rect 474831 274496 474897 274499
rect 341679 274494 474897 274496
rect 341679 274438 341684 274494
rect 341740 274438 474836 274494
rect 474892 274438 474897 274494
rect 341679 274436 474897 274438
rect 341679 274433 341745 274436
rect 474831 274433 474897 274436
rect 42298 273546 42304 273610
rect 42368 273608 42374 273610
rect 669999 273608 670065 273611
rect 42368 273606 670065 273608
rect 42368 273550 670004 273606
rect 670060 273550 670065 273606
rect 42368 273548 670065 273550
rect 42368 273546 42374 273548
rect 669999 273545 670065 273548
rect 62607 273460 62673 273463
rect 672495 273460 672561 273463
rect 62607 273458 672561 273460
rect 62607 273402 62612 273458
rect 62668 273402 672500 273458
rect 672556 273402 672561 273458
rect 62607 273400 672561 273402
rect 62607 273397 62673 273400
rect 672495 273397 672561 273400
rect 378639 273312 378705 273315
rect 565839 273312 565905 273315
rect 378639 273310 565905 273312
rect 378639 273254 378644 273310
rect 378700 273254 565844 273310
rect 565900 273254 565905 273310
rect 378639 273252 565905 273254
rect 378639 273249 378705 273252
rect 565839 273249 565905 273252
rect 382959 273164 383025 273167
rect 576495 273164 576561 273167
rect 382959 273162 576561 273164
rect 382959 273106 382964 273162
rect 383020 273106 576500 273162
rect 576556 273106 576561 273162
rect 382959 273104 576561 273106
rect 382959 273101 383025 273104
rect 576495 273101 576561 273104
rect 41338 272954 41344 273018
rect 41408 273016 41414 273018
rect 41775 273016 41841 273019
rect 41408 273014 41841 273016
rect 41408 272958 41780 273014
rect 41836 272958 41841 273014
rect 41408 272956 41841 272958
rect 41408 272954 41414 272956
rect 41775 272953 41841 272956
rect 390159 273016 390225 273019
rect 594159 273016 594225 273019
rect 390159 273014 594225 273016
rect 390159 272958 390164 273014
rect 390220 272958 594164 273014
rect 594220 272958 594225 273014
rect 390159 272956 594225 272958
rect 390159 272953 390225 272956
rect 594159 272953 594225 272956
rect 392751 272868 392817 272871
rect 601263 272868 601329 272871
rect 392751 272866 601329 272868
rect 392751 272810 392756 272866
rect 392812 272810 601268 272866
rect 601324 272810 601329 272866
rect 392751 272808 601329 272810
rect 392751 272805 392817 272808
rect 601263 272805 601329 272808
rect 91887 272720 91953 272723
rect 200175 272720 200241 272723
rect 91887 272718 200241 272720
rect 91887 272662 91892 272718
rect 91948 272662 200180 272718
rect 200236 272662 200241 272718
rect 91887 272660 200241 272662
rect 91887 272657 91953 272660
rect 200175 272657 200241 272660
rect 398703 272720 398769 272723
rect 615471 272720 615537 272723
rect 398703 272718 615537 272720
rect 398703 272662 398708 272718
rect 398764 272662 615476 272718
rect 615532 272662 615537 272718
rect 398703 272660 615537 272662
rect 398703 272657 398769 272660
rect 615471 272657 615537 272660
rect 88335 272572 88401 272575
rect 199215 272572 199281 272575
rect 88335 272570 199281 272572
rect 88335 272514 88340 272570
rect 88396 272514 199220 272570
rect 199276 272514 199281 272570
rect 88335 272512 199281 272514
rect 88335 272509 88401 272512
rect 199215 272509 199281 272512
rect 404175 272572 404241 272575
rect 629679 272572 629745 272575
rect 404175 272570 629745 272572
rect 404175 272514 404180 272570
rect 404236 272514 629684 272570
rect 629740 272514 629745 272570
rect 404175 272512 629745 272514
rect 404175 272509 404241 272512
rect 629679 272509 629745 272512
rect 41530 272362 41536 272426
rect 41600 272424 41606 272426
rect 41775 272424 41841 272427
rect 41600 272422 41841 272424
rect 41600 272366 41780 272422
rect 41836 272366 41841 272422
rect 41600 272364 41841 272366
rect 41600 272362 41606 272364
rect 41775 272361 41841 272364
rect 78831 272424 78897 272427
rect 196623 272424 196689 272427
rect 78831 272422 196689 272424
rect 78831 272366 78836 272422
rect 78892 272366 196628 272422
rect 196684 272366 196689 272422
rect 78831 272364 196689 272366
rect 78831 272361 78897 272364
rect 196623 272361 196689 272364
rect 407247 272424 407313 272427
rect 636783 272424 636849 272427
rect 407247 272422 636849 272424
rect 407247 272366 407252 272422
rect 407308 272366 636788 272422
rect 636844 272366 636849 272422
rect 407247 272364 636849 272366
rect 407247 272361 407313 272364
rect 636783 272361 636849 272364
rect 72975 272276 73041 272279
rect 194415 272276 194481 272279
rect 72975 272274 194481 272276
rect 72975 272218 72980 272274
rect 73036 272218 194420 272274
rect 194476 272218 194481 272274
rect 72975 272216 194481 272218
rect 72975 272213 73041 272216
rect 194415 272213 194481 272216
rect 410895 272276 410961 272279
rect 646191 272276 646257 272279
rect 410895 272274 646257 272276
rect 410895 272218 410900 272274
rect 410956 272218 646196 272274
rect 646252 272218 646257 272274
rect 410895 272216 646257 272218
rect 410895 272213 410961 272216
rect 646191 272213 646257 272216
rect 70575 272128 70641 272131
rect 193743 272128 193809 272131
rect 70575 272126 193809 272128
rect 70575 272070 70580 272126
rect 70636 272070 193748 272126
rect 193804 272070 193809 272126
rect 70575 272068 193809 272070
rect 70575 272065 70641 272068
rect 193743 272065 193809 272068
rect 411759 272128 411825 272131
rect 648591 272128 648657 272131
rect 411759 272126 648657 272128
rect 411759 272070 411764 272126
rect 411820 272070 648596 272126
rect 648652 272070 648657 272126
rect 411759 272068 648657 272070
rect 411759 272065 411825 272068
rect 648591 272065 648657 272068
rect 375567 271980 375633 271983
rect 558735 271980 558801 271983
rect 375567 271978 558801 271980
rect 375567 271922 375572 271978
rect 375628 271922 558740 271978
rect 558796 271922 558801 271978
rect 375567 271920 558801 271922
rect 375567 271917 375633 271920
rect 558735 271917 558801 271920
rect 370095 271832 370161 271835
rect 544527 271832 544593 271835
rect 370095 271830 544593 271832
rect 370095 271774 370100 271830
rect 370156 271774 544532 271830
rect 544588 271774 544593 271830
rect 370095 271772 544593 271774
rect 370095 271769 370161 271772
rect 544527 271769 544593 271772
rect 369615 271684 369681 271687
rect 543375 271684 543441 271687
rect 369615 271682 543441 271684
rect 369615 271626 369620 271682
rect 369676 271626 543380 271682
rect 543436 271626 543441 271682
rect 369615 271624 543441 271626
rect 369615 271621 369681 271624
rect 543375 271621 543441 271624
rect 40954 270586 40960 270650
rect 41024 270648 41030 270650
rect 41775 270648 41841 270651
rect 41024 270646 41841 270648
rect 41024 270590 41780 270646
rect 41836 270590 41841 270646
rect 41024 270588 41841 270590
rect 41024 270586 41030 270588
rect 41775 270585 41841 270588
rect 62319 270648 62385 270651
rect 674554 270648 674560 270650
rect 62319 270646 674560 270648
rect 62319 270590 62324 270646
rect 62380 270590 674560 270646
rect 62319 270588 674560 270590
rect 62319 270585 62385 270588
rect 674554 270586 674560 270588
rect 674624 270648 674630 270650
rect 679695 270648 679761 270651
rect 674624 270646 679761 270648
rect 674624 270590 679700 270646
rect 679756 270590 679761 270646
rect 674624 270588 679761 270590
rect 674624 270586 674630 270588
rect 679695 270585 679761 270588
rect 374319 270500 374385 270503
rect 555183 270500 555249 270503
rect 374319 270498 555249 270500
rect 374319 270442 374324 270498
rect 374380 270442 555188 270498
rect 555244 270442 555249 270498
rect 374319 270440 555249 270442
rect 374319 270437 374385 270440
rect 555183 270437 555249 270440
rect 284271 270352 284337 270355
rect 284655 270352 284721 270355
rect 284271 270350 284721 270352
rect 284271 270294 284276 270350
rect 284332 270294 284660 270350
rect 284716 270294 284721 270350
rect 284271 270292 284721 270294
rect 284271 270289 284337 270292
rect 284655 270289 284721 270292
rect 377007 270352 377073 270355
rect 562287 270352 562353 270355
rect 377007 270350 562353 270352
rect 377007 270294 377012 270350
rect 377068 270294 562292 270350
rect 562348 270294 562353 270350
rect 377007 270292 562353 270294
rect 377007 270289 377073 270292
rect 562287 270289 562353 270292
rect 388431 270204 388497 270207
rect 590607 270204 590673 270207
rect 388431 270202 590673 270204
rect 388431 270146 388436 270202
rect 388492 270146 590612 270202
rect 590668 270146 590673 270202
rect 388431 270144 590673 270146
rect 388431 270141 388497 270144
rect 590607 270141 590673 270144
rect 41146 269994 41152 270058
rect 41216 270056 41222 270058
rect 41775 270056 41841 270059
rect 41216 270054 41841 270056
rect 41216 269998 41780 270054
rect 41836 269998 41841 270054
rect 41216 269996 41841 269998
rect 41216 269994 41222 269996
rect 41775 269993 41841 269996
rect 391503 270056 391569 270059
rect 597711 270056 597777 270059
rect 391503 270054 597777 270056
rect 391503 269998 391508 270054
rect 391564 269998 597716 270054
rect 597772 269998 597777 270054
rect 391503 269996 597777 269998
rect 391503 269993 391569 269996
rect 597711 269993 597777 269996
rect 139119 269908 139185 269911
rect 213327 269908 213393 269911
rect 139119 269906 213393 269908
rect 139119 269850 139124 269906
rect 139180 269850 213332 269906
rect 213388 269850 213393 269906
rect 139119 269848 213393 269850
rect 139119 269845 139185 269848
rect 213327 269845 213393 269848
rect 397071 269908 397137 269911
rect 611919 269908 611985 269911
rect 397071 269906 611985 269908
rect 397071 269850 397076 269906
rect 397132 269850 611924 269906
rect 611980 269850 611985 269906
rect 397071 269848 611985 269850
rect 397071 269845 397137 269848
rect 611919 269845 611985 269848
rect 77583 269760 77649 269763
rect 196143 269760 196209 269763
rect 77583 269758 196209 269760
rect 77583 269702 77588 269758
rect 77644 269702 196148 269758
rect 196204 269702 196209 269758
rect 77583 269700 196209 269702
rect 77583 269697 77649 269700
rect 196143 269697 196209 269700
rect 403023 269760 403089 269763
rect 626127 269760 626193 269763
rect 403023 269758 626193 269760
rect 403023 269702 403028 269758
rect 403084 269702 626132 269758
rect 626188 269702 626193 269758
rect 403023 269700 626193 269702
rect 403023 269697 403089 269700
rect 626127 269697 626193 269700
rect 69423 269612 69489 269615
rect 193071 269612 193137 269615
rect 69423 269610 193137 269612
rect 69423 269554 69428 269610
rect 69484 269554 193076 269610
rect 193132 269554 193137 269610
rect 69423 269552 193137 269554
rect 69423 269549 69489 269552
rect 193071 269549 193137 269552
rect 405615 269612 405681 269615
rect 633231 269612 633297 269615
rect 405615 269610 633297 269612
rect 405615 269554 405620 269610
rect 405676 269554 633236 269610
rect 633292 269554 633297 269610
rect 405615 269552 633297 269554
rect 405615 269549 405681 269552
rect 633231 269549 633297 269552
rect 71727 269464 71793 269467
rect 194223 269464 194289 269467
rect 71727 269462 194289 269464
rect 71727 269406 71732 269462
rect 71788 269406 194228 269462
rect 194284 269406 194289 269462
rect 71727 269404 194289 269406
rect 71727 269401 71793 269404
rect 194223 269401 194289 269404
rect 410415 269464 410481 269467
rect 645039 269464 645105 269467
rect 410415 269462 645105 269464
rect 410415 269406 410420 269462
rect 410476 269406 645044 269462
rect 645100 269406 645105 269462
rect 410415 269404 645105 269406
rect 410415 269401 410481 269404
rect 645039 269401 645105 269404
rect 65871 269316 65937 269319
rect 192399 269316 192465 269319
rect 65871 269314 192465 269316
rect 65871 269258 65876 269314
rect 65932 269258 192404 269314
rect 192460 269258 192465 269314
rect 65871 269256 192465 269258
rect 65871 269253 65937 269256
rect 192399 269253 192465 269256
rect 411567 269316 411633 269319
rect 647343 269316 647409 269319
rect 411567 269314 647409 269316
rect 411567 269258 411572 269314
rect 411628 269258 647348 269314
rect 647404 269258 647409 269314
rect 411567 269256 647409 269258
rect 411567 269253 411633 269256
rect 647343 269253 647409 269256
rect 40762 269106 40768 269170
rect 40832 269168 40838 269170
rect 41775 269168 41841 269171
rect 40832 269166 41841 269168
rect 40832 269110 41780 269166
rect 41836 269110 41841 269166
rect 40832 269108 41841 269110
rect 40832 269106 40838 269108
rect 41775 269105 41841 269108
rect 368367 269168 368433 269171
rect 540975 269168 541041 269171
rect 368367 269166 541041 269168
rect 368367 269110 368372 269166
rect 368428 269110 540980 269166
rect 541036 269110 541041 269166
rect 368367 269108 541041 269110
rect 368367 269105 368433 269108
rect 540975 269105 541041 269108
rect 367887 269020 367953 269023
rect 539823 269020 539889 269023
rect 367887 269018 539889 269020
rect 367887 268962 367892 269018
rect 367948 268962 539828 269018
rect 539884 268962 539889 269018
rect 367887 268960 539889 268962
rect 367887 268957 367953 268960
rect 539823 268957 539889 268960
rect 385551 268872 385617 268875
rect 523023 268872 523089 268875
rect 385551 268870 523089 268872
rect 385551 268814 385556 268870
rect 385612 268814 523028 268870
rect 523084 268814 523089 268870
rect 385551 268812 523089 268814
rect 385551 268809 385617 268812
rect 523023 268809 523089 268812
rect 209583 268132 209649 268135
rect 214287 268132 214353 268135
rect 209583 268130 214353 268132
rect 209583 268074 209588 268130
rect 209644 268074 214292 268130
rect 214348 268074 214353 268130
rect 209583 268072 214353 268074
rect 209583 268069 209649 268072
rect 214287 268069 214353 268072
rect 44655 267096 44721 267099
rect 646575 267096 646641 267099
rect 44655 267094 646641 267096
rect 44655 267038 44660 267094
rect 44716 267038 646580 267094
rect 646636 267038 646641 267094
rect 44655 267036 646641 267038
rect 44655 267033 44721 267036
rect 646575 267033 646641 267036
rect 43503 266948 43569 266951
rect 652239 266948 652305 266951
rect 43503 266946 652305 266948
rect 43503 266890 43508 266946
rect 43564 266890 652244 266946
rect 652300 266890 652305 266946
rect 43503 266888 652305 266890
rect 43503 266885 43569 266888
rect 652239 266885 652305 266888
rect 676143 266948 676209 266951
rect 676290 266948 676350 267214
rect 676143 266946 676350 266948
rect 676143 266890 676148 266946
rect 676204 266890 676350 266946
rect 676143 266888 676350 266890
rect 676143 266885 676209 266888
rect 62031 266800 62097 266803
rect 672399 266800 672465 266803
rect 62031 266798 672465 266800
rect 62031 266742 62036 266798
rect 62092 266742 672404 266798
rect 672460 266742 672465 266798
rect 62031 266740 672465 266742
rect 62031 266737 62097 266740
rect 672399 266737 672465 266740
rect 61839 266652 61905 266655
rect 672591 266652 672657 266655
rect 61839 266650 672657 266652
rect 61839 266594 61844 266650
rect 61900 266594 672596 266650
rect 672652 266594 672657 266650
rect 61839 266592 672657 266594
rect 61839 266589 61905 266592
rect 672591 266589 672657 266592
rect 676290 266507 676350 266770
rect 62415 266504 62481 266507
rect 675322 266504 675328 266506
rect 62415 266502 675328 266504
rect 62415 266446 62420 266502
rect 62476 266446 675328 266502
rect 62415 266444 675328 266446
rect 62415 266441 62481 266444
rect 675322 266442 675328 266444
rect 675392 266442 675398 266506
rect 676239 266502 676350 266507
rect 676239 266446 676244 266502
rect 676300 266446 676350 266502
rect 676239 266444 676350 266446
rect 676239 266441 676305 266444
rect 62223 266356 62289 266359
rect 674362 266356 674368 266358
rect 62223 266354 674368 266356
rect 62223 266298 62228 266354
rect 62284 266298 674368 266354
rect 62223 266296 674368 266298
rect 62223 266293 62289 266296
rect 674362 266294 674368 266296
rect 674432 266294 674438 266358
rect 676047 266208 676113 266211
rect 676047 266206 676320 266208
rect 676047 266150 676052 266206
rect 676108 266150 676320 266206
rect 676047 266148 676320 266150
rect 676047 266145 676113 266148
rect 673978 265702 673984 265766
rect 674048 265764 674054 265766
rect 674048 265704 676320 265764
rect 674048 265702 674054 265704
rect 674170 264962 674176 265026
rect 674240 265024 674246 265026
rect 676290 265024 676350 265216
rect 674240 264964 676350 265024
rect 674240 264962 674246 264964
rect 679695 264876 679761 264879
rect 679695 264874 679806 264876
rect 679695 264818 679700 264874
rect 679756 264818 679806 264874
rect 679695 264813 679806 264818
rect 679746 264698 679806 264813
rect 676047 264284 676113 264287
rect 676047 264282 676320 264284
rect 676047 264226 676052 264282
rect 676108 264226 676320 264282
rect 676047 264224 676320 264226
rect 676047 264221 676113 264224
rect 679791 264136 679857 264139
rect 679746 264134 679857 264136
rect 679746 264078 679796 264134
rect 679852 264078 679857 264134
rect 679746 264073 679857 264078
rect 679746 263736 679806 264073
rect 649743 263544 649809 263547
rect 180470 263542 649809 263544
rect 180470 263486 649748 263542
rect 649804 263486 649809 263542
rect 180470 263484 649809 263486
rect 43311 261944 43377 261947
rect 180470 261944 180530 263484
rect 649743 263481 649809 263484
rect 674554 263248 674560 263250
rect 659490 263188 674560 263248
rect 659490 263100 659550 263188
rect 674554 263186 674560 263188
rect 674624 263248 674630 263250
rect 674624 263188 676320 263248
rect 674624 263186 674630 263188
rect 43311 261942 180530 261944
rect 43311 261886 43316 261942
rect 43372 261886 180530 261942
rect 43311 261884 180530 261886
rect 43311 261881 43377 261884
rect 180470 261878 180530 261884
rect 180780 263040 659550 263100
rect 44943 261700 45009 261703
rect 180780 261700 180840 263040
rect 676290 262659 676350 262774
rect 676239 262654 676350 262659
rect 676239 262598 676244 262654
rect 676300 262598 676350 262654
rect 676239 262596 676350 262598
rect 676239 262593 676305 262596
rect 420399 262212 420465 262215
rect 412512 262210 420465 262212
rect 412512 262154 420404 262210
rect 420460 262154 420465 262210
rect 412512 262152 420465 262154
rect 420399 262149 420465 262152
rect 674746 262150 674752 262214
rect 674816 262212 674822 262214
rect 674816 262152 676320 262212
rect 674816 262150 674822 262152
rect 44943 261698 180840 261700
rect 44943 261642 44948 261698
rect 45004 261644 180840 261698
rect 45004 261642 180780 261644
rect 44943 261640 180780 261642
rect 44943 261637 45009 261640
rect 676290 261474 676350 261738
rect 676282 261410 676288 261474
rect 676352 261410 676358 261474
rect 676047 261324 676113 261327
rect 676047 261322 676320 261324
rect 676047 261266 676052 261322
rect 676108 261266 676320 261322
rect 676047 261264 676320 261266
rect 676047 261261 676113 261264
rect 675706 260670 675712 260734
rect 675776 260732 675782 260734
rect 675776 260672 676320 260732
rect 675776 260670 675782 260672
rect 676866 259995 676926 260184
rect 676815 259990 676926 259995
rect 676815 259934 676820 259990
rect 676876 259934 676926 259990
rect 676815 259932 676926 259934
rect 676815 259929 676881 259932
rect 420399 259844 420465 259847
rect 412512 259842 420465 259844
rect 412512 259786 420404 259842
rect 420460 259786 420465 259842
rect 412512 259784 420465 259786
rect 420399 259781 420465 259784
rect 675279 259844 675345 259847
rect 675279 259842 676320 259844
rect 675279 259786 675284 259842
rect 675340 259786 676320 259842
rect 675279 259784 676320 259786
rect 675279 259781 675345 259784
rect 191535 259400 191601 259403
rect 191535 259398 191904 259400
rect 191535 259342 191540 259398
rect 191596 259342 191904 259398
rect 191535 259340 191904 259342
rect 191535 259337 191601 259340
rect 676047 259252 676113 259255
rect 676047 259250 676320 259252
rect 676047 259194 676052 259250
rect 676108 259194 676320 259250
rect 676047 259192 676320 259194
rect 676047 259189 676113 259192
rect 676047 258734 676113 258737
rect 676047 258732 676320 258734
rect 676047 258676 676052 258732
rect 676108 258676 676320 258732
rect 676047 258674 676320 258676
rect 676047 258671 676113 258674
rect 675130 258302 675136 258366
rect 675200 258364 675206 258366
rect 675200 258304 676320 258364
rect 675200 258302 675206 258304
rect 674938 257710 674944 257774
rect 675008 257772 675014 257774
rect 675008 257712 676320 257772
rect 675008 257710 675014 257712
rect 412482 257032 412542 257520
rect 676290 257035 676350 257150
rect 420399 257032 420465 257035
rect 412482 257030 420465 257032
rect 412482 256974 420404 257030
rect 420460 256974 420465 257030
rect 412482 256972 420465 256974
rect 420399 256969 420465 256972
rect 676239 257030 676350 257035
rect 676239 256974 676244 257030
rect 676300 256974 676350 257030
rect 676239 256972 676350 256974
rect 676239 256969 676305 256972
rect 676047 256884 676113 256887
rect 676047 256882 676320 256884
rect 676047 256826 676052 256882
rect 676108 256826 676320 256882
rect 676047 256824 676320 256826
rect 676047 256821 676113 256824
rect 40194 256295 40254 256410
rect 40194 256290 40305 256295
rect 40194 256234 40244 256290
rect 40300 256234 40305 256290
rect 40194 256232 40305 256234
rect 40239 256229 40305 256232
rect 676047 256292 676113 256295
rect 676047 256290 676320 256292
rect 676047 256234 676052 256290
rect 676108 256234 676320 256290
rect 676047 256232 676320 256234
rect 676047 256229 676113 256232
rect 41538 255703 41598 255966
rect 41538 255698 41649 255703
rect 41538 255642 41588 255698
rect 41644 255642 41649 255698
rect 41538 255640 41649 255642
rect 41583 255637 41649 255640
rect 679746 255555 679806 255670
rect 679695 255550 679806 255555
rect 679695 255494 679700 255550
rect 679756 255494 679806 255550
rect 679695 255492 679806 255494
rect 679695 255489 679761 255492
rect 41775 255404 41841 255407
rect 41568 255402 41841 255404
rect 41568 255346 41780 255402
rect 41836 255346 41841 255402
rect 41568 255344 41841 255346
rect 41775 255341 41841 255344
rect 420399 255256 420465 255259
rect 412512 255254 420465 255256
rect 412512 255198 420404 255254
rect 420460 255198 420465 255254
rect 412512 255196 420465 255198
rect 420399 255193 420465 255196
rect 685506 254963 685566 255300
rect 41775 254960 41841 254963
rect 41568 254958 41841 254960
rect 41568 254902 41780 254958
rect 41836 254902 41841 254958
rect 41568 254900 41841 254902
rect 41775 254897 41841 254900
rect 679695 254960 679761 254963
rect 679695 254958 679806 254960
rect 679695 254902 679700 254958
rect 679756 254902 679806 254958
rect 679695 254897 679806 254902
rect 685455 254958 685566 254963
rect 685455 254902 685460 254958
rect 685516 254902 685566 254958
rect 685455 254900 685566 254902
rect 685455 254897 685521 254900
rect 679746 254782 679806 254897
rect 41775 254516 41841 254519
rect 41568 254514 41841 254516
rect 41568 254458 41780 254514
rect 41836 254458 41841 254514
rect 41568 254456 41841 254458
rect 41775 254453 41841 254456
rect 685455 254516 685521 254519
rect 685455 254514 685566 254516
rect 685455 254458 685460 254514
rect 685516 254458 685566 254514
rect 685455 254453 685566 254458
rect 23151 254220 23217 254223
rect 23106 254218 23217 254220
rect 23106 254162 23156 254218
rect 23212 254162 23217 254218
rect 685506 254190 685566 254453
rect 23106 254157 23217 254162
rect 23106 253894 23166 254157
rect 23298 253335 23358 253450
rect 23055 253332 23121 253335
rect 23055 253330 23166 253332
rect 23055 253274 23060 253330
rect 23116 253274 23166 253330
rect 23055 253269 23166 253274
rect 23298 253330 23409 253335
rect 23298 253274 23348 253330
rect 23404 253274 23409 253330
rect 23298 253272 23409 253274
rect 23343 253269 23409 253272
rect 675898 253270 675904 253334
rect 675968 253332 675974 253334
rect 676815 253332 676881 253335
rect 675968 253330 676881 253332
rect 675968 253274 676820 253330
rect 676876 253274 676881 253330
rect 675968 253272 676881 253274
rect 675968 253270 675974 253272
rect 676815 253269 676881 253272
rect 23106 252932 23166 253269
rect 420399 252888 420465 252891
rect 412512 252886 420465 252888
rect 412512 252830 420404 252886
rect 420460 252830 420465 252886
rect 412512 252828 420465 252830
rect 420399 252825 420465 252828
rect 23247 252740 23313 252743
rect 23247 252738 23358 252740
rect 23247 252682 23252 252738
rect 23308 252682 23358 252738
rect 23247 252677 23358 252682
rect 23298 252414 23358 252677
rect 40386 251706 40446 251970
rect 40378 251642 40384 251706
rect 40448 251642 40454 251706
rect 190191 251704 190257 251707
rect 190191 251702 191904 251704
rect 190191 251646 190196 251702
rect 190252 251646 191904 251702
rect 190191 251644 191904 251646
rect 190191 251641 190257 251644
rect 40194 251263 40254 251378
rect 40194 251258 40305 251263
rect 40194 251202 40244 251258
rect 40300 251202 40305 251258
rect 40194 251200 40305 251202
rect 40239 251197 40305 251200
rect 40578 250670 40638 250934
rect 675759 250816 675825 250819
rect 676282 250816 676288 250818
rect 675759 250814 676288 250816
rect 675759 250758 675764 250814
rect 675820 250758 676288 250814
rect 675759 250756 676288 250758
rect 675759 250753 675825 250756
rect 676282 250754 676288 250756
rect 676352 250754 676358 250818
rect 40570 250606 40576 250670
rect 40640 250606 40646 250670
rect 420303 250520 420369 250523
rect 412512 250518 420369 250520
rect 41154 250226 41214 250490
rect 412512 250462 420308 250518
rect 420364 250462 420369 250518
rect 412512 250460 420369 250462
rect 420303 250457 420369 250460
rect 41146 250162 41152 250226
rect 41216 250162 41222 250226
rect 34434 249783 34494 249898
rect 34434 249778 34545 249783
rect 34434 249722 34484 249778
rect 34540 249722 34545 249778
rect 34434 249720 34545 249722
rect 34479 249717 34545 249720
rect 41775 249484 41841 249487
rect 41568 249482 41841 249484
rect 41568 249426 41780 249482
rect 41836 249426 41841 249482
rect 41568 249424 41841 249426
rect 41775 249421 41841 249424
rect 40770 248746 40830 249010
rect 40762 248682 40768 248746
rect 40832 248682 40838 248746
rect 40962 248154 41022 248418
rect 40954 248090 40960 248154
rect 41024 248090 41030 248154
rect 420399 248152 420465 248155
rect 412512 248150 420465 248152
rect 412512 248094 420404 248150
rect 420460 248094 420465 248150
rect 412512 248092 420465 248094
rect 420399 248089 420465 248092
rect 41871 247930 41937 247933
rect 41568 247928 41937 247930
rect 41568 247872 41876 247928
rect 41932 247872 41937 247928
rect 41568 247870 41937 247872
rect 41871 247867 41937 247870
rect 42255 247560 42321 247563
rect 41568 247558 42321 247560
rect 41568 247502 42260 247558
rect 42316 247502 42321 247558
rect 41568 247500 42321 247502
rect 42255 247497 42321 247500
rect 41538 246675 41598 246938
rect 41487 246670 41598 246675
rect 41487 246614 41492 246670
rect 41548 246614 41598 246670
rect 41487 246612 41598 246614
rect 41487 246609 41553 246612
rect 41871 246376 41937 246379
rect 41568 246374 41937 246376
rect 41568 246318 41876 246374
rect 41932 246318 41937 246374
rect 41568 246316 41937 246318
rect 41871 246313 41937 246316
rect 41538 245784 41598 246050
rect 41679 245784 41745 245787
rect 41538 245782 41745 245784
rect 41538 245726 41684 245782
rect 41740 245726 41745 245782
rect 41538 245724 41745 245726
rect 41679 245721 41745 245724
rect 42543 245488 42609 245491
rect 41568 245486 42609 245488
rect 41568 245430 42548 245486
rect 42604 245430 42609 245486
rect 41568 245428 42609 245430
rect 42543 245425 42609 245428
rect 412482 245340 412542 245828
rect 420399 245340 420465 245343
rect 412482 245338 420465 245340
rect 412482 245282 420404 245338
rect 420460 245282 420465 245338
rect 412482 245280 420465 245282
rect 420399 245277 420465 245280
rect 41583 245192 41649 245195
rect 41538 245190 41649 245192
rect 41538 245134 41588 245190
rect 41644 245134 41649 245190
rect 41538 245129 41649 245134
rect 41538 244866 41598 245129
rect 41583 244748 41649 244751
rect 41538 244746 41649 244748
rect 41538 244690 41588 244746
rect 41644 244690 41649 244746
rect 41538 244685 41649 244690
rect 41538 244496 41598 244685
rect 148527 244600 148593 244603
rect 143904 244598 148593 244600
rect 143904 244542 148532 244598
rect 148588 244542 148593 244598
rect 143904 244540 148593 244542
rect 148527 244537 148593 244540
rect 41538 243715 41598 243978
rect 41538 243710 41649 243715
rect 41538 243654 41588 243710
rect 41644 243654 41649 243710
rect 41538 243652 41649 243654
rect 41583 243649 41649 243652
rect 148719 243416 148785 243419
rect 143904 243414 148785 243416
rect 143904 243358 148724 243414
rect 148780 243358 148785 243414
rect 143904 243356 148785 243358
rect 148719 243353 148785 243356
rect 187119 243416 187185 243419
rect 191874 243416 191934 243904
rect 420399 243564 420465 243567
rect 412512 243562 420465 243564
rect 412512 243506 420404 243562
rect 420460 243506 420465 243562
rect 412512 243504 420465 243506
rect 420399 243501 420465 243504
rect 675663 243566 675729 243567
rect 675663 243562 675712 243566
rect 675776 243564 675782 243566
rect 675663 243506 675668 243562
rect 675663 243502 675712 243506
rect 675776 243504 675820 243564
rect 675776 243502 675782 243504
rect 675663 243501 675729 243502
rect 187119 243414 191934 243416
rect 187119 243358 187124 243414
rect 187180 243358 191934 243414
rect 187119 243356 191934 243358
rect 187119 243353 187185 243356
rect 143874 242084 143934 242128
rect 148335 242084 148401 242087
rect 143874 242082 148401 242084
rect 143874 242026 148340 242082
rect 148396 242026 148401 242082
rect 143874 242024 148401 242026
rect 148335 242021 148401 242024
rect 674938 241874 674944 241938
rect 675008 241936 675014 241938
rect 675087 241936 675153 241939
rect 675008 241934 675153 241936
rect 675008 241878 675092 241934
rect 675148 241878 675153 241934
rect 675008 241876 675153 241878
rect 675008 241874 675014 241876
rect 675087 241873 675153 241876
rect 420399 241196 420465 241199
rect 412512 241194 420465 241196
rect 412512 241138 420404 241194
rect 420460 241138 420465 241194
rect 412512 241136 420465 241138
rect 420399 241133 420465 241136
rect 675183 241050 675249 241051
rect 675130 241048 675136 241050
rect 675092 240988 675136 241048
rect 675200 241046 675249 241050
rect 675244 240990 675249 241046
rect 675130 240986 675136 240988
rect 675200 240986 675249 240990
rect 675183 240985 675249 240986
rect 149007 240900 149073 240903
rect 143904 240898 149073 240900
rect 143904 240842 149012 240898
rect 149068 240842 149073 240898
rect 143904 240840 149073 240842
rect 149007 240837 149073 240840
rect 412143 240160 412209 240163
rect 627183 240160 627249 240163
rect 412143 240158 627249 240160
rect 412143 240102 412148 240158
rect 412204 240102 627188 240158
rect 627244 240102 627249 240158
rect 412143 240100 627249 240102
rect 412143 240097 412209 240100
rect 627183 240097 627249 240100
rect 412047 240012 412113 240015
rect 569007 240012 569073 240015
rect 412047 240010 569073 240012
rect 412047 239954 412052 240010
rect 412108 239954 569012 240010
rect 569068 239954 569073 240010
rect 412047 239952 569073 239954
rect 412047 239949 412113 239952
rect 569007 239949 569073 239952
rect 148239 239716 148305 239719
rect 143904 239714 148305 239716
rect 143904 239658 148244 239714
rect 148300 239658 148305 239714
rect 143904 239656 148305 239658
rect 148239 239653 148305 239656
rect 413391 238976 413457 238979
rect 555375 238976 555441 238979
rect 413391 238974 555441 238976
rect 413391 238918 413396 238974
rect 413452 238918 555380 238974
rect 555436 238918 555441 238974
rect 413391 238916 555441 238918
rect 413391 238913 413457 238916
rect 555375 238913 555441 238916
rect 414063 238828 414129 238831
rect 581775 238828 581841 238831
rect 414063 238826 581841 238828
rect 414063 238770 414068 238826
rect 414124 238770 581780 238826
rect 581836 238770 581841 238826
rect 414063 238768 581841 238770
rect 414063 238765 414129 238768
rect 581775 238765 581841 238768
rect 413679 238680 413745 238683
rect 550191 238680 550257 238683
rect 413679 238678 550257 238680
rect 413679 238622 413684 238678
rect 413740 238622 550196 238678
rect 550252 238622 550257 238678
rect 413679 238620 550257 238622
rect 413679 238617 413745 238620
rect 550191 238617 550257 238620
rect 148623 238532 148689 238535
rect 143904 238530 148689 238532
rect 143904 238474 148628 238530
rect 148684 238474 148689 238530
rect 143904 238472 148689 238474
rect 148623 238469 148689 238472
rect 413967 238384 414033 238387
rect 544335 238384 544401 238387
rect 413967 238382 544401 238384
rect 413967 238326 413972 238382
rect 414028 238326 544340 238382
rect 544396 238326 544401 238382
rect 413967 238324 544401 238326
rect 413967 238321 414033 238324
rect 544335 238321 544401 238324
rect 415215 238236 415281 238239
rect 559887 238236 559953 238239
rect 415215 238234 559953 238236
rect 415215 238178 415220 238234
rect 415276 238178 559892 238234
rect 559948 238178 559953 238234
rect 415215 238176 559953 238178
rect 415215 238173 415281 238176
rect 559887 238173 559953 238176
rect 674746 238174 674752 238238
rect 674816 238236 674822 238238
rect 675087 238236 675153 238239
rect 674816 238234 675153 238236
rect 674816 238178 675092 238234
rect 675148 238178 675153 238234
rect 674816 238176 675153 238178
rect 674816 238174 674822 238176
rect 675087 238173 675153 238176
rect 414447 238088 414513 238091
rect 537999 238088 538065 238091
rect 414447 238086 538065 238088
rect 414447 238030 414452 238086
rect 414508 238030 538004 238086
rect 538060 238030 538065 238086
rect 414447 238028 538065 238030
rect 414447 238025 414513 238028
rect 537999 238025 538065 238028
rect 143874 236756 143934 237244
rect 372207 237052 372273 237055
rect 386991 237052 387057 237055
rect 387471 237052 387537 237055
rect 372207 237050 387057 237052
rect 372207 236994 372212 237050
rect 372268 236994 386996 237050
rect 387052 236994 387057 237050
rect 372207 236992 387057 236994
rect 372207 236989 372273 236992
rect 386991 236989 387057 236992
rect 387138 237050 387537 237052
rect 387138 236994 387476 237050
rect 387532 236994 387537 237050
rect 387138 236992 387537 236994
rect 373455 236904 373521 236907
rect 387138 236904 387198 236992
rect 387471 236989 387537 236992
rect 387855 237052 387921 237055
rect 397498 237052 397504 237054
rect 387855 237050 397504 237052
rect 387855 236994 387860 237050
rect 387916 236994 397504 237050
rect 387855 236992 397504 236994
rect 387855 236989 387921 236992
rect 397498 236990 397504 236992
rect 397568 236990 397574 237054
rect 397743 237052 397809 237055
rect 573135 237052 573201 237055
rect 397743 237050 573201 237052
rect 397743 236994 397748 237050
rect 397804 236994 573140 237050
rect 573196 236994 573201 237050
rect 397743 236992 573201 236994
rect 397743 236989 397809 236992
rect 573135 236989 573201 236992
rect 397839 236904 397905 236907
rect 373455 236902 387198 236904
rect 373455 236846 373460 236902
rect 373516 236846 387198 236902
rect 373455 236844 387198 236846
rect 387330 236902 397905 236904
rect 387330 236846 397844 236902
rect 397900 236846 397905 236902
rect 387330 236844 397905 236846
rect 373455 236841 373521 236844
rect 148911 236756 148977 236759
rect 143874 236754 148977 236756
rect 143874 236698 148916 236754
rect 148972 236698 148977 236754
rect 143874 236696 148977 236698
rect 148911 236693 148977 236696
rect 370383 236756 370449 236759
rect 387330 236756 387390 236844
rect 397839 236841 397905 236844
rect 398031 236904 398097 236907
rect 567471 236904 567537 236907
rect 398031 236902 567537 236904
rect 398031 236846 398036 236902
rect 398092 236846 567476 236902
rect 567532 236846 567537 236902
rect 398031 236844 567537 236846
rect 398031 236841 398097 236844
rect 567471 236841 567537 236844
rect 675759 236904 675825 236907
rect 675898 236904 675904 236906
rect 675759 236902 675904 236904
rect 675759 236846 675764 236902
rect 675820 236846 675904 236902
rect 675759 236844 675904 236846
rect 675759 236841 675825 236844
rect 675898 236842 675904 236844
rect 675968 236842 675974 236906
rect 370383 236754 387390 236756
rect 370383 236698 370388 236754
rect 370444 236698 387390 236754
rect 370383 236696 387390 236698
rect 387567 236756 387633 236759
rect 397455 236756 397521 236759
rect 387567 236754 397521 236756
rect 387567 236698 387572 236754
rect 387628 236698 397460 236754
rect 397516 236698 397521 236754
rect 387567 236696 397521 236698
rect 370383 236693 370449 236696
rect 387567 236693 387633 236696
rect 397455 236693 397521 236696
rect 397690 236694 397696 236758
rect 397760 236756 397766 236758
rect 407290 236756 407296 236758
rect 397760 236696 407296 236756
rect 397760 236694 397766 236696
rect 407290 236694 407296 236696
rect 407360 236694 407366 236758
rect 407439 236756 407505 236759
rect 565263 236756 565329 236759
rect 407439 236754 565329 236756
rect 407439 236698 407444 236754
rect 407500 236698 565268 236754
rect 565324 236698 565329 236754
rect 407439 236696 565329 236698
rect 407439 236693 407505 236696
rect 565263 236693 565329 236696
rect 379503 236608 379569 236611
rect 382383 236608 382449 236611
rect 379503 236606 382449 236608
rect 379503 236550 379508 236606
rect 379564 236550 382388 236606
rect 382444 236550 382449 236606
rect 379503 236548 382449 236550
rect 379503 236545 379569 236548
rect 382383 236545 382449 236548
rect 382575 236608 382641 236611
rect 387087 236608 387153 236611
rect 559215 236608 559281 236611
rect 382575 236606 387153 236608
rect 382575 236550 382580 236606
rect 382636 236550 387092 236606
rect 387148 236550 387153 236606
rect 382575 236548 387153 236550
rect 382575 236545 382641 236548
rect 387087 236545 387153 236548
rect 387330 236606 559281 236608
rect 387330 236550 559220 236606
rect 559276 236550 559281 236606
rect 387330 236548 559281 236550
rect 368943 236460 369009 236463
rect 387183 236460 387249 236463
rect 368943 236458 387249 236460
rect 368943 236402 368948 236458
rect 369004 236402 387188 236458
rect 387244 236402 387249 236458
rect 368943 236400 387249 236402
rect 368943 236397 369009 236400
rect 387183 236397 387249 236400
rect 374895 236312 374961 236315
rect 387330 236312 387390 236548
rect 559215 236545 559281 236548
rect 387471 236460 387537 236463
rect 558447 236460 558513 236463
rect 387471 236458 558513 236460
rect 387471 236402 387476 236458
rect 387532 236402 558452 236458
rect 558508 236402 558513 236458
rect 387471 236400 558513 236402
rect 387471 236397 387537 236400
rect 558447 236397 558513 236400
rect 374895 236310 387390 236312
rect 374895 236254 374900 236310
rect 374956 236254 387390 236310
rect 374895 236252 387390 236254
rect 387471 236312 387537 236315
rect 397071 236312 397137 236315
rect 387471 236310 397137 236312
rect 387471 236254 387476 236310
rect 387532 236254 397076 236310
rect 397132 236254 397137 236310
rect 387471 236252 397137 236254
rect 374895 236249 374961 236252
rect 387471 236249 387537 236252
rect 397071 236249 397137 236252
rect 397359 236312 397425 236315
rect 407439 236312 407505 236315
rect 397359 236310 407505 236312
rect 397359 236254 397364 236310
rect 397420 236254 407444 236310
rect 407500 236254 407505 236310
rect 397359 236252 407505 236254
rect 397359 236249 397425 236252
rect 407439 236249 407505 236252
rect 407674 236250 407680 236314
rect 407744 236312 407750 236314
rect 413679 236312 413745 236315
rect 415215 236312 415281 236315
rect 407744 236310 413745 236312
rect 407744 236254 413684 236310
rect 413740 236254 413745 236310
rect 407744 236252 413745 236254
rect 407744 236250 407750 236252
rect 413679 236249 413745 236252
rect 413826 236310 415281 236312
rect 413826 236254 415220 236310
rect 415276 236254 415281 236310
rect 413826 236252 415281 236254
rect 413826 236167 413886 236252
rect 415215 236249 415281 236252
rect 415407 236312 415473 236315
rect 621135 236312 621201 236315
rect 415407 236310 621201 236312
rect 415407 236254 415412 236310
rect 415468 236254 621140 236310
rect 621196 236254 621201 236310
rect 415407 236252 621201 236254
rect 415407 236249 415473 236252
rect 621135 236249 621201 236252
rect 356847 236164 356913 236167
rect 406479 236164 406545 236167
rect 356847 236162 406545 236164
rect 356847 236106 356852 236162
rect 356908 236106 406484 236162
rect 406540 236106 406545 236162
rect 356847 236104 406545 236106
rect 356847 236101 356913 236104
rect 406479 236101 406545 236104
rect 409935 236164 410001 236167
rect 413626 236164 413632 236166
rect 409935 236162 413632 236164
rect 409935 236106 409940 236162
rect 409996 236106 413632 236162
rect 409935 236104 413632 236106
rect 409935 236101 410001 236104
rect 413626 236102 413632 236104
rect 413696 236102 413702 236166
rect 413826 236162 413937 236167
rect 413826 236106 413876 236162
rect 413932 236106 413937 236162
rect 413826 236104 413937 236106
rect 413871 236101 413937 236104
rect 414010 236102 414016 236166
rect 414080 236164 414086 236166
rect 590415 236164 590481 236167
rect 414080 236162 590481 236164
rect 414080 236106 590420 236162
rect 590476 236106 590481 236162
rect 414080 236104 590481 236106
rect 414080 236102 414086 236104
rect 590415 236101 590481 236104
rect 149103 236016 149169 236019
rect 143904 236014 149169 236016
rect 143904 235958 149108 236014
rect 149164 235958 149169 236014
rect 143904 235956 149169 235958
rect 149103 235953 149169 235956
rect 385839 236016 385905 236019
rect 580335 236016 580401 236019
rect 385839 236014 580401 236016
rect 385839 235958 385844 236014
rect 385900 235958 580340 236014
rect 580396 235958 580401 236014
rect 385839 235956 580401 235958
rect 385839 235953 385905 235956
rect 580335 235953 580401 235956
rect 389871 235868 389937 235871
rect 587919 235868 587985 235871
rect 389871 235866 587985 235868
rect 389871 235810 389876 235866
rect 389932 235810 587924 235866
rect 587980 235810 587985 235866
rect 389871 235808 587985 235810
rect 389871 235805 389937 235808
rect 587919 235805 587985 235808
rect 342543 235720 342609 235723
rect 390735 235720 390801 235723
rect 342543 235718 390801 235720
rect 342543 235662 342548 235718
rect 342604 235662 390740 235718
rect 390796 235662 390801 235718
rect 342543 235660 390801 235662
rect 342543 235657 342609 235660
rect 390735 235657 390801 235660
rect 393039 235720 393105 235723
rect 591471 235720 591537 235723
rect 393039 235718 591537 235720
rect 393039 235662 393044 235718
rect 393100 235662 591476 235718
rect 591532 235662 591537 235718
rect 393039 235660 591537 235662
rect 393039 235657 393105 235660
rect 591471 235657 591537 235660
rect 367215 235572 367281 235575
rect 397455 235572 397521 235575
rect 367215 235570 397521 235572
rect 367215 235514 367220 235570
rect 367276 235514 397460 235570
rect 397516 235514 397521 235570
rect 367215 235512 397521 235514
rect 367215 235509 367281 235512
rect 397455 235509 397521 235512
rect 399855 235572 399921 235575
rect 608271 235572 608337 235575
rect 399855 235570 608337 235572
rect 399855 235514 399860 235570
rect 399916 235514 608276 235570
rect 608332 235514 608337 235570
rect 399855 235512 608337 235514
rect 399855 235509 399921 235512
rect 608271 235509 608337 235512
rect 401391 235424 401457 235427
rect 611247 235424 611313 235427
rect 401391 235422 611313 235424
rect 401391 235366 401396 235422
rect 401452 235366 611252 235422
rect 611308 235366 611313 235422
rect 401391 235364 611313 235366
rect 401391 235361 401457 235364
rect 611247 235361 611313 235364
rect 402735 235276 402801 235279
rect 614319 235276 614385 235279
rect 402735 235274 614385 235276
rect 402735 235218 402740 235274
rect 402796 235218 614324 235274
rect 614380 235218 614385 235274
rect 402735 235216 614385 235218
rect 402735 235213 402801 235216
rect 614319 235213 614385 235216
rect 405423 235128 405489 235131
rect 618831 235128 618897 235131
rect 405423 235126 618897 235128
rect 405423 235070 405428 235126
rect 405484 235070 618836 235126
rect 618892 235070 618897 235126
rect 405423 235068 618897 235070
rect 405423 235065 405489 235068
rect 618831 235065 618897 235068
rect 299439 234980 299505 234983
rect 355887 234980 355953 234983
rect 299439 234978 355953 234980
rect 299439 234922 299444 234978
rect 299500 234922 355892 234978
rect 355948 234922 355953 234978
rect 299439 234920 355953 234922
rect 299439 234917 299505 234920
rect 355887 234917 355953 234920
rect 356751 234980 356817 234983
rect 403119 234980 403185 234983
rect 356751 234978 403185 234980
rect 356751 234922 356756 234978
rect 356812 234922 403124 234978
rect 403180 234922 403185 234978
rect 356751 234920 403185 234922
rect 356751 234917 356817 234920
rect 403119 234917 403185 234920
rect 403983 234980 404049 234983
rect 616623 234980 616689 234983
rect 403983 234978 616689 234980
rect 403983 234922 403988 234978
rect 404044 234922 616628 234978
rect 616684 234922 616689 234978
rect 403983 234920 616689 234922
rect 403983 234917 404049 234920
rect 616623 234917 616689 234920
rect 148431 234832 148497 234835
rect 143904 234830 148497 234832
rect 143904 234774 148436 234830
rect 148492 234774 148497 234830
rect 143904 234772 148497 234774
rect 148431 234769 148497 234772
rect 347631 234832 347697 234835
rect 405327 234832 405393 234835
rect 347631 234830 405393 234832
rect 347631 234774 347636 234830
rect 347692 234774 405332 234830
rect 405388 234774 405393 234830
rect 347631 234772 405393 234774
rect 347631 234769 347697 234772
rect 405327 234769 405393 234772
rect 405519 234832 405585 234835
rect 619599 234832 619665 234835
rect 405519 234830 619665 234832
rect 405519 234774 405524 234830
rect 405580 234774 619604 234830
rect 619660 234774 619665 234830
rect 405519 234772 619665 234774
rect 405519 234769 405585 234772
rect 619599 234769 619665 234772
rect 299343 234684 299409 234687
rect 405711 234684 405777 234687
rect 299343 234682 405777 234684
rect 299343 234626 299348 234682
rect 299404 234626 405716 234682
rect 405772 234626 405777 234682
rect 299343 234624 405777 234626
rect 299343 234621 299409 234624
rect 405711 234621 405777 234624
rect 408495 234684 408561 234687
rect 625551 234684 625617 234687
rect 408495 234682 625617 234684
rect 408495 234626 408500 234682
rect 408556 234626 625556 234682
rect 625612 234626 625617 234682
rect 408495 234624 625617 234626
rect 408495 234621 408561 234624
rect 625551 234621 625617 234624
rect 379119 234536 379185 234539
rect 409839 234536 409905 234539
rect 379119 234534 409905 234536
rect 379119 234478 379124 234534
rect 379180 234478 409844 234534
rect 409900 234478 409905 234534
rect 379119 234476 409905 234478
rect 379119 234473 379185 234476
rect 409839 234473 409905 234476
rect 411375 234536 411441 234539
rect 590895 234536 590961 234539
rect 411375 234534 590961 234536
rect 411375 234478 411380 234534
rect 411436 234478 590900 234534
rect 590956 234478 590961 234534
rect 411375 234476 590961 234478
rect 411375 234473 411441 234476
rect 590895 234473 590961 234476
rect 382095 234388 382161 234391
rect 410031 234388 410097 234391
rect 382095 234386 410097 234388
rect 382095 234330 382100 234386
rect 382156 234330 410036 234386
rect 410092 234330 410097 234386
rect 382095 234328 410097 234330
rect 382095 234325 382161 234328
rect 410031 234325 410097 234328
rect 410799 234388 410865 234391
rect 587439 234388 587505 234391
rect 410799 234386 587505 234388
rect 410799 234330 410804 234386
rect 410860 234330 587444 234386
rect 587500 234330 587505 234386
rect 410799 234328 587505 234330
rect 410799 234325 410865 234328
rect 587439 234325 587505 234328
rect 341583 234240 341649 234243
rect 490479 234240 490545 234243
rect 341583 234238 490545 234240
rect 341583 234182 341588 234238
rect 341644 234182 490484 234238
rect 490540 234182 490545 234238
rect 341583 234180 490545 234182
rect 341583 234177 341649 234180
rect 490479 234177 490545 234180
rect 332559 234092 332625 234095
rect 472335 234092 472401 234095
rect 332559 234090 472401 234092
rect 332559 234034 332564 234090
rect 332620 234034 472340 234090
rect 472396 234034 472401 234090
rect 332559 234032 472401 234034
rect 332559 234029 332625 234032
rect 472335 234029 472401 234032
rect 400239 233944 400305 233947
rect 480879 233944 480945 233947
rect 400239 233942 480945 233944
rect 400239 233886 400244 233942
rect 400300 233886 480884 233942
rect 480940 233886 480945 233942
rect 400239 233884 480945 233886
rect 400239 233881 400305 233884
rect 480879 233881 480945 233884
rect 364047 233796 364113 233799
rect 405903 233796 405969 233799
rect 364047 233794 405969 233796
rect 364047 233738 364052 233794
rect 364108 233738 405908 233794
rect 405964 233738 405969 233794
rect 364047 233736 405969 233738
rect 364047 233733 364113 233736
rect 405903 233733 405969 233736
rect 148815 233648 148881 233651
rect 143904 233646 148881 233648
rect 143904 233590 148820 233646
rect 148876 233590 148881 233646
rect 143904 233588 148881 233590
rect 148815 233585 148881 233588
rect 365679 233352 365745 233355
rect 380079 233352 380145 233355
rect 365679 233350 380145 233352
rect 365679 233294 365684 233350
rect 365740 233294 380084 233350
rect 380140 233294 380145 233350
rect 365679 233292 380145 233294
rect 365679 233289 365745 233292
rect 380079 233289 380145 233292
rect 343983 233204 344049 233207
rect 495087 233204 495153 233207
rect 343983 233202 495153 233204
rect 343983 233146 343988 233202
rect 344044 233146 495092 233202
rect 495148 233146 495153 233202
rect 343983 233144 495153 233146
rect 343983 233141 344049 233144
rect 495087 233141 495153 233144
rect 371151 233056 371217 233059
rect 549423 233056 549489 233059
rect 371151 233054 549489 233056
rect 371151 232998 371156 233054
rect 371212 232998 549428 233054
rect 549484 232998 549489 233054
rect 371151 232996 549489 232998
rect 371151 232993 371217 232996
rect 549423 232993 549489 232996
rect 370767 232908 370833 232911
rect 551631 232908 551697 232911
rect 370767 232906 551697 232908
rect 370767 232850 370772 232906
rect 370828 232850 551636 232906
rect 551692 232850 551697 232906
rect 370767 232848 551697 232850
rect 370767 232845 370833 232848
rect 551631 232845 551697 232848
rect 374031 232760 374097 232763
rect 557679 232760 557745 232763
rect 374031 232758 557745 232760
rect 374031 232702 374036 232758
rect 374092 232702 557684 232758
rect 557740 232702 557745 232758
rect 374031 232700 557745 232702
rect 374031 232697 374097 232700
rect 557679 232697 557745 232700
rect 375375 232612 375441 232615
rect 560751 232612 560817 232615
rect 375375 232610 560817 232612
rect 375375 232554 375380 232610
rect 375436 232554 560756 232610
rect 560812 232554 560817 232610
rect 375375 232552 560817 232554
rect 375375 232549 375441 232552
rect 560751 232549 560817 232552
rect 381711 232464 381777 232467
rect 570447 232464 570513 232467
rect 381711 232462 570513 232464
rect 381711 232406 381716 232462
rect 381772 232406 570452 232462
rect 570508 232406 570513 232462
rect 381711 232404 570513 232406
rect 381711 232401 381777 232404
rect 570447 232401 570513 232404
rect 147855 232316 147921 232319
rect 143904 232314 147921 232316
rect 143904 232258 147860 232314
rect 147916 232258 147921 232314
rect 143904 232256 147921 232258
rect 147855 232253 147921 232256
rect 384975 232316 385041 232319
rect 576591 232316 576657 232319
rect 384975 232314 576657 232316
rect 384975 232258 384980 232314
rect 385036 232258 576596 232314
rect 576652 232258 576657 232314
rect 384975 232256 576657 232258
rect 384975 232253 385041 232256
rect 576591 232253 576657 232256
rect 382671 232168 382737 232171
rect 575823 232168 575889 232171
rect 382671 232166 575889 232168
rect 382671 232110 382676 232166
rect 382732 232110 575828 232166
rect 575884 232110 575889 232166
rect 382671 232108 575889 232110
rect 382671 232105 382737 232108
rect 575823 232105 575889 232108
rect 385263 232020 385329 232023
rect 578031 232020 578097 232023
rect 385263 232018 578097 232020
rect 385263 231962 385268 232018
rect 385324 231962 578036 232018
rect 578092 231962 578097 232018
rect 385263 231960 578097 231962
rect 385263 231957 385329 231960
rect 578031 231957 578097 231960
rect 333807 231872 333873 231875
rect 368655 231872 368721 231875
rect 333807 231870 368721 231872
rect 333807 231814 333812 231870
rect 333868 231814 368660 231870
rect 368716 231814 368721 231870
rect 333807 231812 368721 231814
rect 333807 231809 333873 231812
rect 368655 231809 368721 231812
rect 405999 231872 406065 231875
rect 604527 231872 604593 231875
rect 405999 231870 604593 231872
rect 405999 231814 406004 231870
rect 406060 231814 604532 231870
rect 604588 231814 604593 231870
rect 405999 231812 604593 231814
rect 405999 231809 406065 231812
rect 604527 231809 604593 231812
rect 330255 231724 330321 231727
rect 470127 231724 470193 231727
rect 330255 231722 470193 231724
rect 330255 231666 330260 231722
rect 330316 231666 470132 231722
rect 470188 231666 470193 231722
rect 330255 231664 470193 231666
rect 330255 231661 330321 231664
rect 470127 231661 470193 231664
rect 322479 231576 322545 231579
rect 455151 231576 455217 231579
rect 322479 231574 455217 231576
rect 322479 231518 322484 231574
rect 322540 231518 455156 231574
rect 455212 231518 455217 231574
rect 322479 231516 455217 231518
rect 322479 231513 322545 231516
rect 455151 231513 455217 231516
rect 319503 231428 319569 231431
rect 448911 231428 448977 231431
rect 319503 231426 448977 231428
rect 319503 231370 319508 231426
rect 319564 231370 448916 231426
rect 448972 231370 448977 231426
rect 319503 231368 448977 231370
rect 319503 231365 319569 231368
rect 448911 231365 448977 231368
rect 316719 231280 316785 231283
rect 442863 231280 442929 231283
rect 316719 231278 442929 231280
rect 316719 231222 316724 231278
rect 316780 231222 442868 231278
rect 442924 231222 442929 231278
rect 316719 231220 442929 231222
rect 316719 231217 316785 231220
rect 442863 231217 442929 231220
rect 149391 231132 149457 231135
rect 143904 231130 149457 231132
rect 143904 231074 149396 231130
rect 149452 231074 149457 231130
rect 143904 231072 149457 231074
rect 149391 231069 149457 231072
rect 307599 231132 307665 231135
rect 424719 231132 424785 231135
rect 307599 231130 424785 231132
rect 307599 231074 307604 231130
rect 307660 231074 424724 231130
rect 424780 231074 424785 231130
rect 307599 231072 424785 231074
rect 307599 231069 307665 231072
rect 424719 231069 424785 231072
rect 408111 230392 408177 230395
rect 575055 230392 575121 230395
rect 408111 230390 575121 230392
rect 408111 230334 408116 230390
rect 408172 230334 575060 230390
rect 575116 230334 575121 230390
rect 408111 230332 575121 230334
rect 408111 230329 408177 230332
rect 575055 230329 575121 230332
rect 363567 230244 363633 230247
rect 534255 230244 534321 230247
rect 363567 230242 534321 230244
rect 363567 230186 363572 230242
rect 363628 230186 534260 230242
rect 534316 230186 534321 230242
rect 363567 230184 534321 230186
rect 363567 230181 363633 230184
rect 534255 230181 534321 230184
rect 358959 230096 359025 230099
rect 527535 230096 527601 230099
rect 358959 230094 527601 230096
rect 358959 230038 358964 230094
rect 359020 230038 527540 230094
rect 527596 230038 527601 230094
rect 358959 230036 527601 230038
rect 358959 230033 359025 230036
rect 527535 230033 527601 230036
rect 146895 229948 146961 229951
rect 143904 229946 146961 229948
rect 143904 229890 146900 229946
rect 146956 229890 146961 229946
rect 143904 229888 146961 229890
rect 146895 229885 146961 229888
rect 366639 229948 366705 229951
rect 540303 229948 540369 229951
rect 366639 229946 540369 229948
rect 366639 229890 366644 229946
rect 366700 229890 540308 229946
rect 540364 229890 540369 229946
rect 366639 229888 540369 229890
rect 366639 229885 366705 229888
rect 540303 229885 540369 229888
rect 40954 229738 40960 229802
rect 41024 229800 41030 229802
rect 41775 229800 41841 229803
rect 41024 229798 41841 229800
rect 41024 229742 41780 229798
rect 41836 229742 41841 229798
rect 41024 229740 41841 229742
rect 41024 229738 41030 229740
rect 41775 229737 41841 229740
rect 373071 229800 373137 229803
rect 553935 229800 554001 229803
rect 373071 229798 554001 229800
rect 373071 229742 373076 229798
rect 373132 229742 553940 229798
rect 553996 229742 554001 229798
rect 373071 229740 554001 229742
rect 373071 229737 373137 229740
rect 553935 229737 554001 229740
rect 379887 229652 379953 229655
rect 569775 229652 569841 229655
rect 379887 229650 569841 229652
rect 379887 229594 379892 229650
rect 379948 229594 569780 229650
rect 569836 229594 569841 229650
rect 379887 229592 569841 229594
rect 379887 229589 379953 229592
rect 569775 229589 569841 229592
rect 381327 229504 381393 229507
rect 572751 229504 572817 229507
rect 381327 229502 572817 229504
rect 381327 229446 381332 229502
rect 381388 229446 572756 229502
rect 572812 229446 572817 229502
rect 381327 229444 572817 229446
rect 381327 229441 381393 229444
rect 572751 229441 572817 229444
rect 383535 229356 383601 229359
rect 573519 229356 573585 229359
rect 383535 229354 573585 229356
rect 383535 229298 383540 229354
rect 383596 229298 573524 229354
rect 573580 229298 573585 229354
rect 383535 229296 573585 229298
rect 383535 229293 383601 229296
rect 573519 229293 573585 229296
rect 41146 229146 41152 229210
rect 41216 229208 41222 229210
rect 41775 229208 41841 229211
rect 41216 229206 41841 229208
rect 41216 229150 41780 229206
rect 41836 229150 41841 229206
rect 41216 229148 41841 229150
rect 41216 229146 41222 229148
rect 41775 229145 41841 229148
rect 296559 229208 296625 229211
rect 362799 229208 362865 229211
rect 296559 229206 362865 229208
rect 296559 229150 296564 229206
rect 296620 229150 362804 229206
rect 362860 229150 362865 229206
rect 296559 229148 362865 229150
rect 296559 229145 296625 229148
rect 362799 229145 362865 229148
rect 384399 229208 384465 229211
rect 578895 229208 578961 229211
rect 384399 229206 578961 229208
rect 384399 229150 384404 229206
rect 384460 229150 578900 229206
rect 578956 229150 578961 229206
rect 384399 229148 578961 229150
rect 384399 229145 384465 229148
rect 578895 229145 578961 229148
rect 292143 229060 292209 229063
rect 359823 229060 359889 229063
rect 292143 229058 359889 229060
rect 292143 229002 292148 229058
rect 292204 229002 359828 229058
rect 359884 229002 359889 229058
rect 292143 229000 359889 229002
rect 292143 228997 292209 229000
rect 359823 228997 359889 229000
rect 400239 229060 400305 229063
rect 599919 229060 599985 229063
rect 400239 229058 599985 229060
rect 400239 229002 400244 229058
rect 400300 229002 599924 229058
rect 599980 229002 599985 229058
rect 400239 229000 599985 229002
rect 400239 228997 400305 229000
rect 599919 228997 599985 229000
rect 293103 228912 293169 228915
rect 365679 228912 365745 228915
rect 293103 228910 365745 228912
rect 293103 228854 293108 228910
rect 293164 228854 365684 228910
rect 365740 228854 365745 228910
rect 293103 228852 365745 228854
rect 293103 228849 293169 228852
rect 365679 228849 365745 228852
rect 399471 228912 399537 228915
rect 607503 228912 607569 228915
rect 399471 228910 607569 228912
rect 399471 228854 399476 228910
rect 399532 228854 607508 228910
rect 607564 228854 607569 228910
rect 399471 228852 607569 228854
rect 399471 228849 399537 228852
rect 607503 228849 607569 228852
rect 360783 228764 360849 228767
rect 528303 228764 528369 228767
rect 360783 228762 528369 228764
rect 360783 228706 360788 228762
rect 360844 228706 528308 228762
rect 528364 228706 528369 228762
rect 360783 228704 528369 228706
rect 360783 228701 360849 228704
rect 528303 228701 528369 228704
rect 143874 228172 143934 228660
rect 345423 228616 345489 228619
rect 497967 228616 498033 228619
rect 345423 228614 498033 228616
rect 345423 228558 345428 228614
rect 345484 228558 497972 228614
rect 498028 228558 498033 228614
rect 345423 228556 498033 228558
rect 345423 228553 345489 228556
rect 497967 228553 498033 228556
rect 342159 228468 342225 228471
rect 494223 228468 494289 228471
rect 342159 228466 494289 228468
rect 342159 228410 342164 228466
rect 342220 228410 494228 228466
rect 494284 228410 494289 228466
rect 342159 228408 494289 228410
rect 342159 228405 342225 228408
rect 494223 228405 494289 228408
rect 339375 228320 339441 228323
rect 488271 228320 488337 228323
rect 339375 228318 488337 228320
rect 339375 228262 339380 228318
rect 339436 228262 488276 228318
rect 488332 228262 488337 228318
rect 339375 228260 488337 228262
rect 339375 228257 339441 228260
rect 488271 228257 488337 228260
rect 149391 228172 149457 228175
rect 143874 228170 149457 228172
rect 143874 228114 149396 228170
rect 149452 228114 149457 228170
rect 143874 228112 149457 228114
rect 149391 228109 149457 228112
rect 333039 228172 333105 228175
rect 476175 228172 476241 228175
rect 333039 228170 476241 228172
rect 333039 228114 333044 228170
rect 333100 228114 476180 228170
rect 476236 228114 476241 228170
rect 333039 228112 476241 228114
rect 333039 228109 333105 228112
rect 476175 228109 476241 228112
rect 40378 227370 40384 227434
rect 40448 227432 40454 227434
rect 41775 227432 41841 227435
rect 149391 227432 149457 227435
rect 40448 227430 41841 227432
rect 40448 227374 41780 227430
rect 41836 227374 41841 227430
rect 40448 227372 41841 227374
rect 143904 227430 149457 227432
rect 143904 227374 149396 227430
rect 149452 227374 149457 227430
rect 143904 227372 149457 227374
rect 40448 227370 40454 227372
rect 41775 227369 41841 227372
rect 149391 227369 149457 227372
rect 336879 227432 336945 227435
rect 481455 227432 481521 227435
rect 336879 227430 481521 227432
rect 336879 227374 336884 227430
rect 336940 227374 481460 227430
rect 481516 227374 481521 227430
rect 336879 227372 481521 227374
rect 336879 227369 336945 227372
rect 481455 227369 481521 227372
rect 343119 227284 343185 227287
rect 493455 227284 493521 227287
rect 343119 227282 493521 227284
rect 343119 227226 343124 227282
rect 343180 227226 493460 227282
rect 493516 227226 493521 227282
rect 343119 227224 493521 227226
rect 343119 227221 343185 227224
rect 493455 227221 493521 227224
rect 344751 227136 344817 227139
rect 498831 227136 498897 227139
rect 344751 227134 498897 227136
rect 344751 227078 344756 227134
rect 344812 227078 498836 227134
rect 498892 227078 498897 227134
rect 344751 227076 498897 227078
rect 344751 227073 344817 227076
rect 498831 227073 498897 227076
rect 391599 226988 391665 226991
rect 591663 226988 591729 226991
rect 391599 226986 591729 226988
rect 391599 226930 391604 226986
rect 391660 226930 591668 226986
rect 591724 226930 591729 226986
rect 391599 226928 591729 226930
rect 391599 226925 391665 226928
rect 591663 226925 591729 226928
rect 40762 226778 40768 226842
rect 40832 226840 40838 226842
rect 41775 226840 41841 226843
rect 40832 226838 41841 226840
rect 40832 226782 41780 226838
rect 41836 226782 41841 226838
rect 40832 226780 41841 226782
rect 40832 226778 40838 226780
rect 41775 226777 41841 226780
rect 391215 226840 391281 226843
rect 590895 226840 590961 226843
rect 391215 226838 590961 226840
rect 391215 226782 391220 226838
rect 391276 226782 590900 226838
rect 590956 226782 590961 226838
rect 391215 226780 590961 226782
rect 391215 226777 391281 226780
rect 590895 226777 590961 226780
rect 394095 226692 394161 226695
rect 596175 226692 596241 226695
rect 394095 226690 596241 226692
rect 394095 226634 394100 226690
rect 394156 226634 596180 226690
rect 596236 226634 596241 226690
rect 394095 226632 596241 226634
rect 394095 226629 394161 226632
rect 596175 226629 596241 226632
rect 394479 226544 394545 226547
rect 596943 226544 597009 226547
rect 394479 226542 597009 226544
rect 394479 226486 394484 226542
rect 394540 226486 596948 226542
rect 597004 226486 597009 226542
rect 394479 226484 597009 226486
rect 394479 226481 394545 226484
rect 596943 226481 597009 226484
rect 147183 226396 147249 226399
rect 143904 226394 147249 226396
rect 143904 226338 147188 226394
rect 147244 226338 147249 226394
rect 143904 226336 147249 226338
rect 147183 226333 147249 226336
rect 404367 226396 404433 226399
rect 617295 226396 617361 226399
rect 404367 226394 617361 226396
rect 404367 226338 404372 226394
rect 404428 226338 617300 226394
rect 617356 226338 617361 226394
rect 404367 226336 617361 226338
rect 404367 226333 404433 226336
rect 617295 226333 617361 226336
rect 405807 226248 405873 226251
rect 620367 226248 620433 226251
rect 405807 226246 620433 226248
rect 405807 226190 405812 226246
rect 405868 226190 620372 226246
rect 620428 226190 620433 226246
rect 405807 226188 620433 226190
rect 405807 226185 405873 226188
rect 620367 226185 620433 226188
rect 407631 226100 407697 226103
rect 623343 226100 623409 226103
rect 407631 226098 623409 226100
rect 407631 226042 407636 226098
rect 407692 226042 623348 226098
rect 623404 226042 623409 226098
rect 407631 226040 623409 226042
rect 407631 226037 407697 226040
rect 623343 226037 623409 226040
rect 40570 225890 40576 225954
rect 40640 225952 40646 225954
rect 41775 225952 41841 225955
rect 40640 225950 41841 225952
rect 40640 225894 41780 225950
rect 41836 225894 41841 225950
rect 40640 225892 41841 225894
rect 40640 225890 40646 225892
rect 41775 225889 41841 225892
rect 340143 225952 340209 225955
rect 487503 225952 487569 225955
rect 340143 225950 487569 225952
rect 340143 225894 340148 225950
rect 340204 225894 487508 225950
rect 487564 225894 487569 225950
rect 340143 225892 487569 225894
rect 340143 225889 340209 225892
rect 487503 225889 487569 225892
rect 330831 225804 330897 225807
rect 469359 225804 469425 225807
rect 330831 225802 469425 225804
rect 330831 225746 330836 225802
rect 330892 225746 469364 225802
rect 469420 225746 469425 225802
rect 330831 225744 469425 225746
rect 330831 225741 330897 225744
rect 469359 225741 469425 225744
rect 328047 225656 328113 225659
rect 463311 225656 463377 225659
rect 328047 225654 463377 225656
rect 328047 225598 328052 225654
rect 328108 225598 463316 225654
rect 463372 225598 463377 225654
rect 328047 225596 463377 225598
rect 328047 225593 328113 225596
rect 463311 225593 463377 225596
rect 327279 225508 327345 225511
rect 457263 225508 457329 225511
rect 327279 225506 457329 225508
rect 327279 225450 327284 225506
rect 327340 225450 457268 225506
rect 457324 225450 457329 225506
rect 327279 225448 457329 225450
rect 327279 225445 327345 225448
rect 457263 225445 457329 225448
rect 318927 225360 318993 225363
rect 445167 225360 445233 225363
rect 318927 225358 445233 225360
rect 318927 225302 318932 225358
rect 318988 225302 445172 225358
rect 445228 225302 445233 225358
rect 318927 225300 445233 225302
rect 318927 225297 318993 225300
rect 445167 225297 445233 225300
rect 149391 225212 149457 225215
rect 143904 225210 149457 225212
rect 143904 225154 149396 225210
rect 149452 225154 149457 225210
rect 143904 225152 149457 225154
rect 149391 225149 149457 225152
rect 368655 225212 368721 225215
rect 475311 225212 475377 225215
rect 368655 225210 475377 225212
rect 368655 225154 368660 225210
rect 368716 225154 475316 225210
rect 475372 225154 475377 225210
rect 368655 225152 475377 225154
rect 368655 225149 368721 225152
rect 475311 225149 475377 225152
rect 354063 224620 354129 224623
rect 518415 224620 518481 224623
rect 354063 224618 518481 224620
rect 354063 224562 354068 224618
rect 354124 224562 518420 224618
rect 518476 224562 518481 224618
rect 354063 224560 518481 224562
rect 354063 224557 354129 224560
rect 518415 224557 518481 224560
rect 357231 224472 357297 224475
rect 524463 224472 524529 224475
rect 357231 224470 524529 224472
rect 357231 224414 357236 224470
rect 357292 224414 524468 224470
rect 524524 224414 524529 224470
rect 357231 224412 524529 224414
rect 357231 224409 357297 224412
rect 524463 224409 524529 224412
rect 360303 224324 360369 224327
rect 530511 224324 530577 224327
rect 360303 224322 530577 224324
rect 360303 224266 360308 224322
rect 360364 224266 530516 224322
rect 530572 224266 530577 224322
rect 360303 224264 530577 224266
rect 360303 224261 360369 224264
rect 530511 224261 530577 224264
rect 361455 224176 361521 224179
rect 532047 224176 532113 224179
rect 361455 224174 532113 224176
rect 361455 224118 361460 224174
rect 361516 224118 532052 224174
rect 532108 224118 532113 224174
rect 361455 224116 532113 224118
rect 361455 224113 361521 224116
rect 532047 224113 532113 224116
rect 359727 224028 359793 224031
rect 528975 224028 529041 224031
rect 359727 224026 529041 224028
rect 359727 223970 359732 224026
rect 359788 223970 528980 224026
rect 529036 223970 529041 224026
rect 359727 223968 529041 223970
rect 359727 223965 359793 223968
rect 528975 223965 529041 223968
rect 149487 223880 149553 223883
rect 143904 223878 149553 223880
rect 143904 223822 149492 223878
rect 149548 223822 149553 223878
rect 143904 223820 149553 223822
rect 149487 223817 149553 223820
rect 363759 223880 363825 223883
rect 536559 223880 536625 223883
rect 363759 223878 536625 223880
rect 363759 223822 363764 223878
rect 363820 223822 536564 223878
rect 536620 223822 536625 223878
rect 363759 223820 536625 223822
rect 363759 223817 363825 223820
rect 536559 223817 536625 223820
rect 367599 223732 367665 223735
rect 544047 223732 544113 223735
rect 367599 223730 544113 223732
rect 367599 223674 367604 223730
rect 367660 223674 544052 223730
rect 544108 223674 544113 223730
rect 367599 223672 544113 223674
rect 367599 223669 367665 223672
rect 544047 223669 544113 223672
rect 377583 223584 377649 223587
rect 562959 223584 563025 223587
rect 377583 223582 563025 223584
rect 377583 223526 377588 223582
rect 377644 223526 562964 223582
rect 563020 223526 563025 223582
rect 377583 223524 563025 223526
rect 377583 223521 377649 223524
rect 562959 223521 563025 223524
rect 376719 223436 376785 223439
rect 562191 223436 562257 223439
rect 376719 223434 562257 223436
rect 376719 223378 376724 223434
rect 376780 223378 562196 223434
rect 562252 223378 562257 223434
rect 376719 223376 562257 223378
rect 376719 223373 376785 223376
rect 562191 223373 562257 223376
rect 381231 223288 381297 223291
rect 571311 223288 571377 223291
rect 381231 223286 571377 223288
rect 381231 223230 381236 223286
rect 381292 223230 571316 223286
rect 571372 223230 571377 223286
rect 381231 223228 571377 223230
rect 381231 223225 381297 223228
rect 571311 223225 571377 223228
rect 384303 223140 384369 223143
rect 577263 223140 577329 223143
rect 384303 223138 577329 223140
rect 384303 223082 384308 223138
rect 384364 223082 577268 223138
rect 577324 223082 577329 223138
rect 384303 223080 577329 223082
rect 384303 223077 384369 223080
rect 577263 223077 577329 223080
rect 358575 222992 358641 222995
rect 525999 222992 526065 222995
rect 358575 222990 526065 222992
rect 358575 222934 358580 222990
rect 358636 222934 526004 222990
rect 526060 222934 526065 222990
rect 358575 222932 526065 222934
rect 358575 222929 358641 222932
rect 525999 222929 526065 222932
rect 359439 222844 359505 222847
rect 526671 222844 526737 222847
rect 359439 222842 526737 222844
rect 359439 222786 359444 222842
rect 359500 222786 526676 222842
rect 526732 222786 526737 222842
rect 359439 222784 526737 222786
rect 359439 222781 359505 222784
rect 526671 222781 526737 222784
rect 149391 222696 149457 222699
rect 143904 222694 149457 222696
rect 143904 222638 149396 222694
rect 149452 222638 149457 222694
rect 143904 222636 149457 222638
rect 149391 222633 149457 222636
rect 355599 222696 355665 222699
rect 519855 222696 519921 222699
rect 355599 222694 519921 222696
rect 355599 222638 355604 222694
rect 355660 222638 519860 222694
rect 519916 222638 519921 222694
rect 355599 222636 519921 222638
rect 355599 222633 355665 222636
rect 519855 222633 519921 222636
rect 406479 222548 406545 222551
rect 522927 222548 522993 222551
rect 406479 222546 522993 222548
rect 406479 222490 406484 222546
rect 406540 222490 522932 222546
rect 522988 222490 522993 222546
rect 406479 222488 522993 222490
rect 406479 222485 406545 222488
rect 522927 222485 522993 222488
rect 676290 221811 676350 222074
rect 676239 221806 676350 221811
rect 676239 221750 676244 221806
rect 676300 221750 676350 221806
rect 676239 221748 676350 221750
rect 676239 221745 676305 221748
rect 146895 221512 146961 221515
rect 143904 221510 146961 221512
rect 143904 221454 146900 221510
rect 146956 221454 146961 221510
rect 143904 221452 146961 221454
rect 146895 221449 146961 221452
rect 676143 221216 676209 221219
rect 676290 221216 676350 221482
rect 676143 221214 676350 221216
rect 676143 221158 676148 221214
rect 676204 221158 676350 221214
rect 676143 221156 676350 221158
rect 676143 221153 676209 221156
rect 186927 221068 186993 221071
rect 186927 221066 190560 221068
rect 186927 221010 186932 221066
rect 186988 221010 190560 221066
rect 186927 221008 190560 221010
rect 186927 221005 186993 221008
rect 676290 220775 676350 221038
rect 676239 220770 676350 220775
rect 676239 220714 676244 220770
rect 676300 220714 676350 220770
rect 676239 220712 676350 220714
rect 676239 220709 676305 220712
rect 185583 220328 185649 220331
rect 185583 220326 190560 220328
rect 185583 220270 185588 220326
rect 185644 220270 190560 220326
rect 185583 220268 190560 220270
rect 185583 220265 185649 220268
rect 143874 219736 143934 220224
rect 149391 219736 149457 219739
rect 143874 219734 149457 219736
rect 143874 219678 149396 219734
rect 149452 219678 149457 219734
rect 143874 219676 149457 219678
rect 149391 219673 149457 219676
rect 184335 219588 184401 219591
rect 184335 219586 190560 219588
rect 184335 219530 184340 219586
rect 184396 219530 190560 219586
rect 184335 219528 190560 219530
rect 184335 219525 184401 219528
rect 147663 218996 147729 218999
rect 143904 218994 147729 218996
rect 143904 218938 147668 218994
rect 147724 218938 147729 218994
rect 143904 218936 147729 218938
rect 147663 218933 147729 218936
rect 184335 218848 184401 218851
rect 184335 218846 190560 218848
rect 184335 218790 184340 218846
rect 184396 218790 190560 218846
rect 184335 218788 190560 218790
rect 184335 218785 184401 218788
rect 639810 218670 639870 220594
rect 674170 220562 674176 220626
rect 674240 220624 674246 220626
rect 674240 220564 676320 220624
rect 674240 220562 674246 220564
rect 674170 219970 674176 220034
rect 674240 220032 674246 220034
rect 674240 219972 676320 220032
rect 674240 219970 674246 219972
rect 676047 219514 676113 219517
rect 676047 219512 676320 219514
rect 676047 219456 676052 219512
rect 676108 219456 676320 219512
rect 676047 219454 676320 219456
rect 676047 219451 676113 219454
rect 673978 219082 673984 219146
rect 674048 219144 674054 219146
rect 674362 219144 674368 219146
rect 674048 219084 674368 219144
rect 674048 219082 674054 219084
rect 674362 219082 674368 219084
rect 674432 219144 674438 219146
rect 674432 219084 676320 219144
rect 674432 219082 674438 219084
rect 674554 218490 674560 218554
rect 674624 218552 674630 218554
rect 674624 218492 676320 218552
rect 674624 218490 674630 218492
rect 186831 218108 186897 218111
rect 186831 218106 190560 218108
rect 186831 218050 186836 218106
rect 186892 218050 190560 218106
rect 186831 218048 190560 218050
rect 186831 218045 186897 218048
rect 149391 217812 149457 217815
rect 143904 217810 149457 217812
rect 143904 217754 149396 217810
rect 149452 217754 149457 217810
rect 143904 217752 149457 217754
rect 149391 217749 149457 217752
rect 190146 217294 190206 218048
rect 674362 217898 674368 217962
rect 674432 217960 674438 217962
rect 675322 217960 675328 217962
rect 674432 217900 675328 217960
rect 674432 217898 674438 217900
rect 675322 217898 675328 217900
rect 675392 217960 675398 217962
rect 675392 217900 676320 217960
rect 675392 217898 675398 217900
rect 675706 217602 675712 217666
rect 675776 217664 675782 217666
rect 675776 217604 676320 217664
rect 675776 217602 675782 217604
rect 190146 217234 190560 217294
rect 676866 216779 676926 217042
rect 676866 216774 676977 216779
rect 149487 216628 149553 216631
rect 143904 216626 149553 216628
rect 143904 216570 149492 216626
rect 149548 216570 149553 216626
rect 143904 216568 149553 216570
rect 149487 216565 149553 216568
rect 187023 216480 187089 216483
rect 187023 216478 190560 216480
rect 187023 216422 187028 216478
rect 187084 216422 190560 216478
rect 187023 216420 190560 216422
rect 187023 216417 187089 216420
rect 190146 215814 190206 216420
rect 190146 215754 190560 215814
rect 143874 214852 143934 215340
rect 186255 215000 186321 215003
rect 186255 214998 190560 215000
rect 186255 214942 186260 214998
rect 186316 214942 190560 214998
rect 186255 214940 190560 214942
rect 186255 214937 186321 214940
rect 149391 214852 149457 214855
rect 143874 214850 149457 214852
rect 143874 214794 149396 214850
rect 149452 214794 149457 214850
rect 143874 214792 149457 214794
rect 149391 214789 149457 214792
rect 190146 214334 190206 214940
rect 640386 214822 640446 216746
rect 676866 216718 676916 216774
rect 676972 216718 676977 216774
rect 676866 216716 676977 216718
rect 676911 216713 676977 216716
rect 675759 216480 675825 216483
rect 675759 216478 676320 216480
rect 675759 216422 675764 216478
rect 675820 216422 676320 216478
rect 675759 216420 676320 216422
rect 675759 216417 675825 216420
rect 676047 216110 676113 216113
rect 676047 216108 676320 216110
rect 676047 216052 676052 216108
rect 676108 216052 676320 216108
rect 676047 216050 676320 216052
rect 676047 216047 676113 216050
rect 675898 215530 675904 215594
rect 675968 215592 675974 215594
rect 675968 215532 676320 215592
rect 675968 215530 675974 215532
rect 676866 214855 676926 214970
rect 676815 214850 676926 214855
rect 676815 214794 676820 214850
rect 676876 214794 676926 214850
rect 676815 214792 676926 214794
rect 676815 214789 676881 214792
rect 676047 214630 676113 214633
rect 676047 214628 676320 214630
rect 676047 214572 676052 214628
rect 676108 214572 676320 214628
rect 676047 214570 676320 214572
rect 676047 214567 676113 214570
rect 190146 214274 190560 214334
rect 147087 214112 147153 214115
rect 143904 214110 147153 214112
rect 143904 214054 147092 214110
rect 147148 214054 147153 214110
rect 143904 214052 147153 214054
rect 147087 214049 147153 214052
rect 675951 214112 676017 214115
rect 675951 214110 676320 214112
rect 675951 214054 675956 214110
rect 676012 214054 676320 214110
rect 675951 214052 676320 214054
rect 675951 214049 676017 214052
rect 186447 213520 186513 213523
rect 186447 213518 190560 213520
rect 186447 213462 186452 213518
rect 186508 213462 190560 213518
rect 186447 213460 190560 213462
rect 186447 213457 186513 213460
rect 41775 213298 41841 213301
rect 41568 213296 41841 213298
rect 41568 213240 41780 213296
rect 41836 213240 41841 213296
rect 41568 213238 41841 213240
rect 41775 213235 41841 213238
rect 41583 212928 41649 212931
rect 146895 212928 146961 212931
rect 41538 212926 41649 212928
rect 41538 212870 41588 212926
rect 41644 212870 41649 212926
rect 41538 212865 41649 212870
rect 143904 212926 146961 212928
rect 143904 212870 146900 212926
rect 146956 212870 146961 212926
rect 143904 212868 146961 212870
rect 146895 212865 146961 212868
rect 41538 212750 41598 212865
rect 190146 212706 190206 213460
rect 676290 213375 676350 213490
rect 676239 213370 676350 213375
rect 676239 213314 676244 213370
rect 676300 213314 676350 213370
rect 676239 213312 676350 213314
rect 676239 213309 676305 213312
rect 674554 213014 674560 213078
rect 674624 213076 674630 213078
rect 674624 213016 676320 213076
rect 674624 213014 674630 213016
rect 190146 212646 190560 212706
rect 640194 212339 640254 212898
rect 676047 212632 676113 212635
rect 676047 212630 676320 212632
rect 676047 212574 676052 212630
rect 676108 212574 676320 212630
rect 676047 212572 676320 212574
rect 676047 212569 676113 212572
rect 640143 212334 640254 212339
rect 640143 212278 640148 212334
rect 640204 212278 640254 212334
rect 640143 212276 640254 212278
rect 640143 212273 640209 212276
rect 41775 212188 41841 212191
rect 41568 212186 41841 212188
rect 41568 212130 41780 212186
rect 41836 212130 41841 212186
rect 41568 212128 41841 212130
rect 41775 212125 41841 212128
rect 186063 212040 186129 212043
rect 676047 212040 676113 212043
rect 186063 212038 190560 212040
rect 186063 211982 186068 212038
rect 186124 211982 190560 212038
rect 186063 211980 190560 211982
rect 676047 212038 676320 212040
rect 676047 211982 676052 212038
rect 676108 211982 676320 212038
rect 676047 211980 676320 211982
rect 186063 211977 186129 211980
rect 41775 211744 41841 211747
rect 147375 211744 147441 211747
rect 41568 211742 41841 211744
rect 41568 211686 41780 211742
rect 41836 211686 41841 211742
rect 41568 211684 41841 211686
rect 143904 211742 147441 211744
rect 143904 211686 147380 211742
rect 147436 211686 147441 211742
rect 143904 211684 147441 211686
rect 41775 211681 41841 211684
rect 147375 211681 147441 211684
rect 41583 211448 41649 211451
rect 41538 211446 41649 211448
rect 41538 211390 41588 211446
rect 41644 211390 41649 211446
rect 41538 211385 41649 211390
rect 41538 211270 41598 211385
rect 190146 211152 190206 211980
rect 676047 211977 676113 211980
rect 640143 211596 640209 211599
rect 640143 211594 640254 211596
rect 640143 211538 640148 211594
rect 640204 211538 640254 211594
rect 640143 211533 640254 211538
rect 190146 211092 190560 211152
rect 640194 210974 640254 211533
rect 676290 211451 676350 211566
rect 676239 211446 676350 211451
rect 676239 211390 676244 211446
rect 676300 211390 676350 211446
rect 676239 211388 676350 211390
rect 676239 211385 676305 211388
rect 675951 211078 676017 211081
rect 675951 211076 676320 211078
rect 675951 211020 675956 211076
rect 676012 211020 676320 211076
rect 675951 211018 676320 211020
rect 675951 211015 676017 211018
rect 41775 210708 41841 210711
rect 679791 210708 679857 210711
rect 41568 210706 41841 210708
rect 41568 210650 41780 210706
rect 41836 210650 41841 210706
rect 41568 210648 41841 210650
rect 41775 210645 41841 210648
rect 679746 210706 679857 210708
rect 679746 210650 679796 210706
rect 679852 210650 679857 210706
rect 679746 210645 679857 210650
rect 186639 210560 186705 210563
rect 186639 210558 190014 210560
rect 186639 210502 186644 210558
rect 186700 210502 190014 210558
rect 679746 210530 679806 210645
rect 186639 210500 190014 210502
rect 186639 210497 186705 210500
rect 189954 210486 190014 210500
rect 189954 210426 190560 210486
rect 147471 210412 147537 210415
rect 143904 210410 147537 210412
rect 143904 210354 147476 210410
rect 147532 210354 147537 210410
rect 143904 210352 147537 210354
rect 147471 210349 147537 210352
rect 41775 210264 41841 210267
rect 41568 210262 41841 210264
rect 41568 210206 41780 210262
rect 41836 210206 41841 210262
rect 41568 210204 41841 210206
rect 41775 210201 41841 210204
rect 41583 209968 41649 209971
rect 41538 209966 41649 209968
rect 41538 209910 41588 209966
rect 41644 209910 41649 209966
rect 41538 209905 41649 209910
rect 41538 209790 41598 209905
rect 190146 209672 190206 210426
rect 685506 209823 685566 210086
rect 679791 209820 679857 209823
rect 679746 209818 679857 209820
rect 679746 209762 679796 209818
rect 679852 209762 679857 209818
rect 679746 209757 679857 209762
rect 685455 209818 685566 209823
rect 685455 209762 685460 209818
rect 685516 209762 685566 209818
rect 685455 209760 685566 209762
rect 685455 209757 685521 209760
rect 190146 209612 190560 209672
rect 679746 209568 679806 209757
rect 41583 209376 41649 209379
rect 41538 209374 41649 209376
rect 41538 209318 41588 209374
rect 41644 209318 41649 209374
rect 41538 209313 41649 209318
rect 685455 209376 685521 209379
rect 685455 209374 685566 209376
rect 685455 209318 685460 209374
rect 685516 209318 685566 209374
rect 685455 209313 685566 209318
rect 41538 209198 41598 209313
rect 146895 209228 146961 209231
rect 143904 209226 146961 209228
rect 143904 209170 146900 209226
rect 146956 209170 146961 209226
rect 143904 209168 146961 209170
rect 146895 209165 146961 209168
rect 186735 209080 186801 209083
rect 186735 209078 190014 209080
rect 186735 209022 186740 209078
rect 186796 209022 190014 209078
rect 186735 209020 190014 209022
rect 186735 209017 186801 209020
rect 189954 209006 190014 209020
rect 189954 208946 190560 209006
rect 40386 208490 40446 208754
rect 40378 208426 40384 208490
rect 40448 208426 40454 208490
rect 41775 208266 41841 208269
rect 41568 208264 41841 208266
rect 41568 208208 41780 208264
rect 41836 208208 41841 208264
rect 41568 208206 41841 208208
rect 41775 208203 41841 208206
rect 190146 208192 190206 208946
rect 190146 208132 190560 208192
rect 147183 208044 147249 208047
rect 143904 208042 147249 208044
rect 143904 207986 147188 208042
rect 147244 207986 147249 208042
rect 143904 207984 147249 207986
rect 147183 207981 147249 207984
rect 40570 207834 40576 207898
rect 40640 207834 40646 207898
rect 40578 207718 40638 207834
rect 189954 207318 190560 207378
rect 186351 207304 186417 207307
rect 189954 207304 190014 207318
rect 186351 207302 190014 207304
rect 40962 207010 41022 207274
rect 186351 207246 186356 207302
rect 186412 207246 190014 207302
rect 639810 207274 639870 209124
rect 685506 209050 685566 209313
rect 676666 207538 676672 207602
rect 676736 207600 676742 207602
rect 676815 207600 676881 207603
rect 676736 207598 676881 207600
rect 676736 207542 676820 207598
rect 676876 207542 676881 207598
rect 676736 207540 676881 207542
rect 676736 207538 676742 207540
rect 676815 207537 676881 207540
rect 676474 207390 676480 207454
rect 676544 207452 676550 207454
rect 676911 207452 676977 207455
rect 676544 207450 676977 207452
rect 676544 207394 676916 207450
rect 676972 207394 676977 207450
rect 676544 207392 676977 207394
rect 676544 207390 676550 207392
rect 676911 207389 676977 207392
rect 186351 207244 190014 207246
rect 186351 207241 186417 207244
rect 40954 206946 40960 207010
rect 41024 206946 41030 207010
rect 34050 206567 34110 206682
rect 34050 206562 34161 206567
rect 34050 206506 34100 206562
rect 34156 206506 34161 206562
rect 34050 206504 34161 206506
rect 34095 206501 34161 206504
rect 143874 206416 143934 206904
rect 189954 206712 190014 207244
rect 189954 206652 190560 206712
rect 147279 206416 147345 206419
rect 143874 206414 147345 206416
rect 143874 206358 147284 206414
rect 147340 206358 147345 206414
rect 143874 206356 147345 206358
rect 147279 206353 147345 206356
rect 42255 206268 42321 206271
rect 41568 206266 42321 206268
rect 41568 206210 42260 206266
rect 42316 206210 42321 206266
rect 41568 206208 42321 206210
rect 42255 206205 42321 206208
rect 186543 205972 186609 205975
rect 186543 205970 190014 205972
rect 186543 205914 186548 205970
rect 186604 205914 190014 205970
rect 186543 205912 190014 205914
rect 186543 205909 186609 205912
rect 189954 205898 190014 205912
rect 189954 205838 190560 205898
rect 40770 205530 40830 205794
rect 149391 205676 149457 205679
rect 143904 205674 149457 205676
rect 143904 205618 149396 205674
rect 149452 205618 149457 205674
rect 143904 205616 149457 205618
rect 149391 205613 149457 205616
rect 40762 205466 40768 205530
rect 40832 205466 40838 205530
rect 190146 205232 190206 205838
rect 41154 204938 41214 205202
rect 190146 205172 190560 205232
rect 41146 204874 41152 204938
rect 41216 204874 41222 204938
rect 34242 204495 34302 204758
rect 34191 204490 34302 204495
rect 149295 204492 149361 204495
rect 34191 204434 34196 204490
rect 34252 204434 34302 204490
rect 34191 204432 34302 204434
rect 143904 204490 149361 204492
rect 143904 204434 149300 204490
rect 149356 204434 149361 204490
rect 143904 204432 149361 204434
rect 34191 204429 34257 204432
rect 149295 204429 149361 204432
rect 185967 204344 186033 204347
rect 185967 204342 190560 204344
rect 34242 204051 34302 204314
rect 185967 204286 185972 204342
rect 186028 204286 190560 204342
rect 185967 204284 190560 204286
rect 185967 204281 186033 204284
rect 34242 204046 34353 204051
rect 34242 203990 34292 204046
rect 34348 203990 34353 204046
rect 34242 203988 34353 203990
rect 34287 203985 34353 203988
rect 41538 203607 41598 203722
rect 41538 203602 41649 203607
rect 41538 203546 41588 203602
rect 41644 203546 41649 203602
rect 41538 203544 41649 203546
rect 190146 203604 190206 204284
rect 190146 203544 190560 203604
rect 41583 203541 41649 203544
rect 639810 203426 639870 205350
rect 675663 204494 675729 204495
rect 675663 204490 675712 204494
rect 675776 204492 675782 204494
rect 675663 204434 675668 204490
rect 675663 204430 675712 204434
rect 675776 204432 675820 204492
rect 675776 204430 675782 204432
rect 675663 204429 675729 204430
rect 149487 203308 149553 203311
rect 143904 203306 149553 203308
rect 143904 203250 149492 203306
rect 149548 203250 149553 203306
rect 143904 203248 149553 203250
rect 149487 203245 149553 203248
rect 34434 203015 34494 203204
rect 34434 203010 34545 203015
rect 34434 202954 34484 203010
rect 34540 202954 34545 203010
rect 34434 202952 34545 202954
rect 34479 202949 34545 202952
rect 41871 202864 41937 202867
rect 41568 202862 41937 202864
rect 41568 202806 41876 202862
rect 41932 202806 41937 202862
rect 41568 202804 41937 202806
rect 41871 202801 41937 202804
rect 186159 202864 186225 202867
rect 186159 202862 190560 202864
rect 186159 202806 186164 202862
rect 186220 202806 190560 202862
rect 186159 202804 190560 202806
rect 186159 202801 186225 202804
rect 34434 201979 34494 202242
rect 190146 202124 190206 202804
rect 190146 202064 190560 202124
rect 34383 201974 34494 201979
rect 34383 201918 34388 201974
rect 34444 201918 34494 201974
rect 34383 201916 34494 201918
rect 143874 201976 143934 202020
rect 149391 201976 149457 201979
rect 143874 201974 149457 201976
rect 143874 201918 149396 201974
rect 149452 201918 149457 201974
rect 143874 201916 149457 201918
rect 34383 201913 34449 201916
rect 149391 201913 149457 201916
rect 41967 201680 42033 201683
rect 41568 201678 42033 201680
rect 41568 201622 41972 201678
rect 42028 201622 42033 201678
rect 41568 201620 42033 201622
rect 41967 201617 42033 201620
rect 41583 201532 41649 201535
rect 41538 201530 41649 201532
rect 41538 201474 41588 201530
rect 41644 201474 41649 201530
rect 41538 201469 41649 201474
rect 41538 201354 41598 201469
rect 190287 201384 190353 201387
rect 190287 201382 190560 201384
rect 190287 201326 190292 201382
rect 190348 201326 190560 201382
rect 190287 201324 190560 201326
rect 190287 201321 190353 201324
rect 640194 200943 640254 201502
rect 41583 200940 41649 200943
rect 41538 200938 41649 200940
rect 41538 200882 41588 200938
rect 41644 200882 41649 200938
rect 41538 200877 41649 200882
rect 640143 200938 640254 200943
rect 640143 200882 640148 200938
rect 640204 200882 640254 200938
rect 640143 200880 640254 200882
rect 640143 200877 640209 200880
rect 41538 200762 41598 200877
rect 149391 200792 149457 200795
rect 143904 200790 149457 200792
rect 143904 200734 149396 200790
rect 149452 200734 149457 200790
rect 143904 200732 149457 200734
rect 149391 200729 149457 200732
rect 190287 200570 190353 200573
rect 190287 200568 190560 200570
rect 190287 200512 190292 200568
rect 190348 200512 190560 200568
rect 190287 200510 190560 200512
rect 190287 200507 190353 200510
rect 640143 200200 640209 200203
rect 640143 200198 640254 200200
rect 640143 200142 640148 200198
rect 640204 200142 640254 200198
rect 640143 200137 640254 200142
rect 185967 199756 186033 199759
rect 185967 199754 190560 199756
rect 185967 199698 185972 199754
rect 186028 199698 190560 199754
rect 185967 199696 190560 199698
rect 185967 199693 186033 199696
rect 147471 199608 147537 199611
rect 143904 199606 147537 199608
rect 143904 199550 147476 199606
rect 147532 199550 147537 199606
rect 640194 199578 640254 200137
rect 143904 199548 147537 199550
rect 147471 199545 147537 199548
rect 187215 199164 187281 199167
rect 187215 199162 190014 199164
rect 187215 199106 187220 199162
rect 187276 199106 190014 199162
rect 187215 199104 190014 199106
rect 187215 199101 187281 199104
rect 189954 199090 190014 199104
rect 189954 199030 190560 199090
rect 149487 198424 149553 198427
rect 143904 198422 149553 198424
rect 143904 198366 149492 198422
rect 149548 198366 149553 198422
rect 143904 198364 149553 198366
rect 149487 198361 149553 198364
rect 675759 198424 675825 198427
rect 675898 198424 675904 198426
rect 675759 198422 675904 198424
rect 675759 198366 675764 198422
rect 675820 198366 675904 198422
rect 675759 198364 675904 198366
rect 675759 198361 675825 198364
rect 675898 198362 675904 198364
rect 675968 198362 675974 198426
rect 185487 198276 185553 198279
rect 185487 198274 190560 198276
rect 185487 198218 185492 198274
rect 185548 198218 190560 198274
rect 185487 198216 190560 198218
rect 185487 198213 185553 198216
rect 184239 197684 184305 197687
rect 184239 197682 190014 197684
rect 184239 197626 184244 197682
rect 184300 197626 190014 197682
rect 184239 197624 190014 197626
rect 184239 197621 184305 197624
rect 189954 197610 190014 197624
rect 189954 197550 190560 197610
rect 149391 197092 149457 197095
rect 143904 197090 149457 197092
rect 143904 197034 149396 197090
rect 149452 197034 149457 197090
rect 143904 197032 149457 197034
rect 149391 197029 149457 197032
rect 185967 196796 186033 196799
rect 185967 196794 190560 196796
rect 185967 196738 185972 196794
rect 186028 196738 190560 196794
rect 185967 196736 190560 196738
rect 185967 196733 186033 196736
rect 186063 196056 186129 196059
rect 186063 196054 190560 196056
rect 186063 195998 186068 196054
rect 186124 195998 190560 196054
rect 186063 195996 190560 195998
rect 186063 195993 186129 195996
rect 149391 195908 149457 195911
rect 143904 195906 149457 195908
rect 143904 195850 149396 195906
rect 149452 195850 149457 195906
rect 143904 195848 149457 195850
rect 149391 195845 149457 195848
rect 639810 195730 639870 197654
rect 184335 195316 184401 195319
rect 184335 195314 190560 195316
rect 184335 195258 184340 195314
rect 184396 195258 190560 195314
rect 184335 195256 190560 195258
rect 184335 195253 184401 195256
rect 674554 194810 674560 194874
rect 674624 194872 674630 194874
rect 675087 194872 675153 194875
rect 674624 194870 675153 194872
rect 674624 194814 675092 194870
rect 675148 194814 675153 194870
rect 674624 194812 675153 194814
rect 674624 194810 674630 194812
rect 675087 194809 675153 194812
rect 149487 194724 149553 194727
rect 143904 194722 149553 194724
rect 143904 194666 149492 194722
rect 149548 194666 149553 194722
rect 143904 194664 149553 194666
rect 149487 194661 149553 194664
rect 184431 194428 184497 194431
rect 184431 194426 190560 194428
rect 184431 194370 184436 194426
rect 184492 194370 190560 194426
rect 184431 194368 190560 194370
rect 184431 194365 184497 194368
rect 184527 193836 184593 193839
rect 184527 193834 190014 193836
rect 184527 193778 184532 193834
rect 184588 193778 190014 193834
rect 184527 193776 190014 193778
rect 184527 193773 184593 193776
rect 189954 193762 190014 193776
rect 189954 193702 190560 193762
rect 143874 193392 143934 193436
rect 149391 193392 149457 193395
rect 143874 193390 149457 193392
rect 143874 193334 149396 193390
rect 149452 193334 149457 193390
rect 143874 193332 149457 193334
rect 149391 193329 149457 193332
rect 184431 192948 184497 192951
rect 184431 192946 190560 192948
rect 184431 192890 184436 192946
rect 184492 192890 190560 192946
rect 184431 192888 190560 192890
rect 184431 192885 184497 192888
rect 184335 192356 184401 192359
rect 184335 192354 190014 192356
rect 184335 192298 184340 192354
rect 184396 192298 190014 192354
rect 184335 192296 190014 192298
rect 184335 192293 184401 192296
rect 189954 192282 190014 192296
rect 189954 192222 190560 192282
rect 149391 192208 149457 192211
rect 143904 192206 149457 192208
rect 143904 192150 149396 192206
rect 149452 192150 149457 192206
rect 143904 192148 149457 192150
rect 149391 192145 149457 192148
rect 639810 192030 639870 193880
rect 675759 193540 675825 193543
rect 676474 193540 676480 193542
rect 675759 193538 676480 193540
rect 675759 193482 675764 193538
rect 675820 193482 676480 193538
rect 675759 193480 676480 193482
rect 675759 193477 675825 193480
rect 676474 193478 676480 193480
rect 676544 193478 676550 193542
rect 675759 191616 675825 191619
rect 676666 191616 676672 191618
rect 675759 191614 676672 191616
rect 675759 191558 675764 191614
rect 675820 191558 676672 191614
rect 675759 191556 676672 191558
rect 675759 191553 675825 191556
rect 676666 191554 676672 191556
rect 676736 191554 676742 191618
rect 184527 191468 184593 191471
rect 184527 191466 190560 191468
rect 184527 191410 184532 191466
rect 184588 191410 190560 191466
rect 184527 191408 190560 191410
rect 184527 191405 184593 191408
rect 147375 191024 147441 191027
rect 143904 191022 147441 191024
rect 143904 190966 147380 191022
rect 147436 190966 147441 191022
rect 143904 190964 147441 190966
rect 147375 190961 147441 190964
rect 184623 190728 184689 190731
rect 184623 190726 190014 190728
rect 184623 190670 184628 190726
rect 184684 190670 190014 190726
rect 184623 190668 190014 190670
rect 184623 190665 184689 190668
rect 189954 190654 190014 190668
rect 189954 190594 190560 190654
rect 184335 189988 184401 189991
rect 184335 189986 190560 189988
rect 184335 189930 184340 189986
rect 184396 189930 190560 189986
rect 184335 189928 190560 189930
rect 184335 189925 184401 189928
rect 149391 189840 149457 189843
rect 143904 189838 149457 189840
rect 143904 189782 149396 189838
rect 149452 189782 149457 189838
rect 143904 189780 149457 189782
rect 149391 189777 149457 189780
rect 184527 189248 184593 189251
rect 184527 189246 190014 189248
rect 184527 189190 184532 189246
rect 184588 189190 190014 189246
rect 184527 189188 190014 189190
rect 184527 189185 184593 189188
rect 189954 189174 190014 189188
rect 189954 189114 190560 189174
rect 143874 188064 143934 188552
rect 184335 188508 184401 188511
rect 184335 188506 190560 188508
rect 184335 188450 184340 188506
rect 184396 188450 190560 188506
rect 184335 188448 190560 188450
rect 184335 188445 184401 188448
rect 639810 188182 639870 190106
rect 149487 188064 149553 188067
rect 143874 188062 149553 188064
rect 143874 188006 149492 188062
rect 149548 188006 149553 188062
rect 143874 188004 149553 188006
rect 149487 188001 149553 188004
rect 184431 187620 184497 187623
rect 184431 187618 190560 187620
rect 184431 187562 184436 187618
rect 184492 187562 190560 187618
rect 184431 187560 190560 187562
rect 184431 187557 184497 187560
rect 149295 187472 149361 187475
rect 143904 187470 149361 187472
rect 143904 187414 149300 187470
rect 149356 187414 149361 187470
rect 143904 187412 149361 187414
rect 149295 187409 149361 187412
rect 184335 186880 184401 186883
rect 184335 186878 190560 186880
rect 184335 186822 184340 186878
rect 184396 186822 190560 186878
rect 184335 186820 190560 186822
rect 184335 186817 184401 186820
rect 41146 186670 41152 186734
rect 41216 186732 41222 186734
rect 41775 186732 41841 186735
rect 41216 186730 41841 186732
rect 41216 186674 41780 186730
rect 41836 186674 41841 186730
rect 41216 186672 41841 186674
rect 41216 186670 41222 186672
rect 41775 186669 41841 186672
rect 149199 186288 149265 186291
rect 143904 186286 149265 186288
rect 143904 186230 149204 186286
rect 149260 186230 149265 186286
rect 143904 186228 149265 186230
rect 149199 186225 149265 186228
rect 184431 186140 184497 186143
rect 184431 186138 190560 186140
rect 184431 186082 184436 186138
rect 184492 186082 190560 186138
rect 184431 186080 190560 186082
rect 184431 186077 184497 186080
rect 40954 185782 40960 185846
rect 41024 185844 41030 185846
rect 41775 185844 41841 185847
rect 41024 185842 41841 185844
rect 41024 185786 41780 185842
rect 41836 185786 41841 185842
rect 41024 185784 41841 185786
rect 41024 185782 41030 185784
rect 41775 185781 41841 185784
rect 640194 185699 640254 186258
rect 640194 185694 640305 185699
rect 640194 185638 640244 185694
rect 640300 185638 640305 185694
rect 640194 185636 640305 185638
rect 640239 185633 640305 185636
rect 184623 185400 184689 185403
rect 184623 185398 190014 185400
rect 184623 185342 184628 185398
rect 184684 185342 190014 185398
rect 184623 185340 190014 185342
rect 184623 185337 184689 185340
rect 189954 185326 190014 185340
rect 189954 185266 190560 185326
rect 143874 184512 143934 185000
rect 640239 184956 640305 184959
rect 640194 184954 640305 184956
rect 640194 184898 640244 184954
rect 640300 184898 640305 184954
rect 640194 184893 640305 184898
rect 184527 184660 184593 184663
rect 184527 184658 190560 184660
rect 184527 184602 184532 184658
rect 184588 184602 190560 184658
rect 184527 184600 190560 184602
rect 184527 184597 184593 184600
rect 149583 184512 149649 184515
rect 143874 184510 149649 184512
rect 143874 184454 149588 184510
rect 149644 184454 149649 184510
rect 143874 184452 149649 184454
rect 149583 184449 149649 184452
rect 640194 184334 640254 184893
rect 40378 184154 40384 184218
rect 40448 184216 40454 184218
rect 41775 184216 41841 184219
rect 40448 184214 41841 184216
rect 40448 184158 41780 184214
rect 41836 184158 41841 184214
rect 40448 184156 41841 184158
rect 40448 184154 40454 184156
rect 41775 184153 41841 184156
rect 184335 183920 184401 183923
rect 184335 183918 190014 183920
rect 184335 183862 184340 183918
rect 184396 183862 190014 183918
rect 184335 183860 190014 183862
rect 184335 183857 184401 183860
rect 189954 183846 190014 183860
rect 189954 183786 190560 183846
rect 149391 183772 149457 183775
rect 143904 183770 149457 183772
rect 143904 183714 149396 183770
rect 149452 183714 149457 183770
rect 143904 183712 149457 183714
rect 149391 183709 149457 183712
rect 40762 183562 40768 183626
rect 40832 183624 40838 183626
rect 41775 183624 41841 183627
rect 40832 183622 41841 183624
rect 40832 183566 41780 183622
rect 41836 183566 41841 183622
rect 40832 183564 41841 183566
rect 40832 183562 40838 183564
rect 41775 183561 41841 183564
rect 186735 183180 186801 183183
rect 186735 183178 190560 183180
rect 186735 183122 186740 183178
rect 186796 183122 190560 183178
rect 186735 183120 190560 183122
rect 186735 183117 186801 183120
rect 645135 183032 645201 183035
rect 640386 183030 645201 183032
rect 640386 182974 645140 183030
rect 645196 182974 645201 183030
rect 640386 182972 645201 182974
rect 40570 182822 40576 182886
rect 40640 182884 40646 182886
rect 41775 182884 41841 182887
rect 40640 182882 41841 182884
rect 40640 182826 41780 182882
rect 41836 182826 41841 182882
rect 40640 182824 41841 182826
rect 40640 182822 40646 182824
rect 41775 182821 41841 182824
rect 149487 182588 149553 182591
rect 143904 182586 149553 182588
rect 143904 182530 149492 182586
rect 149548 182530 149553 182586
rect 143904 182528 149553 182530
rect 149487 182525 149553 182528
rect 185775 182440 185841 182443
rect 640386 182440 640446 182972
rect 645135 182969 645201 182972
rect 185775 182438 190014 182440
rect 185775 182382 185780 182438
rect 185836 182382 190014 182438
rect 640224 182410 640446 182440
rect 185775 182380 190014 182382
rect 185775 182377 185841 182380
rect 189954 182366 190014 182380
rect 640194 182380 640416 182410
rect 189954 182306 190560 182366
rect 184431 181552 184497 181555
rect 184431 181550 190560 181552
rect 184431 181494 184436 181550
rect 184492 181494 190560 181550
rect 184431 181492 190560 181494
rect 184431 181489 184497 181492
rect 149295 181404 149361 181407
rect 143904 181402 149361 181404
rect 143904 181346 149300 181402
rect 149356 181346 149361 181402
rect 143904 181344 149361 181346
rect 149295 181341 149361 181344
rect 184335 180812 184401 180815
rect 184335 180810 190560 180812
rect 184335 180754 184340 180810
rect 184396 180754 190560 180810
rect 184335 180752 190560 180754
rect 184335 180749 184401 180752
rect 640194 180560 640254 182380
rect 143874 179628 143934 180116
rect 184431 180072 184497 180075
rect 184431 180070 190560 180072
rect 184431 180014 184436 180070
rect 184492 180014 190560 180070
rect 184431 180012 190560 180014
rect 184431 180009 184497 180012
rect 149487 179628 149553 179631
rect 143874 179626 149553 179628
rect 143874 179570 149492 179626
rect 149548 179570 149553 179626
rect 143874 179568 149553 179570
rect 149487 179565 149553 179568
rect 184623 179332 184689 179335
rect 645135 179332 645201 179335
rect 184623 179330 190560 179332
rect 184623 179274 184628 179330
rect 184684 179274 190560 179330
rect 184623 179272 190560 179274
rect 640194 179330 645201 179332
rect 640194 179274 645140 179330
rect 645196 179274 645201 179330
rect 640194 179272 645201 179274
rect 184623 179269 184689 179272
rect 149391 178888 149457 178891
rect 143904 178886 149457 178888
rect 143904 178830 149396 178886
rect 149452 178830 149457 178886
rect 143904 178828 149457 178830
rect 149391 178825 149457 178828
rect 184527 178592 184593 178595
rect 184527 178590 190560 178592
rect 184527 178534 184532 178590
rect 184588 178534 190560 178590
rect 184527 178532 190560 178534
rect 184527 178529 184593 178532
rect 149391 177704 149457 177707
rect 143904 177702 149457 177704
rect 143904 177646 149396 177702
rect 149452 177646 149457 177702
rect 143904 177644 149457 177646
rect 149391 177641 149457 177644
rect 184431 177704 184497 177707
rect 184431 177702 190560 177704
rect 184431 177646 184436 177702
rect 184492 177646 190560 177702
rect 184431 177644 190560 177646
rect 184431 177641 184497 177644
rect 184335 177112 184401 177115
rect 184335 177110 190014 177112
rect 184335 177054 184340 177110
rect 184396 177054 190014 177110
rect 184335 177052 190014 177054
rect 184335 177049 184401 177052
rect 189954 177038 190014 177052
rect 189954 176978 190560 177038
rect 640194 176786 640254 179272
rect 645135 179269 645201 179272
rect 676143 177408 676209 177411
rect 676290 177408 676350 177674
rect 676143 177406 676350 177408
rect 676143 177350 676148 177406
rect 676204 177350 676350 177406
rect 676143 177348 676350 177350
rect 676143 177345 676209 177348
rect 676290 176819 676350 177082
rect 676290 176814 676401 176819
rect 676290 176758 676340 176814
rect 676396 176758 676401 176814
rect 676290 176756 676401 176758
rect 676335 176753 676401 176756
rect 147759 176520 147825 176523
rect 143904 176518 147825 176520
rect 143904 176462 147764 176518
rect 147820 176462 147825 176518
rect 143904 176460 147825 176462
rect 147759 176457 147825 176460
rect 676290 176375 676350 176638
rect 676239 176370 676350 176375
rect 676239 176314 676244 176370
rect 676300 176314 676350 176370
rect 676239 176312 676350 176314
rect 676239 176309 676305 176312
rect 184527 176224 184593 176227
rect 184527 176222 190560 176224
rect 184527 176166 184532 176222
rect 184588 176166 190560 176222
rect 184527 176164 190560 176166
rect 184527 176161 184593 176164
rect 674170 176162 674176 176226
rect 674240 176224 674246 176226
rect 674240 176164 676320 176224
rect 674240 176162 674246 176164
rect 184335 175632 184401 175635
rect 184335 175630 190014 175632
rect 184335 175574 184340 175630
rect 184396 175574 190014 175630
rect 184335 175572 190014 175574
rect 184335 175569 184401 175572
rect 189954 175558 190014 175572
rect 674554 175570 674560 175634
rect 674624 175632 674630 175634
rect 674624 175572 676320 175632
rect 674624 175570 674630 175572
rect 189954 175498 190560 175558
rect 673978 175422 673984 175486
rect 674048 175484 674054 175486
rect 674048 175424 676350 175484
rect 674048 175422 674054 175424
rect 149391 175188 149457 175191
rect 143904 175186 149457 175188
rect 143904 175130 149396 175186
rect 149452 175130 149457 175186
rect 143904 175128 149457 175130
rect 149391 175125 149457 175128
rect 676290 175084 676350 175424
rect 645135 174892 645201 174895
rect 640416 174890 645201 174892
rect 640416 174862 645140 174890
rect 640386 174834 645140 174862
rect 645196 174834 645201 174890
rect 640386 174832 645201 174834
rect 186255 174744 186321 174747
rect 186255 174742 190560 174744
rect 186255 174686 186260 174742
rect 186316 174686 190560 174742
rect 186255 174684 190560 174686
rect 186255 174681 186321 174684
rect 148911 174004 148977 174007
rect 143904 174002 148977 174004
rect 143904 173946 148916 174002
rect 148972 173946 148977 174002
rect 143904 173944 148977 173946
rect 148911 173941 148977 173944
rect 184431 174004 184497 174007
rect 184431 174002 190014 174004
rect 184431 173946 184436 174002
rect 184492 173946 190014 174002
rect 184431 173944 190014 173946
rect 184431 173941 184497 173944
rect 189954 173930 190014 173944
rect 189954 173870 190560 173930
rect 185583 173264 185649 173267
rect 185583 173262 190560 173264
rect 185583 173206 185588 173262
rect 185644 173206 190560 173262
rect 185583 173204 190560 173206
rect 185583 173201 185649 173204
rect 640386 172938 640446 174832
rect 645135 174829 645201 174832
rect 672399 174744 672465 174747
rect 673978 174744 673984 174746
rect 672399 174742 673984 174744
rect 672399 174686 672404 174742
rect 672460 174686 673984 174742
rect 672399 174684 673984 174686
rect 672399 174681 672465 174684
rect 673978 174682 673984 174684
rect 674048 174744 674054 174746
rect 674048 174684 676320 174744
rect 674048 174682 674054 174684
rect 674362 174090 674368 174154
rect 674432 174152 674438 174154
rect 674432 174092 676320 174152
rect 674432 174090 674438 174092
rect 672591 173560 672657 173563
rect 674170 173560 674176 173562
rect 672591 173558 674176 173560
rect 672591 173502 672596 173558
rect 672652 173502 674176 173558
rect 672591 173500 674176 173502
rect 672591 173497 672657 173500
rect 674170 173498 674176 173500
rect 674240 173560 674246 173562
rect 674240 173500 676320 173560
rect 674240 173498 674246 173500
rect 676482 172970 676542 173234
rect 676474 172906 676480 172970
rect 676544 172906 676550 172970
rect 149295 172820 149361 172823
rect 143904 172818 149361 172820
rect 143904 172762 149300 172818
rect 149356 172762 149361 172818
rect 143904 172760 149361 172762
rect 149295 172757 149361 172760
rect 674746 172610 674752 172674
rect 674816 172672 674822 172674
rect 674816 172612 676320 172672
rect 674816 172610 674822 172612
rect 184335 172524 184401 172527
rect 184335 172522 190014 172524
rect 184335 172466 184340 172522
rect 184396 172466 190014 172522
rect 184335 172464 190014 172466
rect 184335 172461 184401 172464
rect 189954 172450 190014 172464
rect 189954 172390 190560 172450
rect 675567 172080 675633 172083
rect 675567 172078 676320 172080
rect 675567 172022 675572 172078
rect 675628 172022 676320 172078
rect 675567 172020 676320 172022
rect 675567 172017 675633 172020
rect 184431 171784 184497 171787
rect 184431 171782 190560 171784
rect 184431 171726 184436 171782
rect 184492 171726 190560 171782
rect 184431 171724 190560 171726
rect 184431 171721 184497 171724
rect 143874 171044 143934 171532
rect 675514 171278 675520 171342
rect 675584 171340 675590 171342
rect 676290 171340 676350 171680
rect 675584 171280 676350 171340
rect 675584 171278 675590 171280
rect 674938 171130 674944 171194
rect 675008 171192 675014 171194
rect 675008 171132 676320 171192
rect 675008 171130 675014 171132
rect 149583 171044 149649 171047
rect 645135 171044 645201 171047
rect 143874 171042 149649 171044
rect 143874 170986 149588 171042
rect 149644 170986 149649 171042
rect 640416 171042 645201 171044
rect 640416 171014 645140 171042
rect 143874 170984 149649 170986
rect 149583 170981 149649 170984
rect 640386 170986 645140 171014
rect 645196 170986 645201 171042
rect 640386 170984 645201 170986
rect 184623 170896 184689 170899
rect 184623 170894 190560 170896
rect 184623 170838 184628 170894
rect 184684 170838 190560 170894
rect 184623 170836 190560 170838
rect 184623 170833 184689 170836
rect 149199 170304 149265 170307
rect 143904 170302 149265 170304
rect 143904 170246 149204 170302
rect 149260 170246 149265 170302
rect 143904 170244 149265 170246
rect 149199 170241 149265 170244
rect 184527 170304 184593 170307
rect 184527 170302 190014 170304
rect 184527 170246 184532 170302
rect 184588 170246 190014 170302
rect 184527 170244 190014 170246
rect 184527 170241 184593 170244
rect 189954 170230 190014 170244
rect 189954 170170 190560 170230
rect 184431 169416 184497 169419
rect 184431 169414 190560 169416
rect 184431 169358 184436 169414
rect 184492 169358 190560 169414
rect 184431 169356 190560 169358
rect 184431 169353 184497 169356
rect 149487 169120 149553 169123
rect 143904 169118 149553 169120
rect 143904 169062 149492 169118
rect 149548 169062 149553 169118
rect 640386 169090 640446 170984
rect 645135 170981 645201 170984
rect 676290 170454 676350 170570
rect 676282 170390 676288 170454
rect 676352 170390 676358 170454
rect 676047 170230 676113 170233
rect 676047 170228 676320 170230
rect 676047 170172 676052 170228
rect 676108 170172 676320 170228
rect 676047 170170 676320 170172
rect 676047 170167 676113 170170
rect 676047 169712 676113 169715
rect 676047 169710 676320 169712
rect 676047 169654 676052 169710
rect 676108 169654 676320 169710
rect 676047 169652 676320 169654
rect 676047 169649 676113 169652
rect 143904 169060 149553 169062
rect 149487 169057 149553 169060
rect 676290 168975 676350 169090
rect 676239 168970 676350 168975
rect 676239 168914 676244 168970
rect 676300 168914 676350 168970
rect 676239 168912 676350 168914
rect 676239 168909 676305 168912
rect 184335 168676 184401 168679
rect 184335 168674 190014 168676
rect 184335 168618 184340 168674
rect 184396 168618 190014 168674
rect 184335 168616 190014 168618
rect 184335 168613 184401 168616
rect 189954 168602 190014 168616
rect 675322 168614 675328 168678
rect 675392 168676 675398 168678
rect 675392 168616 676320 168676
rect 675392 168614 675398 168616
rect 189954 168542 190560 168602
rect 675130 168170 675136 168234
rect 675200 168232 675206 168234
rect 675200 168172 676320 168232
rect 675200 168170 675206 168172
rect 148911 168084 148977 168087
rect 143904 168082 148977 168084
rect 143904 168026 148916 168082
rect 148972 168026 148977 168082
rect 143904 168024 148977 168026
rect 148911 168021 148977 168024
rect 184623 167936 184689 167939
rect 184623 167934 190560 167936
rect 184623 167878 184628 167934
rect 184684 167878 190560 167934
rect 184623 167876 190560 167878
rect 184623 167873 184689 167876
rect 645135 167788 645201 167791
rect 640386 167786 645201 167788
rect 640386 167730 645140 167786
rect 645196 167730 645201 167786
rect 640386 167728 645201 167730
rect 184527 167196 184593 167199
rect 184527 167194 190014 167196
rect 184527 167138 184532 167194
rect 184588 167138 190014 167194
rect 184527 167136 190014 167138
rect 184527 167133 184593 167136
rect 189954 167122 190014 167136
rect 189954 167062 190560 167122
rect 143874 166308 143934 166796
rect 184335 166456 184401 166459
rect 184335 166454 190560 166456
rect 184335 166398 184340 166454
rect 184396 166398 190560 166454
rect 184335 166396 190560 166398
rect 184335 166393 184401 166396
rect 148527 166308 148593 166311
rect 143874 166306 148593 166308
rect 143874 166250 148532 166306
rect 148588 166250 148593 166306
rect 143874 166248 148593 166250
rect 148527 166245 148593 166248
rect 640386 166012 640446 167728
rect 645135 167725 645201 167728
rect 675898 167578 675904 167642
rect 675968 167640 675974 167642
rect 675968 167580 676320 167640
rect 675968 167578 675974 167580
rect 675706 167134 675712 167198
rect 675776 167196 675782 167198
rect 675776 167136 676320 167196
rect 675776 167134 675782 167136
rect 676090 166246 676096 166310
rect 676160 166308 676166 166310
rect 676290 166308 676350 166648
rect 676160 166248 676350 166308
rect 676160 166246 676166 166248
rect 676047 166160 676113 166163
rect 676047 166158 676320 166160
rect 676047 166102 676052 166158
rect 676108 166102 676320 166158
rect 676047 166100 676320 166102
rect 676047 166097 676113 166100
rect 640194 165952 640446 166012
rect 184431 165716 184497 165719
rect 184431 165714 190014 165716
rect 184431 165658 184436 165714
rect 184492 165658 190014 165714
rect 184431 165656 190014 165658
rect 184431 165653 184497 165656
rect 189954 165642 190014 165656
rect 189954 165582 190560 165642
rect 148335 165568 148401 165571
rect 143904 165566 148401 165568
rect 143904 165510 148340 165566
rect 148396 165510 148401 165566
rect 143904 165508 148401 165510
rect 148335 165505 148401 165508
rect 640194 165242 640254 165952
rect 676143 165420 676209 165423
rect 676290 165420 676350 165686
rect 676143 165418 676350 165420
rect 676143 165362 676148 165418
rect 676204 165362 676350 165418
rect 676143 165360 676350 165362
rect 676143 165357 676209 165360
rect 676290 164831 676350 165168
rect 184527 164828 184593 164831
rect 184527 164826 190560 164828
rect 184527 164770 184532 164826
rect 184588 164770 190560 164826
rect 184527 164768 190560 164770
rect 676239 164826 676350 164831
rect 676239 164770 676244 164826
rect 676300 164770 676350 164826
rect 676239 164768 676350 164770
rect 184527 164765 184593 164768
rect 676239 164765 676305 164768
rect 148719 164384 148785 164387
rect 143904 164382 148785 164384
rect 143904 164326 148724 164382
rect 148780 164326 148785 164382
rect 143904 164324 148785 164326
rect 148719 164321 148785 164324
rect 184335 164088 184401 164091
rect 184335 164086 190560 164088
rect 184335 164030 184340 164086
rect 184396 164030 190560 164086
rect 184335 164028 190560 164030
rect 184335 164025 184401 164028
rect 184527 163348 184593 163351
rect 645135 163348 645201 163351
rect 184527 163346 190560 163348
rect 184527 163290 184532 163346
rect 184588 163290 190560 163346
rect 640416 163346 645201 163348
rect 640416 163318 645140 163346
rect 184527 163288 190560 163290
rect 640386 163290 645140 163318
rect 645196 163290 645201 163346
rect 640386 163288 645201 163290
rect 184527 163285 184593 163288
rect 148431 163200 148497 163203
rect 143904 163198 148497 163200
rect 143904 163142 148436 163198
rect 148492 163142 148497 163198
rect 143904 163140 148497 163142
rect 148431 163137 148497 163140
rect 184335 162608 184401 162611
rect 184335 162606 190560 162608
rect 184335 162550 184340 162606
rect 184396 162550 190560 162606
rect 184335 162548 190560 162550
rect 184335 162545 184401 162548
rect 148239 161868 148305 161871
rect 143904 161866 148305 161868
rect 143904 161810 148244 161866
rect 148300 161810 148305 161866
rect 143904 161808 148305 161810
rect 148239 161805 148305 161808
rect 184431 161868 184497 161871
rect 184431 161866 190560 161868
rect 184431 161810 184436 161866
rect 184492 161810 190560 161866
rect 184431 161808 190560 161810
rect 184431 161805 184497 161808
rect 640386 161394 640446 163288
rect 645135 163285 645201 163288
rect 184431 160980 184497 160983
rect 184431 160978 190560 160980
rect 184431 160922 184436 160978
rect 184492 160922 190560 160978
rect 184431 160920 190560 160922
rect 184431 160917 184497 160920
rect 148623 160684 148689 160687
rect 143904 160682 148689 160684
rect 143904 160626 148628 160682
rect 148684 160626 148689 160682
rect 143904 160624 148689 160626
rect 148623 160621 148689 160624
rect 184527 160388 184593 160391
rect 184527 160386 190014 160388
rect 184527 160330 184532 160386
rect 184588 160330 190014 160386
rect 184527 160328 190014 160330
rect 184527 160325 184593 160328
rect 189954 160314 190014 160328
rect 189954 160254 190560 160314
rect 147087 159500 147153 159503
rect 143904 159498 147153 159500
rect 143904 159442 147092 159498
rect 147148 159442 147153 159498
rect 143904 159440 147153 159442
rect 147087 159437 147153 159440
rect 184335 159500 184401 159503
rect 645135 159500 645201 159503
rect 184335 159498 190560 159500
rect 184335 159442 184340 159498
rect 184396 159442 190560 159498
rect 640416 159498 645201 159500
rect 640416 159470 645140 159498
rect 184335 159440 190560 159442
rect 640386 159442 645140 159470
rect 645196 159442 645201 159498
rect 640386 159440 645201 159442
rect 184335 159437 184401 159440
rect 184623 158908 184689 158911
rect 184623 158906 190014 158908
rect 184623 158850 184628 158906
rect 184684 158850 190014 158906
rect 184623 158848 190014 158850
rect 184623 158845 184689 158848
rect 189954 158834 190014 158848
rect 189954 158774 190560 158834
rect 143874 157724 143934 158212
rect 184335 158020 184401 158023
rect 184335 158018 190560 158020
rect 184335 157962 184340 158018
rect 184396 157962 190560 158018
rect 184335 157960 190560 157962
rect 184335 157957 184401 157960
rect 148815 157724 148881 157727
rect 143874 157722 148881 157724
rect 143874 157666 148820 157722
rect 148876 157666 148881 157722
rect 143874 157664 148881 157666
rect 148815 157661 148881 157664
rect 640386 157546 640446 159440
rect 645135 159437 645201 159440
rect 675759 159352 675825 159355
rect 676474 159352 676480 159354
rect 675759 159350 676480 159352
rect 675759 159294 675764 159350
rect 675820 159294 676480 159350
rect 675759 159292 676480 159294
rect 675759 159289 675825 159292
rect 676474 159290 676480 159292
rect 676544 159290 676550 159354
rect 675471 157726 675537 157727
rect 675471 157722 675520 157726
rect 675584 157724 675590 157726
rect 675471 157666 675476 157722
rect 675471 157662 675520 157666
rect 675584 157664 675628 157724
rect 675584 157662 675590 157664
rect 675471 157661 675537 157662
rect 184431 157428 184497 157431
rect 184431 157426 190014 157428
rect 184431 157370 184436 157426
rect 184492 157370 190014 157426
rect 184431 157368 190014 157370
rect 184431 157365 184497 157368
rect 189954 157354 190014 157368
rect 189954 157294 190560 157354
rect 146895 156984 146961 156987
rect 143904 156982 146961 156984
rect 143904 156926 146900 156982
rect 146956 156926 146961 156982
rect 143904 156924 146961 156926
rect 146895 156921 146961 156924
rect 184527 156540 184593 156543
rect 184527 156538 190560 156540
rect 184527 156482 184532 156538
rect 184588 156482 190560 156538
rect 184527 156480 190560 156482
rect 184527 156477 184593 156480
rect 149679 155800 149745 155803
rect 143904 155798 149745 155800
rect 143904 155742 149684 155798
rect 149740 155742 149745 155798
rect 143904 155740 149745 155742
rect 149679 155737 149745 155740
rect 184623 155652 184689 155655
rect 184623 155650 190560 155652
rect 184623 155594 184628 155650
rect 184684 155594 190560 155650
rect 184623 155592 190560 155594
rect 184623 155589 184689 155592
rect 640194 155504 640254 155622
rect 645135 155504 645201 155507
rect 640194 155502 645201 155504
rect 640194 155446 645140 155502
rect 645196 155446 645201 155502
rect 640194 155444 645201 155446
rect 184335 155060 184401 155063
rect 184335 155058 190560 155060
rect 184335 155002 184340 155058
rect 184396 155002 190560 155058
rect 184335 155000 190560 155002
rect 184335 154997 184401 155000
rect 149295 154616 149361 154619
rect 143904 154614 149361 154616
rect 143904 154558 149300 154614
rect 149356 154558 149361 154614
rect 143904 154556 149361 154558
rect 149295 154553 149361 154556
rect 184431 154172 184497 154175
rect 184431 154170 190560 154172
rect 184431 154114 184436 154170
rect 184492 154114 190560 154170
rect 184431 154112 190560 154114
rect 184431 154109 184497 154112
rect 640386 153772 640446 155444
rect 645135 155441 645201 155444
rect 675759 155504 675825 155507
rect 675898 155504 675904 155506
rect 675759 155502 675904 155504
rect 675759 155446 675764 155502
rect 675820 155446 675904 155502
rect 675759 155444 675904 155446
rect 675759 155441 675825 155444
rect 675898 155442 675904 155444
rect 675968 155442 675974 155506
rect 674938 155294 674944 155358
rect 675008 155356 675014 155358
rect 675087 155356 675153 155359
rect 675008 155354 675153 155356
rect 675008 155298 675092 155354
rect 675148 155298 675153 155354
rect 675008 155296 675153 155298
rect 675008 155294 675014 155296
rect 675087 155293 675153 155296
rect 184527 153580 184593 153583
rect 184527 153578 190014 153580
rect 184527 153522 184532 153578
rect 184588 153522 190014 153578
rect 184527 153520 190014 153522
rect 184527 153517 184593 153520
rect 189954 153506 190014 153520
rect 189954 153446 190560 153506
rect 143874 153136 143934 153328
rect 149487 153136 149553 153139
rect 143874 153134 149553 153136
rect 143874 153078 149492 153134
rect 149548 153078 149553 153134
rect 143874 153076 149553 153078
rect 149487 153073 149553 153076
rect 184623 152692 184689 152695
rect 184623 152690 190560 152692
rect 184623 152634 184628 152690
rect 184684 152634 190560 152690
rect 184623 152632 190560 152634
rect 184623 152629 184689 152632
rect 645135 152544 645201 152547
rect 675183 152546 675249 152547
rect 675130 152544 675136 152546
rect 640194 152542 645201 152544
rect 640194 152486 645140 152542
rect 645196 152486 645201 152542
rect 640194 152484 645201 152486
rect 675092 152484 675136 152544
rect 675200 152542 675249 152546
rect 675244 152486 675249 152542
rect 149679 152100 149745 152103
rect 143904 152098 149745 152100
rect 143904 152042 149684 152098
rect 149740 152042 149745 152098
rect 143904 152040 149745 152042
rect 149679 152037 149745 152040
rect 184335 151952 184401 151955
rect 184335 151950 190014 151952
rect 184335 151894 184340 151950
rect 184396 151894 190014 151950
rect 184335 151892 190014 151894
rect 184335 151889 184401 151892
rect 189954 151878 190014 151892
rect 189954 151818 190560 151878
rect 184431 151212 184497 151215
rect 184431 151210 190560 151212
rect 184431 151154 184436 151210
rect 184492 151154 190560 151210
rect 184431 151152 190560 151154
rect 184431 151149 184497 151152
rect 149487 150916 149553 150919
rect 143904 150914 149553 150916
rect 143904 150858 149492 150914
rect 149548 150858 149553 150914
rect 143904 150856 149553 150858
rect 149487 150853 149553 150856
rect 184527 150472 184593 150475
rect 184527 150470 190014 150472
rect 184527 150414 184532 150470
rect 184588 150414 190014 150470
rect 184527 150412 190014 150414
rect 184527 150409 184593 150412
rect 189954 150398 190014 150412
rect 189954 150338 190560 150398
rect 640194 149998 640254 152484
rect 645135 152481 645201 152484
rect 675130 152482 675136 152484
rect 675200 152482 675249 152486
rect 675183 152481 675249 152482
rect 675663 152546 675729 152547
rect 675663 152542 675712 152546
rect 675776 152544 675782 152546
rect 675663 152486 675668 152542
rect 675663 152482 675712 152486
rect 675776 152484 675820 152544
rect 675776 152482 675782 152484
rect 675663 152481 675729 152482
rect 675759 151360 675825 151363
rect 676090 151360 676096 151362
rect 675759 151358 676096 151360
rect 675759 151302 675764 151358
rect 675820 151302 676096 151358
rect 675759 151300 676096 151302
rect 675759 151297 675825 151300
rect 676090 151298 676096 151300
rect 676160 151298 676166 151362
rect 675322 150262 675328 150326
rect 675392 150324 675398 150326
rect 675471 150324 675537 150327
rect 675392 150322 675537 150324
rect 675392 150266 675476 150322
rect 675532 150266 675537 150322
rect 675392 150264 675537 150266
rect 675392 150262 675398 150264
rect 675471 150261 675537 150264
rect 149295 149880 149361 149883
rect 143874 149878 149361 149880
rect 143874 149822 149300 149878
rect 149356 149822 149361 149878
rect 143874 149820 149361 149822
rect 143874 149776 143934 149820
rect 149295 149817 149361 149820
rect 184335 149732 184401 149735
rect 184335 149730 190560 149732
rect 184335 149674 184340 149730
rect 184396 149674 190560 149730
rect 184335 149672 190560 149674
rect 184335 149669 184401 149672
rect 674746 149670 674752 149734
rect 674816 149732 674822 149734
rect 675087 149732 675153 149735
rect 674816 149730 675153 149732
rect 674816 149674 675092 149730
rect 675148 149674 675153 149730
rect 674816 149672 675153 149674
rect 674816 149670 674822 149672
rect 675087 149669 675153 149672
rect 184431 148992 184497 148995
rect 184431 148990 190014 148992
rect 184431 148934 184436 148990
rect 184492 148934 190014 148990
rect 184431 148932 190014 148934
rect 184431 148929 184497 148932
rect 189954 148918 190014 148932
rect 189954 148858 190560 148918
rect 149295 148548 149361 148551
rect 143904 148546 149361 148548
rect 143904 148490 149300 148546
rect 149356 148490 149361 148546
rect 143904 148488 149361 148490
rect 149295 148485 149361 148488
rect 186735 148104 186801 148107
rect 645135 148104 645201 148107
rect 186735 148102 190560 148104
rect 186735 148046 186740 148102
rect 186796 148046 190560 148102
rect 640416 148102 645201 148104
rect 640416 148074 645140 148102
rect 186735 148044 190560 148046
rect 640386 148046 645140 148074
rect 645196 148046 645201 148102
rect 640386 148044 645201 148046
rect 186735 148041 186801 148044
rect 149487 147364 149553 147367
rect 143904 147362 149553 147364
rect 143904 147306 149492 147362
rect 149548 147306 149553 147362
rect 143904 147304 149553 147306
rect 149487 147301 149553 147304
rect 184527 147364 184593 147367
rect 184527 147362 190560 147364
rect 184527 147306 184532 147362
rect 184588 147306 190560 147362
rect 184527 147304 190560 147306
rect 184527 147301 184593 147304
rect 184623 146624 184689 146627
rect 184623 146622 190560 146624
rect 184623 146566 184628 146622
rect 184684 146566 190560 146622
rect 184623 146564 190560 146566
rect 184623 146561 184689 146564
rect 147663 146180 147729 146183
rect 143904 146178 147729 146180
rect 143904 146122 147668 146178
rect 147724 146122 147729 146178
rect 640386 146150 640446 148044
rect 645135 148041 645201 148044
rect 675759 146624 675825 146627
rect 676282 146624 676288 146626
rect 675759 146622 676288 146624
rect 675759 146566 675764 146622
rect 675820 146566 676288 146622
rect 675759 146564 676288 146566
rect 675759 146561 675825 146564
rect 676282 146562 676288 146564
rect 676352 146562 676358 146626
rect 143904 146120 147729 146122
rect 147663 146117 147729 146120
rect 184335 145884 184401 145887
rect 184335 145882 190560 145884
rect 184335 145826 184340 145882
rect 184396 145826 190560 145882
rect 184335 145824 190560 145826
rect 184335 145821 184401 145824
rect 184431 145144 184497 145147
rect 184431 145142 190014 145144
rect 184431 145086 184436 145142
rect 184492 145086 190014 145142
rect 184431 145084 190014 145086
rect 184431 145081 184497 145084
rect 189954 145070 190014 145084
rect 189954 145010 190560 145070
rect 143874 144552 143934 144892
rect 147663 144552 147729 144555
rect 143874 144550 147729 144552
rect 143874 144494 147668 144550
rect 147724 144494 147729 144550
rect 143874 144492 147729 144494
rect 147663 144489 147729 144492
rect 184527 144404 184593 144407
rect 184527 144402 190560 144404
rect 184527 144346 184532 144402
rect 184588 144346 190560 144402
rect 184527 144344 190560 144346
rect 184527 144341 184593 144344
rect 646671 144256 646737 144259
rect 640416 144254 646737 144256
rect 640416 144226 646676 144254
rect 640386 144198 646676 144226
rect 646732 144198 646737 144254
rect 640386 144196 646737 144198
rect 147279 143664 147345 143667
rect 143904 143662 147345 143664
rect 143904 143606 147284 143662
rect 147340 143606 147345 143662
rect 143904 143604 147345 143606
rect 147279 143601 147345 143604
rect 184335 143664 184401 143667
rect 184335 143662 190014 143664
rect 184335 143606 184340 143662
rect 184396 143606 190014 143662
rect 184335 143604 190014 143606
rect 184335 143601 184401 143604
rect 189954 143590 190014 143604
rect 189954 143530 190560 143590
rect 184431 142776 184497 142779
rect 184431 142774 190560 142776
rect 184431 142718 184436 142774
rect 184492 142718 190560 142774
rect 184431 142716 190560 142718
rect 184431 142713 184497 142716
rect 147471 142480 147537 142483
rect 143904 142478 147537 142480
rect 143904 142422 147476 142478
rect 147532 142422 147537 142478
rect 143904 142420 147537 142422
rect 147471 142417 147537 142420
rect 640386 142302 640446 144196
rect 646671 144193 646737 144196
rect 184623 142184 184689 142187
rect 184623 142182 190014 142184
rect 184623 142126 184628 142182
rect 184684 142126 190014 142182
rect 184623 142124 190014 142126
rect 184623 142121 184689 142124
rect 189954 142110 190014 142124
rect 189954 142050 190560 142110
rect 149679 141296 149745 141299
rect 143904 141294 149745 141296
rect 143904 141238 149684 141294
rect 149740 141238 149745 141294
rect 143904 141236 149745 141238
rect 149679 141233 149745 141236
rect 184527 141296 184593 141299
rect 184527 141294 190560 141296
rect 184527 141238 184532 141294
rect 184588 141238 190560 141294
rect 184527 141236 190560 141238
rect 184527 141233 184593 141236
rect 646767 141000 646833 141003
rect 640386 140998 646833 141000
rect 640386 140942 646772 140998
rect 646828 140942 646833 140998
rect 640386 140940 646833 140942
rect 184335 140556 184401 140559
rect 184335 140554 190560 140556
rect 184335 140498 184340 140554
rect 184396 140498 190560 140554
rect 184335 140496 190560 140498
rect 184335 140493 184401 140496
rect 640386 140408 640446 140940
rect 646767 140937 646833 140940
rect 640224 140378 640446 140408
rect 640194 140348 640416 140378
rect 147471 139964 147537 139967
rect 143904 139962 147537 139964
rect 143904 139906 147476 139962
rect 147532 139906 147537 139962
rect 143904 139904 147537 139906
rect 147471 139901 147537 139904
rect 184431 139816 184497 139819
rect 184431 139814 190560 139816
rect 184431 139758 184436 139814
rect 184492 139758 190560 139814
rect 184431 139756 190560 139758
rect 184431 139753 184497 139756
rect 184527 138928 184593 138931
rect 184527 138926 190560 138928
rect 184527 138870 184532 138926
rect 184588 138870 190560 138926
rect 184527 138868 190560 138870
rect 184527 138865 184593 138868
rect 147663 138780 147729 138783
rect 143904 138778 147729 138780
rect 143904 138722 147668 138778
rect 147724 138722 147729 138778
rect 143904 138720 147729 138722
rect 147663 138717 147729 138720
rect 640194 138528 640254 140348
rect 186063 138336 186129 138339
rect 186063 138334 190560 138336
rect 186063 138278 186068 138334
rect 186124 138278 190560 138334
rect 186063 138276 190560 138278
rect 186063 138273 186129 138276
rect 149583 137596 149649 137599
rect 143904 137594 149649 137596
rect 143904 137538 149588 137594
rect 149644 137538 149649 137594
rect 143904 137536 149649 137538
rect 149583 137533 149649 137536
rect 185967 137448 186033 137451
rect 185967 137446 190560 137448
rect 185967 137390 185972 137446
rect 186028 137390 190560 137446
rect 185967 137388 190560 137390
rect 185967 137385 186033 137388
rect 186159 136856 186225 136859
rect 186159 136854 190014 136856
rect 186159 136798 186164 136854
rect 186220 136798 190014 136854
rect 186159 136796 190014 136798
rect 186159 136793 186225 136796
rect 189954 136782 190014 136796
rect 189954 136722 190560 136782
rect 143874 135968 143934 136308
rect 149679 135968 149745 135971
rect 143874 135966 149745 135968
rect 143874 135910 149684 135966
rect 149740 135910 149745 135966
rect 143874 135908 149745 135910
rect 149679 135905 149745 135908
rect 186447 135968 186513 135971
rect 186447 135966 190560 135968
rect 186447 135910 186452 135966
rect 186508 135910 190560 135966
rect 186447 135908 190560 135910
rect 186447 135905 186513 135908
rect 185775 135228 185841 135231
rect 185775 135226 190014 135228
rect 185775 135170 185780 135226
rect 185836 135170 190014 135226
rect 185775 135168 190014 135170
rect 185775 135165 185841 135168
rect 189954 135154 190014 135168
rect 189954 135094 190560 135154
rect 149679 135080 149745 135083
rect 143904 135078 149745 135080
rect 143904 135022 149684 135078
rect 149740 135022 149745 135078
rect 143904 135020 149745 135022
rect 149679 135017 149745 135020
rect 647055 134784 647121 134787
rect 640416 134782 647121 134784
rect 640416 134726 647060 134782
rect 647116 134726 647121 134782
rect 640416 134724 647121 134726
rect 647055 134721 647121 134724
rect 184335 134488 184401 134491
rect 184335 134486 190560 134488
rect 184335 134430 184340 134486
rect 184396 134430 190560 134486
rect 184335 134428 190560 134430
rect 184335 134425 184401 134428
rect 148911 133896 148977 133899
rect 143904 133894 148977 133896
rect 143904 133838 148916 133894
rect 148972 133838 148977 133894
rect 143904 133836 148977 133838
rect 148911 133833 148977 133836
rect 186255 133748 186321 133751
rect 186255 133746 190014 133748
rect 186255 133690 186260 133746
rect 186316 133690 190014 133746
rect 186255 133688 190014 133690
rect 186255 133685 186321 133688
rect 189954 133674 190014 133688
rect 189954 133614 190560 133674
rect 184431 133008 184497 133011
rect 184431 133006 190560 133008
rect 184431 132950 184436 133006
rect 184492 132950 190560 133006
rect 184431 132948 190560 132950
rect 184431 132945 184497 132948
rect 148815 132712 148881 132715
rect 143904 132710 148881 132712
rect 143904 132654 148820 132710
rect 148876 132654 148881 132710
rect 143904 132652 148881 132654
rect 148815 132649 148881 132652
rect 184335 132268 184401 132271
rect 184335 132266 190014 132268
rect 184335 132210 184340 132266
rect 184396 132210 190014 132266
rect 184335 132208 190014 132210
rect 184335 132205 184401 132208
rect 189954 132194 190014 132208
rect 189954 132134 190560 132194
rect 676143 131824 676209 131827
rect 676290 131824 676350 132090
rect 676143 131822 676350 131824
rect 676143 131766 676148 131822
rect 676204 131766 676350 131822
rect 676143 131764 676350 131766
rect 676143 131761 676209 131764
rect 184431 131528 184497 131531
rect 184431 131526 190560 131528
rect 184431 131470 184436 131526
rect 184492 131470 190560 131526
rect 184431 131468 190560 131470
rect 184431 131465 184497 131468
rect 143874 130936 143934 131424
rect 676290 131235 676350 131498
rect 676290 131230 676401 131235
rect 676290 131174 676340 131230
rect 676396 131174 676401 131230
rect 676290 131172 676401 131174
rect 676335 131169 676401 131172
rect 149679 130936 149745 130939
rect 647823 130936 647889 130939
rect 143874 130934 149745 130936
rect 143874 130878 149684 130934
rect 149740 130878 149745 130934
rect 143874 130876 149745 130878
rect 640416 130934 647889 130936
rect 640416 130878 647828 130934
rect 647884 130878 647889 130934
rect 640416 130876 647889 130878
rect 149679 130873 149745 130876
rect 647823 130873 647889 130876
rect 676290 130791 676350 130980
rect 676239 130786 676350 130791
rect 676239 130730 676244 130786
rect 676300 130730 676350 130786
rect 676239 130728 676350 130730
rect 676239 130725 676305 130728
rect 184527 130640 184593 130643
rect 184527 130638 190560 130640
rect 184527 130582 184532 130638
rect 184588 130582 190560 130638
rect 184527 130580 190560 130582
rect 184527 130577 184593 130580
rect 674362 130578 674368 130642
rect 674432 130640 674438 130642
rect 674432 130580 676320 130640
rect 674432 130578 674438 130580
rect 147471 130344 147537 130347
rect 143904 130342 147537 130344
rect 143904 130286 147476 130342
rect 147532 130286 147537 130342
rect 143904 130284 147537 130286
rect 147471 130281 147537 130284
rect 184623 129900 184689 129903
rect 184623 129898 190560 129900
rect 184623 129842 184628 129898
rect 184684 129842 190560 129898
rect 184623 129840 190560 129842
rect 184623 129837 184689 129840
rect 676290 129755 676350 130018
rect 676239 129750 676350 129755
rect 676239 129694 676244 129750
rect 676300 129694 676350 129750
rect 676239 129692 676350 129694
rect 676239 129689 676305 129692
rect 673978 129394 673984 129458
rect 674048 129456 674054 129458
rect 674048 129396 676320 129456
rect 674048 129394 674054 129396
rect 149103 129160 149169 129163
rect 143904 129158 149169 129160
rect 143904 129102 149108 129158
rect 149164 129102 149169 129158
rect 143904 129100 149169 129102
rect 149103 129097 149169 129100
rect 186735 129160 186801 129163
rect 186735 129158 190560 129160
rect 186735 129102 186740 129158
rect 186796 129102 190560 129158
rect 186735 129100 190560 129102
rect 186735 129097 186801 129100
rect 645711 129012 645777 129015
rect 640416 129010 645777 129012
rect 640416 128954 645716 129010
rect 645772 128954 645777 129010
rect 640416 128952 645777 128954
rect 645711 128949 645777 128952
rect 676143 128864 676209 128867
rect 676290 128864 676350 129130
rect 676143 128862 676350 128864
rect 676143 128806 676148 128862
rect 676204 128806 676350 128862
rect 676143 128804 676350 128806
rect 676143 128801 676209 128804
rect 674170 128506 674176 128570
rect 674240 128568 674246 128570
rect 674240 128508 676320 128568
rect 674240 128506 674246 128508
rect 184335 128420 184401 128423
rect 184335 128418 190014 128420
rect 184335 128362 184340 128418
rect 184396 128362 190014 128418
rect 184335 128360 190014 128362
rect 184335 128357 184401 128360
rect 189954 128346 190014 128360
rect 189954 128286 190560 128346
rect 147663 127976 147729 127979
rect 143904 127974 147729 127976
rect 143904 127918 147668 127974
rect 147724 127918 147729 127974
rect 143904 127916 147729 127918
rect 147663 127913 147729 127916
rect 676290 127831 676350 127946
rect 676239 127826 676350 127831
rect 676239 127770 676244 127826
rect 676300 127770 676350 127826
rect 676239 127768 676350 127770
rect 676239 127765 676305 127768
rect 184431 127680 184497 127683
rect 646959 127680 647025 127683
rect 184431 127678 190560 127680
rect 184431 127622 184436 127678
rect 184492 127622 190560 127678
rect 184431 127620 190560 127622
rect 640386 127678 647025 127680
rect 640386 127622 646964 127678
rect 647020 127622 647025 127678
rect 640386 127620 647025 127622
rect 184431 127617 184497 127620
rect 640386 127058 640446 127620
rect 646959 127617 647025 127620
rect 676047 127606 676113 127609
rect 676047 127604 676320 127606
rect 676047 127548 676052 127604
rect 676108 127548 676320 127604
rect 676047 127546 676320 127548
rect 676047 127543 676113 127546
rect 184527 126940 184593 126943
rect 184527 126938 190014 126940
rect 184527 126882 184532 126938
rect 184588 126882 190014 126938
rect 184527 126880 190014 126882
rect 184527 126877 184593 126880
rect 189954 126866 190014 126880
rect 189954 126806 190560 126866
rect 676866 126795 676926 127058
rect 676866 126790 676977 126795
rect 676866 126734 676916 126790
rect 676972 126734 676977 126790
rect 676866 126732 676977 126734
rect 676911 126729 676977 126732
rect 149295 126644 149361 126647
rect 143904 126642 149361 126644
rect 143904 126586 149300 126642
rect 149356 126586 149361 126642
rect 143904 126584 149361 126586
rect 149295 126581 149361 126584
rect 676290 126351 676350 126466
rect 676239 126346 676350 126351
rect 676239 126290 676244 126346
rect 676300 126290 676350 126346
rect 676239 126288 676350 126290
rect 676239 126285 676305 126288
rect 676047 126126 676113 126129
rect 676047 126124 676320 126126
rect 676047 126068 676052 126124
rect 676108 126068 676320 126124
rect 676047 126066 676320 126068
rect 676047 126063 676113 126066
rect 184431 126052 184497 126055
rect 184431 126050 190560 126052
rect 184431 125994 184436 126050
rect 184492 125994 190560 126050
rect 184431 125992 190560 125994
rect 184431 125989 184497 125992
rect 646863 125756 646929 125759
rect 640386 125754 646929 125756
rect 640386 125698 646868 125754
rect 646924 125698 646929 125754
rect 640386 125696 646929 125698
rect 149583 125460 149649 125463
rect 143904 125458 149649 125460
rect 143904 125402 149588 125458
rect 149644 125402 149649 125458
rect 143904 125400 149649 125402
rect 149583 125397 149649 125400
rect 184335 125460 184401 125463
rect 184335 125458 190014 125460
rect 184335 125402 184340 125458
rect 184396 125402 190014 125458
rect 184335 125400 190014 125402
rect 184335 125397 184401 125400
rect 189954 125386 190014 125400
rect 189954 125326 190560 125386
rect 640386 125208 640446 125696
rect 646863 125693 646929 125696
rect 673978 125546 673984 125610
rect 674048 125608 674054 125610
rect 674048 125548 676320 125608
rect 674048 125546 674054 125548
rect 676866 124871 676926 124986
rect 676815 124866 676926 124871
rect 676815 124810 676820 124866
rect 676876 124810 676926 124866
rect 676815 124808 676926 124810
rect 676815 124805 676881 124808
rect 184527 124572 184593 124575
rect 676047 124572 676113 124575
rect 184527 124570 190560 124572
rect 184527 124514 184532 124570
rect 184588 124514 190560 124570
rect 184527 124512 190560 124514
rect 676047 124570 676320 124572
rect 676047 124514 676052 124570
rect 676108 124514 676320 124570
rect 676047 124512 676320 124514
rect 184527 124509 184593 124512
rect 676047 124509 676113 124512
rect 149391 124276 149457 124279
rect 143904 124274 149457 124276
rect 143904 124218 149396 124274
rect 149452 124218 149457 124274
rect 143904 124216 149457 124218
rect 149391 124213 149457 124216
rect 675951 124128 676017 124131
rect 675951 124126 676320 124128
rect 675951 124070 675956 124126
rect 676012 124070 676320 124126
rect 675951 124068 676320 124070
rect 675951 124065 676017 124068
rect 184335 123832 184401 123835
rect 646575 123832 646641 123835
rect 184335 123830 190560 123832
rect 184335 123774 184340 123830
rect 184396 123774 190560 123830
rect 184335 123772 190560 123774
rect 640194 123830 646641 123832
rect 640194 123774 646580 123830
rect 646636 123774 646641 123830
rect 640194 123772 646641 123774
rect 184335 123769 184401 123772
rect 640194 123358 640254 123772
rect 646575 123769 646641 123772
rect 676047 123536 676113 123539
rect 676047 123534 676320 123536
rect 676047 123478 676052 123534
rect 676108 123478 676320 123534
rect 676047 123476 676320 123478
rect 676047 123473 676113 123476
rect 184431 123092 184497 123095
rect 184431 123090 190560 123092
rect 184431 123034 184436 123090
rect 184492 123034 190560 123090
rect 184431 123032 190560 123034
rect 184431 123029 184497 123032
rect 674170 123030 674176 123094
rect 674240 123092 674246 123094
rect 674240 123032 676320 123092
rect 674240 123030 674246 123032
rect 143874 122500 143934 122988
rect 149199 122500 149265 122503
rect 143874 122498 149265 122500
rect 143874 122442 149204 122498
rect 149260 122442 149265 122498
rect 143874 122440 149265 122442
rect 149199 122437 149265 122440
rect 184335 122204 184401 122207
rect 184335 122202 190560 122204
rect 184335 122146 184340 122202
rect 184396 122146 190560 122202
rect 184335 122144 190560 122146
rect 184335 122141 184401 122144
rect 674362 122142 674368 122206
rect 674432 122204 674438 122206
rect 676290 122204 676350 122544
rect 674432 122144 676350 122204
rect 674432 122142 674438 122144
rect 646479 122056 646545 122059
rect 640194 122054 646545 122056
rect 640194 121998 646484 122054
rect 646540 121998 646545 122054
rect 640194 121996 646545 121998
rect 148911 121760 148977 121763
rect 143904 121758 148977 121760
rect 143904 121702 148916 121758
rect 148972 121702 148977 121758
rect 143904 121700 148977 121702
rect 148911 121697 148977 121700
rect 184527 121612 184593 121615
rect 184527 121610 190560 121612
rect 184527 121554 184532 121610
rect 184588 121554 190560 121610
rect 184527 121552 190560 121554
rect 184527 121549 184593 121552
rect 640194 121434 640254 121996
rect 646479 121993 646545 121996
rect 676047 122056 676113 122059
rect 676047 122054 676320 122056
rect 676047 121998 676052 122054
rect 676108 121998 676320 122054
rect 676047 121996 676320 121998
rect 676047 121993 676113 121996
rect 676290 121467 676350 121582
rect 676239 121462 676350 121467
rect 676239 121406 676244 121462
rect 676300 121406 676350 121462
rect 676239 121404 676350 121406
rect 676239 121401 676305 121404
rect 676047 121094 676113 121097
rect 676047 121092 676320 121094
rect 676047 121036 676052 121092
rect 676108 121036 676320 121092
rect 676047 121034 676320 121036
rect 676047 121031 676113 121034
rect 184335 120724 184401 120727
rect 184335 120722 190560 120724
rect 184335 120666 184340 120722
rect 184396 120666 190560 120722
rect 184335 120664 190560 120666
rect 184335 120661 184401 120664
rect 147471 120576 147537 120579
rect 143904 120574 147537 120576
rect 143904 120518 147476 120574
rect 147532 120518 147537 120574
rect 143904 120516 147537 120518
rect 147471 120513 147537 120516
rect 676047 120576 676113 120579
rect 676047 120574 676320 120576
rect 676047 120518 676052 120574
rect 676108 120518 676320 120574
rect 676047 120516 676320 120518
rect 676047 120513 676113 120516
rect 184431 120132 184497 120135
rect 184431 120130 190014 120132
rect 184431 120074 184436 120130
rect 184492 120074 190014 120130
rect 184431 120072 190014 120074
rect 184431 120069 184497 120072
rect 189954 120058 190014 120072
rect 189954 119998 190560 120058
rect 676143 119836 676209 119839
rect 676290 119836 676350 120102
rect 676143 119834 676350 119836
rect 676143 119778 676148 119834
rect 676204 119778 676350 119834
rect 676143 119776 676350 119778
rect 676143 119773 676209 119776
rect 647919 119540 647985 119543
rect 640416 119538 647985 119540
rect 640416 119482 647924 119538
rect 647980 119482 647985 119538
rect 640416 119480 647985 119482
rect 647919 119477 647985 119480
rect 149487 119392 149553 119395
rect 143904 119390 149553 119392
rect 143904 119334 149492 119390
rect 149548 119334 149553 119390
rect 143904 119332 149553 119334
rect 149487 119329 149553 119332
rect 676290 119247 676350 119510
rect 184527 119244 184593 119247
rect 184527 119242 190560 119244
rect 184527 119186 184532 119242
rect 184588 119186 190560 119242
rect 184527 119184 190560 119186
rect 676239 119242 676350 119247
rect 676239 119186 676244 119242
rect 676300 119186 676350 119242
rect 676239 119184 676350 119186
rect 184527 119181 184593 119184
rect 676239 119181 676305 119184
rect 184719 118652 184785 118655
rect 184719 118650 190014 118652
rect 184719 118594 184724 118650
rect 184780 118594 190014 118650
rect 184719 118592 190014 118594
rect 184719 118589 184785 118592
rect 189954 118578 190014 118592
rect 189954 118518 190560 118578
rect 149391 118208 149457 118211
rect 143874 118206 149457 118208
rect 143874 118150 149396 118206
rect 149452 118150 149457 118206
rect 143874 118148 149457 118150
rect 143874 118104 143934 118148
rect 149391 118145 149457 118148
rect 676666 117998 676672 118062
rect 676736 118060 676742 118062
rect 676815 118060 676881 118063
rect 676736 118058 676881 118060
rect 676736 118002 676820 118058
rect 676876 118002 676881 118058
rect 676736 118000 676881 118002
rect 676736 117998 676742 118000
rect 676815 117997 676881 118000
rect 675898 117850 675904 117914
rect 675968 117912 675974 117914
rect 676911 117912 676977 117915
rect 675968 117910 676977 117912
rect 675968 117854 676916 117910
rect 676972 117854 676977 117910
rect 675968 117852 676977 117854
rect 675968 117850 675974 117852
rect 676911 117849 676977 117852
rect 184335 117764 184401 117767
rect 184335 117762 190560 117764
rect 184335 117706 184340 117762
rect 184396 117706 190560 117762
rect 184335 117704 190560 117706
rect 184335 117701 184401 117704
rect 645231 117616 645297 117619
rect 640416 117614 645297 117616
rect 640416 117558 645236 117614
rect 645292 117558 645297 117614
rect 640416 117556 645297 117558
rect 645231 117553 645297 117556
rect 184431 117024 184497 117027
rect 184431 117022 190014 117024
rect 184431 116966 184436 117022
rect 184492 116966 190014 117022
rect 184431 116964 190014 116966
rect 184431 116961 184497 116964
rect 189954 116950 190014 116964
rect 189954 116890 190560 116950
rect 149487 116876 149553 116879
rect 143904 116874 149553 116876
rect 143904 116818 149492 116874
rect 149548 116818 149553 116874
rect 143904 116816 149553 116818
rect 149487 116813 149553 116816
rect 184527 116284 184593 116287
rect 184527 116282 190560 116284
rect 184527 116226 184532 116282
rect 184588 116226 190560 116282
rect 184527 116224 190560 116226
rect 184527 116221 184593 116224
rect 149391 115692 149457 115695
rect 647919 115692 647985 115695
rect 143904 115690 149457 115692
rect 143904 115634 149396 115690
rect 149452 115634 149457 115690
rect 143904 115632 149457 115634
rect 640416 115690 647985 115692
rect 640416 115634 647924 115690
rect 647980 115634 647985 115690
rect 640416 115632 647985 115634
rect 149391 115629 149457 115632
rect 647919 115629 647985 115632
rect 184623 115396 184689 115399
rect 184623 115394 190560 115396
rect 184623 115338 184628 115394
rect 184684 115338 190560 115394
rect 184623 115336 190560 115338
rect 184623 115333 184689 115336
rect 149103 115248 149169 115251
rect 149391 115248 149457 115251
rect 149103 115246 149457 115248
rect 149103 115190 149108 115246
rect 149164 115190 149396 115246
rect 149452 115190 149457 115246
rect 149103 115188 149457 115190
rect 149103 115185 149169 115188
rect 149391 115185 149457 115188
rect 184335 114804 184401 114807
rect 184335 114802 190560 114804
rect 184335 114746 184340 114802
rect 184396 114746 190560 114802
rect 184335 114744 190560 114746
rect 184335 114741 184401 114744
rect 149487 114508 149553 114511
rect 143904 114506 149553 114508
rect 143904 114450 149492 114506
rect 149548 114450 149553 114506
rect 143904 114448 149553 114450
rect 149487 114445 149553 114448
rect 184431 113916 184497 113919
rect 184431 113914 190560 113916
rect 184431 113858 184436 113914
rect 184492 113858 190560 113914
rect 184431 113856 190560 113858
rect 184431 113853 184497 113856
rect 149391 113176 149457 113179
rect 143904 113174 149457 113176
rect 143904 113118 149396 113174
rect 149452 113118 149457 113174
rect 143904 113116 149457 113118
rect 149391 113113 149457 113116
rect 184527 113176 184593 113179
rect 640194 113176 640254 113738
rect 646479 113176 646545 113179
rect 184527 113174 190560 113176
rect 184527 113118 184532 113174
rect 184588 113118 190560 113174
rect 184527 113116 190560 113118
rect 640194 113174 646545 113176
rect 640194 113118 646484 113174
rect 646540 113118 646545 113174
rect 640194 113116 646545 113118
rect 184527 113113 184593 113116
rect 646479 113113 646545 113116
rect 184623 112436 184689 112439
rect 184623 112434 190560 112436
rect 184623 112378 184628 112434
rect 184684 112378 190560 112434
rect 184623 112376 190560 112378
rect 184623 112373 184689 112376
rect 148431 111992 148497 111995
rect 143904 111990 148497 111992
rect 143904 111934 148436 111990
rect 148492 111934 148497 111990
rect 143904 111932 148497 111934
rect 148431 111929 148497 111932
rect 184335 111696 184401 111699
rect 184335 111694 190014 111696
rect 184335 111638 184340 111694
rect 184396 111638 190014 111694
rect 184335 111636 190014 111638
rect 184335 111633 184401 111636
rect 189954 111622 190014 111636
rect 189954 111562 190560 111622
rect 640386 111400 640446 111888
rect 647151 111400 647217 111403
rect 640386 111398 647217 111400
rect 640386 111342 647156 111398
rect 647212 111342 647217 111398
rect 640386 111340 647217 111342
rect 647151 111337 647217 111340
rect 149391 110956 149457 110959
rect 143904 110954 149457 110956
rect 143904 110898 149396 110954
rect 149452 110898 149457 110954
rect 143904 110896 149457 110898
rect 149391 110893 149457 110896
rect 184431 110956 184497 110959
rect 184431 110954 190560 110956
rect 184431 110898 184436 110954
rect 184492 110898 190560 110954
rect 184431 110896 190560 110898
rect 184431 110893 184497 110896
rect 184527 110216 184593 110219
rect 184527 110214 190014 110216
rect 184527 110158 184532 110214
rect 184588 110158 190014 110214
rect 184527 110156 190014 110158
rect 184527 110153 184593 110156
rect 189954 110142 190014 110156
rect 189954 110082 190560 110142
rect 143874 109624 143934 109668
rect 148623 109624 148689 109627
rect 143874 109622 148689 109624
rect 143874 109566 148628 109622
rect 148684 109566 148689 109622
rect 143874 109564 148689 109566
rect 148623 109561 148689 109564
rect 640386 109476 640446 109890
rect 646671 109476 646737 109479
rect 640386 109474 646737 109476
rect 640386 109418 646676 109474
rect 646732 109418 646737 109474
rect 640386 109416 646737 109418
rect 646671 109413 646737 109416
rect 184335 109328 184401 109331
rect 184335 109326 190560 109328
rect 184335 109270 184340 109326
rect 184396 109270 190560 109326
rect 184335 109268 190560 109270
rect 184335 109265 184401 109268
rect 185679 108736 185745 108739
rect 185679 108734 190014 108736
rect 185679 108678 185684 108734
rect 185740 108678 190014 108734
rect 185679 108676 190014 108678
rect 185679 108673 185745 108676
rect 189954 108662 190014 108676
rect 189954 108602 190560 108662
rect 147183 108440 147249 108443
rect 143904 108438 147249 108440
rect 143904 108382 147188 108438
rect 147244 108382 147249 108438
rect 143904 108380 147249 108382
rect 147183 108377 147249 108380
rect 646767 107996 646833 107999
rect 640416 107994 646833 107996
rect 640416 107938 646772 107994
rect 646828 107938 646833 107994
rect 640416 107936 646833 107938
rect 646767 107933 646833 107936
rect 186159 107848 186225 107851
rect 186159 107846 190560 107848
rect 186159 107790 186164 107846
rect 186220 107790 190560 107846
rect 186159 107788 190560 107790
rect 186159 107785 186225 107788
rect 673978 107638 673984 107702
rect 674048 107700 674054 107702
rect 675183 107700 675249 107703
rect 674048 107698 675249 107700
rect 674048 107642 675188 107698
rect 675244 107642 675249 107698
rect 674048 107640 675249 107642
rect 674048 107638 674054 107640
rect 675183 107637 675249 107640
rect 148335 107256 148401 107259
rect 143904 107254 148401 107256
rect 143904 107198 148340 107254
rect 148396 107198 148401 107254
rect 143904 107196 148401 107198
rect 148335 107193 148401 107196
rect 184431 107108 184497 107111
rect 184431 107106 190560 107108
rect 184431 107050 184436 107106
rect 184492 107050 190560 107106
rect 184431 107048 190560 107050
rect 184431 107045 184497 107048
rect 674362 106454 674368 106518
rect 674432 106516 674438 106518
rect 675087 106516 675153 106519
rect 674432 106514 675153 106516
rect 674432 106458 675092 106514
rect 675148 106458 675153 106514
rect 674432 106456 675153 106458
rect 674432 106454 674438 106456
rect 675087 106453 675153 106456
rect 185295 106368 185361 106371
rect 185295 106366 190560 106368
rect 185295 106310 185300 106366
rect 185356 106310 190560 106366
rect 185295 106308 190560 106310
rect 185295 106305 185361 106308
rect 148623 106072 148689 106075
rect 646095 106072 646161 106075
rect 143904 106070 148689 106072
rect 143904 106014 148628 106070
rect 148684 106014 148689 106070
rect 143904 106012 148689 106014
rect 640416 106070 646161 106072
rect 640416 106014 646100 106070
rect 646156 106014 646161 106070
rect 640416 106012 646161 106014
rect 148623 106009 148689 106012
rect 646095 106009 646161 106012
rect 665154 105631 665214 106082
rect 184335 105628 184401 105631
rect 184335 105626 190560 105628
rect 184335 105570 184340 105626
rect 184396 105570 190560 105626
rect 184335 105568 190560 105570
rect 665154 105626 665265 105631
rect 665154 105570 665204 105626
rect 665260 105570 665265 105626
rect 665154 105568 665265 105570
rect 184335 105565 184401 105568
rect 665199 105565 665265 105568
rect 674170 105566 674176 105630
rect 674240 105628 674246 105630
rect 675087 105628 675153 105631
rect 674240 105626 675153 105628
rect 674240 105570 675092 105626
rect 675148 105570 675153 105626
rect 674240 105568 675153 105570
rect 674240 105566 674246 105568
rect 675087 105565 675153 105568
rect 665346 105332 665406 105361
rect 665583 105332 665649 105335
rect 665346 105330 665649 105332
rect 665346 105274 665588 105330
rect 665644 105274 665649 105330
rect 665346 105272 665649 105274
rect 665583 105269 665649 105272
rect 665295 105184 665361 105187
rect 665295 105182 665406 105184
rect 665295 105126 665300 105182
rect 665356 105126 665406 105182
rect 665295 105121 665406 105126
rect 665346 104996 665406 105121
rect 184527 104888 184593 104891
rect 184527 104886 190014 104888
rect 184527 104830 184532 104886
rect 184588 104830 190014 104886
rect 184527 104828 190014 104830
rect 184527 104825 184593 104828
rect 189954 104814 190014 104828
rect 189954 104754 190560 104814
rect 148239 104740 148305 104743
rect 143904 104738 148305 104740
rect 143904 104682 148244 104738
rect 148300 104682 148305 104738
rect 143904 104680 148305 104682
rect 148239 104677 148305 104680
rect 647919 104148 647985 104151
rect 640416 104146 647985 104148
rect 640416 104090 647924 104146
rect 647980 104090 647985 104146
rect 640416 104088 647985 104090
rect 647919 104085 647985 104088
rect 184431 104000 184497 104003
rect 184431 103998 190560 104000
rect 184431 103942 184436 103998
rect 184492 103942 190560 103998
rect 184431 103940 190560 103942
rect 184431 103937 184497 103940
rect 148719 103556 148785 103559
rect 143904 103554 148785 103556
rect 143904 103498 148724 103554
rect 148780 103498 148785 103554
rect 143904 103496 148785 103498
rect 148719 103493 148785 103496
rect 184431 103408 184497 103411
rect 184431 103406 190014 103408
rect 184431 103350 184436 103406
rect 184492 103350 190014 103406
rect 184431 103348 190014 103350
rect 184431 103345 184497 103348
rect 189954 103334 190014 103348
rect 189954 103274 190560 103334
rect 675759 103260 675825 103263
rect 675898 103260 675904 103262
rect 675759 103258 675904 103260
rect 675759 103202 675764 103258
rect 675820 103202 675904 103258
rect 675759 103200 675904 103202
rect 675759 103197 675825 103200
rect 675898 103198 675904 103200
rect 675968 103198 675974 103262
rect 184335 102520 184401 102523
rect 184335 102518 190560 102520
rect 184335 102462 184340 102518
rect 184396 102462 190560 102518
rect 184335 102460 190560 102462
rect 184335 102457 184401 102460
rect 148527 102372 148593 102375
rect 143904 102370 148593 102372
rect 143904 102314 148532 102370
rect 148588 102314 148593 102370
rect 143904 102312 148593 102314
rect 148527 102309 148593 102312
rect 645135 102224 645201 102227
rect 640416 102222 645201 102224
rect 640416 102166 645140 102222
rect 645196 102166 645201 102222
rect 640416 102164 645201 102166
rect 645135 102161 645201 102164
rect 184527 101928 184593 101931
rect 184527 101926 190014 101928
rect 184527 101870 184532 101926
rect 184588 101870 190014 101926
rect 184527 101868 190014 101870
rect 184527 101865 184593 101868
rect 189954 101854 190014 101868
rect 189954 101794 190560 101854
rect 675759 101484 675825 101487
rect 676666 101484 676672 101486
rect 675759 101482 676672 101484
rect 675759 101426 675764 101482
rect 675820 101426 676672 101482
rect 675759 101424 676672 101426
rect 675759 101421 675825 101424
rect 676666 101422 676672 101424
rect 676736 101422 676742 101486
rect 143874 100892 143934 101084
rect 184623 101040 184689 101043
rect 184623 101038 190560 101040
rect 184623 100982 184628 101038
rect 184684 100982 190560 101038
rect 184623 100980 190560 100982
rect 184623 100977 184689 100980
rect 149391 100892 149457 100895
rect 143874 100890 149457 100892
rect 143874 100834 149396 100890
rect 149452 100834 149457 100890
rect 143874 100832 149457 100834
rect 149391 100829 149457 100832
rect 184335 100300 184401 100303
rect 184335 100298 190014 100300
rect 184335 100242 184340 100298
rect 184396 100242 190014 100298
rect 184335 100240 190014 100242
rect 184335 100237 184401 100240
rect 189954 100226 190014 100240
rect 189954 100166 190560 100226
rect 149487 99856 149553 99859
rect 143904 99854 149553 99856
rect 143904 99798 149492 99854
rect 149548 99798 149553 99854
rect 143904 99796 149553 99798
rect 149487 99793 149553 99796
rect 640194 99708 640254 100270
rect 647919 99708 647985 99711
rect 640194 99706 647985 99708
rect 640194 99650 647924 99706
rect 647980 99650 647985 99706
rect 640194 99648 647985 99650
rect 647919 99645 647985 99648
rect 184431 99560 184497 99563
rect 184431 99558 190560 99560
rect 184431 99502 184436 99558
rect 184492 99502 190560 99558
rect 184431 99500 190560 99502
rect 184431 99497 184497 99500
rect 149391 98672 149457 98675
rect 143904 98670 149457 98672
rect 143904 98614 149396 98670
rect 149452 98614 149457 98670
rect 143904 98612 149457 98614
rect 149391 98609 149457 98612
rect 184527 98672 184593 98675
rect 184527 98670 190560 98672
rect 184527 98614 184532 98670
rect 184588 98614 190560 98670
rect 184527 98612 190560 98614
rect 184527 98609 184593 98612
rect 184623 98080 184689 98083
rect 640386 98080 640446 98420
rect 647055 98080 647121 98083
rect 184623 98078 190560 98080
rect 184623 98022 184628 98078
rect 184684 98022 190560 98078
rect 184623 98020 190560 98022
rect 640386 98078 647121 98080
rect 640386 98022 647060 98078
rect 647116 98022 647121 98078
rect 640386 98020 647121 98022
rect 184623 98017 184689 98020
rect 647055 98017 647121 98020
rect 149487 97488 149553 97491
rect 143904 97486 149553 97488
rect 143904 97430 149492 97486
rect 149548 97430 149553 97486
rect 143904 97428 149553 97430
rect 149487 97425 149553 97428
rect 184335 97192 184401 97195
rect 184335 97190 190560 97192
rect 184335 97134 184340 97190
rect 184396 97134 190560 97190
rect 184335 97132 190560 97134
rect 184335 97129 184401 97132
rect 184431 96452 184497 96455
rect 184431 96450 190560 96452
rect 184431 96394 184436 96450
rect 184492 96394 190560 96450
rect 184431 96392 190560 96394
rect 184431 96389 184497 96392
rect 143874 95712 143934 96200
rect 640386 96008 640446 96570
rect 645423 96008 645489 96011
rect 640386 96006 645489 96008
rect 640386 95950 645428 96006
rect 645484 95950 645489 96006
rect 640386 95948 645489 95950
rect 645423 95945 645489 95948
rect 149391 95712 149457 95715
rect 143874 95710 149457 95712
rect 143874 95654 149396 95710
rect 149452 95654 149457 95710
rect 143874 95652 149457 95654
rect 149391 95649 149457 95652
rect 184719 95712 184785 95715
rect 184719 95710 190560 95712
rect 184719 95654 184724 95710
rect 184780 95654 190560 95710
rect 184719 95652 190560 95654
rect 184719 95649 184785 95652
rect 149295 94972 149361 94975
rect 143904 94970 149361 94972
rect 143904 94914 149300 94970
rect 149356 94914 149361 94970
rect 143904 94912 149361 94914
rect 149295 94909 149361 94912
rect 189954 94838 190560 94898
rect 184335 94824 184401 94827
rect 189954 94824 190014 94838
rect 184335 94822 190014 94824
rect 184335 94766 184340 94822
rect 184396 94766 190014 94822
rect 184335 94764 190014 94766
rect 184335 94761 184401 94764
rect 184431 94232 184497 94235
rect 184431 94230 190560 94232
rect 184431 94174 184436 94230
rect 184492 94174 190560 94230
rect 184431 94172 190560 94174
rect 184431 94169 184497 94172
rect 640386 94084 640446 94646
rect 647727 94084 647793 94087
rect 640386 94082 647793 94084
rect 640386 94026 647732 94082
rect 647788 94026 647793 94082
rect 640386 94024 647793 94026
rect 647727 94021 647793 94024
rect 149487 93788 149553 93791
rect 143904 93786 149553 93788
rect 143904 93730 149492 93786
rect 149548 93730 149553 93786
rect 143904 93728 149553 93730
rect 149487 93725 149553 93728
rect 184527 93492 184593 93495
rect 184527 93490 190014 93492
rect 184527 93434 184532 93490
rect 184588 93434 190014 93490
rect 184527 93432 190014 93434
rect 184527 93429 184593 93432
rect 189954 93418 190014 93432
rect 189954 93358 190560 93418
rect 184623 92752 184689 92755
rect 647823 92752 647889 92755
rect 184623 92750 190560 92752
rect 184623 92694 184628 92750
rect 184684 92694 190560 92750
rect 184623 92692 190560 92694
rect 640416 92750 647889 92752
rect 640416 92694 647828 92750
rect 647884 92694 647889 92750
rect 640416 92692 647889 92694
rect 184623 92689 184689 92692
rect 647823 92689 647889 92692
rect 149391 92604 149457 92607
rect 143904 92602 149457 92604
rect 143904 92546 149396 92602
rect 149452 92546 149457 92602
rect 143904 92544 149457 92546
rect 149391 92541 149457 92544
rect 184335 92012 184401 92015
rect 184335 92010 190014 92012
rect 184335 91954 184340 92010
rect 184396 91954 190014 92010
rect 184335 91952 190014 91954
rect 184335 91949 184401 91952
rect 189954 91938 190014 91952
rect 189954 91878 190560 91938
rect 149679 91420 149745 91423
rect 143904 91418 149745 91420
rect 143904 91362 149684 91418
rect 149740 91362 149745 91418
rect 143904 91360 149745 91362
rect 149679 91357 149745 91360
rect 184623 91124 184689 91127
rect 184623 91122 190560 91124
rect 184623 91066 184628 91122
rect 184684 91066 190560 91122
rect 184623 91064 190560 91066
rect 184623 91061 184689 91064
rect 659343 90828 659409 90831
rect 640416 90826 659409 90828
rect 640416 90770 659348 90826
rect 659404 90770 659409 90826
rect 640416 90768 659409 90770
rect 659343 90765 659409 90768
rect 184431 90384 184497 90387
rect 184431 90382 190560 90384
rect 184431 90326 184436 90382
rect 184492 90326 190560 90382
rect 184431 90324 190560 90326
rect 184431 90321 184497 90324
rect 149391 90236 149457 90239
rect 143904 90234 149457 90236
rect 143904 90178 149396 90234
rect 149452 90178 149457 90234
rect 143904 90176 149457 90178
rect 149391 90173 149457 90176
rect 184527 89644 184593 89647
rect 184527 89642 190560 89644
rect 184527 89586 184532 89642
rect 184588 89586 190560 89642
rect 184527 89584 190560 89586
rect 184527 89581 184593 89584
rect 149391 89052 149457 89055
rect 143904 89050 149457 89052
rect 143904 88994 149396 89050
rect 149452 88994 149457 89050
rect 143904 88992 149457 88994
rect 149391 88989 149457 88992
rect 184335 88904 184401 88907
rect 645903 88904 645969 88907
rect 184335 88902 190560 88904
rect 184335 88846 184340 88902
rect 184396 88846 190560 88902
rect 184335 88844 190560 88846
rect 640416 88902 645969 88904
rect 640416 88846 645908 88902
rect 645964 88846 645969 88902
rect 640416 88844 645969 88846
rect 184335 88841 184401 88844
rect 645903 88841 645969 88844
rect 184431 88164 184497 88167
rect 184431 88162 190014 88164
rect 184431 88106 184436 88162
rect 184492 88106 190014 88162
rect 184431 88104 190014 88106
rect 184431 88101 184497 88104
rect 189954 88090 190014 88104
rect 189954 88030 190560 88090
rect 143874 87276 143934 87764
rect 149487 87276 149553 87279
rect 143874 87274 149553 87276
rect 143874 87218 149492 87274
rect 149548 87218 149553 87274
rect 143874 87216 149553 87218
rect 149487 87213 149553 87216
rect 184527 87276 184593 87279
rect 184527 87274 190560 87276
rect 184527 87218 184532 87274
rect 184588 87218 190560 87274
rect 184527 87216 190560 87218
rect 184527 87213 184593 87216
rect 647919 87128 647985 87131
rect 640386 87126 647985 87128
rect 640386 87070 647924 87126
rect 647980 87070 647985 87126
rect 640386 87068 647985 87070
rect 640386 86950 640446 87068
rect 647919 87065 647985 87068
rect 653679 86980 653745 86983
rect 653679 86978 656736 86980
rect 653679 86922 653684 86978
rect 653740 86922 656736 86978
rect 653679 86920 656736 86922
rect 653679 86917 653745 86920
rect 184623 86684 184689 86687
rect 184623 86682 190014 86684
rect 184623 86626 184628 86682
rect 184684 86626 190014 86682
rect 184623 86624 190014 86626
rect 184623 86621 184689 86624
rect 189954 86610 190014 86624
rect 189954 86550 190560 86610
rect 148623 86536 148689 86539
rect 143904 86534 148689 86536
rect 143904 86478 148628 86534
rect 148684 86478 148689 86534
rect 143904 86476 148689 86478
rect 148623 86473 148689 86476
rect 663279 86388 663345 86391
rect 663234 86386 663345 86388
rect 663234 86330 663284 86386
rect 663340 86330 663345 86386
rect 663234 86325 663345 86330
rect 650895 86240 650961 86243
rect 650895 86238 656736 86240
rect 650895 86182 650900 86238
rect 650956 86182 656736 86238
rect 663234 86210 663294 86325
rect 650895 86180 656736 86182
rect 650895 86177 650961 86180
rect 184431 85796 184497 85799
rect 184431 85794 190560 85796
rect 184431 85738 184436 85794
rect 184492 85738 190560 85794
rect 184431 85736 190560 85738
rect 184431 85733 184497 85736
rect 148431 85352 148497 85355
rect 143904 85350 148497 85352
rect 143904 85294 148436 85350
rect 148492 85294 148497 85350
rect 143904 85292 148497 85294
rect 148431 85289 148497 85292
rect 652335 85352 652401 85355
rect 652335 85350 656736 85352
rect 652335 85294 652340 85350
rect 652396 85294 656736 85350
rect 652335 85292 656736 85294
rect 652335 85289 652401 85292
rect 184335 85204 184401 85207
rect 184335 85202 190014 85204
rect 184335 85146 184340 85202
rect 184396 85146 190014 85202
rect 184335 85144 190014 85146
rect 184335 85141 184401 85144
rect 189954 85130 190014 85144
rect 189954 85070 190560 85130
rect 640194 84464 640254 85026
rect 663234 84763 663294 85322
rect 663234 84758 663345 84763
rect 663234 84702 663284 84758
rect 663340 84702 663345 84758
rect 663234 84700 663345 84702
rect 663279 84697 663345 84700
rect 645711 84464 645777 84467
rect 640194 84462 645777 84464
rect 640194 84406 645716 84462
rect 645772 84406 645777 84462
rect 640194 84404 645777 84406
rect 645711 84401 645777 84404
rect 184527 84316 184593 84319
rect 653679 84316 653745 84319
rect 184527 84314 190560 84316
rect 184527 84258 184532 84314
rect 184588 84258 190560 84314
rect 184527 84256 190560 84258
rect 653679 84314 656736 84316
rect 653679 84258 653684 84314
rect 653740 84258 656736 84314
rect 653679 84256 656736 84258
rect 184527 84253 184593 84256
rect 653679 84253 653745 84256
rect 146991 84168 147057 84171
rect 143904 84166 147057 84168
rect 143904 84110 146996 84166
rect 147052 84110 147057 84166
rect 143904 84108 147057 84110
rect 146991 84105 147057 84108
rect 663426 84023 663486 84582
rect 663426 84018 663537 84023
rect 663426 83962 663476 84018
rect 663532 83962 663537 84018
rect 663426 83960 663537 83962
rect 663471 83957 663537 83960
rect 189954 83442 190560 83502
rect 184335 83428 184401 83431
rect 189954 83428 190014 83442
rect 184335 83426 190014 83428
rect 184335 83370 184340 83426
rect 184396 83370 190014 83426
rect 184335 83368 190014 83370
rect 652239 83428 652305 83431
rect 652239 83426 656736 83428
rect 652239 83370 652244 83426
rect 652300 83370 656736 83426
rect 652239 83368 656736 83370
rect 184335 83365 184401 83368
rect 652239 83365 652305 83368
rect 143874 82392 143934 82880
rect 186159 82836 186225 82839
rect 186159 82834 190560 82836
rect 186159 82778 186164 82834
rect 186220 82778 190560 82834
rect 186159 82776 190560 82778
rect 186159 82773 186225 82776
rect 640386 82688 640446 83176
rect 663426 82839 663486 83398
rect 663375 82834 663486 82839
rect 663375 82778 663380 82834
rect 663436 82778 663486 82834
rect 663375 82776 663486 82778
rect 663375 82773 663441 82776
rect 647919 82688 647985 82691
rect 640386 82686 647985 82688
rect 640386 82630 647924 82686
rect 647980 82630 647985 82686
rect 640386 82628 647985 82630
rect 647919 82625 647985 82628
rect 652431 82688 652497 82691
rect 652431 82686 656736 82688
rect 652431 82630 652436 82686
rect 652492 82630 656736 82686
rect 652431 82628 656736 82630
rect 652431 82625 652497 82628
rect 149199 82392 149265 82395
rect 143874 82390 149265 82392
rect 143874 82334 149204 82390
rect 149260 82334 149265 82390
rect 143874 82332 149265 82334
rect 149199 82329 149265 82332
rect 663234 82099 663294 82658
rect 663234 82094 663345 82099
rect 663234 82038 663284 82094
rect 663340 82038 663345 82094
rect 663234 82036 663345 82038
rect 663279 82033 663345 82036
rect 184239 81948 184305 81951
rect 184239 81946 190560 81948
rect 184239 81890 184244 81946
rect 184300 81890 190560 81946
rect 184239 81888 190560 81890
rect 184239 81885 184305 81888
rect 148335 81652 148401 81655
rect 143904 81650 148401 81652
rect 143904 81594 148340 81650
rect 148396 81594 148401 81650
rect 143904 81592 148401 81594
rect 148335 81589 148401 81592
rect 662415 81652 662481 81655
rect 663042 81652 663102 81770
rect 662415 81650 663102 81652
rect 662415 81594 662420 81650
rect 662476 81594 663102 81650
rect 662415 81592 663102 81594
rect 662415 81589 662481 81592
rect 184431 81356 184497 81359
rect 184431 81354 190560 81356
rect 184431 81298 184436 81354
rect 184492 81298 190560 81354
rect 184431 81296 190560 81298
rect 184431 81293 184497 81296
rect 640386 81060 640446 81326
rect 647919 81060 647985 81063
rect 640386 81058 647985 81060
rect 640386 81002 647924 81058
rect 647980 81002 647985 81058
rect 640386 81000 647985 81002
rect 647919 80997 647985 81000
rect 149295 80468 149361 80471
rect 143904 80466 149361 80468
rect 143904 80410 149300 80466
rect 149356 80410 149361 80466
rect 143904 80408 149361 80410
rect 149295 80405 149361 80408
rect 184623 80468 184689 80471
rect 184623 80466 190560 80468
rect 184623 80410 184628 80466
rect 184684 80410 190560 80466
rect 184623 80408 190560 80410
rect 184623 80405 184689 80408
rect 184431 79876 184497 79879
rect 184431 79874 190014 79876
rect 184431 79818 184436 79874
rect 184492 79818 190014 79874
rect 184431 79816 190014 79818
rect 184431 79813 184497 79816
rect 189954 79802 190014 79816
rect 189954 79742 190560 79802
rect 646671 79432 646737 79435
rect 640416 79430 646737 79432
rect 640416 79374 646676 79430
rect 646732 79374 646737 79430
rect 640416 79372 646737 79374
rect 646671 79369 646737 79372
rect 149583 79284 149649 79287
rect 143904 79282 149649 79284
rect 143904 79226 149588 79282
rect 149644 79226 149649 79282
rect 143904 79224 149649 79226
rect 149583 79221 149649 79224
rect 184335 78988 184401 78991
rect 184335 78986 190560 78988
rect 184335 78930 184340 78986
rect 184396 78930 190560 78986
rect 184335 78928 190560 78930
rect 184335 78925 184401 78928
rect 184527 78248 184593 78251
rect 184527 78246 190014 78248
rect 184527 78190 184532 78246
rect 184588 78190 190014 78246
rect 184527 78188 190014 78190
rect 184527 78185 184593 78188
rect 189954 78174 190014 78188
rect 189954 78114 190560 78174
rect 148815 77952 148881 77955
rect 143904 77950 148881 77952
rect 143904 77894 148820 77950
rect 148876 77894 148881 77950
rect 143904 77892 148881 77894
rect 148815 77889 148881 77892
rect 184431 77508 184497 77511
rect 647919 77508 647985 77511
rect 184431 77506 190560 77508
rect 184431 77450 184436 77506
rect 184492 77450 190560 77506
rect 184431 77448 190560 77450
rect 640416 77506 647985 77508
rect 640416 77450 647924 77506
rect 647980 77450 647985 77506
rect 640416 77448 647985 77450
rect 184431 77445 184497 77448
rect 647919 77445 647985 77448
rect 149391 76768 149457 76771
rect 143904 76766 149457 76768
rect 143904 76710 149396 76766
rect 149452 76710 149457 76766
rect 143904 76708 149457 76710
rect 149391 76705 149457 76708
rect 184335 76768 184401 76771
rect 184335 76766 190014 76768
rect 184335 76710 184340 76766
rect 184396 76710 190014 76766
rect 184335 76708 190014 76710
rect 184335 76705 184401 76708
rect 189954 76694 190014 76708
rect 189954 76634 190560 76694
rect 184623 76028 184689 76031
rect 184623 76026 190560 76028
rect 184623 75970 184628 76026
rect 184684 75970 190560 76026
rect 184623 75968 190560 75970
rect 184623 75965 184689 75968
rect 149487 75584 149553 75587
rect 646287 75584 646353 75587
rect 143904 75582 149553 75584
rect 143904 75526 149492 75582
rect 149548 75526 149553 75582
rect 143904 75524 149553 75526
rect 640416 75582 646353 75584
rect 640416 75526 646292 75582
rect 646348 75526 646353 75582
rect 640416 75524 646353 75526
rect 149487 75521 149553 75524
rect 646287 75521 646353 75524
rect 184527 75140 184593 75143
rect 184527 75138 190560 75140
rect 184527 75082 184532 75138
rect 184588 75082 190560 75138
rect 184527 75080 190560 75082
rect 184527 75077 184593 75080
rect 184335 74400 184401 74403
rect 184335 74398 190560 74400
rect 184335 74342 184340 74398
rect 184396 74342 190560 74398
rect 184335 74340 190560 74342
rect 184335 74337 184401 74340
rect 143874 73808 143934 74296
rect 149295 73808 149361 73811
rect 143874 73806 149361 73808
rect 143874 73750 149300 73806
rect 149356 73750 149361 73806
rect 143874 73748 149361 73750
rect 149295 73745 149361 73748
rect 184527 73660 184593 73663
rect 647919 73660 647985 73663
rect 184527 73658 190560 73660
rect 184527 73602 184532 73658
rect 184588 73602 190560 73658
rect 184527 73600 190560 73602
rect 640416 73658 647985 73660
rect 640416 73602 647924 73658
rect 647980 73602 647985 73658
rect 640416 73600 647985 73602
rect 184527 73597 184593 73600
rect 647919 73597 647985 73600
rect 149679 73068 149745 73071
rect 143904 73066 149745 73068
rect 143904 73010 149684 73066
rect 149740 73010 149745 73066
rect 143904 73008 149745 73010
rect 149679 73005 149745 73008
rect 184431 72920 184497 72923
rect 184431 72918 190560 72920
rect 184431 72862 184436 72918
rect 184492 72862 190560 72918
rect 184431 72860 190560 72862
rect 184431 72857 184497 72860
rect 184623 72180 184689 72183
rect 184623 72178 190560 72180
rect 184623 72122 184628 72178
rect 184684 72122 190560 72178
rect 184623 72120 190560 72122
rect 184623 72117 184689 72120
rect 149103 72032 149169 72035
rect 143904 72030 149169 72032
rect 143904 71974 149108 72030
rect 149164 71974 149169 72030
rect 143904 71972 149169 71974
rect 149103 71969 149169 71972
rect 646959 71884 647025 71887
rect 640386 71882 647025 71884
rect 640386 71826 646964 71882
rect 647020 71826 647025 71882
rect 640386 71824 647025 71826
rect 640386 71706 640446 71824
rect 646959 71821 647025 71824
rect 184335 71440 184401 71443
rect 184335 71438 190014 71440
rect 184335 71382 184340 71438
rect 184396 71382 190014 71438
rect 184335 71380 190014 71382
rect 184335 71377 184401 71380
rect 189954 71366 190014 71380
rect 189954 71306 190560 71366
rect 149487 70848 149553 70851
rect 143904 70846 149553 70848
rect 143904 70790 149492 70846
rect 149548 70790 149553 70846
rect 143904 70788 149553 70790
rect 149487 70785 149553 70788
rect 184431 70552 184497 70555
rect 184431 70550 190560 70552
rect 184431 70494 184436 70550
rect 184492 70494 190560 70550
rect 184431 70492 190560 70494
rect 184431 70489 184497 70492
rect 184527 69960 184593 69963
rect 184527 69958 190014 69960
rect 184527 69902 184532 69958
rect 184588 69902 190014 69958
rect 184527 69900 190014 69902
rect 184527 69897 184593 69900
rect 189954 69886 190014 69900
rect 189954 69826 190560 69886
rect 640386 69664 640446 69856
rect 647919 69664 647985 69667
rect 640386 69662 647985 69664
rect 640386 69606 647924 69662
rect 647980 69606 647985 69662
rect 640386 69604 647985 69606
rect 647919 69601 647985 69604
rect 149391 69516 149457 69519
rect 143904 69514 149457 69516
rect 143904 69458 149396 69514
rect 149452 69458 149457 69514
rect 143904 69456 149457 69458
rect 149391 69453 149457 69456
rect 184335 69072 184401 69075
rect 184335 69070 190560 69072
rect 184335 69014 184340 69070
rect 184396 69014 190560 69070
rect 184335 69012 190560 69014
rect 184335 69009 184401 69012
rect 646863 68628 646929 68631
rect 640194 68626 646929 68628
rect 640194 68570 646868 68626
rect 646924 68570 646929 68626
rect 640194 68568 646929 68570
rect 184335 68480 184401 68483
rect 184335 68478 190014 68480
rect 184335 68422 184340 68478
rect 184396 68422 190014 68478
rect 184335 68420 190014 68422
rect 184335 68417 184401 68420
rect 189954 68406 190014 68420
rect 189954 68346 190560 68406
rect 149295 68332 149361 68335
rect 143904 68330 149361 68332
rect 143904 68274 149300 68330
rect 149356 68274 149361 68330
rect 143904 68272 149361 68274
rect 149295 68269 149361 68272
rect 640194 68006 640254 68568
rect 646863 68565 646929 68568
rect 184527 67592 184593 67595
rect 184527 67590 190560 67592
rect 184527 67534 184532 67590
rect 184588 67534 190560 67590
rect 184527 67532 190560 67534
rect 184527 67529 184593 67532
rect 149199 67148 149265 67151
rect 143904 67146 149265 67148
rect 143904 67090 149204 67146
rect 149260 67090 149265 67146
rect 143904 67088 149265 67090
rect 149199 67085 149265 67088
rect 184431 66852 184497 66855
rect 184431 66850 190560 66852
rect 184431 66794 184436 66850
rect 184492 66794 190560 66850
rect 184431 66792 190560 66794
rect 184431 66789 184497 66792
rect 645999 66260 646065 66263
rect 640194 66258 646065 66260
rect 640194 66202 646004 66258
rect 646060 66202 646065 66258
rect 640194 66200 646065 66202
rect 184335 66112 184401 66115
rect 184335 66110 190560 66112
rect 184335 66054 184340 66110
rect 184396 66054 190560 66110
rect 640194 66082 640254 66200
rect 645999 66197 646065 66200
rect 184335 66052 190560 66054
rect 184335 66049 184401 66052
rect 143874 65372 143934 65860
rect 149391 65372 149457 65375
rect 143874 65370 149457 65372
rect 143874 65314 149396 65370
rect 149452 65314 149457 65370
rect 143874 65312 149457 65314
rect 149391 65309 149457 65312
rect 184527 65224 184593 65227
rect 184527 65222 190560 65224
rect 184527 65166 184532 65222
rect 184588 65166 190560 65222
rect 184527 65164 190560 65166
rect 184527 65161 184593 65164
rect 149487 64632 149553 64635
rect 143904 64630 149553 64632
rect 143904 64574 149492 64630
rect 149548 64574 149553 64630
rect 143904 64572 149553 64574
rect 149487 64569 149553 64572
rect 184431 64632 184497 64635
rect 184431 64630 190014 64632
rect 184431 64574 184436 64630
rect 184492 64574 190014 64630
rect 184431 64572 190014 64574
rect 184431 64569 184497 64572
rect 189954 64558 190014 64572
rect 189954 64498 190560 64558
rect 647919 64188 647985 64191
rect 640416 64186 647985 64188
rect 640416 64130 647924 64186
rect 647980 64130 647985 64186
rect 640416 64128 647985 64130
rect 647919 64125 647985 64128
rect 184335 63744 184401 63747
rect 184335 63742 190560 63744
rect 184335 63686 184340 63742
rect 184396 63686 190560 63742
rect 184335 63684 190560 63686
rect 184335 63681 184401 63684
rect 149583 63448 149649 63451
rect 143904 63446 149649 63448
rect 143904 63390 149588 63446
rect 149644 63390 149649 63446
rect 143904 63388 149649 63390
rect 149583 63385 149649 63388
rect 184431 63152 184497 63155
rect 184431 63150 190014 63152
rect 184431 63094 184436 63150
rect 184492 63094 190014 63150
rect 184431 63092 190014 63094
rect 184431 63089 184497 63092
rect 189954 63078 190014 63092
rect 189954 63018 190560 63078
rect 149391 62264 149457 62267
rect 143904 62262 149457 62264
rect 143904 62206 149396 62262
rect 149452 62206 149457 62262
rect 143904 62204 149457 62206
rect 149391 62201 149457 62204
rect 184335 62264 184401 62267
rect 647919 62264 647985 62267
rect 184335 62262 190560 62264
rect 184335 62206 184340 62262
rect 184396 62206 190560 62262
rect 184335 62204 190560 62206
rect 640416 62262 647985 62264
rect 640416 62206 647924 62262
rect 647980 62206 647985 62262
rect 640416 62204 647985 62206
rect 184335 62201 184401 62204
rect 647919 62201 647985 62204
rect 184623 61524 184689 61527
rect 184623 61522 190014 61524
rect 184623 61466 184628 61522
rect 184684 61466 190014 61522
rect 184623 61464 190014 61466
rect 184623 61461 184689 61464
rect 189954 61450 190014 61464
rect 189954 61390 190560 61450
rect 143874 60636 143934 60976
rect 184527 60784 184593 60787
rect 184527 60782 190560 60784
rect 184527 60726 184532 60782
rect 184588 60726 190560 60782
rect 184527 60724 190560 60726
rect 184527 60721 184593 60724
rect 149295 60636 149361 60639
rect 143874 60634 149361 60636
rect 143874 60578 149300 60634
rect 149356 60578 149361 60634
rect 143874 60576 149361 60578
rect 149295 60573 149361 60576
rect 647151 60340 647217 60343
rect 640416 60338 647217 60340
rect 640416 60282 647156 60338
rect 647212 60282 647217 60338
rect 640416 60280 647217 60282
rect 647151 60277 647217 60280
rect 184335 60044 184401 60047
rect 184335 60042 190014 60044
rect 184335 59986 184340 60042
rect 184396 59986 190014 60042
rect 184335 59984 190014 59986
rect 184335 59981 184401 59984
rect 189954 59970 190014 59984
rect 189954 59910 190560 59970
rect 149391 59748 149457 59751
rect 143904 59746 149457 59748
rect 143904 59690 149396 59746
rect 149452 59690 149457 59746
rect 143904 59688 149457 59690
rect 149391 59685 149457 59688
rect 184431 59304 184497 59307
rect 184431 59302 190560 59304
rect 184431 59246 184436 59302
rect 184492 59246 190560 59302
rect 184431 59244 190560 59246
rect 184431 59241 184497 59244
rect 645999 59008 646065 59011
rect 640386 59006 646065 59008
rect 640386 58950 646004 59006
rect 646060 58950 646065 59006
rect 640386 58948 646065 58950
rect 149391 58564 149457 58567
rect 143904 58562 149457 58564
rect 143904 58506 149396 58562
rect 149452 58506 149457 58562
rect 143904 58504 149457 58506
rect 149391 58501 149457 58504
rect 184527 58416 184593 58419
rect 184527 58414 190560 58416
rect 184527 58358 184532 58414
rect 184588 58358 190560 58414
rect 640386 58386 640446 58948
rect 645999 58945 646065 58948
rect 184527 58356 190560 58358
rect 184527 58353 184593 58356
rect 184335 57676 184401 57679
rect 184335 57674 190560 57676
rect 184335 57618 184340 57674
rect 184396 57618 190560 57674
rect 184335 57616 190560 57618
rect 184335 57613 184401 57616
rect 149487 57380 149553 57383
rect 143904 57378 149553 57380
rect 143904 57322 149492 57378
rect 149548 57322 149553 57378
rect 143904 57320 149553 57322
rect 149487 57317 149553 57320
rect 646767 57084 646833 57087
rect 640386 57082 646833 57084
rect 640386 57026 646772 57082
rect 646828 57026 646833 57082
rect 640386 57024 646833 57026
rect 184335 56936 184401 56939
rect 184335 56934 190560 56936
rect 184335 56878 184340 56934
rect 184396 56878 190560 56934
rect 184335 56876 190560 56878
rect 184335 56873 184401 56876
rect 640386 56536 640446 57024
rect 646767 57021 646833 57024
rect 149391 56196 149457 56199
rect 143874 56194 149457 56196
rect 143874 56138 149396 56194
rect 149452 56138 149457 56194
rect 143874 56136 149457 56138
rect 143874 56092 143934 56136
rect 149391 56133 149457 56136
rect 184335 56196 184401 56199
rect 184335 56194 190560 56196
rect 184335 56138 184340 56194
rect 184396 56138 190560 56194
rect 184335 56136 190560 56138
rect 184335 56133 184401 56136
rect 184431 55456 184497 55459
rect 184431 55454 190560 55456
rect 184431 55398 184436 55454
rect 184492 55398 190560 55454
rect 184431 55396 190560 55398
rect 184431 55393 184497 55396
rect 149679 54864 149745 54867
rect 143904 54862 149745 54864
rect 143904 54806 149684 54862
rect 149740 54806 149745 54862
rect 143904 54804 149745 54806
rect 149679 54801 149745 54804
rect 184335 54716 184401 54719
rect 646479 54716 646545 54719
rect 184335 54714 190014 54716
rect 184335 54658 184340 54714
rect 184396 54658 190014 54714
rect 184335 54656 190014 54658
rect 184335 54653 184401 54656
rect 189954 54642 190014 54656
rect 640386 54714 646545 54716
rect 640386 54658 646484 54714
rect 646540 54658 646545 54714
rect 640386 54656 646545 54658
rect 189954 54582 190560 54642
rect 640386 54612 640446 54656
rect 646479 54653 646545 54656
rect 184335 53976 184401 53979
rect 184335 53974 190560 53976
rect 184335 53918 184340 53974
rect 184396 53918 190560 53974
rect 184335 53916 190560 53918
rect 184335 53913 184401 53916
rect 149391 53828 149457 53831
rect 143904 53826 149457 53828
rect 143904 53770 149396 53826
rect 149452 53770 149457 53826
rect 143904 53768 149457 53770
rect 149391 53765 149457 53768
rect 302895 42136 302961 42139
rect 311151 42136 311217 42139
rect 302895 42134 311217 42136
rect 302895 42078 302900 42134
rect 302956 42078 311156 42134
rect 311212 42078 311217 42134
rect 302895 42076 311217 42078
rect 302895 42073 302961 42076
rect 311151 42073 311217 42076
rect 412527 42136 412593 42139
rect 412527 42134 437790 42136
rect 412527 42078 412532 42134
rect 412588 42078 437790 42134
rect 412527 42076 437790 42078
rect 412527 42073 412593 42076
rect 416847 41988 416913 41991
rect 416847 41986 417630 41988
rect 416847 41930 416852 41986
rect 416908 41930 417630 41986
rect 416847 41928 417630 41930
rect 416847 41925 416913 41928
rect 357711 41840 357777 41843
rect 362031 41840 362097 41843
rect 389199 41840 389265 41843
rect 357711 41838 361854 41840
rect 357711 41782 357716 41838
rect 357772 41782 361854 41838
rect 357711 41780 361854 41782
rect 357711 41777 357777 41780
rect 361794 40508 361854 41780
rect 362031 41838 389265 41840
rect 362031 41782 362036 41838
rect 362092 41782 389204 41838
rect 389260 41782 389265 41838
rect 362031 41780 389265 41782
rect 362031 41777 362097 41780
rect 389199 41777 389265 41780
rect 403215 40508 403281 40511
rect 361794 40506 403281 40508
rect 361794 40450 403220 40506
rect 403276 40450 403281 40506
rect 361794 40448 403281 40450
rect 417570 40508 417630 41928
rect 437730 40656 437790 42076
rect 467343 41840 467409 41843
rect 471663 41840 471729 41843
rect 522831 41840 522897 41843
rect 467343 41838 471486 41840
rect 467343 41782 467348 41838
rect 467404 41782 471486 41838
rect 467343 41780 471486 41782
rect 467343 41777 467409 41780
rect 471426 40804 471486 41780
rect 471663 41838 478110 41840
rect 471663 41782 471668 41838
rect 471724 41782 478110 41838
rect 471663 41780 478110 41782
rect 471663 41777 471729 41780
rect 478050 40804 478110 41780
rect 498210 41838 522897 41840
rect 498210 41782 522836 41838
rect 522892 41782 522897 41838
rect 498210 41780 522897 41782
rect 498210 40804 498270 41780
rect 522831 41777 522897 41780
rect 471426 40744 475902 40804
rect 478050 40744 498270 40804
rect 475695 40656 475761 40659
rect 437730 40654 475761 40656
rect 437730 40598 475700 40654
rect 475756 40598 475761 40654
rect 437730 40596 475761 40598
rect 475695 40593 475761 40596
rect 458607 40508 458673 40511
rect 417570 40506 458673 40508
rect 417570 40450 458612 40506
rect 458668 40450 458673 40506
rect 417570 40448 458673 40450
rect 475842 40508 475902 40744
rect 541455 40508 541521 40511
rect 475842 40506 541521 40508
rect 475842 40450 541460 40506
rect 541516 40450 541521 40506
rect 475842 40448 541521 40450
rect 403215 40445 403281 40448
rect 458607 40445 458673 40448
rect 541455 40445 541521 40448
rect 142095 40360 142161 40363
rect 141762 40358 142161 40360
rect 141762 40302 142100 40358
rect 142156 40302 142161 40358
rect 141762 40300 142161 40302
rect 141762 39886 141822 40300
rect 142095 40297 142161 40300
rect 311055 37252 311121 37255
rect 334095 37252 334161 37255
rect 311055 37250 334161 37252
rect 311055 37194 311060 37250
rect 311116 37194 334100 37250
rect 334156 37194 334161 37250
rect 311055 37192 334161 37194
rect 311055 37189 311121 37192
rect 334095 37189 334161 37192
<< via3 >>
rect 40384 815078 40448 815142
rect 40576 814042 40640 814106
rect 41344 810194 41408 810258
rect 41536 802254 41600 802318
rect 41728 800426 41792 800490
rect 42496 800426 42560 800490
rect 42304 800278 42368 800342
rect 42304 796726 42368 796790
rect 42496 794358 42560 794422
rect 41728 792878 41792 792942
rect 41536 791842 41600 791906
rect 41344 791694 41408 791758
rect 674944 788290 675008 788354
rect 675520 787166 675584 787170
rect 675532 787110 675584 787166
rect 675520 787106 675584 787110
rect 674752 786218 674816 786282
rect 675328 784798 675392 784802
rect 675328 784742 675380 784798
rect 675328 784738 675392 784742
rect 674176 784294 674240 784358
rect 673984 783406 674048 783470
rect 676672 782962 676736 783026
rect 676096 780594 676160 780658
rect 676480 780002 676544 780066
rect 676288 778818 676352 778882
rect 40576 772306 40640 772370
rect 40192 771862 40256 771926
rect 40384 771862 40448 771926
rect 675520 771862 675584 771926
rect 40576 770826 40640 770890
rect 40768 758838 40832 758902
rect 40960 757506 41024 757570
rect 40768 746258 40832 746322
rect 40960 745962 41024 746026
rect 676288 745370 676352 745434
rect 676864 745370 676928 745434
rect 674368 742410 674432 742474
rect 675712 741730 675776 741734
rect 675724 741674 675776 741730
rect 675712 741670 675776 741674
rect 676480 741522 676544 741586
rect 677056 741522 677120 741586
rect 675136 740042 675200 740106
rect 675904 739154 675968 739218
rect 674560 738562 674624 738626
rect 676480 735010 676544 735074
rect 675520 734478 675584 734482
rect 675532 734422 675584 734478
rect 675520 734418 675584 734422
rect 676288 734270 676352 734334
rect 40576 729238 40640 729302
rect 40384 728706 40448 728710
rect 40384 728650 40436 728706
rect 40436 728650 40448 728706
rect 40384 728646 40448 728650
rect 676864 728054 676928 728118
rect 677440 728054 677504 728118
rect 40576 727610 40640 727674
rect 40576 717304 40640 717368
rect 40384 715770 40448 715834
rect 42688 711626 42752 711690
rect 42688 711182 42752 711246
rect 674752 711182 674816 711246
rect 674944 710442 675008 710506
rect 675328 709702 675392 709766
rect 676096 709406 676160 709470
rect 674176 707630 674240 707694
rect 673984 707038 674048 707102
rect 677440 705854 677504 705918
rect 677248 705410 677312 705474
rect 677056 704966 677120 705030
rect 40576 702894 40640 702958
rect 40384 702746 40448 702810
rect 675328 697922 675392 697926
rect 675328 697866 675380 697922
rect 675328 697862 675392 697866
rect 674176 697122 674240 697186
rect 674752 696974 674816 697038
rect 676288 694902 676352 694966
rect 674944 694606 675008 694670
rect 673984 693422 674048 693486
rect 677056 686762 677120 686826
rect 40384 685430 40448 685494
rect 40576 684394 40640 684458
rect 40768 672856 40832 672920
rect 42496 671282 42560 671286
rect 42496 671226 42508 671282
rect 42508 671226 42560 671282
rect 42496 671222 42560 671226
rect 42304 671074 42368 671138
rect 42112 670630 42176 670694
rect 42112 668410 42176 668474
rect 42496 667730 42560 667734
rect 42496 667674 42508 667730
rect 42508 667674 42560 667730
rect 42496 667670 42560 667674
rect 675712 666190 675776 666254
rect 676480 665302 676544 665366
rect 675136 664710 675200 664774
rect 674368 663378 674432 663442
rect 675904 662638 675968 662702
rect 674560 662046 674624 662110
rect 40768 660862 40832 660926
rect 675520 661158 675584 661222
rect 676864 660418 676928 660482
rect 42304 659530 42368 659594
rect 674368 652130 674432 652194
rect 675520 651450 675584 651454
rect 675532 651394 675584 651450
rect 675520 651390 675584 651394
rect 674560 650946 674624 651010
rect 675712 649822 675776 649826
rect 675724 649766 675776 649822
rect 675712 649762 675776 649766
rect 675136 648342 675200 648346
rect 675136 648286 675188 648342
rect 675136 648282 675200 648286
rect 676480 648282 676544 648346
rect 676096 645322 676160 645386
rect 40576 644730 40640 644794
rect 41728 642510 41792 642574
rect 40384 642214 40448 642278
rect 43072 642214 43136 642278
rect 40576 628006 40640 628070
rect 40384 627858 40448 627922
rect 674752 620902 674816 620966
rect 675328 619866 675392 619930
rect 676288 619274 676352 619338
rect 674176 617942 674240 618006
rect 674944 617794 675008 617858
rect 673984 616906 674048 616970
rect 40576 616462 40640 616526
rect 40384 616314 40448 616378
rect 677056 615130 677120 615194
rect 674176 607730 674240 607794
rect 674944 607434 675008 607498
rect 675904 606398 675968 606462
rect 674752 604770 674816 604834
rect 41728 602166 41792 602170
rect 41728 602110 41740 602166
rect 41740 602110 41792 602166
rect 41728 602106 41792 602110
rect 675328 602018 675392 602022
rect 675340 601962 675392 602018
rect 675328 601958 675392 601962
rect 676288 600182 676352 600246
rect 42880 587514 42944 587518
rect 42880 587458 42932 587514
rect 42932 587458 42944 587514
rect 42880 587454 42944 587458
rect 40384 586212 40448 586276
rect 40576 585916 40640 585980
rect 42880 577302 42944 577306
rect 42880 577246 42892 577302
rect 42892 577246 42944 577302
rect 42880 577242 42944 577246
rect 40384 573986 40448 574050
rect 675520 573986 675584 574050
rect 40576 573838 40640 573902
rect 674560 572802 674624 572866
rect 675712 572506 675776 572570
rect 676096 572210 676160 572274
rect 674368 571174 674432 571238
rect 675136 570434 675200 570498
rect 676480 570138 676544 570202
rect 674368 562886 674432 562950
rect 675520 561762 675584 561766
rect 675532 561706 675584 561762
rect 675520 561702 675584 561706
rect 675136 561406 675200 561470
rect 674560 558890 674624 558954
rect 677056 554598 677120 554662
rect 676864 553266 676928 553330
rect 40384 539798 40448 539862
rect 41536 538022 41600 538086
rect 43072 536986 43136 537050
rect 40960 536246 41024 536310
rect 40768 535062 40832 535126
rect 41344 534174 41408 534238
rect 40576 533878 40640 533942
rect 41920 533050 41984 533054
rect 41920 532994 41932 533050
rect 41932 532994 41984 533050
rect 41920 532990 41984 532994
rect 41152 530770 41216 530834
rect 675904 530770 675968 530834
rect 41728 530090 41792 530094
rect 41728 530034 41780 530090
rect 41780 530034 41792 530090
rect 41728 530030 41792 530034
rect 674176 529882 674240 529946
rect 42112 529350 42176 529354
rect 42112 529294 42164 529350
rect 42164 529294 42176 529350
rect 42112 529290 42176 529294
rect 674752 529290 674816 529354
rect 676288 528994 676352 529058
rect 674944 527810 675008 527874
rect 42496 527218 42560 527282
rect 42304 527130 42368 527134
rect 675328 527218 675392 527282
rect 42304 527074 42316 527130
rect 42316 527074 42368 527130
rect 42304 527070 42368 527074
rect 675136 486370 675200 486434
rect 674368 485630 674432 485694
rect 675520 483410 675584 483474
rect 674560 482818 674624 482882
rect 676864 481042 676928 481106
rect 40768 480746 40832 480810
rect 42688 480746 42752 480810
rect 677056 480598 677120 480662
rect 40576 478082 40640 478146
rect 40576 473198 40640 473262
rect 43072 473050 43136 473114
rect 42496 471570 42560 471634
rect 41536 471274 41600 471338
rect 42304 470090 42368 470154
rect 42304 470002 42368 470006
rect 42304 469946 42316 470002
rect 42316 469946 42368 470002
rect 42304 469942 42368 469946
rect 41920 469498 41984 469562
rect 40576 469350 40640 469414
rect 42112 468018 42176 468082
rect 41728 467426 41792 467490
rect 40960 467278 41024 467342
rect 41344 466834 41408 466898
rect 41152 466242 41216 466306
rect 40768 465798 40832 465862
rect 42688 465058 42752 465122
rect 40576 423886 40640 423950
rect 41728 423442 41792 423506
rect 40768 422850 40832 422914
rect 40960 422406 41024 422470
rect 42112 422110 42176 422174
rect 41152 420926 41216 420990
rect 41920 420778 41984 420842
rect 42112 406066 42176 406070
rect 42112 406010 42124 406066
rect 42124 406010 42176 406066
rect 42112 406006 42176 406010
rect 40960 402010 41024 402074
rect 40576 400086 40640 400150
rect 673984 399642 674048 399706
rect 41152 399494 41216 399558
rect 40768 398754 40832 398818
rect 675712 398606 675776 398670
rect 676288 397866 676352 397930
rect 674368 397570 674432 397634
rect 676288 396386 676352 396450
rect 676672 395794 676736 395858
rect 676096 395350 676160 395414
rect 675328 394610 675392 394674
rect 674752 393278 674816 393342
rect 675520 393130 675584 393194
rect 675904 392168 675968 392232
rect 675136 391650 675200 391714
rect 41920 388080 41984 388144
rect 676480 384694 676544 384758
rect 41728 383214 41792 383278
rect 676288 382918 676352 382982
rect 675328 382326 675392 382390
rect 40576 381290 40640 381354
rect 40768 380254 40832 380318
rect 41344 379662 41408 379726
rect 41728 378774 41792 378838
rect 676672 378774 676736 378838
rect 40960 378182 41024 378246
rect 675904 378034 675968 378098
rect 41152 377738 41216 377802
rect 675520 377206 675584 377210
rect 675532 377150 675584 377206
rect 675520 377146 675584 377150
rect 675136 376466 675200 376470
rect 675136 376410 675188 376466
rect 675136 376406 675200 376410
rect 674752 375666 674816 375730
rect 674368 374334 674432 374398
rect 676096 371966 676160 372030
rect 41152 359238 41216 359302
rect 41344 358794 41408 358858
rect 40576 356870 40640 356934
rect 40960 356426 41024 356490
rect 40768 355538 40832 355602
rect 673984 355982 674048 356046
rect 673984 355834 674048 355898
rect 674176 355242 674240 355306
rect 675712 354650 675776 354714
rect 674368 354206 674432 354270
rect 674560 353170 674624 353234
rect 674752 350950 674816 351014
rect 674944 348730 675008 348794
rect 41728 343166 41792 343170
rect 41728 343110 41740 343166
rect 41740 343110 41792 343166
rect 41728 343106 41792 343110
rect 675904 342958 675968 343022
rect 675712 342810 675776 342874
rect 40576 338518 40640 338582
rect 40768 338074 40832 338138
rect 40960 337038 41024 337102
rect 41344 336594 41408 336658
rect 41152 334966 41216 335030
rect 41536 334522 41600 334586
rect 675712 333546 675776 333550
rect 675712 333490 675764 333546
rect 675712 333486 675776 333490
rect 674944 332302 675008 332366
rect 675904 330526 675968 330590
rect 674560 328158 674624 328222
rect 674752 326826 674816 326890
rect 41536 316170 41600 316234
rect 41344 315430 41408 315494
rect 40768 313654 40832 313718
rect 41152 313210 41216 313274
rect 40960 312322 41024 312386
rect 673984 310990 674048 311054
rect 673984 310398 674048 310462
rect 674176 309806 674240 309870
rect 676864 309658 676928 309722
rect 674560 309066 674624 309130
rect 674368 308918 674432 308982
rect 675904 308326 675968 308390
rect 676288 307586 676352 307650
rect 674752 307438 674816 307502
rect 675328 306402 675392 306466
rect 675712 305958 675776 306022
rect 674176 305366 674240 305430
rect 674944 303442 675008 303506
rect 675136 302702 675200 302766
rect 676096 302554 676160 302618
rect 675520 301962 675584 302026
rect 676480 301074 676544 301138
rect 40960 294858 41024 294922
rect 676288 294562 676352 294626
rect 40768 293822 40832 293886
rect 41536 293378 41600 293442
rect 675328 292846 675392 292850
rect 675328 292790 675380 292846
rect 675328 292786 675392 292790
rect 41152 291898 41216 291962
rect 41344 291306 41408 291370
rect 676096 290714 676160 290778
rect 675712 288554 675776 288558
rect 675724 288498 675776 288554
rect 675712 288494 675776 288498
rect 675520 287814 675584 287818
rect 675520 287758 675572 287814
rect 675520 287754 675584 287758
rect 675136 287162 675200 287226
rect 676480 286570 676544 286634
rect 674944 285534 675008 285598
rect 674752 283166 674816 283230
rect 674176 282130 674240 282194
rect 40576 278578 40640 278642
rect 676864 278430 676928 278494
rect 675904 278282 675968 278346
rect 43072 276358 43136 276422
rect 42304 273546 42368 273610
rect 41344 272954 41408 273018
rect 41536 272362 41600 272426
rect 40960 270586 41024 270650
rect 674560 270586 674624 270650
rect 41152 269994 41216 270058
rect 40768 269106 40832 269170
rect 675328 266442 675392 266506
rect 674368 266294 674432 266358
rect 673984 265702 674048 265766
rect 674176 264962 674240 265026
rect 674560 263186 674624 263250
rect 674752 262150 674816 262214
rect 676288 261410 676352 261474
rect 675712 260670 675776 260734
rect 675136 258302 675200 258366
rect 674944 257710 675008 257774
rect 675904 253270 675968 253334
rect 40384 251642 40448 251706
rect 676288 250754 676352 250818
rect 40576 250606 40640 250670
rect 41152 250162 41216 250226
rect 40768 248682 40832 248746
rect 40960 248090 41024 248154
rect 675712 243562 675776 243566
rect 675724 243506 675776 243562
rect 675712 243502 675776 243506
rect 674944 241874 675008 241938
rect 675136 241046 675200 241050
rect 675136 240990 675188 241046
rect 675136 240986 675200 240990
rect 674752 238174 674816 238238
rect 397504 236990 397568 237054
rect 675904 236842 675968 236906
rect 397696 236694 397760 236758
rect 407296 236694 407360 236758
rect 407680 236250 407744 236314
rect 413632 236102 413696 236166
rect 414016 236102 414080 236166
rect 40960 229738 41024 229802
rect 41152 229146 41216 229210
rect 40384 227370 40448 227434
rect 40768 226778 40832 226842
rect 40576 225890 40640 225954
rect 674176 220562 674240 220626
rect 674176 219970 674240 220034
rect 673984 219082 674048 219146
rect 674368 219082 674432 219146
rect 674560 218490 674624 218554
rect 674368 217898 674432 217962
rect 675328 217898 675392 217962
rect 675712 217602 675776 217666
rect 675904 215530 675968 215594
rect 674560 213014 674624 213078
rect 40384 208426 40448 208490
rect 40576 207834 40640 207898
rect 676672 207538 676736 207602
rect 676480 207390 676544 207454
rect 40960 206946 41024 207010
rect 40768 205466 40832 205530
rect 41152 204874 41216 204938
rect 675712 204490 675776 204494
rect 675724 204434 675776 204490
rect 675712 204430 675776 204434
rect 675904 198362 675968 198426
rect 674560 194810 674624 194874
rect 676480 193478 676544 193542
rect 676672 191554 676736 191618
rect 41152 186670 41216 186734
rect 40960 185782 41024 185846
rect 40384 184154 40448 184218
rect 40768 183562 40832 183626
rect 40576 182822 40640 182886
rect 674176 176162 674240 176226
rect 674560 175570 674624 175634
rect 673984 175422 674048 175486
rect 673984 174682 674048 174746
rect 674368 174090 674432 174154
rect 674176 173498 674240 173562
rect 676480 172906 676544 172970
rect 674752 172610 674816 172674
rect 675520 171278 675584 171342
rect 674944 171130 675008 171194
rect 676288 170390 676352 170454
rect 675328 168614 675392 168678
rect 675136 168170 675200 168234
rect 675904 167578 675968 167642
rect 675712 167134 675776 167198
rect 676096 166246 676160 166310
rect 676480 159290 676544 159354
rect 675520 157722 675584 157726
rect 675532 157666 675584 157722
rect 675520 157662 675584 157666
rect 675904 155442 675968 155506
rect 674944 155294 675008 155358
rect 675136 152542 675200 152546
rect 675136 152486 675188 152542
rect 675136 152482 675200 152486
rect 675712 152542 675776 152546
rect 675724 152486 675776 152542
rect 675712 152482 675776 152486
rect 676096 151298 676160 151362
rect 675328 150262 675392 150326
rect 674752 149670 674816 149734
rect 676288 146562 676352 146626
rect 674368 130578 674432 130642
rect 673984 129394 674048 129458
rect 674176 128506 674240 128570
rect 673984 125546 674048 125610
rect 674176 123030 674240 123094
rect 674368 122142 674432 122206
rect 676672 117998 676736 118062
rect 675904 117850 675968 117914
rect 673984 107638 674048 107702
rect 674368 106454 674432 106518
rect 674176 105566 674240 105630
rect 675904 103198 675968 103262
rect 676672 101422 676736 101486
<< metal4 >>
rect 40383 815142 40449 815143
rect 40383 815078 40384 815142
rect 40448 815078 40449 815142
rect 40383 815077 40449 815078
rect 40386 779004 40446 815077
rect 40575 814106 40641 814107
rect 40575 814042 40576 814106
rect 40640 814042 40641 814106
rect 40575 814041 40641 814042
rect 39938 778944 40446 779004
rect 40578 779046 40638 814041
rect 41343 810258 41409 810259
rect 41343 810194 41344 810258
rect 41408 810194 41409 810258
rect 41343 810193 41409 810194
rect 41346 791759 41406 810193
rect 41535 802318 41601 802319
rect 41535 802254 41536 802318
rect 41600 802254 41601 802318
rect 41535 802253 41601 802254
rect 41538 791907 41598 802253
rect 41727 800490 41793 800491
rect 41727 800426 41728 800490
rect 41792 800426 41793 800490
rect 41727 800425 41793 800426
rect 42495 800490 42561 800491
rect 42495 800426 42496 800490
rect 42560 800426 42561 800490
rect 42495 800425 42561 800426
rect 41730 792943 41790 800425
rect 42303 800342 42369 800343
rect 42303 800278 42304 800342
rect 42368 800278 42369 800342
rect 42303 800277 42369 800278
rect 42306 796791 42366 800277
rect 42303 796790 42369 796791
rect 42303 796726 42304 796790
rect 42368 796726 42369 796790
rect 42303 796725 42369 796726
rect 42498 794423 42558 800425
rect 42495 794422 42561 794423
rect 42495 794358 42496 794422
rect 42560 794358 42561 794422
rect 42495 794357 42561 794358
rect 41727 792942 41793 792943
rect 41727 792878 41728 792942
rect 41792 792878 41793 792942
rect 41727 792877 41793 792878
rect 41535 791906 41601 791907
rect 41535 791842 41536 791906
rect 41600 791842 41601 791906
rect 41535 791841 41601 791842
rect 41343 791758 41409 791759
rect 41343 791694 41344 791758
rect 41408 791694 41409 791758
rect 41343 791693 41409 791694
rect 674943 788354 675009 788355
rect 674943 788290 674944 788354
rect 675008 788290 675009 788354
rect 674943 788289 675009 788290
rect 674751 786282 674817 786283
rect 674751 786218 674752 786282
rect 674816 786218 674817 786282
rect 674751 786217 674817 786218
rect 674175 784358 674241 784359
rect 674175 784294 674176 784358
rect 674240 784294 674241 784358
rect 674175 784293 674241 784294
rect 673983 783470 674049 783471
rect 673983 783406 673984 783470
rect 674048 783406 674049 783470
rect 673983 783405 674049 783406
rect 40578 778986 41271 779046
rect 39938 777498 39998 778944
rect 41211 777498 41271 778986
rect 39938 777438 40446 777498
rect 40386 771927 40446 777438
rect 40578 777438 41271 777498
rect 40578 772371 40638 777438
rect 40575 772370 40641 772371
rect 40575 772306 40576 772370
rect 40640 772306 40641 772370
rect 40575 772305 40641 772306
rect 40191 771926 40257 771927
rect 40191 771862 40192 771926
rect 40256 771862 40257 771926
rect 40191 771861 40257 771862
rect 40383 771926 40449 771927
rect 40383 771862 40384 771926
rect 40448 771862 40449 771926
rect 40383 771861 40449 771862
rect 40194 771591 40254 771861
rect 40194 771531 40446 771591
rect 40386 736026 40446 771531
rect 40575 770890 40641 770891
rect 40575 770826 40576 770890
rect 40640 770826 40641 770890
rect 40575 770825 40641 770826
rect 39901 735966 40446 736026
rect 40578 736079 40638 770825
rect 40767 758902 40833 758903
rect 40767 758838 40768 758902
rect 40832 758838 40833 758902
rect 40767 758837 40833 758838
rect 40770 746323 40830 758837
rect 40959 757570 41025 757571
rect 40959 757506 40960 757570
rect 41024 757506 41025 757570
rect 40959 757505 41025 757506
rect 40767 746322 40833 746323
rect 40767 746258 40768 746322
rect 40832 746258 40833 746322
rect 40767 746257 40833 746258
rect 40962 746027 41022 757505
rect 40959 746026 41025 746027
rect 40959 745962 40960 746026
rect 41024 745962 41025 746026
rect 40959 745961 41025 745962
rect 40578 736019 41279 736079
rect 39901 734331 39961 735966
rect 41219 734331 41279 736019
rect 39901 734271 40446 734331
rect 40386 728711 40446 734271
rect 40578 734271 41279 734331
rect 40578 729303 40638 734271
rect 40575 729302 40641 729303
rect 40575 729238 40576 729302
rect 40640 729238 40641 729302
rect 40575 729237 40641 729238
rect 40383 728710 40449 728711
rect 40383 728646 40384 728710
rect 40448 728646 40449 728710
rect 40383 728645 40449 728646
rect 40578 727675 40638 729237
rect 40575 727674 40641 727675
rect 40575 727610 40576 727674
rect 40640 727610 40641 727674
rect 40575 727609 40641 727610
rect 673986 725634 674046 783405
rect 669711 725574 674046 725634
rect 40575 717368 40641 717369
rect 40575 717304 40576 717368
rect 40640 717304 40641 717368
rect 40575 717303 40641 717304
rect 40383 715834 40449 715835
rect 40383 715770 40384 715834
rect 40448 715770 40449 715834
rect 40383 715769 40449 715770
rect 40386 702811 40446 715769
rect 40578 702959 40638 717303
rect 669711 714927 669771 725574
rect 674178 725442 674238 784293
rect 674367 742474 674433 742475
rect 674367 742410 674368 742474
rect 674432 742410 674433 742474
rect 674367 742409 674433 742410
rect 669903 725382 674238 725442
rect 669903 715119 669963 725382
rect 674370 725250 674430 742409
rect 674559 738626 674625 738627
rect 674559 738562 674560 738626
rect 674624 738562 674625 738626
rect 674559 738561 674625 738562
rect 670095 725190 674430 725250
rect 670095 715311 670155 725190
rect 674562 725058 674622 738561
rect 670287 724998 674622 725058
rect 670287 715503 670347 724998
rect 674754 724866 674814 786217
rect 670479 724806 674814 724866
rect 670479 715695 670539 724806
rect 674946 724674 675006 788289
rect 675519 787170 675585 787171
rect 675519 787166 675520 787170
rect 675519 787110 675532 787166
rect 675519 787106 675520 787110
rect 675584 787106 675585 787170
rect 675519 787105 675585 787106
rect 675327 784802 675393 784803
rect 675327 784738 675328 784802
rect 675392 784798 675393 784802
rect 675380 784742 675393 784798
rect 675392 784738 675393 784742
rect 675327 784737 675393 784738
rect 675135 740106 675201 740107
rect 675135 740042 675136 740106
rect 675200 740042 675201 740106
rect 675135 740041 675201 740042
rect 670671 724614 675006 724674
rect 670671 715887 670731 724614
rect 675138 724482 675198 740041
rect 670863 724422 675198 724482
rect 670863 716079 670923 724422
rect 675330 724290 675390 784737
rect 675522 771927 675582 787105
rect 676671 783026 676737 783027
rect 676671 782962 676672 783026
rect 676736 782962 676737 783026
rect 676671 782961 676737 782962
rect 676095 780658 676161 780659
rect 676095 780594 676096 780658
rect 676160 780594 676161 780658
rect 676095 780593 676161 780594
rect 675519 771926 675585 771927
rect 675519 771862 675520 771926
rect 675584 771862 675585 771926
rect 675519 771861 675585 771862
rect 675711 741734 675777 741735
rect 675711 741730 675712 741734
rect 675711 741674 675724 741730
rect 675711 741670 675712 741674
rect 675776 741670 675777 741734
rect 675711 741669 675777 741670
rect 675519 734482 675585 734483
rect 675519 734478 675520 734482
rect 675519 734422 675532 734478
rect 675519 734418 675520 734422
rect 675584 734418 675585 734482
rect 675519 734417 675585 734418
rect 671055 724230 675390 724290
rect 671055 716271 671115 724230
rect 675522 724098 675582 734417
rect 671247 724038 675582 724098
rect 671247 716463 671307 724038
rect 675714 723906 675774 741669
rect 675903 739218 675969 739219
rect 675903 739154 675904 739218
rect 675968 739154 675969 739218
rect 675903 739153 675969 739154
rect 671439 723846 675774 723906
rect 671439 716655 671499 723846
rect 675906 723714 675966 739153
rect 671631 723654 675966 723714
rect 671631 716847 671691 723654
rect 676098 723522 676158 780593
rect 676479 780066 676545 780067
rect 676479 780002 676480 780066
rect 676544 780002 676545 780066
rect 676479 780001 676545 780002
rect 676287 778882 676353 778883
rect 676287 778818 676288 778882
rect 676352 778818 676353 778882
rect 676287 778817 676353 778818
rect 676290 745435 676350 778817
rect 676287 745434 676353 745435
rect 676287 745370 676288 745434
rect 676352 745370 676353 745434
rect 676287 745369 676353 745370
rect 676482 741587 676542 780001
rect 676479 741586 676545 741587
rect 676479 741522 676480 741586
rect 676544 741522 676545 741586
rect 676479 741521 676545 741522
rect 676479 735074 676545 735075
rect 676479 735010 676480 735074
rect 676544 735010 676545 735074
rect 676479 735009 676545 735010
rect 676287 734334 676353 734335
rect 676287 734270 676288 734334
rect 676352 734270 676353 734334
rect 676287 734269 676353 734270
rect 671823 723462 676158 723522
rect 671823 717039 671883 723462
rect 676290 723138 676350 734269
rect 676482 727635 676542 735009
rect 676674 731550 676734 782961
rect 676863 745434 676929 745435
rect 676863 745370 676864 745434
rect 676928 745370 676929 745434
rect 676863 745369 676929 745370
rect 676866 740289 676926 745369
rect 677055 741586 677121 741587
rect 677055 741522 677056 741586
rect 677120 741522 677121 741586
rect 677055 741521 677121 741522
rect 677058 740955 677118 741521
rect 677058 740895 677310 740955
rect 676866 740229 677118 740289
rect 676674 731490 676926 731550
rect 676866 728119 676926 731490
rect 676863 728118 676929 728119
rect 676863 728054 676864 728118
rect 676928 728054 676929 728118
rect 676863 728053 676929 728054
rect 676482 727575 676926 727635
rect 672207 723078 676350 723138
rect 672207 717423 672267 723078
rect 676866 722754 676926 727575
rect 672591 722694 676926 722754
rect 672591 717807 672651 722694
rect 677058 722562 677118 740229
rect 672783 722502 677118 722562
rect 672783 717999 672843 722502
rect 677250 722370 677310 740895
rect 677439 728118 677505 728119
rect 677439 728054 677440 728118
rect 677504 728054 677505 728118
rect 677439 728053 677505 728054
rect 672975 722310 677310 722370
rect 672975 718191 673035 722310
rect 677442 722178 677502 728053
rect 673167 722118 677502 722178
rect 673167 718383 673227 722118
rect 673167 718323 677502 718383
rect 672975 718131 677310 718191
rect 672783 717939 677118 717999
rect 672591 717747 676926 717807
rect 672207 717363 676542 717423
rect 671823 716979 676158 717039
rect 671631 716787 675966 716847
rect 671439 716595 675774 716655
rect 671247 716403 675582 716463
rect 671055 716211 675390 716271
rect 670863 716019 675198 716079
rect 670671 715827 675006 715887
rect 670479 715635 674814 715695
rect 670287 715443 674622 715503
rect 670095 715251 674430 715311
rect 669903 715059 674238 715119
rect 669711 714867 674046 714927
rect 42687 711690 42753 711691
rect 42687 711626 42688 711690
rect 42752 711626 42753 711690
rect 42687 711625 42753 711626
rect 42690 711247 42750 711625
rect 42687 711246 42753 711247
rect 42687 711182 42688 711246
rect 42752 711182 42753 711246
rect 42687 711181 42753 711182
rect 673986 707103 674046 714867
rect 674178 707695 674238 715059
rect 674175 707694 674241 707695
rect 674175 707630 674176 707694
rect 674240 707630 674241 707694
rect 674175 707629 674241 707630
rect 673983 707102 674049 707103
rect 673983 707038 673984 707102
rect 674048 707038 674049 707102
rect 673983 707037 674049 707038
rect 40575 702958 40641 702959
rect 40575 702894 40576 702958
rect 40640 702894 40641 702958
rect 40575 702893 40641 702894
rect 40383 702810 40449 702811
rect 40383 702746 40384 702810
rect 40448 702746 40449 702810
rect 40383 702745 40449 702746
rect 674175 697186 674241 697187
rect 674175 697122 674176 697186
rect 674240 697122 674241 697186
rect 674175 697121 674241 697122
rect 673983 693486 674049 693487
rect 673983 693422 673984 693486
rect 674048 693422 674049 693486
rect 673983 693421 674049 693422
rect 40383 685494 40449 685495
rect 40383 685430 40384 685494
rect 40448 685430 40449 685494
rect 40383 685429 40449 685430
rect 40386 649363 40446 685429
rect 40575 684458 40641 684459
rect 40575 684394 40576 684458
rect 40640 684394 40641 684458
rect 40575 684393 40641 684394
rect 39954 649303 40446 649363
rect 40578 649367 40638 684393
rect 673986 679840 674046 693421
rect 669777 679780 674046 679840
rect 40767 672920 40833 672921
rect 40767 672856 40768 672920
rect 40832 672856 40833 672920
rect 40767 672855 40833 672856
rect 40770 660927 40830 672855
rect 42495 671286 42561 671287
rect 42495 671222 42496 671286
rect 42560 671222 42561 671286
rect 42495 671221 42561 671222
rect 42303 671138 42369 671139
rect 42303 671074 42304 671138
rect 42368 671074 42369 671138
rect 42303 671073 42369 671074
rect 42111 670694 42177 670695
rect 42111 670630 42112 670694
rect 42176 670630 42177 670694
rect 42111 670629 42177 670630
rect 42114 668475 42174 670629
rect 42111 668474 42177 668475
rect 42111 668410 42112 668474
rect 42176 668410 42177 668474
rect 42111 668409 42177 668410
rect 40767 660926 40833 660927
rect 40767 660862 40768 660926
rect 40832 660862 40833 660926
rect 40767 660861 40833 660862
rect 42306 659595 42366 671073
rect 42498 667735 42558 671221
rect 669777 670459 669837 679780
rect 674178 679648 674238 697121
rect 669969 679588 674238 679648
rect 669969 670651 670029 679588
rect 674370 679456 674430 715251
rect 670161 679396 674430 679456
rect 670161 670843 670221 679396
rect 674562 679264 674622 715443
rect 674754 711247 674814 715635
rect 674751 711246 674817 711247
rect 674751 711182 674752 711246
rect 674816 711182 674817 711246
rect 674751 711181 674817 711182
rect 674946 710507 675006 715827
rect 674943 710506 675009 710507
rect 674943 710442 674944 710506
rect 675008 710442 675009 710506
rect 674943 710441 675009 710442
rect 674751 697038 674817 697039
rect 674751 696974 674752 697038
rect 674816 696974 674817 697038
rect 674751 696973 674817 696974
rect 670353 679204 674622 679264
rect 670353 671035 670413 679204
rect 674754 679072 674814 696973
rect 674943 694670 675009 694671
rect 674943 694606 674944 694670
rect 675008 694606 675009 694670
rect 674943 694605 675009 694606
rect 670545 679012 674814 679072
rect 670545 671227 670605 679012
rect 674946 678880 675006 694605
rect 670737 678820 675006 678880
rect 670737 671419 670797 678820
rect 675138 678688 675198 716019
rect 675330 709767 675390 716211
rect 675327 709766 675393 709767
rect 675327 709702 675328 709766
rect 675392 709702 675393 709766
rect 675327 709701 675393 709702
rect 675327 697926 675393 697927
rect 675327 697862 675328 697926
rect 675392 697922 675393 697926
rect 675380 697866 675393 697922
rect 675392 697862 675393 697866
rect 675327 697861 675393 697862
rect 670929 678628 675198 678688
rect 670929 671611 670989 678628
rect 675330 678496 675390 697861
rect 671121 678436 675390 678496
rect 671121 671803 671181 678436
rect 675522 678304 675582 716403
rect 671313 678244 675582 678304
rect 671313 671995 671373 678244
rect 675714 678112 675774 716595
rect 671505 678052 675774 678112
rect 671505 672187 671565 678052
rect 675906 677920 675966 716787
rect 676098 709471 676158 716979
rect 676095 709470 676161 709471
rect 676095 709406 676096 709470
rect 676160 709406 676161 709470
rect 676095 709405 676161 709406
rect 676287 694966 676353 694967
rect 676287 694902 676288 694966
rect 676352 694902 676353 694966
rect 676287 694901 676353 694902
rect 671697 677860 675966 677920
rect 671697 672379 671757 677860
rect 676290 677536 676350 694901
rect 672081 677476 676350 677536
rect 672081 672763 672141 677476
rect 676482 677344 676542 717363
rect 672273 677284 676542 677344
rect 672273 672955 672333 677284
rect 676866 676960 676926 717747
rect 677058 705031 677118 717939
rect 677250 705475 677310 718131
rect 677442 705919 677502 718323
rect 677439 705918 677505 705919
rect 677439 705854 677440 705918
rect 677504 705854 677505 705918
rect 677439 705853 677505 705854
rect 677247 705474 677313 705475
rect 677247 705410 677248 705474
rect 677312 705410 677313 705474
rect 677247 705409 677313 705410
rect 677055 705030 677121 705031
rect 677055 704966 677056 705030
rect 677120 704966 677121 705030
rect 677055 704965 677121 704966
rect 677055 686826 677121 686827
rect 677055 686762 677056 686826
rect 677120 686762 677121 686826
rect 677055 686761 677121 686762
rect 672657 676900 676926 676960
rect 672657 673339 672717 676900
rect 677058 676768 677118 686761
rect 672849 676708 677118 676768
rect 672849 673531 672909 676708
rect 672849 673471 677118 673531
rect 672657 673279 676926 673339
rect 672273 672895 676542 672955
rect 672081 672703 676350 672763
rect 671697 672319 675966 672379
rect 671505 672127 675774 672187
rect 671313 671935 675582 671995
rect 671121 671743 675390 671803
rect 670929 671551 675198 671611
rect 670737 671359 675006 671419
rect 670545 671167 674814 671227
rect 670353 670975 674622 671035
rect 670161 670783 674430 670843
rect 669969 670591 674238 670651
rect 669777 670399 674046 670459
rect 42495 667734 42561 667735
rect 42495 667670 42496 667734
rect 42560 667670 42561 667734
rect 42495 667669 42561 667670
rect 42303 659594 42369 659595
rect 42303 659530 42304 659594
rect 42368 659530 42369 659594
rect 42303 659529 42369 659530
rect 40578 649307 41286 649367
rect 39954 648068 40014 649303
rect 41226 648070 41286 649307
rect 40386 648068 40446 648070
rect 39954 648008 40446 648068
rect 40386 642279 40446 648008
rect 40578 648010 41286 648070
rect 40578 644795 40638 648010
rect 40575 644794 40641 644795
rect 40575 644730 40576 644794
rect 40640 644730 40641 644794
rect 40575 644729 40641 644730
rect 41727 642574 41793 642575
rect 41727 642510 41728 642574
rect 41792 642510 41793 642574
rect 41727 642509 41793 642510
rect 40383 642278 40449 642279
rect 40383 642214 40384 642278
rect 40448 642214 40449 642278
rect 40383 642213 40449 642214
rect 40575 628070 40641 628071
rect 40575 628006 40576 628070
rect 40640 628006 40641 628070
rect 40575 628005 40641 628006
rect 40383 627922 40449 627923
rect 40383 627858 40384 627922
rect 40448 627858 40449 627922
rect 40383 627857 40449 627858
rect 40386 616379 40446 627857
rect 40578 616527 40638 628005
rect 40575 616526 40641 616527
rect 40575 616462 40576 616526
rect 40640 616462 40641 616526
rect 40575 616461 40641 616462
rect 40383 616378 40449 616379
rect 40383 616314 40384 616378
rect 40448 616314 40449 616378
rect 40383 616313 40449 616314
rect 41730 604917 41790 642509
rect 43071 642278 43137 642279
rect 43071 642214 43072 642278
rect 43136 642214 43137 642278
rect 43071 642213 43137 642214
rect 41730 604857 42537 604917
rect 42477 603532 42537 604857
rect 41730 603472 42537 603532
rect 41730 602171 41790 603472
rect 41727 602170 41793 602171
rect 41727 602106 41728 602170
rect 41792 602106 41793 602170
rect 41727 602105 41793 602106
rect 42879 587518 42945 587519
rect 42879 587454 42880 587518
rect 42944 587454 42945 587518
rect 42879 587453 42945 587454
rect 40383 586276 40449 586277
rect 40383 586212 40384 586276
rect 40448 586212 40449 586276
rect 40383 586211 40449 586212
rect 40386 574051 40446 586211
rect 40575 585980 40641 585981
rect 40575 585916 40576 585980
rect 40640 585916 40641 585980
rect 40575 585915 40641 585916
rect 40383 574050 40449 574051
rect 40383 573986 40384 574050
rect 40448 573986 40449 574050
rect 40383 573985 40449 573986
rect 40578 573903 40638 585915
rect 42882 577307 42942 587453
rect 42879 577306 42945 577307
rect 42879 577242 42880 577306
rect 42944 577242 42945 577306
rect 42879 577241 42945 577242
rect 40575 573902 40641 573903
rect 40575 573838 40576 573902
rect 40640 573838 40641 573902
rect 40575 573837 40641 573838
rect 40383 539862 40449 539863
rect 40383 539798 40384 539862
rect 40448 539798 40449 539862
rect 40383 539797 40449 539798
rect 40386 479329 40446 539797
rect 41535 538086 41601 538087
rect 41535 538022 41536 538086
rect 41600 538022 41601 538086
rect 41535 538021 41601 538022
rect 40959 536310 41025 536311
rect 40959 536246 40960 536310
rect 41024 536246 41025 536310
rect 40959 536245 41025 536246
rect 40767 535126 40833 535127
rect 40767 535062 40768 535126
rect 40832 535062 40833 535126
rect 40767 535061 40833 535062
rect 40575 533942 40641 533943
rect 40575 533878 40576 533942
rect 40640 533878 40641 533942
rect 40575 533877 40641 533878
rect 40578 480549 40638 533877
rect 40770 480811 40830 535061
rect 40767 480810 40833 480811
rect 40767 480746 40768 480810
rect 40832 480746 40833 480810
rect 40767 480745 40833 480746
rect 40578 480489 40830 480549
rect 39982 479269 40446 479329
rect 39982 478038 40042 479269
rect 40770 479199 40830 480489
rect 40962 479375 41022 536245
rect 41343 534238 41409 534239
rect 41343 534174 41344 534238
rect 41408 534174 41409 534238
rect 41343 534173 41409 534174
rect 41151 530834 41217 530835
rect 41151 530770 41152 530834
rect 41216 530770 41217 530834
rect 41151 530769 41217 530770
rect 41154 479503 41214 530769
rect 41346 479673 41406 534173
rect 41538 479815 41598 538021
rect 43074 537051 43134 642213
rect 673986 633270 674046 670399
rect 671687 633210 674046 633270
rect 671687 627746 671747 633210
rect 674178 633078 674238 670591
rect 674370 663443 674430 670783
rect 674367 663442 674433 663443
rect 674367 663378 674368 663442
rect 674432 663378 674433 663442
rect 674367 663377 674433 663378
rect 674562 662111 674622 670975
rect 674559 662110 674625 662111
rect 674559 662046 674560 662110
rect 674624 662046 674625 662110
rect 674559 662045 674625 662046
rect 674367 652194 674433 652195
rect 674367 652130 674368 652194
rect 674432 652130 674433 652194
rect 674367 652129 674433 652130
rect 671879 633018 674238 633078
rect 671879 627938 671939 633018
rect 674370 632886 674430 652129
rect 674559 651010 674625 651011
rect 674559 650946 674560 651010
rect 674624 650946 674625 651010
rect 674559 650945 674625 650946
rect 672071 632826 674430 632886
rect 672071 628130 672131 632826
rect 674562 632694 674622 650945
rect 672263 632634 674622 632694
rect 672263 628322 672323 632634
rect 674754 632502 674814 671167
rect 672455 632442 674814 632502
rect 672455 628514 672515 632442
rect 674946 632310 675006 671359
rect 675138 664775 675198 671551
rect 675135 664774 675201 664775
rect 675135 664710 675136 664774
rect 675200 664710 675201 664774
rect 675135 664709 675201 664710
rect 675135 648346 675201 648347
rect 675135 648282 675136 648346
rect 675200 648342 675201 648346
rect 675188 648286 675201 648342
rect 675200 648282 675201 648286
rect 675135 648281 675201 648282
rect 672647 632250 675006 632310
rect 672647 628706 672707 632250
rect 675138 632118 675198 648281
rect 672839 632058 675198 632118
rect 672839 628898 672899 632058
rect 675330 631926 675390 671743
rect 675522 661223 675582 671935
rect 675714 666255 675774 672127
rect 675711 666254 675777 666255
rect 675711 666190 675712 666254
rect 675776 666190 675777 666254
rect 675711 666189 675777 666190
rect 675906 662703 675966 672319
rect 675903 662702 675969 662703
rect 675903 662638 675904 662702
rect 675968 662638 675969 662702
rect 675903 662637 675969 662638
rect 675519 661222 675585 661223
rect 675519 661158 675520 661222
rect 675584 661158 675585 661222
rect 675519 661157 675585 661158
rect 675519 651454 675585 651455
rect 675519 651450 675520 651454
rect 675519 651394 675532 651450
rect 675519 651390 675520 651394
rect 675584 651390 675585 651454
rect 675519 651389 675585 651390
rect 673031 631866 675390 631926
rect 673031 629090 673091 631866
rect 675522 631734 675582 651389
rect 675711 649826 675777 649827
rect 675711 649822 675712 649826
rect 675711 649766 675724 649822
rect 675711 649762 675712 649766
rect 675776 649762 675777 649826
rect 675711 649761 675777 649762
rect 673223 631674 675582 631734
rect 673223 629282 673283 631674
rect 675714 631542 675774 649761
rect 676095 645386 676161 645387
rect 676095 645322 676096 645386
rect 676160 645322 676161 645386
rect 676095 645321 676161 645322
rect 673415 631482 675774 631542
rect 673415 629474 673475 631482
rect 676098 630257 676158 645321
rect 675954 630197 676158 630257
rect 673415 629414 675774 629474
rect 673223 629222 675582 629282
rect 673031 629030 675390 629090
rect 672839 628838 675198 628898
rect 672647 628646 675006 628706
rect 672455 628454 674814 628514
rect 672263 628262 674622 628322
rect 672071 628070 674430 628130
rect 671879 627878 674238 627938
rect 671687 627686 674046 627746
rect 673986 616971 674046 627686
rect 674178 618007 674238 627878
rect 674175 618006 674241 618007
rect 674175 617942 674176 618006
rect 674240 617942 674241 618006
rect 674175 617941 674241 617942
rect 673983 616970 674049 616971
rect 673983 616906 673984 616970
rect 674048 616906 674049 616970
rect 673983 616905 674049 616906
rect 674175 607794 674241 607795
rect 674175 607730 674176 607794
rect 674240 607730 674241 607794
rect 674175 607729 674241 607730
rect 674178 589071 674238 607729
rect 670595 589011 674238 589071
rect 670595 580018 670655 589011
rect 674370 588879 674430 628070
rect 670787 588819 674430 588879
rect 670787 580210 670847 588819
rect 674562 588687 674622 628262
rect 674754 620967 674814 628454
rect 674751 620966 674817 620967
rect 674751 620902 674752 620966
rect 674816 620902 674817 620966
rect 674751 620901 674817 620902
rect 674946 617859 675006 628646
rect 674943 617858 675009 617859
rect 674943 617794 674944 617858
rect 675008 617794 675009 617858
rect 674943 617793 675009 617794
rect 674943 607498 675009 607499
rect 674943 607434 674944 607498
rect 675008 607434 675009 607498
rect 674943 607433 675009 607434
rect 674751 604834 674817 604835
rect 674751 604770 674752 604834
rect 674816 604770 674817 604834
rect 674751 604769 674817 604770
rect 670979 588627 674622 588687
rect 670979 580402 671039 588627
rect 674754 588495 674814 604769
rect 671171 588435 674814 588495
rect 671171 580594 671231 588435
rect 674946 588303 675006 607433
rect 671363 588243 675006 588303
rect 671363 580786 671423 588243
rect 675138 588111 675198 628838
rect 675330 619931 675390 629030
rect 675327 619930 675393 619931
rect 675327 619866 675328 619930
rect 675392 619866 675393 619930
rect 675327 619865 675393 619866
rect 675327 602022 675393 602023
rect 675327 602018 675328 602022
rect 675327 601962 675340 602018
rect 675327 601958 675328 601962
rect 675392 601958 675393 602022
rect 675327 601957 675393 601958
rect 671555 588051 675198 588111
rect 671555 580978 671615 588051
rect 675330 587919 675390 601957
rect 671747 587859 675390 587919
rect 671747 581170 671807 587859
rect 675522 587727 675582 629222
rect 671939 587667 675582 587727
rect 671939 581362 671999 587667
rect 675714 587535 675774 629414
rect 675954 628407 676014 630197
rect 676290 630096 676350 672703
rect 676482 665367 676542 672895
rect 676479 665366 676545 665367
rect 676479 665302 676480 665366
rect 676544 665302 676545 665366
rect 676479 665301 676545 665302
rect 676866 660483 676926 673279
rect 676863 660482 676929 660483
rect 676863 660418 676864 660482
rect 676928 660418 676929 660482
rect 676863 660417 676929 660418
rect 676479 648346 676545 648347
rect 676479 648282 676480 648346
rect 676544 648282 676545 648346
rect 676479 648281 676545 648282
rect 676160 630036 676350 630096
rect 676482 630096 676542 648281
rect 677058 630319 677118 673471
rect 677058 630259 677631 630319
rect 676482 630036 677391 630096
rect 676160 628786 676220 630036
rect 676160 628726 676350 628786
rect 675954 628347 676158 628407
rect 675903 606462 675969 606463
rect 675903 606398 675904 606462
rect 675968 606398 675969 606462
rect 675903 606397 675969 606398
rect 672131 587475 675774 587535
rect 672131 581554 672191 587475
rect 675906 587343 675966 606397
rect 672323 587283 675966 587343
rect 672323 581746 672383 587283
rect 676098 587151 676158 628347
rect 676290 619339 676350 628726
rect 677331 628518 677391 630036
rect 676482 628458 677391 628518
rect 676287 619338 676353 619339
rect 676287 619274 676288 619338
rect 676352 619274 676353 619338
rect 676287 619273 676353 619274
rect 676287 600246 676353 600247
rect 676287 600182 676288 600246
rect 676352 600182 676353 600246
rect 676287 600181 676353 600182
rect 672515 587091 676158 587151
rect 672515 581938 672575 587091
rect 676290 586959 676350 600181
rect 672707 586899 676350 586959
rect 672707 582130 672767 586899
rect 676482 586767 676542 628458
rect 677571 628337 677631 630259
rect 677058 628277 677631 628337
rect 677058 615195 677118 628277
rect 677055 615194 677121 615195
rect 677055 615130 677056 615194
rect 677120 615130 677121 615194
rect 677055 615129 677121 615130
rect 672899 586707 676542 586767
rect 672899 582322 672959 586707
rect 672899 582262 676542 582322
rect 672707 582070 676350 582130
rect 672515 581878 676158 581938
rect 672323 581686 675966 581746
rect 672131 581494 675774 581554
rect 671939 581302 675582 581362
rect 671747 581110 675390 581170
rect 671555 580918 675198 580978
rect 671363 580726 675006 580786
rect 671171 580534 674814 580594
rect 670979 580342 674622 580402
rect 670787 580150 674430 580210
rect 670595 579958 674238 580018
rect 674178 542465 674238 579958
rect 674370 571239 674430 580150
rect 674562 572867 674622 580342
rect 674559 572866 674625 572867
rect 674559 572802 674560 572866
rect 674624 572802 674625 572866
rect 674559 572801 674625 572802
rect 674367 571238 674433 571239
rect 674367 571174 674368 571238
rect 674432 571174 674433 571238
rect 674367 571173 674433 571174
rect 674367 562950 674433 562951
rect 674367 562886 674368 562950
rect 674432 562886 674433 562950
rect 674367 562885 674433 562886
rect 672301 542405 674238 542465
rect 672301 537329 672361 542405
rect 674370 542273 674430 562885
rect 674559 558954 674625 558955
rect 674559 558890 674560 558954
rect 674624 558890 674625 558954
rect 674559 558889 674625 558890
rect 672493 542213 674430 542273
rect 672493 537521 672553 542213
rect 674562 542081 674622 558889
rect 672685 542021 674622 542081
rect 672685 537713 672745 542021
rect 674754 541889 674814 580534
rect 672877 541829 674814 541889
rect 672877 537905 672937 541829
rect 674946 541697 675006 580726
rect 675138 570499 675198 580918
rect 675135 570498 675201 570499
rect 675135 570434 675136 570498
rect 675200 570434 675201 570498
rect 675135 570433 675201 570434
rect 675135 561470 675201 561471
rect 675135 561406 675136 561470
rect 675200 561406 675201 561470
rect 675135 561405 675201 561406
rect 673069 541637 675006 541697
rect 673069 538097 673129 541637
rect 675138 541505 675198 561405
rect 673261 541445 675198 541505
rect 673261 538289 673321 541445
rect 675330 541313 675390 581110
rect 675522 574051 675582 581302
rect 675519 574050 675585 574051
rect 675519 573986 675520 574050
rect 675584 573986 675585 574050
rect 675519 573985 675585 573986
rect 675714 572571 675774 581494
rect 675711 572570 675777 572571
rect 675711 572506 675712 572570
rect 675776 572506 675777 572570
rect 675711 572505 675777 572506
rect 675519 561766 675585 561767
rect 675519 561762 675520 561766
rect 675519 561706 675532 561762
rect 675519 561702 675520 561706
rect 675584 561702 675585 561766
rect 675519 561701 675585 561702
rect 673453 541253 675390 541313
rect 673453 538481 673513 541253
rect 675522 541121 675582 561701
rect 673645 541061 675582 541121
rect 673645 538673 673705 541061
rect 673645 538613 675582 538673
rect 673453 538421 675390 538481
rect 673261 538229 675198 538289
rect 673069 538037 675006 538097
rect 672877 537845 674814 537905
rect 672685 537653 674622 537713
rect 672493 537461 674430 537521
rect 672301 537269 674238 537329
rect 43071 537050 43137 537051
rect 43071 536986 43072 537050
rect 43136 536986 43137 537050
rect 43071 536985 43137 536986
rect 41919 533054 41985 533055
rect 41919 532990 41920 533054
rect 41984 532990 41985 533054
rect 41919 532989 41985 532990
rect 41727 530094 41793 530095
rect 41727 530030 41728 530094
rect 41792 530030 41793 530094
rect 41727 530029 41793 530030
rect 41730 479957 41790 530029
rect 41922 480099 41982 532989
rect 674178 529947 674238 537269
rect 674175 529946 674241 529947
rect 674175 529882 674176 529946
rect 674240 529882 674241 529946
rect 674175 529881 674241 529882
rect 42111 529354 42177 529355
rect 42111 529290 42112 529354
rect 42176 529290 42177 529354
rect 42111 529289 42177 529290
rect 42114 480241 42174 529289
rect 42495 527282 42561 527283
rect 42495 527218 42496 527282
rect 42560 527218 42561 527282
rect 42495 527217 42561 527218
rect 42303 527134 42369 527135
rect 42303 527070 42304 527134
rect 42368 527070 42369 527134
rect 42303 527069 42369 527070
rect 42306 480383 42366 527069
rect 42498 480525 42558 527217
rect 674370 485695 674430 537461
rect 674367 485694 674433 485695
rect 674367 485630 674368 485694
rect 674432 485630 674433 485694
rect 674367 485629 674433 485630
rect 674562 482883 674622 537653
rect 674754 529355 674814 537845
rect 674751 529354 674817 529355
rect 674751 529290 674752 529354
rect 674816 529290 674817 529354
rect 674751 529289 674817 529290
rect 674946 527875 675006 538037
rect 674943 527874 675009 527875
rect 674943 527810 674944 527874
rect 675008 527810 675009 527874
rect 674943 527809 675009 527810
rect 675138 497551 675198 538229
rect 675330 527283 675390 538421
rect 675327 527282 675393 527283
rect 675327 527218 675328 527282
rect 675392 527218 675393 527282
rect 675327 527217 675393 527218
rect 674832 497491 675198 497551
rect 675522 497541 675582 538613
rect 675906 530835 675966 581686
rect 676098 572275 676158 581878
rect 676095 572274 676161 572275
rect 676095 572210 676096 572274
rect 676160 572210 676161 572274
rect 676095 572209 676161 572210
rect 675903 530834 675969 530835
rect 675903 530770 675904 530834
rect 675968 530770 675969 530834
rect 675903 530769 675969 530770
rect 676290 529059 676350 582070
rect 676482 570203 676542 582262
rect 676479 570202 676545 570203
rect 676479 570138 676480 570202
rect 676544 570138 676545 570202
rect 676479 570137 676545 570138
rect 677055 554662 677121 554663
rect 677055 554598 677056 554662
rect 677120 554598 677121 554662
rect 677055 554597 677121 554598
rect 676863 553330 676929 553331
rect 676863 553266 676864 553330
rect 676928 553266 676929 553330
rect 676863 553265 676929 553266
rect 676866 539735 676926 553265
rect 677058 539991 677118 554597
rect 677058 539931 677692 539991
rect 676866 539675 677416 539735
rect 676866 539674 676926 539675
rect 677356 538472 677416 539675
rect 676866 538412 677416 538472
rect 676287 529058 676353 529059
rect 676287 528994 676288 529058
rect 676352 528994 676353 529058
rect 676287 528993 676353 528994
rect 674832 496191 674892 497491
rect 675522 497481 675992 497541
rect 675932 496246 675992 497481
rect 674832 496131 675198 496191
rect 675138 486435 675198 496131
rect 675522 496186 675992 496246
rect 675135 486434 675201 486435
rect 675135 486370 675136 486434
rect 675200 486370 675201 486434
rect 675135 486369 675201 486370
rect 675522 483475 675582 496186
rect 676866 496113 676926 538412
rect 676176 496053 676926 496113
rect 677058 538266 677118 538271
rect 677632 538266 677692 539931
rect 677058 538206 677692 538266
rect 677058 496090 677118 538206
rect 676176 494803 676236 496053
rect 677058 496030 677515 496090
rect 676176 494743 676926 494803
rect 677455 494777 677515 496030
rect 675519 483474 675585 483475
rect 675519 483410 675520 483474
rect 675584 483410 675585 483474
rect 675519 483409 675585 483410
rect 674559 482882 674625 482883
rect 674559 482818 674560 482882
rect 674624 482818 674625 482882
rect 674559 482817 674625 482818
rect 676866 481107 676926 494743
rect 677058 494717 677515 494777
rect 676863 481106 676929 481107
rect 676863 481042 676864 481106
rect 676928 481042 676929 481106
rect 676863 481041 676929 481042
rect 42687 480810 42753 480811
rect 42687 480746 42688 480810
rect 42752 480746 42753 480810
rect 42687 480745 42753 480746
rect 42690 480667 42750 480745
rect 42690 480607 44945 480667
rect 677058 480663 677118 494717
rect 42498 480465 44753 480525
rect 42306 480323 44561 480383
rect 42114 480181 44369 480241
rect 41922 480039 44177 480099
rect 41730 479897 43985 479957
rect 41538 479755 43793 479815
rect 41346 479613 43601 479673
rect 41154 479443 41477 479503
rect 40962 479315 41307 479375
rect 40770 479139 41157 479199
rect 40575 478146 40641 478147
rect 40575 478082 40576 478146
rect 40640 478082 40641 478146
rect 41097 478125 41157 479139
rect 40575 478081 40641 478082
rect 39982 477978 40446 478038
rect 40386 469470 40446 477978
rect 40578 473263 40638 478081
rect 40770 478065 41157 478125
rect 40575 473262 40641 473263
rect 40575 473198 40576 473262
rect 40640 473198 40641 473262
rect 40575 473197 40641 473198
rect 40386 469415 40638 469470
rect 40386 469414 40641 469415
rect 40386 469410 40576 469414
rect 40575 469350 40576 469410
rect 40640 469350 40641 469414
rect 40575 469349 40641 469350
rect 40770 465863 40830 478065
rect 41247 477961 41307 479315
rect 40962 477901 41307 477961
rect 40962 467343 41022 477901
rect 41417 477827 41477 479443
rect 41154 477767 41477 477827
rect 40959 467342 41025 467343
rect 40959 467278 40960 467342
rect 41024 467278 41025 467342
rect 40959 467277 41025 467278
rect 41154 466307 41214 477767
rect 43541 476486 43601 479613
rect 41346 476426 43601 476486
rect 41346 466899 41406 476426
rect 43733 476294 43793 479755
rect 41538 476234 43793 476294
rect 41538 471339 41598 476234
rect 43925 476102 43985 479897
rect 41730 476042 43985 476102
rect 41535 471338 41601 471339
rect 41535 471274 41536 471338
rect 41600 471274 41601 471338
rect 41535 471273 41601 471274
rect 41730 467491 41790 476042
rect 44117 475910 44177 480039
rect 41922 475850 44177 475910
rect 41922 469563 41982 475850
rect 44309 475718 44369 480181
rect 42114 475658 44369 475718
rect 41919 469562 41985 469563
rect 41919 469498 41920 469562
rect 41984 469498 41985 469562
rect 41919 469497 41985 469498
rect 42114 468083 42174 475658
rect 44501 475526 44561 480323
rect 42306 475466 44561 475526
rect 42306 470155 42366 475466
rect 44693 475334 44753 480465
rect 42498 475274 44753 475334
rect 42498 471635 42558 475274
rect 44885 475142 44945 480607
rect 677055 480662 677121 480663
rect 677055 480598 677056 480662
rect 677120 480598 677121 480662
rect 677055 480597 677121 480598
rect 42690 475082 44945 475142
rect 42495 471634 42561 471635
rect 42495 471570 42496 471634
rect 42560 471570 42561 471634
rect 42495 471569 42561 471570
rect 42303 470154 42369 470155
rect 42303 470090 42304 470154
rect 42368 470090 42369 470154
rect 42303 470089 42369 470090
rect 42303 470006 42369 470007
rect 42303 469942 42304 470006
rect 42368 469942 42369 470006
rect 42303 469941 42369 469942
rect 42111 468082 42177 468083
rect 42111 468018 42112 468082
rect 42176 468018 42177 468082
rect 42111 468017 42177 468018
rect 41727 467490 41793 467491
rect 41727 467426 41728 467490
rect 41792 467426 41793 467490
rect 41727 467425 41793 467426
rect 41343 466898 41409 466899
rect 41343 466834 41344 466898
rect 41408 466834 41409 466898
rect 41343 466833 41409 466834
rect 41151 466306 41217 466307
rect 41151 466242 41152 466306
rect 41216 466242 41217 466306
rect 41151 466241 41217 466242
rect 40767 465862 40833 465863
rect 40767 465798 40768 465862
rect 40832 465798 40833 465862
rect 40767 465797 40833 465798
rect 40575 423950 40641 423951
rect 40575 423886 40576 423950
rect 40640 423886 40641 423950
rect 40575 423885 40641 423886
rect 40578 400151 40638 423885
rect 41727 423506 41793 423507
rect 41727 423442 41728 423506
rect 41792 423442 41793 423506
rect 41727 423441 41793 423442
rect 40767 422914 40833 422915
rect 40767 422850 40768 422914
rect 40832 422850 40833 422914
rect 40767 422849 40833 422850
rect 40575 400150 40641 400151
rect 40575 400086 40576 400150
rect 40640 400086 40641 400150
rect 40575 400085 40641 400086
rect 40770 398819 40830 422849
rect 40959 422470 41025 422471
rect 40959 422406 40960 422470
rect 41024 422406 41025 422470
rect 40959 422405 41025 422406
rect 40962 402075 41022 422405
rect 41151 420990 41217 420991
rect 41151 420926 41152 420990
rect 41216 420926 41217 420990
rect 41151 420925 41217 420926
rect 40959 402074 41025 402075
rect 40959 402010 40960 402074
rect 41024 402010 41025 402074
rect 40959 402009 41025 402010
rect 41154 399559 41214 420925
rect 41151 399558 41217 399559
rect 41151 399494 41152 399558
rect 41216 399494 41217 399558
rect 41151 399493 41217 399494
rect 40767 398818 40833 398819
rect 40767 398754 40768 398818
rect 40832 398754 40833 398818
rect 40767 398753 40833 398754
rect 41730 391092 41790 423441
rect 42111 422174 42177 422175
rect 42111 422110 42112 422174
rect 42176 422110 42177 422174
rect 42111 422109 42177 422110
rect 41919 420842 41985 420843
rect 41919 420778 41920 420842
rect 41984 420778 41985 420842
rect 41919 420777 41985 420778
rect 40784 391032 41790 391092
rect 40784 389414 40844 391032
rect 41922 390917 41982 420777
rect 42114 406071 42174 422109
rect 42111 406070 42177 406071
rect 42111 406006 42112 406070
rect 42176 406006 42177 406070
rect 42111 406005 42177 406006
rect 40988 390857 41982 390917
rect 40988 389633 41048 390857
rect 40988 389573 41982 389633
rect 40784 389354 41790 389414
rect 41730 383279 41790 389354
rect 41922 388145 41982 389573
rect 41919 388144 41985 388145
rect 41919 388080 41920 388144
rect 41984 388080 41985 388144
rect 41919 388079 41985 388080
rect 41727 383278 41793 383279
rect 41727 383214 41728 383278
rect 41792 383214 41793 383278
rect 41727 383213 41793 383214
rect 40575 381354 40641 381355
rect 40575 381290 40576 381354
rect 40640 381290 40641 381354
rect 40575 381289 40641 381290
rect 40578 356935 40638 381289
rect 40767 380318 40833 380319
rect 40767 380254 40768 380318
rect 40832 380254 40833 380318
rect 40767 380253 40833 380254
rect 40575 356934 40641 356935
rect 40575 356870 40576 356934
rect 40640 356870 40641 356934
rect 40575 356869 40641 356870
rect 40770 355603 40830 380253
rect 41343 379726 41409 379727
rect 41343 379662 41344 379726
rect 41408 379662 41409 379726
rect 41343 379661 41409 379662
rect 40959 378246 41025 378247
rect 40959 378182 40960 378246
rect 41024 378182 41025 378246
rect 40959 378181 41025 378182
rect 40962 356491 41022 378181
rect 41151 377802 41217 377803
rect 41151 377738 41152 377802
rect 41216 377738 41217 377802
rect 41151 377737 41217 377738
rect 41154 359303 41214 377737
rect 41151 359302 41217 359303
rect 41151 359238 41152 359302
rect 41216 359238 41217 359302
rect 41151 359237 41217 359238
rect 41346 358859 41406 379661
rect 41727 378838 41793 378839
rect 41727 378774 41728 378838
rect 41792 378774 41793 378838
rect 41727 378773 41793 378774
rect 41343 358858 41409 358859
rect 41343 358794 41344 358858
rect 41408 358794 41409 358858
rect 41343 358793 41409 358794
rect 40959 356490 41025 356491
rect 40959 356426 40960 356490
rect 41024 356426 41025 356490
rect 40959 356425 41025 356426
rect 40767 355602 40833 355603
rect 40767 355538 40768 355602
rect 40832 355538 40833 355602
rect 40767 355537 40833 355538
rect 41730 347996 41790 378773
rect 41048 347936 41790 347996
rect 41048 346427 41108 347936
rect 41048 346367 41790 346427
rect 41730 343171 41790 346367
rect 41727 343170 41793 343171
rect 41727 343106 41728 343170
rect 41792 343106 41793 343170
rect 41727 343105 41793 343106
rect 40575 338582 40641 338583
rect 40575 338518 40576 338582
rect 40640 338518 40641 338582
rect 40575 338517 40641 338518
rect 40578 306566 40638 338517
rect 40767 338138 40833 338139
rect 40767 338074 40768 338138
rect 40832 338074 40833 338138
rect 40767 338073 40833 338074
rect 40770 313719 40830 338073
rect 40959 337102 41025 337103
rect 40959 337038 40960 337102
rect 41024 337038 41025 337102
rect 40959 337037 41025 337038
rect 40767 313718 40833 313719
rect 40767 313654 40768 313718
rect 40832 313654 40833 313718
rect 40767 313653 40833 313654
rect 40962 312387 41022 337037
rect 41343 336658 41409 336659
rect 41343 336594 41344 336658
rect 41408 336594 41409 336658
rect 41343 336593 41409 336594
rect 41151 335030 41217 335031
rect 41151 334966 41152 335030
rect 41216 334966 41217 335030
rect 41151 334965 41217 334966
rect 41154 313275 41214 334965
rect 41346 315495 41406 336593
rect 41535 334586 41601 334587
rect 41535 334522 41536 334586
rect 41600 334522 41601 334586
rect 41535 334521 41601 334522
rect 41538 316235 41598 334521
rect 41535 316234 41601 316235
rect 41535 316170 41536 316234
rect 41600 316170 41601 316234
rect 41535 316169 41601 316170
rect 41343 315494 41409 315495
rect 41343 315430 41344 315494
rect 41408 315430 41409 315494
rect 41343 315429 41409 315430
rect 41151 313274 41217 313275
rect 41151 313210 41152 313274
rect 41216 313210 41217 313274
rect 41151 313209 41217 313210
rect 40959 312386 41025 312387
rect 40959 312322 40960 312386
rect 41024 312322 41025 312386
rect 40959 312321 41025 312322
rect 40578 306506 41226 306566
rect 41166 304969 41226 306506
rect 40578 304909 41226 304969
rect 40578 278643 40638 304909
rect 40959 294922 41025 294923
rect 40959 294858 40960 294922
rect 41024 294858 41025 294922
rect 40959 294857 41025 294858
rect 40767 293886 40833 293887
rect 40767 293822 40768 293886
rect 40832 293822 40833 293886
rect 40767 293821 40833 293822
rect 40575 278642 40641 278643
rect 40575 278578 40576 278642
rect 40640 278578 40641 278642
rect 40575 278577 40641 278578
rect 40770 269171 40830 293821
rect 40962 270651 41022 294857
rect 41535 293442 41601 293443
rect 41535 293378 41536 293442
rect 41600 293378 41601 293442
rect 41535 293377 41601 293378
rect 41151 291962 41217 291963
rect 41151 291898 41152 291962
rect 41216 291898 41217 291962
rect 41151 291897 41217 291898
rect 40959 270650 41025 270651
rect 40959 270586 40960 270650
rect 41024 270586 41025 270650
rect 40959 270585 41025 270586
rect 41154 270059 41214 291897
rect 41343 291370 41409 291371
rect 41343 291306 41344 291370
rect 41408 291306 41409 291370
rect 41343 291305 41409 291306
rect 41346 273019 41406 291305
rect 41343 273018 41409 273019
rect 41343 272954 41344 273018
rect 41408 272954 41409 273018
rect 41343 272953 41409 272954
rect 41538 272427 41598 293377
rect 42306 273611 42366 469941
rect 42690 465123 42750 475082
rect 43071 473114 43137 473115
rect 43071 473050 43072 473114
rect 43136 473050 43137 473114
rect 43071 473049 43137 473050
rect 42687 465122 42753 465123
rect 42687 465058 42688 465122
rect 42752 465058 42753 465122
rect 42687 465057 42753 465058
rect 43074 276423 43134 473049
rect 673983 399706 674049 399707
rect 673983 399642 673984 399706
rect 674048 399642 674049 399706
rect 673983 399641 674049 399642
rect 673986 356047 674046 399641
rect 675711 398670 675777 398671
rect 675711 398606 675712 398670
rect 675776 398606 675777 398670
rect 675711 398605 675777 398606
rect 674367 397634 674433 397635
rect 674367 397570 674368 397634
rect 674432 397570 674433 397634
rect 674367 397569 674433 397570
rect 674370 374399 674430 397569
rect 675327 394674 675393 394675
rect 675327 394610 675328 394674
rect 675392 394610 675393 394674
rect 675327 394609 675393 394610
rect 674751 393342 674817 393343
rect 674751 393278 674752 393342
rect 674816 393278 674817 393342
rect 674751 393277 674817 393278
rect 674754 375731 674814 393277
rect 675135 391714 675201 391715
rect 675135 391650 675136 391714
rect 675200 391650 675201 391714
rect 675135 391649 675201 391650
rect 675138 376471 675198 391649
rect 675330 382391 675390 394609
rect 675519 393194 675585 393195
rect 675519 393130 675520 393194
rect 675584 393130 675585 393194
rect 675519 393129 675585 393130
rect 675327 382390 675393 382391
rect 675327 382326 675328 382390
rect 675392 382326 675393 382390
rect 675327 382325 675393 382326
rect 675522 377211 675582 393129
rect 675519 377210 675585 377211
rect 675519 377206 675520 377210
rect 675519 377150 675532 377206
rect 675519 377146 675520 377150
rect 675584 377146 675585 377210
rect 675519 377145 675585 377146
rect 675135 376470 675201 376471
rect 675135 376406 675136 376470
rect 675200 376466 675201 376470
rect 675188 376410 675201 376466
rect 675200 376406 675201 376410
rect 675135 376405 675201 376406
rect 674751 375730 674817 375731
rect 674751 375666 674752 375730
rect 674816 375666 674817 375730
rect 674751 375665 674817 375666
rect 674367 374398 674433 374399
rect 674367 374334 674368 374398
rect 674432 374334 674433 374398
rect 674367 374333 674433 374334
rect 675714 364554 675774 398605
rect 676287 397930 676353 397931
rect 676287 397866 676288 397930
rect 676352 397866 676353 397930
rect 676287 397865 676353 397866
rect 676290 397470 676350 397865
rect 676290 397410 676542 397470
rect 676287 396450 676353 396451
rect 676287 396386 676288 396450
rect 676352 396386 676353 396450
rect 676287 396385 676353 396386
rect 676095 395414 676161 395415
rect 676095 395350 676096 395414
rect 676160 395350 676161 395414
rect 676095 395349 676161 395350
rect 675903 392232 675969 392233
rect 675903 392168 675904 392232
rect 675968 392168 675969 392232
rect 675903 392167 675969 392168
rect 675906 378099 675966 392167
rect 675903 378098 675969 378099
rect 675903 378034 675904 378098
rect 675968 378034 675969 378098
rect 675903 378033 675969 378034
rect 676098 372031 676158 395349
rect 676290 382983 676350 396385
rect 676482 384759 676542 397410
rect 676671 395858 676737 395859
rect 676671 395794 676672 395858
rect 676736 395794 676737 395858
rect 676671 395793 676737 395794
rect 676479 384758 676545 384759
rect 676479 384694 676480 384758
rect 676544 384694 676545 384758
rect 676479 384693 676545 384694
rect 676287 382982 676353 382983
rect 676287 382918 676288 382982
rect 676352 382918 676353 382982
rect 676287 382917 676353 382918
rect 676674 378839 676734 395793
rect 676671 378838 676737 378839
rect 676671 378774 676672 378838
rect 676736 378774 676737 378838
rect 676671 378773 676737 378774
rect 676095 372030 676161 372031
rect 676095 371966 676096 372030
rect 676160 371966 676161 372030
rect 676095 371965 676161 371966
rect 675714 364494 676106 364554
rect 676046 362907 676106 364494
rect 675714 362847 676106 362907
rect 673983 356046 674049 356047
rect 673983 355982 673984 356046
rect 674048 355982 674049 356046
rect 673983 355981 674049 355982
rect 673983 355898 674049 355899
rect 673983 355834 673984 355898
rect 674048 355834 674049 355898
rect 673983 355833 674049 355834
rect 673986 311055 674046 355833
rect 674175 355306 674241 355307
rect 674175 355242 674176 355306
rect 674240 355242 674241 355306
rect 674175 355241 674241 355242
rect 673983 311054 674049 311055
rect 673983 310990 673984 311054
rect 674048 310990 674049 311054
rect 673983 310989 674049 310990
rect 673983 310462 674049 310463
rect 673983 310398 673984 310462
rect 674048 310398 674049 310462
rect 673983 310397 674049 310398
rect 43071 276422 43137 276423
rect 43071 276358 43072 276422
rect 43136 276358 43137 276422
rect 43071 276357 43137 276358
rect 42303 273610 42369 273611
rect 42303 273546 42304 273610
rect 42368 273546 42369 273610
rect 42303 273545 42369 273546
rect 41535 272426 41601 272427
rect 41535 272362 41536 272426
rect 41600 272362 41601 272426
rect 41535 272361 41601 272362
rect 41151 270058 41217 270059
rect 41151 269994 41152 270058
rect 41216 269994 41217 270058
rect 41151 269993 41217 269994
rect 40767 269170 40833 269171
rect 40767 269106 40768 269170
rect 40832 269106 40833 269170
rect 40767 269105 40833 269106
rect 673986 265767 674046 310397
rect 674178 309871 674238 355241
rect 675714 354715 675774 362847
rect 675711 354714 675777 354715
rect 675711 354650 675712 354714
rect 675776 354650 675777 354714
rect 675711 354649 675777 354650
rect 674367 354270 674433 354271
rect 674367 354206 674368 354270
rect 674432 354206 674433 354270
rect 674367 354205 674433 354206
rect 674175 309870 674241 309871
rect 674175 309806 674176 309870
rect 674240 309806 674241 309870
rect 674175 309805 674241 309806
rect 674370 308983 674430 354205
rect 674559 353234 674625 353235
rect 674559 353170 674560 353234
rect 674624 353170 674625 353234
rect 674559 353169 674625 353170
rect 674562 328223 674622 353169
rect 674751 351014 674817 351015
rect 674751 350950 674752 351014
rect 674816 350950 674817 351014
rect 674751 350949 674817 350950
rect 674559 328222 674625 328223
rect 674559 328158 674560 328222
rect 674624 328158 674625 328222
rect 674559 328157 674625 328158
rect 674754 326891 674814 350949
rect 674943 348794 675009 348795
rect 674943 348730 674944 348794
rect 675008 348730 675009 348794
rect 674943 348729 675009 348730
rect 674946 332367 675006 348729
rect 675903 343022 675969 343023
rect 675903 342958 675904 343022
rect 675968 342958 675969 343022
rect 675903 342957 675969 342958
rect 675711 342874 675777 342875
rect 675711 342810 675712 342874
rect 675776 342810 675777 342874
rect 675711 342809 675777 342810
rect 675714 333551 675774 342809
rect 675711 333550 675777 333551
rect 675711 333486 675712 333550
rect 675776 333546 675777 333550
rect 675764 333490 675777 333546
rect 675776 333486 675777 333490
rect 675711 333485 675777 333486
rect 674943 332366 675009 332367
rect 674943 332302 674944 332366
rect 675008 332302 675009 332366
rect 674943 332301 675009 332302
rect 675906 330591 675966 342957
rect 675903 330590 675969 330591
rect 675903 330526 675904 330590
rect 675968 330526 675969 330590
rect 675903 330525 675969 330526
rect 674751 326890 674817 326891
rect 674751 326826 674752 326890
rect 674816 326826 674817 326890
rect 674751 326825 674817 326826
rect 676863 309722 676929 309723
rect 676863 309658 676864 309722
rect 676928 309658 676929 309722
rect 676863 309657 676929 309658
rect 674559 309130 674625 309131
rect 674559 309066 674560 309130
rect 674624 309066 674625 309130
rect 674559 309065 674625 309066
rect 674367 308982 674433 308983
rect 674367 308918 674368 308982
rect 674432 308918 674433 308982
rect 674367 308917 674433 308918
rect 674175 305430 674241 305431
rect 674175 305366 674176 305430
rect 674240 305366 674241 305430
rect 674175 305365 674241 305366
rect 674178 282195 674238 305365
rect 674175 282194 674241 282195
rect 674175 282130 674176 282194
rect 674240 282130 674241 282194
rect 674175 282129 674241 282130
rect 674562 270651 674622 309065
rect 675903 308390 675969 308391
rect 675903 308326 675904 308390
rect 675968 308326 675969 308390
rect 675903 308325 675969 308326
rect 674751 307502 674817 307503
rect 674751 307438 674752 307502
rect 674816 307438 674817 307502
rect 674751 307437 674817 307438
rect 674754 283231 674814 307437
rect 675327 306466 675393 306467
rect 675327 306402 675328 306466
rect 675392 306402 675393 306466
rect 675327 306401 675393 306402
rect 674943 303506 675009 303507
rect 674943 303442 674944 303506
rect 675008 303442 675009 303506
rect 674943 303441 675009 303442
rect 674946 285599 675006 303441
rect 675135 302766 675201 302767
rect 675135 302702 675136 302766
rect 675200 302702 675201 302766
rect 675135 302701 675201 302702
rect 675138 287227 675198 302701
rect 675330 292851 675390 306401
rect 675711 306022 675777 306023
rect 675711 305958 675712 306022
rect 675776 305958 675777 306022
rect 675711 305957 675777 305958
rect 675519 302026 675585 302027
rect 675519 301962 675520 302026
rect 675584 301962 675585 302026
rect 675519 301961 675585 301962
rect 675327 292850 675393 292851
rect 675327 292786 675328 292850
rect 675392 292846 675393 292850
rect 675380 292790 675393 292846
rect 675392 292786 675393 292790
rect 675327 292785 675393 292786
rect 675522 287819 675582 301961
rect 675714 288559 675774 305957
rect 675711 288558 675777 288559
rect 675711 288554 675712 288558
rect 675711 288498 675724 288554
rect 675711 288494 675712 288498
rect 675776 288494 675777 288558
rect 675711 288493 675777 288494
rect 675519 287818 675585 287819
rect 675519 287754 675520 287818
rect 675584 287814 675585 287818
rect 675572 287758 675585 287814
rect 675584 287754 675585 287758
rect 675519 287753 675585 287754
rect 675135 287226 675201 287227
rect 675135 287162 675136 287226
rect 675200 287162 675201 287226
rect 675135 287161 675201 287162
rect 674943 285598 675009 285599
rect 674943 285534 674944 285598
rect 675008 285534 675009 285598
rect 674943 285533 675009 285534
rect 674751 283230 674817 283231
rect 674751 283166 674752 283230
rect 674816 283166 674817 283230
rect 674751 283165 674817 283166
rect 675906 278347 675966 308325
rect 676287 307650 676353 307651
rect 676287 307586 676288 307650
rect 676352 307586 676353 307650
rect 676287 307585 676353 307586
rect 676095 302618 676161 302619
rect 676095 302554 676096 302618
rect 676160 302554 676161 302618
rect 676095 302553 676161 302554
rect 676098 290779 676158 302553
rect 676290 294627 676350 307585
rect 676479 301138 676545 301139
rect 676479 301074 676480 301138
rect 676544 301074 676545 301138
rect 676479 301073 676545 301074
rect 676287 294626 676353 294627
rect 676287 294562 676288 294626
rect 676352 294562 676353 294626
rect 676287 294561 676353 294562
rect 676095 290778 676161 290779
rect 676095 290714 676096 290778
rect 676160 290714 676161 290778
rect 676095 290713 676161 290714
rect 676482 286635 676542 301073
rect 676479 286634 676545 286635
rect 676479 286570 676480 286634
rect 676544 286570 676545 286634
rect 676479 286569 676545 286570
rect 676866 278495 676926 309657
rect 676863 278494 676929 278495
rect 676863 278430 676864 278494
rect 676928 278430 676929 278494
rect 676863 278429 676929 278430
rect 675903 278346 675969 278347
rect 675903 278282 675904 278346
rect 675968 278282 675969 278346
rect 675903 278281 675969 278282
rect 674559 270650 674625 270651
rect 674559 270586 674560 270650
rect 674624 270586 674625 270650
rect 674559 270585 674625 270586
rect 675327 266506 675393 266507
rect 675327 266442 675328 266506
rect 675392 266442 675393 266506
rect 675327 266441 675393 266442
rect 674367 266358 674433 266359
rect 674367 266294 674368 266358
rect 674432 266294 674433 266358
rect 674367 266293 674433 266294
rect 673983 265766 674049 265767
rect 673983 265702 673984 265766
rect 674048 265702 674049 265766
rect 673983 265701 674049 265702
rect 674175 265026 674241 265027
rect 674175 264962 674176 265026
rect 674240 264962 674241 265026
rect 674175 264961 674241 264962
rect 40383 251706 40449 251707
rect 40383 251642 40384 251706
rect 40448 251642 40449 251706
rect 40383 251641 40449 251642
rect 40386 227435 40446 251641
rect 40575 250670 40641 250671
rect 40575 250606 40576 250670
rect 40640 250606 40641 250670
rect 40575 250605 40641 250606
rect 40383 227434 40449 227435
rect 40383 227370 40384 227434
rect 40448 227370 40449 227434
rect 40383 227369 40449 227370
rect 40578 225955 40638 250605
rect 41151 250226 41217 250227
rect 41151 250162 41152 250226
rect 41216 250162 41217 250226
rect 41151 250161 41217 250162
rect 40767 248746 40833 248747
rect 40767 248682 40768 248746
rect 40832 248682 40833 248746
rect 40767 248681 40833 248682
rect 40770 226843 40830 248681
rect 40959 248154 41025 248155
rect 40959 248090 40960 248154
rect 41024 248090 41025 248154
rect 40959 248089 41025 248090
rect 40962 229803 41022 248089
rect 40959 229802 41025 229803
rect 40959 229738 40960 229802
rect 41024 229738 41025 229802
rect 40959 229737 41025 229738
rect 41154 229211 41214 250161
rect 397503 237054 397569 237055
rect 397503 236990 397504 237054
rect 397568 236990 397569 237054
rect 397503 236989 397569 236990
rect 397506 236793 397566 236989
rect 397506 236759 397758 236793
rect 407298 236759 407742 236793
rect 397506 236758 397761 236759
rect 397506 236733 397696 236758
rect 397695 236694 397696 236733
rect 397760 236694 397761 236758
rect 397695 236693 397761 236694
rect 407295 236758 407742 236759
rect 407295 236694 407296 236758
rect 407360 236733 407742 236758
rect 407360 236694 407361 236733
rect 407295 236693 407361 236694
rect 407682 236315 407742 236733
rect 407679 236314 407745 236315
rect 407679 236250 407680 236314
rect 407744 236250 407745 236314
rect 407679 236249 407745 236250
rect 413631 236166 413697 236167
rect 413631 236102 413632 236166
rect 413696 236127 413697 236166
rect 414015 236166 414081 236167
rect 414015 236127 414016 236166
rect 413696 236102 414016 236127
rect 414080 236102 414081 236166
rect 413631 236101 414081 236102
rect 413634 236067 414078 236101
rect 674178 231599 674238 264961
rect 674370 231791 674430 266293
rect 674559 263250 674625 263251
rect 674559 263186 674560 263250
rect 674624 263186 674625 263250
rect 674559 263185 674625 263186
rect 674562 231983 674622 263185
rect 674751 262214 674817 262215
rect 674751 262150 674752 262214
rect 674816 262150 674817 262214
rect 674751 262149 674817 262150
rect 674754 238239 674814 262149
rect 675135 258366 675201 258367
rect 675135 258302 675136 258366
rect 675200 258302 675201 258366
rect 675135 258301 675201 258302
rect 674943 257774 675009 257775
rect 674943 257710 674944 257774
rect 675008 257710 675009 257774
rect 674943 257709 675009 257710
rect 674946 241939 675006 257709
rect 674943 241938 675009 241939
rect 674943 241874 674944 241938
rect 675008 241874 675009 241938
rect 674943 241873 675009 241874
rect 675138 241051 675198 258301
rect 675135 241050 675201 241051
rect 675135 240986 675136 241050
rect 675200 241046 675201 241050
rect 675188 240990 675201 241046
rect 675200 240986 675201 240990
rect 675135 240985 675201 240986
rect 674751 238238 674817 238239
rect 674751 238174 674752 238238
rect 674816 238174 674817 238238
rect 674751 238173 674817 238174
rect 675330 232839 675390 266441
rect 676287 261474 676353 261475
rect 676287 261410 676288 261474
rect 676352 261410 676353 261474
rect 676287 261409 676353 261410
rect 675711 260734 675777 260735
rect 675711 260670 675712 260734
rect 675776 260670 675777 260734
rect 675711 260669 675777 260670
rect 675714 243567 675774 260669
rect 675903 253334 675969 253335
rect 675903 253270 675904 253334
rect 675968 253270 675969 253334
rect 675903 253269 675969 253270
rect 675711 243566 675777 243567
rect 675711 243562 675712 243566
rect 675711 243506 675724 243562
rect 675711 243502 675712 243506
rect 675776 243502 675777 243566
rect 675711 243501 675777 243502
rect 675906 236907 675966 253269
rect 676290 250819 676350 261409
rect 676287 250818 676353 250819
rect 676287 250754 676288 250818
rect 676352 250754 676353 250818
rect 676287 250753 676353 250754
rect 675903 236906 675969 236907
rect 675903 236842 675904 236906
rect 675968 236842 675969 236906
rect 675903 236841 675969 236842
rect 675330 232779 676170 232839
rect 674562 231923 675389 231983
rect 674370 231731 675197 231791
rect 674178 231539 675005 231599
rect 674945 230163 675005 231539
rect 674178 230103 675005 230163
rect 41151 229210 41217 229211
rect 41151 229146 41152 229210
rect 41216 229146 41217 229210
rect 41151 229145 41217 229146
rect 40767 226842 40833 226843
rect 40767 226778 40768 226842
rect 40832 226778 40833 226842
rect 40767 226777 40833 226778
rect 40575 225954 40641 225955
rect 40575 225890 40576 225954
rect 40640 225890 40641 225954
rect 40575 225889 40641 225890
rect 674178 220627 674238 230103
rect 675137 229971 675197 231731
rect 674370 229911 675197 229971
rect 674175 220626 674241 220627
rect 674175 220562 674176 220626
rect 674240 220562 674241 220626
rect 674175 220561 674241 220562
rect 674175 220034 674241 220035
rect 674175 219970 674176 220034
rect 674240 219970 674241 220034
rect 674175 219969 674241 219970
rect 673983 219146 674049 219147
rect 673983 219082 673984 219146
rect 674048 219082 674049 219146
rect 673983 219081 674049 219082
rect 40383 208490 40449 208491
rect 40383 208426 40384 208490
rect 40448 208426 40449 208490
rect 40383 208425 40449 208426
rect 40386 184219 40446 208425
rect 40575 207898 40641 207899
rect 40575 207834 40576 207898
rect 40640 207834 40641 207898
rect 40575 207833 40641 207834
rect 40383 184218 40449 184219
rect 40383 184154 40384 184218
rect 40448 184154 40449 184218
rect 40383 184153 40449 184154
rect 40578 182887 40638 207833
rect 40959 207010 41025 207011
rect 40959 206946 40960 207010
rect 41024 206946 41025 207010
rect 40959 206945 41025 206946
rect 40767 205530 40833 205531
rect 40767 205466 40768 205530
rect 40832 205466 40833 205530
rect 40767 205465 40833 205466
rect 40770 183627 40830 205465
rect 40962 185847 41022 206945
rect 41151 204938 41217 204939
rect 41151 204874 41152 204938
rect 41216 204874 41217 204938
rect 41151 204873 41217 204874
rect 41154 186735 41214 204873
rect 41151 186734 41217 186735
rect 41151 186670 41152 186734
rect 41216 186670 41217 186734
rect 41151 186669 41217 186670
rect 673986 186411 674046 219081
rect 674178 186603 674238 219969
rect 674370 219147 674430 229911
rect 675329 229779 675389 231923
rect 674562 229719 675389 229779
rect 674367 219146 674433 219147
rect 674367 219082 674368 219146
rect 674432 219082 674433 219146
rect 674367 219081 674433 219082
rect 674562 218555 674622 229719
rect 675330 225553 675390 225554
rect 676110 225553 676170 232779
rect 675330 225493 676170 225553
rect 674559 218554 674625 218555
rect 674559 218490 674560 218554
rect 674624 218490 674625 218554
rect 674559 218489 674625 218490
rect 675330 217963 675390 225493
rect 674367 217962 674433 217963
rect 674367 217898 674368 217962
rect 674432 217898 674433 217962
rect 674367 217897 674433 217898
rect 675327 217962 675393 217963
rect 675327 217898 675328 217962
rect 675392 217898 675393 217962
rect 675327 217897 675393 217898
rect 674370 186795 674430 217897
rect 675711 217666 675777 217667
rect 675711 217602 675712 217666
rect 675776 217602 675777 217666
rect 675711 217601 675777 217602
rect 674559 213078 674625 213079
rect 674559 213014 674560 213078
rect 674624 213014 674625 213078
rect 674559 213013 674625 213014
rect 674562 194875 674622 213013
rect 675714 204495 675774 217601
rect 675903 215594 675969 215595
rect 675903 215530 675904 215594
rect 675968 215530 675969 215594
rect 675903 215529 675969 215530
rect 675711 204494 675777 204495
rect 675711 204490 675712 204494
rect 675711 204434 675724 204490
rect 675711 204430 675712 204434
rect 675776 204430 675777 204494
rect 675711 204429 675777 204430
rect 675906 198427 675966 215529
rect 676671 207602 676737 207603
rect 676671 207538 676672 207602
rect 676736 207538 676737 207602
rect 676671 207537 676737 207538
rect 676479 207454 676545 207455
rect 676479 207390 676480 207454
rect 676544 207390 676545 207454
rect 676479 207389 676545 207390
rect 675903 198426 675969 198427
rect 675903 198362 675904 198426
rect 675968 198362 675969 198426
rect 675903 198361 675969 198362
rect 674559 194874 674625 194875
rect 674559 194810 674560 194874
rect 674624 194810 674625 194874
rect 674559 194809 674625 194810
rect 676482 193543 676542 207389
rect 676479 193542 676545 193543
rect 676479 193478 676480 193542
rect 676544 193478 676545 193542
rect 676479 193477 676545 193478
rect 676674 191619 676734 207537
rect 676671 191618 676737 191619
rect 676671 191554 676672 191618
rect 676736 191554 676737 191618
rect 676671 191553 676737 191554
rect 674370 186735 675545 186795
rect 674178 186543 675353 186603
rect 673986 186351 675161 186411
rect 40959 185846 41025 185847
rect 40959 185782 40960 185846
rect 41024 185782 41025 185846
rect 40959 185781 41025 185782
rect 675101 184731 675161 186351
rect 673986 184671 675161 184731
rect 40767 183626 40833 183627
rect 40767 183562 40768 183626
rect 40832 183562 40833 183626
rect 40767 183561 40833 183562
rect 40575 182886 40641 182887
rect 40575 182822 40576 182886
rect 40640 182822 40641 182886
rect 40575 182821 40641 182822
rect 673986 175487 674046 184671
rect 675293 184539 675353 186543
rect 674178 184479 675353 184539
rect 674178 176227 674238 184479
rect 675485 184347 675545 186735
rect 674370 184287 675545 184347
rect 674175 176226 674241 176227
rect 674175 176162 674176 176226
rect 674240 176162 674241 176226
rect 674175 176161 674241 176162
rect 673983 175486 674049 175487
rect 673983 175422 673984 175486
rect 674048 175422 674049 175486
rect 673983 175421 674049 175422
rect 673983 174746 674049 174747
rect 673983 174682 673984 174746
rect 674048 174682 674049 174746
rect 673983 174681 674049 174682
rect 673986 140845 674046 174681
rect 674370 174155 674430 184287
rect 674559 175634 674625 175635
rect 674559 175570 674560 175634
rect 674624 175570 674625 175634
rect 674559 175569 674625 175570
rect 674367 174154 674433 174155
rect 674367 174090 674368 174154
rect 674432 174090 674433 174154
rect 674367 174089 674433 174090
rect 674175 173562 674241 173563
rect 674175 173498 674176 173562
rect 674240 173498 674241 173562
rect 674175 173497 674241 173498
rect 673158 140785 674046 140845
rect 673158 139119 673218 140785
rect 674178 140653 674238 173497
rect 673350 140593 674238 140653
rect 673350 139311 673410 140593
rect 673350 139251 674238 139311
rect 673158 139059 674046 139119
rect 673986 129459 674046 139059
rect 673983 129458 674049 129459
rect 673983 129394 673984 129458
rect 674048 129394 674049 129458
rect 673983 129393 674049 129394
rect 674178 128571 674238 139251
rect 674562 135390 674622 175569
rect 676479 172970 676545 172971
rect 676479 172906 676480 172970
rect 676544 172906 676545 172970
rect 676479 172905 676545 172906
rect 674751 172674 674817 172675
rect 674751 172610 674752 172674
rect 674816 172610 674817 172674
rect 674751 172609 674817 172610
rect 674754 149735 674814 172609
rect 675519 171342 675585 171343
rect 675519 171278 675520 171342
rect 675584 171278 675585 171342
rect 675519 171277 675585 171278
rect 674943 171194 675009 171195
rect 674943 171130 674944 171194
rect 675008 171130 675009 171194
rect 674943 171129 675009 171130
rect 674946 155359 675006 171129
rect 675327 168678 675393 168679
rect 675327 168614 675328 168678
rect 675392 168614 675393 168678
rect 675327 168613 675393 168614
rect 675135 168234 675201 168235
rect 675135 168170 675136 168234
rect 675200 168170 675201 168234
rect 675135 168169 675201 168170
rect 674943 155358 675009 155359
rect 674943 155294 674944 155358
rect 675008 155294 675009 155358
rect 674943 155293 675009 155294
rect 675138 152547 675198 168169
rect 675135 152546 675201 152547
rect 675135 152482 675136 152546
rect 675200 152542 675201 152546
rect 675188 152486 675201 152542
rect 675200 152482 675201 152486
rect 675135 152481 675201 152482
rect 675330 150327 675390 168613
rect 675522 157727 675582 171277
rect 676287 170454 676353 170455
rect 676287 170390 676288 170454
rect 676352 170390 676353 170454
rect 676287 170389 676353 170390
rect 675903 167642 675969 167643
rect 675903 167578 675904 167642
rect 675968 167578 675969 167642
rect 675903 167577 675969 167578
rect 675711 167198 675777 167199
rect 675711 167134 675712 167198
rect 675776 167134 675777 167198
rect 675711 167133 675777 167134
rect 675519 157726 675585 157727
rect 675519 157722 675520 157726
rect 675519 157666 675532 157722
rect 675519 157662 675520 157666
rect 675584 157662 675585 157726
rect 675519 157661 675585 157662
rect 675714 152547 675774 167133
rect 675906 155507 675966 167577
rect 676095 166310 676161 166311
rect 676095 166246 676096 166310
rect 676160 166246 676161 166310
rect 676095 166245 676161 166246
rect 675903 155506 675969 155507
rect 675903 155442 675904 155506
rect 675968 155442 675969 155506
rect 675903 155441 675969 155442
rect 675711 152546 675777 152547
rect 675711 152542 675712 152546
rect 675711 152486 675724 152542
rect 675711 152482 675712 152486
rect 675776 152482 675777 152546
rect 675711 152481 675777 152482
rect 676098 151363 676158 166245
rect 676095 151362 676161 151363
rect 676095 151298 676096 151362
rect 676160 151298 676161 151362
rect 676095 151297 676161 151298
rect 675327 150326 675393 150327
rect 675327 150262 675328 150326
rect 675392 150262 675393 150326
rect 675327 150261 675393 150262
rect 674751 149734 674817 149735
rect 674751 149670 674752 149734
rect 674816 149670 674817 149734
rect 674751 149669 674817 149670
rect 676290 146627 676350 170389
rect 676482 159355 676542 172905
rect 676479 159354 676545 159355
rect 676479 159290 676480 159354
rect 676544 159290 676545 159354
rect 676479 159289 676545 159290
rect 676287 146626 676353 146627
rect 676287 146562 676288 146626
rect 676352 146562 676353 146626
rect 676287 146561 676353 146562
rect 674370 135330 674622 135390
rect 674370 130643 674430 135330
rect 674367 130642 674433 130643
rect 674367 130578 674368 130642
rect 674432 130578 674433 130642
rect 674367 130577 674433 130578
rect 674175 128570 674241 128571
rect 674175 128506 674176 128570
rect 674240 128506 674241 128570
rect 674175 128505 674241 128506
rect 673983 125610 674049 125611
rect 673983 125546 673984 125610
rect 674048 125546 674049 125610
rect 673983 125545 674049 125546
rect 673986 107703 674046 125545
rect 674175 123094 674241 123095
rect 674175 123030 674176 123094
rect 674240 123030 674241 123094
rect 674175 123029 674241 123030
rect 673983 107702 674049 107703
rect 673983 107638 673984 107702
rect 674048 107638 674049 107702
rect 673983 107637 674049 107638
rect 674178 105631 674238 123029
rect 674367 122206 674433 122207
rect 674367 122142 674368 122206
rect 674432 122142 674433 122206
rect 674367 122141 674433 122142
rect 674370 106519 674430 122141
rect 676671 118062 676737 118063
rect 676671 117998 676672 118062
rect 676736 117998 676737 118062
rect 676671 117997 676737 117998
rect 675903 117914 675969 117915
rect 675903 117850 675904 117914
rect 675968 117850 675969 117914
rect 675903 117849 675969 117850
rect 674367 106518 674433 106519
rect 674367 106454 674368 106518
rect 674432 106454 674433 106518
rect 674367 106453 674433 106454
rect 674175 105630 674241 105631
rect 674175 105566 674176 105630
rect 674240 105566 674241 105630
rect 674175 105565 674241 105566
rect 675906 103263 675966 117849
rect 675903 103262 675969 103263
rect 675903 103198 675904 103262
rect 675968 103198 675969 103262
rect 675903 103197 675969 103198
rect 676674 101487 676734 117997
rect 676671 101486 676737 101487
rect 676671 101422 676672 101486
rect 676736 101422 676737 101486
rect 676671 101421 676737 101422
<< metal5 >>
rect 78610 1018624 90778 1030788
rect 130010 1018624 142178 1030788
rect 181410 1018624 193578 1030788
rect 231810 1018624 243978 1030788
rect 284410 1018624 296578 1030788
rect 334810 1018624 346978 1030788
rect 386210 1018624 398378 1030788
rect 475210 1018624 487378 1030788
rect 526610 1018624 538778 1030788
rect 577010 1018624 589178 1030788
rect 628410 1018624 640578 1030788
rect 6811 956610 18975 968778
rect 698624 953022 710788 965190
rect 6167 914054 19619 924934
rect 697980 909666 711432 920546
rect 6811 871210 18975 883378
rect 698512 863640 711002 876180
rect 6811 829010 18975 841178
rect 698624 819822 710788 831990
rect 6598 786620 19088 799160
rect 698512 774440 711002 786980
rect 6598 743420 19088 755960
rect 698512 729440 711002 741980
rect 6598 700220 19088 712760
rect 698512 684440 711002 696980
rect 6598 657020 19088 669560
rect 698512 639240 711002 651780
rect 6598 613820 19088 626360
rect 698512 594240 711002 606780
rect 6598 570620 19088 583160
rect 698512 549040 711002 561580
rect 6598 527420 19088 539960
rect 698624 505222 710788 517390
rect 6811 484410 18975 496578
rect 697980 461866 711432 472746
rect 6167 442854 19619 453734
rect 698624 417022 710788 429190
rect 6598 399820 19088 412360
rect 698512 371840 711002 384380
rect 6598 356620 19088 369160
rect 698512 326640 711002 339180
rect 6598 313420 19088 325960
rect 6598 270220 19088 282760
rect 698512 281640 711002 294180
rect 182164 262913 189643 264077
rect 179295 260388 186774 261552
rect 179546 257823 187025 258987
rect 180260 255444 187739 256608
rect 413512 252916 420991 254080
rect 413752 250339 421231 251503
rect 414135 247866 421614 249030
rect 414519 245406 421998 246570
rect 183287 242831 190766 243995
rect 414666 240372 422145 241536
rect 6598 227020 19088 239560
rect 698512 236640 711002 249180
rect 6598 183820 19088 196360
rect 698512 191440 711002 203980
rect 698512 146440 711002 158980
rect 6811 111610 18975 123778
rect 698512 101240 711002 113780
rect 6167 70054 19619 80934
rect 667805 67044 669486 74622
rect 671570 67513 673251 75091
rect 80222 6811 92390 18975
rect 136713 7143 144149 18309
rect 187640 6598 200180 19088
rect 243266 6167 254146 19619
rect 296240 6598 308780 19088
rect 351040 6598 363580 19088
rect 405840 6598 418380 19088
rect 460640 6598 473180 19088
rect 515440 6598 527980 19088
rect 570422 6811 582590 18975
rect 624222 6811 636390 18975
use gpio_control_block  gpio_control_bidir_1\[0\] ../maglef
timestamp 1624273664
transform -1 0 710203 0 1 118400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1624273664
transform -1 0 710203 0 1 164000
box -1620 -364 34000 13964
use simple_por  por ../maglef
timestamp 1606790297
transform 1 0 654146 0 -1 112882
box 25 11 11344 8291
use sky130_fd_sc_hvl__lsbufhv2lv_1_wrapped  rstb_level
timestamp 1608587411
transform -1 0 145710 0 -1 50488
box 414 -400 3522 3800
use mgmt_core  soc ../maglef
timestamp 1624566096
transform 1 0 190434 0 1 53602
box 0 0 450000 168026
use storage  storage ../maglef
timestamp 1624446576
transform 1 0 52032 0 1 53156
box 1066 70 92000 191480
use user_id_programming  user_id_value ../maglef
timestamp 1607107372
transform 1 0 656624 0 1 80926
box 0 0 7109 7077
use gpio_control_block  gpio_control_in_2\[10\]
timestamp 1624273664
transform 1 0 7631 0 1 286000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1624273664
transform 1 0 7631 0 1 199600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1624273664
transform 1 0 7631 0 1 242800
box -1620 -364 34000 13964
use mgmt_protect  mgmt_buffers ../maglef
timestamp 1624984707
transform 1 0 192180 0 1 240036
box -2762 -2778 222734 26170
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1624273664
transform -1 0 710203 0 1 253600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1624273664
transform -1 0 710203 0 1 208400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1624273664
transform 1 0 7631 0 1 329200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1624273664
transform 1 0 7631 0 1 372400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1624273664
transform -1 0 710203 0 1 344600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1624273664
transform -1 0 710203 0 1 298800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1624273664
transform -1 0 710203 0 1 389000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1624273664
transform -1 0 710203 0 1 477200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1624273664
transform 1 0 7631 0 1 462400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1624273664
transform 1 0 7631 0 1 415000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1624273664
transform 1 0 7631 0 1 674600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1624273664
transform 1 0 7631 0 1 631400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1624273664
transform 1 0 7631 0 1 588224
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[10\]
timestamp 1624273664
transform -1 0 710203 0 1 702000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[6\]
timestamp 1624273664
transform -1 0 710203 0 1 521600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[7\]
timestamp 1624273664
transform -1 0 710203 0 1 564800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[8\]
timestamp 1624273664
transform -1 0 710203 0 1 611800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[9\]
timestamp 1624273664
transform -1 0 710203 0 1 657000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1624273664
transform 1 0 7631 0 1 804200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1624273664
transform 1 0 7631 0 1 761000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1624273664
transform 1 0 7631 0 1 717800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[11\]
timestamp 1624273664
transform -1 0 710203 0 1 880800
box -1620 -364 34000 13964
use chip_io_alt  padframe
timestamp 1625169553
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use user_analog_project_wrapper  mprj
timestamp 1620244087
transform 1 0 65308 0 1 278718
box -800 -800 584800 704800
use caravan_power_routing  caravan_power_routing_0
timestamp 1625173552
transform 1 0 38561 0 1 38708
box -33118 599 673272 959285
<< labels >>
flabel metal5 s 187640 6598 200180 19088 0 FreeSans 16000 0 0 0 clock
port 0 nsew signal input
flabel metal5 s 351040 6598 363580 19088 0 FreeSans 16000 0 0 0 flash_clk
port 1 nsew signal tristate
flabel metal5 s 296240 6598 308780 19088 0 FreeSans 16000 0 0 0 flash_csb
port 2 nsew signal tristate
flabel metal5 s 405840 6598 418380 19088 0 FreeSans 16000 0 0 0 flash_io0
port 3 nsew signal tristate
flabel metal5 s 460640 6598 473180 19088 0 FreeSans 16000 0 0 0 flash_io1
port 4 nsew signal tristate
flabel metal5 s 515440 6598 527980 19088 0 FreeSans 16000 0 0 0 gpio
port 5 nsew signal bidirectional
flabel metal5 s 698512 101240 711002 113780 0 FreeSans 16000 0 0 0 mprj_io[0]
port 6 nsew signal bidirectional
flabel metal5 s 698512 684440 711002 696980 0 FreeSans 16000 0 0 0 mprj_io[10]
port 7 nsew signal bidirectional
flabel metal5 s 698512 729440 711002 741980 0 FreeSans 16000 0 0 0 mprj_io[11]
port 8 nsew signal bidirectional
flabel metal5 s 698512 774440 711002 786980 0 FreeSans 16000 0 0 0 mprj_io[12]
port 9 nsew signal bidirectional
flabel metal5 s 698512 863640 711002 876180 0 FreeSans 16000 0 0 0 mprj_io[13]
port 10 nsew signal bidirectional
flabel metal5 s 628410 1018624 640578 1030788 0 FreeSans 16000 0 0 0 mprj_io[15]
port 12 nsew signal bidirectional
flabel metal5 s 526610 1018624 538778 1030788 0 FreeSans 16000 0 0 0 mprj_io[16]
port 13 nsew signal bidirectional
flabel metal5 s 475210 1018624 487378 1030788 0 FreeSans 16000 0 0 0 mprj_io[17]
port 14 nsew signal bidirectional
flabel metal5 s 698512 146440 711002 158980 0 FreeSans 16000 0 0 0 mprj_io[1]
port 17 nsew signal bidirectional
flabel metal5 s 231810 1018624 243978 1030788 0 FreeSans 16000 0 0 0 mprj_io[20]
port 18 nsew signal bidirectional
flabel metal5 s 181410 1018624 193578 1030788 0 FreeSans 16000 0 0 0 mprj_io[21]
port 19 nsew signal bidirectional
flabel metal5 s 130010 1018624 142178 1030788 0 FreeSans 16000 0 0 0 mprj_io[22]
port 20 nsew signal bidirectional
flabel metal5 s 78610 1018624 90778 1030788 0 FreeSans 16000 0 0 0 mprj_io[23]
port 21 nsew signal bidirectional
flabel metal5 s 6811 956610 18975 968778 0 FreeSans 16000 0 0 0 mprj_io[24]
port 22 nsew signal bidirectional
flabel metal5 s 6598 786620 19088 799160 0 FreeSans 16000 0 0 0 mprj_io[25]
port 23 nsew signal bidirectional
flabel metal5 s 6598 743420 19088 755960 0 FreeSans 16000 0 0 0 mprj_io[26]
port 24 nsew signal bidirectional
flabel metal5 s 6598 700220 19088 712760 0 FreeSans 16000 0 0 0 mprj_io[27]
port 25 nsew signal bidirectional
flabel metal5 s 6598 657020 19088 669560 0 FreeSans 16000 0 0 0 mprj_io[28]
port 26 nsew signal bidirectional
flabel metal5 s 6598 613820 19088 626360 0 FreeSans 16000 0 0 0 mprj_io[29]
port 27 nsew signal bidirectional
flabel metal5 s 698512 191440 711002 203980 0 FreeSans 16000 0 0 0 mprj_io[2]
port 28 nsew signal bidirectional
flabel metal5 s 6598 570620 19088 583160 0 FreeSans 16000 0 0 0 mprj_io[30]
port 29 nsew signal bidirectional
flabel metal5 s 6598 527420 19088 539960 0 FreeSans 16000 0 0 0 mprj_io[31]
port 30 nsew signal bidirectional
flabel metal5 s 6598 399820 19088 412360 0 FreeSans 16000 0 0 0 mprj_io[32]
port 31 nsew signal bidirectional
flabel metal5 s 6598 356620 19088 369160 0 FreeSans 16000 0 0 0 mprj_io[33]
port 32 nsew signal bidirectional
flabel metal5 s 6598 313420 19088 325960 0 FreeSans 16000 0 0 0 mprj_io[34]
port 33 nsew signal bidirectional
flabel metal5 s 6598 270220 19088 282760 0 FreeSans 16000 0 0 0 mprj_io[35]
port 34 nsew signal bidirectional
flabel metal5 s 6598 227020 19088 239560 0 FreeSans 16000 0 0 0 mprj_io[36]
port 35 nsew signal bidirectional
flabel metal5 s 6598 183820 19088 196360 0 FreeSans 16000 0 0 0 mprj_io[37]
port 36 nsew signal bidirectional
flabel metal5 s 698512 236640 711002 249180 0 FreeSans 16000 0 0 0 mprj_io[3]
port 37 nsew signal bidirectional
flabel metal5 s 698512 281640 711002 294180 0 FreeSans 16000 0 0 0 mprj_io[4]
port 38 nsew signal bidirectional
flabel metal5 s 698512 326640 711002 339180 0 FreeSans 16000 0 0 0 mprj_io[5]
port 39 nsew signal bidirectional
flabel metal5 s 698512 371840 711002 384380 0 FreeSans 16000 0 0 0 mprj_io[6]
port 40 nsew signal bidirectional
flabel metal5 s 698512 549040 711002 561580 0 FreeSans 16000 0 0 0 mprj_io[7]
port 41 nsew signal bidirectional
flabel metal5 s 698512 594240 711002 606780 0 FreeSans 16000 0 0 0 mprj_io[8]
port 42 nsew signal bidirectional
flabel metal5 s 698512 639240 711002 651780 0 FreeSans 16000 0 0 0 mprj_io[9]
port 43 nsew signal bidirectional
flabel metal5 s 136713 7143 144149 18309 0 FreeSans 16000 0 0 0 resetb
port 44 nsew signal input
flabel metal5 s 697980 909666 711432 920546 0 FreeSans 16000 0 0 0 vccd1
port 45 nsew signal bidirectional
flabel metal5 s 6167 914054 19619 924934 0 FreeSans 16000 0 0 0 vccd2
port 46 nsew signal bidirectional
flabel metal5 s 624222 6811 636390 18975 0 FreeSans 16000 0 0 0 vdda
port 47 nsew signal bidirectional
flabel metal5 s 698624 819822 710788 831990 0 FreeSans 16000 0 0 0 vdda1
port 48 nsew signal bidirectional
flabel metal5 s 698624 505222 710788 517390 0 FreeSans 16000 0 0 0 vdda1_2
port 49 nsew signal bidirectional
flabel metal5 s 6811 484410 18975 496578 0 FreeSans 16000 0 0 0 vdda2
port 50 nsew signal bidirectional
flabel metal5 s 6811 871210 18975 883378 0 FreeSans 16000 0 0 0 vddio_2
port 51 nsew signal bidirectional
flabel metal5 s 577010 1018624 589178 1030788 0 FreeSans 16000 0 0 0 vssa1
port 52 nsew signal bidirectional
flabel metal5 s 698624 417022 710788 429190 0 FreeSans 16000 0 0 0 vssa1_2
port 53 nsew signal bidirectional
flabel metal5 s 6811 829010 18975 841178 0 FreeSans 16000 0 0 0 vssa2
port 54 nsew signal bidirectional
flabel metal5 s 697980 461866 711432 472746 0 FreeSans 16000 0 0 0 vssd1
port 55 nsew signal bidirectional
flabel metal5 s 6167 442854 19619 453734 0 FreeSans 16000 0 0 0 vssd2
port 56 nsew signal bidirectional
flabel metal5 s 334810 1018624 346978 1030788 0 FreeSans 16000 0 0 0 vssio_2
port 57 nsew signal bidirectional
flabel metal5 s 6811 111610 18975 123778 0 FreeSans 16000 0 0 0 vddio
port 58 nsew signal bidirectional
flabel metal5 s 570422 6811 582590 18975 0 FreeSans 16000 0 0 0 vssio
port 59 nsew signal bidirectional
flabel metal5 s 80222 6811 92390 18975 0 FreeSans 16000 0 0 0 vssa
port 60 nsew signal bidirectional
flabel metal5 s 6167 70054 19619 80934 0 FreeSans 16000 0 0 0 vccd
port 61 nsew signal bidirectional
flabel metal5 s 243266 6167 254146 19619 0 FreeSans 16000 0 0 0 vssd
port 62 nsew signal bidirectional
flabel metal2 s 579796 53602 579852 54402 0 FreeSans 16000 0 0 0 pwr_ctrl_out[0]
port 63 nsew signal tristate
flabel metal2 s 597092 53602 597148 54402 0 FreeSans 16000 0 0 0 pwr_ctrl_out[1]
port 64 nsew signal tristate
flabel metal2 s 614388 53602 614444 54402 0 FreeSans 16000 0 0 0 pwr_ctrl_out[2]
port 65 nsew signal tristate
flabel metal2 s 631684 53602 631740 54402 0 FreeSans 16000 0 0 0 pwr_ctrl_out[3]
port 66 nsew signal tristate
flabel metal5 417118 253512 417118 253512 0 FreeSans 8000 0 0 0 vccd1_core
flabel metal5 417486 250996 417486 250996 0 FreeSans 8000 0 0 0 vssd1_core
flabel metal5 417793 248603 417793 248603 0 FreeSans 8000 0 0 0 vdda1_core
flabel metal5 418100 245964 418100 245964 0 FreeSans 8000 0 0 0 vssa1_core
flabel metal5 417916 240932 417916 240932 0 FreeSans 8000 0 0 0 vssd_core
flabel metal5 186454 243448 186454 243448 0 FreeSans 8000 0 0 0 vccd_core
flabel metal5 183999 256028 183999 256028 0 FreeSans 8000 0 0 0 vssa2_core
flabel metal5 183201 258482 183201 258482 0 FreeSans 8000 0 0 0 vdda2_core
flabel metal5 182956 261182 182956 261182 0 FreeSans 8000 0 0 0 vssd2_core
flabel metal5 184920 263575 184920 263575 0 FreeSans 8000 0 0 0 vccd2_core
flabel metal5 668612 70870 668612 70870 0 FreeSans 8000 90 0 0 vddio_core
flabel metal5 672443 71154 672443 71154 0 FreeSans 8000 90 0 0 vssio_core
flabel metal5 s 698624 953022 710788 965190 0 FreeSans 16000 0 0 0 mprj_io[14]
port 15 nsew signal bidirectional
flabel metal5 s 284410 1018624 296578 1030788 0 FreeSans 16000 0 0 0 mprj_io[19]
port 16 nsew signal bidirectional
flabel metal5 s 386210 1018624 398378 1030788 0 FreeSans 16000 0 0 0 mprj_io[18]
port 11 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
