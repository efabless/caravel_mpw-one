.SUBCKT sky130_fd_io__gnd2gnd_sub_dnwl 1 2
**
X0 1 2 sky130_fd_pr__model__parasitic__diode_ps2nw a=283.052 p=67.56 m=1
.ENDS
