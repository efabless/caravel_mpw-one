* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param
+ sky130_fd_pr__nfet_g5v0d16v0__mm_mult = 0.8
.param sky130_fd_pr__nfet_g5v0d16v0__toxe_slope_spectre = 0.0
.param sky130_fd_pr__nfet_g5v0d16v0__wint_slope_spectre = 0.0
.param sky130_fd_pr__nfet_g5v0d16v0__lint_slope_spectre = 0.0
.param sky130_fd_pr__nfet_g5v0d16v0__vth0_slope_spectre = 0.0
.param sky130_fd_pr__nfet_g5v0d16v0__voff_slope_spectre = 0.0
.param sky130_fd_pr__nfet_g5v0d16v0__nfactor_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__nfet_g5v0d16v0__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_g5v0d16v0__wint_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_g5v0d16v0__lint_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_g5v0d16v0__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_g5v0d16v0__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_g5v0d16v0__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__nfet_g5v0d16v0__base d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1 delvto = 0.0
msky130_fd_pr__nfet_g5v0d16v0__base d g s b sky130_fd_pr__nfet_g5v0d16v0__model_base l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} 
.model sky130_fd_pr__nfet_g5v0d16v0__model_base.0 nmos
* Model Flag Parameters
+ lmin = 6.95e-007 lmax = 7.05e-007 wmin = 1.9995e-005 wmax = 2.00005e-5
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 1.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d16v0__toxe_mult}
+ toxm = 1.16e-8
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d16v0__wint_diff}
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d16v0__lint_diff}
+ vth0 = {0.77216+sky130_fd_pr__nfet_g5v0d16v0__vth0_diff_0}
+ k1 = 0.82559
+ k2 = {-0.047197+1.7195e-02+sky130_fd_pr__nfet_g5v0d16v0__k2_diff_0}
+ k3 = -0.884
+ k3b = 0.43
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ dsub = {0.504+sky130_fd_pr__nfet_g5v0d16v0__dsub_diff_0}
+ minv = 0.0
+ voffl = -4.257949e-7
+ lpe0 = 0.0
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -0.0008
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d16v0__voff_diff_0}
+ nfactor = {0.83837+sky130_fd_pr__nfet_g5v0d16v0__nfactor_diff_0}
+ eta0 = {0.016128+sky130_fd_pr__nfet_g5v0d16v0__eta0_diff_0}
+ etab = -0.02983
+ u0 = {0.041428+sky130_fd_pr__nfet_g5v0d16v0__u0_diff_0}
+ ua = {2.3635e-009+sky130_fd_pr__nfet_g5v0d16v0__ua_diff_0}
+ ub = {1.1377e-018+sky130_fd_pr__nfet_g5v0d16v0__ub_diff_0}
+ uc = 2.241e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {73440+sky130_fd_pr__nfet_g5v0d16v0__vsat_diff_0}
+ a0 = {0.73473+sky130_fd_pr__nfet_g5v0d16v0__a0_diff_0}
+ ags = {1.0424+sky130_fd_pr__nfet_g5v0d16v0__ags_diff_0}
+ a1 = 0.0
+ a2 = 0.6597262
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d16v0__b0_diff_0}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d16v0__b1_diff_0}
+ keta = {-0.19104+sky130_fd_pr__nfet_g5v0d16v0__keta_diff_0}
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
+ pclm = 0.82741
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36652
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.005
+ fprout = 10.125
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 724.62
+ rsw = 0.0
+ rdw = 1.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0279e-5
+ alpha1 = 1.1218
+ beta0 = 75.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {0.00e-011+sky130_fd_pr__nfet_g5v0d16v0__agidl_diff_0}
+ bgidl = {1.058e+009+sky130_fd_pr__nfet_g5v0d16v0__bgidl_diff_0}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d16v0__cgidl_diff_0}
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 1.16e-8
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
* Charge AND Capacitance Model Parameters
+ dlc = {-3.5995e-008+sky130_fd_pr__nfet_g5v0d16v0__dlc_diff}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d16v0__dwc_diff}
+ xpart = 0.0
+ cgso = {1.5674e-010*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ cgbo = 0.0
+ cgdl = {4.49025e-011*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ cgsl = {4.49025e-011*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = {0*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.2104
* High-Speed/RF Model Parameters
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.89
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ lintnoi = 0.0
+ tnoia = 7.5e+6
+ tnoib = 7.2e+6
+ rnoia = 0.794
+ rnoib = 0.38
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.000375
+ jsws = 5.84e-11
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.636
+ xjbvs = 1.0
+ pbs = 0.72468
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d16v0__ajunction_mult}
+ mjs = 0.295
+ pbsws = 0.29067
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d16v0__pjunction_mult}
+ mjsws = 0.037586
+ pbswgs = 0.54958
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d16v0__pjunction_mult}
+ mjswgs = 0.78692
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.37073+sky130_fd_pr__nfet_g5v0d16v0__kt1_diff_0}
+ kt2 = {-0.019151+sky130_fd_pr__nfet_g5v0d16v0__kt2_diff_0}
+ at = 29000.0
+ ute = {-1.2471+sky130_fd_pr__nfet_g5v0d16v0__ute_diff_0}
+ ua1 = 2.0117e-9
+ ub1 = -2.2981e-18
+ uc1 = -5.5992e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d16v0__tvoff_diff_0}
+ njs = 1.0773
+ tpb = 0.001344
+ tcj = 0.00067434
+ tpbsw = 0.00099005
+ tcjsw = 0.0002493
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 0.76
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = .28e-6
+ sbref = 1.585e-6
+ kvth0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__kvth0_diff}
+ lkvth0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__lkvth0_diff}
+ wkvth0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 1.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__ku0_diff}
+ lku0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__lku0_diff}
+ wku0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__wku0_diff}
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 1.0
+ wlodku0 = 1.0
+ kvsat = {0.0+sky130_fd_pr__nfet_g5v0d16v0__kvsat_diff}
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_g5v0d16v0__model_base.1 nmos
* Model Flag Parameters
+ lmin = 6.95e-007 lmax = 7.05e-007 wmin = 4.995e-006 wmax = 5.0005e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 1.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d16v0__toxe_mult}
+ toxm = 1.16e-8
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d16v0__wint_diff}
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d16v0__lint_diff}
+ vth0 = {0.78433+sky130_fd_pr__nfet_g5v0d16v0__vth0_diff_1}
+ k1 = 0.89738
+ k2 = {-0.047197+sky130_fd_pr__nfet_g5v0d16v0__k2_diff_1}
+ k3 = -0.884
+ k3b = 0.43
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ dsub = {0.504+sky130_fd_pr__nfet_g5v0d16v0__dsub_diff_1}
+ minv = 0.0
+ voffl = -4.257949e-7
+ lpe0 = 0.0
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -0.0008
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d16v0__voff_diff_1}
+ nfactor = {0.83837+sky130_fd_pr__nfet_g5v0d16v0__nfactor_diff_1}
+ eta0 = {0.016128+sky130_fd_pr__nfet_g5v0d16v0__eta0_diff_1}
+ etab = -0.02983
+ u0 = {0.034999+sky130_fd_pr__nfet_g5v0d16v0__u0_diff_1}
+ ua = {6.84e-010+sky130_fd_pr__nfet_g5v0d16v0__ua_diff_1}
+ ub = {1.5447e-018+sky130_fd_pr__nfet_g5v0d16v0__ub_diff_1}
+ uc = -1.5747e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {73440+sky130_fd_pr__nfet_g5v0d16v0__vsat_diff_1}
+ a0 = {0.73473+sky130_fd_pr__nfet_g5v0d16v0__a0_diff_1}
+ ags = {1.0424+sky130_fd_pr__nfet_g5v0d16v0__ags_diff_1}
+ a1 = 0.0
+ a2 = 0.6597262
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d16v0__b0_diff_1}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d16v0__b1_diff_1}
+ keta = {-0.19104+sky130_fd_pr__nfet_g5v0d16v0__keta_diff_1}
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
+ pclm = 0.82741
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36652
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.005
+ fprout = 10.125
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 724.62
+ rsw = 0.0
+ rdw = 1.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0279e-5
+ alpha1 = 1.1218
+ beta0 = 75.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {0.00e-011+sky130_fd_pr__nfet_g5v0d16v0__agidl_diff_1}
+ bgidl = {1.058e+009+sky130_fd_pr__nfet_g5v0d16v0__bgidl_diff_1}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d16v0__cgidl_diff_1}
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 1.16e-8
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
* Charge AND Capacitance Model Parameters
+ dlc = {-3.5995e-008+sky130_fd_pr__nfet_g5v0d16v0__dlc_diff}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d16v0__dwc_diff}
+ xpart = 0.0
+ cgso = {1.5674e-010*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ cgbo = 0.0
+ cgdl = {4.49025e-011*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ cgsl = {4.49025e-011*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = {0*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.2104
* High-Speed/RF Model Parameters
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.89
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ lintnoi = 0.0
+ tnoia = 7.5e+6
+ tnoib = 7.2e+6
+ rnoia = 0.794
+ rnoib = 0.38
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.000375
+ jsws = 5.84e-11
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.636
+ xjbvs = 1.0
+ pbs = 0.72468
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d16v0__ajunction_mult}
+ mjs = 0.295
+ pbsws = 0.29067
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d16v0__pjunction_mult}
+ mjsws = 0.037586
+ pbswgs = 0.54958
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d16v0__pjunction_mult}
+ mjswgs = 0.78692
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.37073+sky130_fd_pr__nfet_g5v0d16v0__kt1_diff_1}
+ kt2 = {-0.019151+sky130_fd_pr__nfet_g5v0d16v0__kt2_diff_1}
+ at = 29000.0
+ ute = {-1.2471+sky130_fd_pr__nfet_g5v0d16v0__ute_diff_1}
+ ua1 = 2.0117e-9
+ ub1 = -2.2981e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d16v0__tvoff_diff_1}
+ njs = 1.0773
+ tpb = 0.001344
+ tcj = 0.00067434
+ tpbsw = 0.00099005
+ tcjsw = 0.0002493
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 0.76
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = .28e-6
+ sbref = 1.585e-6
+ kvth0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__kvth0_diff}
+ lkvth0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__lkvth0_diff}
+ wkvth0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 1.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__ku0_diff}
+ lku0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__lku0_diff}
+ wku0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__wku0_diff}
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 1.0
+ wlodku0 = 1.0
+ kvsat = {0.0+sky130_fd_pr__nfet_g5v0d16v0__kvsat_diff}
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_g5v0d16v0__model_base.2 nmos
* Model Flag Parameters
+ lmin = 6.95e-007 lmax = 7.05e-007 wmin = 4.995e-005 wmax = 6.0005e-5
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 1.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d16v0__toxe_mult}
+ toxm = 1.16e-8
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d16v0__wint_diff}
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d16v0__lint_diff}
+ vth0 = {0.77216+sky130_fd_pr__nfet_g5v0d16v0__vth0_diff_2}
+ k1 = 0.82559
+ k2 = {-0.047197+1.6900e-02+sky130_fd_pr__nfet_g5v0d16v0__k2_diff_2}
+ k3 = -0.884
+ k3b = 0.43
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ dsub = {0.504+sky130_fd_pr__nfet_g5v0d16v0__dsub_diff_2}
+ minv = 0.0
+ voffl = -4.257949e-7
+ lpe0 = 0.0
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -0.0008
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d16v0__voff_diff_2}
+ nfactor = {0.83837+sky130_fd_pr__nfet_g5v0d16v0__nfactor_diff_2}
+ eta0 = {0.016128+sky130_fd_pr__nfet_g5v0d16v0__eta0_diff_2}
+ etab = -0.02983
+ u0 = {0.041428+sky130_fd_pr__nfet_g5v0d16v0__u0_diff_2}
+ ua = {2.9307e-009+sky130_fd_pr__nfet_g5v0d16v0__ua_diff_2}
+ ub = {7.5689e-019+sky130_fd_pr__nfet_g5v0d16v0__ub_diff_2}
+ uc = 3.33389e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {73440+sky130_fd_pr__nfet_g5v0d16v0__vsat_diff_2}
+ a0 = {0.73473+sky130_fd_pr__nfet_g5v0d16v0__a0_diff_2}
+ ags = {1.0424+sky130_fd_pr__nfet_g5v0d16v0__ags_diff_2}
+ a1 = 0.0
+ a2 = 0.6597262
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d16v0__b0_diff_2}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d16v0__b1_diff_2}
+ keta = {-0.19104+sky130_fd_pr__nfet_g5v0d16v0__keta_diff_2}
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
+ pclm = 0.82741
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36652
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.005
+ fprout = 10.125
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 724.62
+ rsw = 0.0
+ rdw = 1.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0279e-5
+ alpha1 = 1.1218
+ beta0 = 75.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {0.00e-011+sky130_fd_pr__nfet_g5v0d16v0__agidl_diff_2}
+ bgidl = {1.058e+009+sky130_fd_pr__nfet_g5v0d16v0__bgidl_diff_2}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d16v0__cgidl_diff_2}
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 1.16e-8
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
* Charge AND Capacitance Model Parameters
+ dlc = {-3.5995e-008+sky130_fd_pr__nfet_g5v0d16v0__dlc_diff}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d16v0__dwc_diff}
+ xpart = 0.0
+ cgso = {1.5674e-010*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ cgbo = 0.0
+ cgdl = {4.49025e-011*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ cgsl = {4.49025e-011*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = {0*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.2104
* High-Speed/RF Model Parameters
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.89
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ lintnoi = 0.0
+ tnoia = 7.5e+6
+ tnoib = 7.2e+6
+ rnoia = 0.794
+ rnoib = 0.38
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.000375
+ jsws = 5.84e-11
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.636
+ xjbvs = 1.0
+ pbs = 0.72468
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d16v0__ajunction_mult}
+ mjs = 0.295
+ pbsws = 0.29067
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d16v0__pjunction_mult}
+ mjsws = 0.037586
+ pbswgs = 0.54958
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d16v0__pjunction_mult}
+ mjswgs = 0.78692
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.37073+sky130_fd_pr__nfet_g5v0d16v0__kt1_diff_2}
+ kt2 = {-0.062945+sky130_fd_pr__nfet_g5v0d16v0__kt2_diff_2}
+ at = 29000.0
+ ute = {-1.4726+sky130_fd_pr__nfet_g5v0d16v0__ute_diff_2}
+ ua1 = 2.0117e-9
+ ub1 = -2.2981e-18
+ uc1 = -2.2901e-12
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d16v0__tvoff_diff_2}
+ njs = 1.0773
+ tpb = 0.001344
+ tcj = 0.00067434
+ tpbsw = 0.00099005
+ tcjsw = 0.0002493
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 0.76
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = .28e-6
+ sbref = 1.585e-6
+ kvth0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__kvth0_diff}
+ lkvth0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__lkvth0_diff}
+ wkvth0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 1.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__ku0_diff}
+ lku0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__lku0_diff}
+ wku0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__wku0_diff}
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 1.0
+ wlodku0 = 1.0
+ kvsat = {0.0+sky130_fd_pr__nfet_g5v0d16v0__kvsat_diff}
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_g5v0d16v0__model_base.3 nmos
* Model Flag Parameters
+ lmin = 2.195e-006 lmax = 2.25e-006 wmin = 1.9995e-005 wmax = 2.0005e-5
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 1.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d16v0__toxe_mult}
+ toxm = 1.16e-8
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d16v0__wint_diff}
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d16v0__lint_diff}
+ vth0 = {0.78433+sky130_fd_pr__nfet_g5v0d16v0__vth0_diff_3}
+ k1 = 0.89738
+ k2 = {-0.044197+sky130_fd_pr__nfet_g5v0d16v0__k2_diff_3}
+ k3 = -0.884
+ k3b = 0.43
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ dsub = {0.504+sky130_fd_pr__nfet_g5v0d16v0__dsub_diff_3}
+ minv = 0.0
+ voffl = -4.257949e-7
+ lpe0 = 0.0
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -0.0008
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d16v0__voff_diff_3}
+ nfactor = {0.83837+sky130_fd_pr__nfet_g5v0d16v0__nfactor_diff_3}
+ eta0 = {0.016128+sky130_fd_pr__nfet_g5v0d16v0__eta0_diff_3}
+ etab = -0.02983
+ u0 = {0.036814+sky130_fd_pr__nfet_g5v0d16v0__u0_diff_3}
+ ua = {8e-011+sky130_fd_pr__nfet_g5v0d16v0__ua_diff_3}
+ ub = {2.1405e-018+sky130_fd_pr__nfet_g5v0d16v0__ub_diff_3}
+ uc = 6.0747e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {100550+sky130_fd_pr__nfet_g5v0d16v0__vsat_diff_3}
+ a0 = {0.3+sky130_fd_pr__nfet_g5v0d16v0__a0_diff_3}
+ ags = {0.13326+sky130_fd_pr__nfet_g5v0d16v0__ags_diff_3}
+ a1 = 0.0
+ a2 = 0.6597262
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d16v0__b0_diff_3}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d16v0__b1_diff_3}
+ keta = {-0.05+sky130_fd_pr__nfet_g5v0d16v0__keta_diff_3}
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
+ pclm = 0.16548
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36652
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.001
+ fprout = 10.125
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 724.62
+ rsw = 0.0
+ rdw = 1.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0448e-7
+ alpha1 = 0.72
+ beta0 = 37.72
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {0.00e-011+sky130_fd_pr__nfet_g5v0d16v0__agidl_diff_3}
+ bgidl = {1.058e+009+sky130_fd_pr__nfet_g5v0d16v0__bgidl_diff_3}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d16v0__cgidl_diff_3}
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 1.16e-8
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
* Charge AND Capacitance Model Parameters
+ dlc = {-3.5995e-008+sky130_fd_pr__nfet_g5v0d16v0__dlc_diff}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d16v0__dwc_diff}
+ xpart = 0.0
+ cgso = {1.5674e-010*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ cgbo = 0.0
+ cgdl = {4.49025e-011*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ cgsl = {4.49025e-011*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = {0*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.2104
* High-Speed/RF Model Parameters
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.89
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ lintnoi = 0.0
+ tnoia = 7.5e+6
+ tnoib = 7.2e+6
+ rnoia = 0.794
+ rnoib = 0.38
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.000375
+ jsws = 5.84e-11
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.636
+ xjbvs = 1.0
+ pbs = 0.72468
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d16v0__ajunction_mult}
+ mjs = 0.295
+ pbsws = 0.29067
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d16v0__pjunction_mult}
+ mjsws = 0.037586
+ pbswgs = 0.54958
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d16v0__pjunction_mult}
+ mjswgs = 0.78692
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.37073+sky130_fd_pr__nfet_g5v0d16v0__kt1_diff_3}
+ kt2 = {-0.019151+sky130_fd_pr__nfet_g5v0d16v0__kt2_diff_3}
+ at = 29000.0
+ ute = {-1.4324+sky130_fd_pr__nfet_g5v0d16v0__ute_diff_3}
+ ua1 = 2.0117e-9
+ ub1 = -2.9862e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d16v0__tvoff_diff_3}
+ njs = 1.0773
+ tpb = 0.001344
+ tcj = 0.00067434
+ tpbsw = 0.00099005
+ tcjsw = 0.0002493
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 0.76
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = .28e-6
+ sbref = 1.585e-6
+ kvth0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__kvth0_diff}
+ lkvth0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__lkvth0_diff}
+ wkvth0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 1.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__ku0_diff}
+ lku0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__lku0_diff}
+ wku0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__wku0_diff}
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 1.0
+ wlodku0 = 1.0
+ kvsat = {0.0+sky130_fd_pr__nfet_g5v0d16v0__kvsat_diff}
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_g5v0d16v0__model_base.4 nmos
* Model Flag Parameters
+ lmin = 2.195e-006 lmax = 2.25e-006 wmin = 4.995e-006 wmax = 5.005e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 1.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d16v0__toxe_mult}
+ toxm = 1.16e-8
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d16v0__wint_diff}
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d16v0__lint_diff}
+ vth0 = {0.78433+sky130_fd_pr__nfet_g5v0d16v0__vth0_diff_4}
+ k1 = 0.89738
+ k2 = {-0.044197+sky130_fd_pr__nfet_g5v0d16v0__k2_diff_4}
+ k3 = -0.884
+ k3b = 0.43
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ dsub = {0.504+sky130_fd_pr__nfet_g5v0d16v0__dsub_diff_4}
+ minv = 0.0
+ voffl = -4.257949e-7
+ lpe0 = 0.0
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -0.0008
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d16v0__voff_diff_4}
+ nfactor = {0.83837+sky130_fd_pr__nfet_g5v0d16v0__nfactor_diff_4}
+ eta0 = {0.016128+sky130_fd_pr__nfet_g5v0d16v0__eta0_diff_4}
+ etab = -0.02983
+ u0 = {0.036814+sky130_fd_pr__nfet_g5v0d16v0__u0_diff_4}
+ ua = {8e-011+sky130_fd_pr__nfet_g5v0d16v0__ua_diff_4}
+ ub = {1.7638e-018+sky130_fd_pr__nfet_g5v0d16v0__ub_diff_4}
+ uc = 2.6729e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {100550+sky130_fd_pr__nfet_g5v0d16v0__vsat_diff_4}
+ a0 = {0.3+sky130_fd_pr__nfet_g5v0d16v0__a0_diff_4}
+ ags = {0.13326+sky130_fd_pr__nfet_g5v0d16v0__ags_diff_4}
+ a1 = 0.0
+ a2 = 0.6597262
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d16v0__b0_diff_4}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d16v0__b1_diff_4}
+ keta = {-0.05+sky130_fd_pr__nfet_g5v0d16v0__keta_diff_4}
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
+ pclm = 0.16548
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36652
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.001
+ fprout = 10.125
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 724.62
+ rsw = 0.0
+ rdw = 1.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0448e-7
+ alpha1 = 0.72
+ beta0 = 37.72
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {0.00e-011+sky130_fd_pr__nfet_g5v0d16v0__agidl_diff_4}
+ bgidl = {1.058e+009+sky130_fd_pr__nfet_g5v0d16v0__bgidl_diff_4}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d16v0__cgidl_diff_4}
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 1.16e-8
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
* Charge AND Capacitance Model Parameters
+ dlc = {-3.5995e-008+sky130_fd_pr__nfet_g5v0d16v0__dlc_diff}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d16v0__dwc_diff}
+ xpart = 0.0
+ cgso = {1.5674e-010*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ cgbo = 0.0
+ cgdl = {4.49025e-011*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ cgsl = {4.49025e-011*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = {0*sky130_fd_pr__nfet_g5v0d16v0__overlap_mult}
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.2104
* High-Speed/RF Model Parameters
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.89
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ lintnoi = 0.0
+ tnoia = 7.5e+6
+ tnoib = 7.2e+6
+ rnoia = 0.794
+ rnoib = 0.38
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.000375
+ jsws = 5.84e-11
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.636
+ xjbvs = 1.0
+ pbs = 0.72468
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d16v0__ajunction_mult}
+ mjs = 0.295
+ pbsws = 0.29067
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d16v0__pjunction_mult}
+ mjsws = 0.037586
+ pbswgs = 0.54958
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d16v0__pjunction_mult}
+ mjswgs = 0.78692
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.37073+sky130_fd_pr__nfet_g5v0d16v0__kt1_diff_4}
+ kt2 = {-0.019151+sky130_fd_pr__nfet_g5v0d16v0__kt2_diff_4}
+ at = 29000.0
+ ute = {-1.4324+sky130_fd_pr__nfet_g5v0d16v0__ute_diff_4}
+ ua1 = 2.0117e-9
+ ub1 = -2.9309e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d16v0__tvoff_diff_4}
+ njs = 1.0773
+ tpb = 0.001344
+ tcj = 0.00067434
+ tpbsw = 0.00099005
+ tcjsw = 0.0002493
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 0.76
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = .28e-6
+ sbref = 1.585e-6
+ kvth0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__kvth0_diff}
+ lkvth0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__lkvth0_diff}
+ wkvth0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 1.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__ku0_diff}
+ lku0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__lku0_diff}
+ wku0 = {0.0+sky130_fd_pr__nfet_g5v0d16v0__wku0_diff}
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 1.0
+ wlodku0 = 1.0
+ kvsat = {0.0+sky130_fd_pr__nfet_g5v0d16v0__kvsat_diff}
+ steta0 = 0.0
.ends sky130_fd_pr__nfet_g5v0d16v0__base
* Well Proximity Effect Parameters
