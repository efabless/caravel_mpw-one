magic
tech sky130A
magscale 1 2
timestamp 1606855431
<< obsli1 >>
rect 38 559 87806 188001
<< obsm1 >>
rect 38 6 87806 188554
<< obsm2 >>
rect 890 0 87186 189211
<< metal3 >>
rect 88454 189114 88934 189234
rect 88454 187890 88934 188010
rect 88454 186666 88934 186786
rect 88454 185442 88934 185562
rect 88454 184218 88934 184338
rect 88454 182994 88934 183114
rect 88454 181906 88934 182026
rect 88454 180682 88934 180802
rect 88454 179458 88934 179578
rect 88454 178234 88934 178354
rect 88454 177010 88934 177130
rect 88454 175786 88934 175906
rect 88454 174698 88934 174818
rect 88454 173474 88934 173594
rect 88454 172250 88934 172370
rect 88454 171026 88934 171146
rect 88454 169802 88934 169922
rect 88454 168578 88934 168698
rect 88454 167490 88934 167610
rect 88454 166266 88934 166386
rect 88454 165042 88934 165162
rect 88454 163818 88934 163938
rect 88454 162594 88934 162714
rect 88454 161370 88934 161490
rect 88454 160146 88934 160266
rect 88454 159058 88934 159178
rect 88454 157834 88934 157954
rect 88454 156610 88934 156730
rect 88454 155386 88934 155506
rect 88454 154162 88934 154282
rect 88454 152938 88934 153058
rect 88454 151850 88934 151970
rect 88454 150626 88934 150746
rect 88454 149402 88934 149522
rect 88454 148178 88934 148298
rect 88454 146954 88934 147074
rect 88454 145730 88934 145850
rect 88454 144642 88934 144762
rect 88454 143418 88934 143538
rect 88454 142194 88934 142314
rect 88454 140970 88934 141090
rect 88454 139746 88934 139866
rect 88454 138522 88934 138642
rect 88454 137298 88934 137418
rect 88454 136210 88934 136330
rect 88454 134986 88934 135106
rect 88454 133762 88934 133882
rect 88454 132538 88934 132658
rect 88454 131314 88934 131434
rect 88454 130090 88934 130210
rect 88454 129002 88934 129122
rect 88454 127778 88934 127898
rect 88454 126554 88934 126674
rect 88454 125330 88934 125450
rect 88454 124106 88934 124226
rect 88454 122882 88934 123002
rect 88454 121794 88934 121914
rect 88454 120570 88934 120690
rect 88454 119346 88934 119466
rect 88454 118122 88934 118242
rect 88454 116898 88934 117018
rect 88454 115674 88934 115794
rect 88454 114450 88934 114570
rect 88454 113362 88934 113482
rect 88454 112138 88934 112258
rect 88454 110914 88934 111034
rect 88454 109690 88934 109810
rect 88454 108466 88934 108586
rect 88454 107242 88934 107362
rect 88454 106154 88934 106274
rect 88454 104930 88934 105050
rect 88454 103706 88934 103826
rect 88454 102482 88934 102602
rect 88454 101258 88934 101378
rect 88454 100034 88934 100154
rect 88454 98946 88934 99066
rect 88454 97722 88934 97842
rect 88454 96498 88934 96618
rect 88454 95274 88934 95394
rect 88454 94050 88934 94170
rect 88454 92826 88934 92946
rect 88454 91602 88934 91722
rect 88454 90514 88934 90634
rect 88454 89290 88934 89410
rect 88454 88066 88934 88186
rect 88454 86842 88934 86962
rect 88454 85618 88934 85738
rect 88454 84394 88934 84514
rect 88454 83306 88934 83426
rect 88454 82082 88934 82202
rect 88454 80858 88934 80978
rect 88454 79634 88934 79754
rect 88454 78410 88934 78530
rect 88454 77186 88934 77306
rect 88454 76098 88934 76218
rect 88454 74874 88934 74994
rect 88454 73650 88934 73770
rect 88454 72426 88934 72546
rect 88454 71202 88934 71322
rect 88454 69978 88934 70098
rect 88454 68754 88934 68874
rect 88454 67666 88934 67786
rect 88454 66442 88934 66562
rect 88454 65218 88934 65338
rect 88454 63994 88934 64114
rect 88454 62770 88934 62890
rect 88454 61546 88934 61666
rect 88454 60458 88934 60578
rect 88454 59234 88934 59354
rect 88454 58010 88934 58130
rect 88454 56786 88934 56906
rect 88454 55562 88934 55682
rect 88454 54338 88934 54458
rect 88454 53250 88934 53370
rect 88454 52026 88934 52146
rect 88454 50802 88934 50922
rect 88454 49578 88934 49698
rect 88454 48354 88934 48474
rect 88454 47130 88934 47250
rect 88454 45906 88934 46026
rect 88454 44818 88934 44938
rect 88454 43594 88934 43714
rect 88454 42370 88934 42490
rect 88454 41146 88934 41266
rect 88454 39922 88934 40042
rect 88454 38698 88934 38818
rect 88454 37610 88934 37730
rect 88454 36386 88934 36506
rect 88454 35162 88934 35282
rect 88454 33938 88934 34058
rect 88454 32714 88934 32834
rect 88454 31490 88934 31610
rect 88454 30402 88934 30522
rect 88454 29178 88934 29298
rect 88454 27954 88934 28074
rect 88454 26730 88934 26850
rect 88454 25506 88934 25626
rect 88454 24282 88934 24402
rect 88454 23058 88934 23178
rect 88454 21970 88934 22090
rect 88454 20746 88934 20866
rect 88454 19522 88934 19642
rect 88454 18298 88934 18418
rect 88454 17074 88934 17194
rect 88454 15850 88934 15970
rect 88454 14762 88934 14882
rect 88454 13538 88934 13658
rect 88454 12314 88934 12434
rect 88454 11090 88934 11210
rect 88454 9866 88934 9986
rect 88454 8642 88934 8762
rect 88454 7554 88934 7674
rect 88454 6330 88934 6450
rect 88454 5106 88934 5226
rect 88454 3882 88934 4002
rect 88454 2658 88934 2778
rect 88454 1434 88934 1554
rect 88454 346 88934 466
<< obsm3 >>
rect 878 189034 88374 189207
rect 878 188090 88454 189034
rect 878 187810 88374 188090
rect 878 186866 88454 187810
rect 878 186586 88374 186866
rect 878 185642 88454 186586
rect 878 185362 88374 185642
rect 878 184418 88454 185362
rect 878 184138 88374 184418
rect 878 183194 88454 184138
rect 878 182914 88374 183194
rect 878 182106 88454 182914
rect 878 181826 88374 182106
rect 878 180882 88454 181826
rect 878 180602 88374 180882
rect 878 179658 88454 180602
rect 878 179378 88374 179658
rect 878 178434 88454 179378
rect 878 178154 88374 178434
rect 878 177210 88454 178154
rect 878 176930 88374 177210
rect 878 175986 88454 176930
rect 878 175706 88374 175986
rect 878 174898 88454 175706
rect 878 174618 88374 174898
rect 878 173674 88454 174618
rect 878 173394 88374 173674
rect 878 172450 88454 173394
rect 878 172170 88374 172450
rect 878 171226 88454 172170
rect 878 170946 88374 171226
rect 878 170002 88454 170946
rect 878 169722 88374 170002
rect 878 168778 88454 169722
rect 878 168498 88374 168778
rect 878 167690 88454 168498
rect 878 167410 88374 167690
rect 878 166466 88454 167410
rect 878 166186 88374 166466
rect 878 165242 88454 166186
rect 878 164962 88374 165242
rect 878 164018 88454 164962
rect 878 163738 88374 164018
rect 878 162794 88454 163738
rect 878 162514 88374 162794
rect 878 161570 88454 162514
rect 878 161290 88374 161570
rect 878 160346 88454 161290
rect 878 160066 88374 160346
rect 878 159258 88454 160066
rect 878 158978 88374 159258
rect 878 158034 88454 158978
rect 878 157754 88374 158034
rect 878 156810 88454 157754
rect 878 156530 88374 156810
rect 878 155586 88454 156530
rect 878 155306 88374 155586
rect 878 154362 88454 155306
rect 878 154082 88374 154362
rect 878 153138 88454 154082
rect 878 152858 88374 153138
rect 878 152050 88454 152858
rect 878 151770 88374 152050
rect 878 150826 88454 151770
rect 878 150546 88374 150826
rect 878 149602 88454 150546
rect 878 149322 88374 149602
rect 878 148378 88454 149322
rect 878 148098 88374 148378
rect 878 147154 88454 148098
rect 878 146874 88374 147154
rect 878 145930 88454 146874
rect 878 145650 88374 145930
rect 878 144842 88454 145650
rect 878 144562 88374 144842
rect 878 143618 88454 144562
rect 878 143338 88374 143618
rect 878 142394 88454 143338
rect 878 142114 88374 142394
rect 878 141170 88454 142114
rect 878 140890 88374 141170
rect 878 139946 88454 140890
rect 878 139666 88374 139946
rect 878 138722 88454 139666
rect 878 138442 88374 138722
rect 878 137498 88454 138442
rect 878 137218 88374 137498
rect 878 136410 88454 137218
rect 878 136130 88374 136410
rect 878 135186 88454 136130
rect 878 134906 88374 135186
rect 878 133962 88454 134906
rect 878 133682 88374 133962
rect 878 132738 88454 133682
rect 878 132458 88374 132738
rect 878 131514 88454 132458
rect 878 131234 88374 131514
rect 878 130290 88454 131234
rect 878 130010 88374 130290
rect 878 129202 88454 130010
rect 878 128922 88374 129202
rect 878 127978 88454 128922
rect 878 127698 88374 127978
rect 878 126754 88454 127698
rect 878 126474 88374 126754
rect 878 125530 88454 126474
rect 878 125250 88374 125530
rect 878 124306 88454 125250
rect 878 124026 88374 124306
rect 878 123082 88454 124026
rect 878 122802 88374 123082
rect 878 121994 88454 122802
rect 878 121714 88374 121994
rect 878 120770 88454 121714
rect 878 120490 88374 120770
rect 878 119546 88454 120490
rect 878 119266 88374 119546
rect 878 118322 88454 119266
rect 878 118042 88374 118322
rect 878 117098 88454 118042
rect 878 116818 88374 117098
rect 878 115874 88454 116818
rect 878 115594 88374 115874
rect 878 114650 88454 115594
rect 878 114370 88374 114650
rect 878 113562 88454 114370
rect 878 113282 88374 113562
rect 878 112338 88454 113282
rect 878 112058 88374 112338
rect 878 111114 88454 112058
rect 878 110834 88374 111114
rect 878 109890 88454 110834
rect 878 109610 88374 109890
rect 878 108666 88454 109610
rect 878 108386 88374 108666
rect 878 107442 88454 108386
rect 878 107162 88374 107442
rect 878 106354 88454 107162
rect 878 106074 88374 106354
rect 878 105130 88454 106074
rect 878 104850 88374 105130
rect 878 103906 88454 104850
rect 878 103626 88374 103906
rect 878 102682 88454 103626
rect 878 102402 88374 102682
rect 878 101458 88454 102402
rect 878 101178 88374 101458
rect 878 100234 88454 101178
rect 878 99954 88374 100234
rect 878 99146 88454 99954
rect 878 98866 88374 99146
rect 878 97922 88454 98866
rect 878 97642 88374 97922
rect 878 96698 88454 97642
rect 878 96418 88374 96698
rect 878 95474 88454 96418
rect 878 95194 88374 95474
rect 878 94250 88454 95194
rect 878 93970 88374 94250
rect 878 93026 88454 93970
rect 878 92746 88374 93026
rect 878 91802 88454 92746
rect 878 91522 88374 91802
rect 878 90714 88454 91522
rect 878 90434 88374 90714
rect 878 89490 88454 90434
rect 878 89210 88374 89490
rect 878 88266 88454 89210
rect 878 87986 88374 88266
rect 878 87042 88454 87986
rect 878 86762 88374 87042
rect 878 85818 88454 86762
rect 878 85538 88374 85818
rect 878 84594 88454 85538
rect 878 84314 88374 84594
rect 878 83506 88454 84314
rect 878 83226 88374 83506
rect 878 82282 88454 83226
rect 878 82002 88374 82282
rect 878 81058 88454 82002
rect 878 80778 88374 81058
rect 878 79834 88454 80778
rect 878 79554 88374 79834
rect 878 78610 88454 79554
rect 878 78330 88374 78610
rect 878 77386 88454 78330
rect 878 77106 88374 77386
rect 878 76298 88454 77106
rect 878 76018 88374 76298
rect 878 75074 88454 76018
rect 878 74794 88374 75074
rect 878 73850 88454 74794
rect 878 73570 88374 73850
rect 878 72626 88454 73570
rect 878 72346 88374 72626
rect 878 71402 88454 72346
rect 878 71122 88374 71402
rect 878 70178 88454 71122
rect 878 69898 88374 70178
rect 878 68954 88454 69898
rect 878 68674 88374 68954
rect 878 67866 88454 68674
rect 878 67586 88374 67866
rect 878 66642 88454 67586
rect 878 66362 88374 66642
rect 878 65418 88454 66362
rect 878 65138 88374 65418
rect 878 64194 88454 65138
rect 878 63914 88374 64194
rect 878 62970 88454 63914
rect 878 62690 88374 62970
rect 878 61746 88454 62690
rect 878 61466 88374 61746
rect 878 60658 88454 61466
rect 878 60378 88374 60658
rect 878 59434 88454 60378
rect 878 59154 88374 59434
rect 878 58210 88454 59154
rect 878 57930 88374 58210
rect 878 56986 88454 57930
rect 878 56706 88374 56986
rect 878 55762 88454 56706
rect 878 55482 88374 55762
rect 878 54538 88454 55482
rect 878 54258 88374 54538
rect 878 53450 88454 54258
rect 878 53170 88374 53450
rect 878 52226 88454 53170
rect 878 51946 88374 52226
rect 878 51002 88454 51946
rect 878 50722 88374 51002
rect 878 49778 88454 50722
rect 878 49498 88374 49778
rect 878 48554 88454 49498
rect 878 48274 88374 48554
rect 878 47330 88454 48274
rect 878 47050 88374 47330
rect 878 46106 88454 47050
rect 878 45826 88374 46106
rect 878 45018 88454 45826
rect 878 44738 88374 45018
rect 878 43794 88454 44738
rect 878 43514 88374 43794
rect 878 42570 88454 43514
rect 878 42290 88374 42570
rect 878 41346 88454 42290
rect 878 41066 88374 41346
rect 878 40122 88454 41066
rect 878 39842 88374 40122
rect 878 38898 88454 39842
rect 878 38618 88374 38898
rect 878 37810 88454 38618
rect 878 37530 88374 37810
rect 878 36586 88454 37530
rect 878 36306 88374 36586
rect 878 35362 88454 36306
rect 878 35082 88374 35362
rect 878 34138 88454 35082
rect 878 33858 88374 34138
rect 878 32914 88454 33858
rect 878 32634 88374 32914
rect 878 31690 88454 32634
rect 878 31410 88374 31690
rect 878 30602 88454 31410
rect 878 30322 88374 30602
rect 878 29378 88454 30322
rect 878 29098 88374 29378
rect 878 28154 88454 29098
rect 878 27874 88374 28154
rect 878 26930 88454 27874
rect 878 26650 88374 26930
rect 878 25706 88454 26650
rect 878 25426 88374 25706
rect 878 24482 88454 25426
rect 878 24202 88374 24482
rect 878 23258 88454 24202
rect 878 22978 88374 23258
rect 878 22170 88454 22978
rect 878 21890 88374 22170
rect 878 20946 88454 21890
rect 878 20666 88374 20946
rect 878 19722 88454 20666
rect 878 19442 88374 19722
rect 878 18498 88454 19442
rect 878 18218 88374 18498
rect 878 17274 88454 18218
rect 878 16994 88374 17274
rect 878 16050 88454 16994
rect 878 15770 88374 16050
rect 878 14962 88454 15770
rect 878 14682 88374 14962
rect 878 13738 88454 14682
rect 878 13458 88374 13738
rect 878 12514 88454 13458
rect 878 12234 88374 12514
rect 878 11290 88454 12234
rect 878 11010 88374 11290
rect 878 10066 88454 11010
rect 878 9786 88374 10066
rect 878 8842 88454 9786
rect 878 8562 88374 8842
rect 878 7754 88454 8562
rect 878 7474 88374 7754
rect 878 6530 88454 7474
rect 878 6250 88374 6530
rect 878 5306 88454 6250
rect 878 5026 88374 5306
rect 878 4082 88454 5026
rect 878 3802 88374 4082
rect 878 2858 88454 3802
rect 878 2578 88374 2858
rect 878 1634 88454 2578
rect 878 1354 88374 1634
rect 878 546 88454 1354
rect 878 266 88374 546
rect 878 101 88454 266
<< obsm4 >>
rect 878 101 87198 187983
<< metal5 >>
rect 38 10092 87806 10412
rect 38 5092 87806 5412
<< obsm5 >>
rect 38 15092 87806 185412
<< labels >>
rlabel metal3 s 88454 346 88934 466 6 mgmt_addr[0]
port 1 nsew default input
rlabel metal3 s 88454 1434 88934 1554 6 mgmt_addr[1]
port 2 nsew default input
rlabel metal3 s 88454 2658 88934 2778 6 mgmt_addr[2]
port 3 nsew default input
rlabel metal3 s 88454 3882 88934 4002 6 mgmt_addr[3]
port 4 nsew default input
rlabel metal3 s 88454 5106 88934 5226 6 mgmt_addr[4]
port 5 nsew default input
rlabel metal3 s 88454 6330 88934 6450 6 mgmt_addr[5]
port 6 nsew default input
rlabel metal3 s 88454 7554 88934 7674 6 mgmt_addr[6]
port 7 nsew default input
rlabel metal3 s 88454 8642 88934 8762 6 mgmt_addr[7]
port 8 nsew default input
rlabel metal3 s 88454 9866 88934 9986 6 mgmt_addr_ro[0]
port 9 nsew default input
rlabel metal3 s 88454 11090 88934 11210 6 mgmt_addr_ro[1]
port 10 nsew default input
rlabel metal3 s 88454 12314 88934 12434 6 mgmt_addr_ro[2]
port 11 nsew default input
rlabel metal3 s 88454 13538 88934 13658 6 mgmt_addr_ro[3]
port 12 nsew default input
rlabel metal3 s 88454 14762 88934 14882 6 mgmt_addr_ro[4]
port 13 nsew default input
rlabel metal3 s 88454 15850 88934 15970 6 mgmt_addr_ro[5]
port 14 nsew default input
rlabel metal3 s 88454 17074 88934 17194 6 mgmt_addr_ro[6]
port 15 nsew default input
rlabel metal3 s 88454 18298 88934 18418 6 mgmt_addr_ro[7]
port 16 nsew default input
rlabel metal3 s 88454 19522 88934 19642 6 mgmt_clk
port 17 nsew default input
rlabel metal3 s 88454 20746 88934 20866 6 mgmt_ena[0]
port 18 nsew default input
rlabel metal3 s 88454 21970 88934 22090 6 mgmt_ena[1]
port 19 nsew default input
rlabel metal3 s 88454 23058 88934 23178 6 mgmt_ena_ro
port 20 nsew default input
rlabel metal3 s 88454 24282 88934 24402 6 mgmt_rdata[0]
port 21 nsew default output
rlabel metal3 s 88454 36386 88934 36506 6 mgmt_rdata[10]
port 22 nsew default output
rlabel metal3 s 88454 37610 88934 37730 6 mgmt_rdata[11]
port 23 nsew default output
rlabel metal3 s 88454 38698 88934 38818 6 mgmt_rdata[12]
port 24 nsew default output
rlabel metal3 s 88454 39922 88934 40042 6 mgmt_rdata[13]
port 25 nsew default output
rlabel metal3 s 88454 41146 88934 41266 6 mgmt_rdata[14]
port 26 nsew default output
rlabel metal3 s 88454 42370 88934 42490 6 mgmt_rdata[15]
port 27 nsew default output
rlabel metal3 s 88454 43594 88934 43714 6 mgmt_rdata[16]
port 28 nsew default output
rlabel metal3 s 88454 44818 88934 44938 6 mgmt_rdata[17]
port 29 nsew default output
rlabel metal3 s 88454 45906 88934 46026 6 mgmt_rdata[18]
port 30 nsew default output
rlabel metal3 s 88454 47130 88934 47250 6 mgmt_rdata[19]
port 31 nsew default output
rlabel metal3 s 88454 25506 88934 25626 6 mgmt_rdata[1]
port 32 nsew default output
rlabel metal3 s 88454 48354 88934 48474 6 mgmt_rdata[20]
port 33 nsew default output
rlabel metal3 s 88454 49578 88934 49698 6 mgmt_rdata[21]
port 34 nsew default output
rlabel metal3 s 88454 50802 88934 50922 6 mgmt_rdata[22]
port 35 nsew default output
rlabel metal3 s 88454 52026 88934 52146 6 mgmt_rdata[23]
port 36 nsew default output
rlabel metal3 s 88454 53250 88934 53370 6 mgmt_rdata[24]
port 37 nsew default output
rlabel metal3 s 88454 54338 88934 54458 6 mgmt_rdata[25]
port 38 nsew default output
rlabel metal3 s 88454 55562 88934 55682 6 mgmt_rdata[26]
port 39 nsew default output
rlabel metal3 s 88454 56786 88934 56906 6 mgmt_rdata[27]
port 40 nsew default output
rlabel metal3 s 88454 58010 88934 58130 6 mgmt_rdata[28]
port 41 nsew default output
rlabel metal3 s 88454 59234 88934 59354 6 mgmt_rdata[29]
port 42 nsew default output
rlabel metal3 s 88454 26730 88934 26850 6 mgmt_rdata[2]
port 43 nsew default output
rlabel metal3 s 88454 60458 88934 60578 6 mgmt_rdata[30]
port 44 nsew default output
rlabel metal3 s 88454 61546 88934 61666 6 mgmt_rdata[31]
port 45 nsew default output
rlabel metal3 s 88454 62770 88934 62890 6 mgmt_rdata[32]
port 46 nsew default output
rlabel metal3 s 88454 63994 88934 64114 6 mgmt_rdata[33]
port 47 nsew default output
rlabel metal3 s 88454 65218 88934 65338 6 mgmt_rdata[34]
port 48 nsew default output
rlabel metal3 s 88454 66442 88934 66562 6 mgmt_rdata[35]
port 49 nsew default output
rlabel metal3 s 88454 67666 88934 67786 6 mgmt_rdata[36]
port 50 nsew default output
rlabel metal3 s 88454 68754 88934 68874 6 mgmt_rdata[37]
port 51 nsew default output
rlabel metal3 s 88454 69978 88934 70098 6 mgmt_rdata[38]
port 52 nsew default output
rlabel metal3 s 88454 71202 88934 71322 6 mgmt_rdata[39]
port 53 nsew default output
rlabel metal3 s 88454 27954 88934 28074 6 mgmt_rdata[3]
port 54 nsew default output
rlabel metal3 s 88454 72426 88934 72546 6 mgmt_rdata[40]
port 55 nsew default output
rlabel metal3 s 88454 73650 88934 73770 6 mgmt_rdata[41]
port 56 nsew default output
rlabel metal3 s 88454 74874 88934 74994 6 mgmt_rdata[42]
port 57 nsew default output
rlabel metal3 s 88454 76098 88934 76218 6 mgmt_rdata[43]
port 58 nsew default output
rlabel metal3 s 88454 77186 88934 77306 6 mgmt_rdata[44]
port 59 nsew default output
rlabel metal3 s 88454 78410 88934 78530 6 mgmt_rdata[45]
port 60 nsew default output
rlabel metal3 s 88454 79634 88934 79754 6 mgmt_rdata[46]
port 61 nsew default output
rlabel metal3 s 88454 80858 88934 80978 6 mgmt_rdata[47]
port 62 nsew default output
rlabel metal3 s 88454 82082 88934 82202 6 mgmt_rdata[48]
port 63 nsew default output
rlabel metal3 s 88454 83306 88934 83426 6 mgmt_rdata[49]
port 64 nsew default output
rlabel metal3 s 88454 29178 88934 29298 6 mgmt_rdata[4]
port 65 nsew default output
rlabel metal3 s 88454 84394 88934 84514 6 mgmt_rdata[50]
port 66 nsew default output
rlabel metal3 s 88454 85618 88934 85738 6 mgmt_rdata[51]
port 67 nsew default output
rlabel metal3 s 88454 86842 88934 86962 6 mgmt_rdata[52]
port 68 nsew default output
rlabel metal3 s 88454 88066 88934 88186 6 mgmt_rdata[53]
port 69 nsew default output
rlabel metal3 s 88454 89290 88934 89410 6 mgmt_rdata[54]
port 70 nsew default output
rlabel metal3 s 88454 90514 88934 90634 6 mgmt_rdata[55]
port 71 nsew default output
rlabel metal3 s 88454 91602 88934 91722 6 mgmt_rdata[56]
port 72 nsew default output
rlabel metal3 s 88454 92826 88934 92946 6 mgmt_rdata[57]
port 73 nsew default output
rlabel metal3 s 88454 94050 88934 94170 6 mgmt_rdata[58]
port 74 nsew default output
rlabel metal3 s 88454 95274 88934 95394 6 mgmt_rdata[59]
port 75 nsew default output
rlabel metal3 s 88454 30402 88934 30522 6 mgmt_rdata[5]
port 76 nsew default output
rlabel metal3 s 88454 96498 88934 96618 6 mgmt_rdata[60]
port 77 nsew default output
rlabel metal3 s 88454 97722 88934 97842 6 mgmt_rdata[61]
port 78 nsew default output
rlabel metal3 s 88454 98946 88934 99066 6 mgmt_rdata[62]
port 79 nsew default output
rlabel metal3 s 88454 100034 88934 100154 6 mgmt_rdata[63]
port 80 nsew default output
rlabel metal3 s 88454 31490 88934 31610 6 mgmt_rdata[6]
port 81 nsew default output
rlabel metal3 s 88454 32714 88934 32834 6 mgmt_rdata[7]
port 82 nsew default output
rlabel metal3 s 88454 33938 88934 34058 6 mgmt_rdata[8]
port 83 nsew default output
rlabel metal3 s 88454 35162 88934 35282 6 mgmt_rdata[9]
port 84 nsew default output
rlabel metal3 s 88454 101258 88934 101378 6 mgmt_rdata_ro[0]
port 85 nsew default output
rlabel metal3 s 88454 113362 88934 113482 6 mgmt_rdata_ro[10]
port 86 nsew default output
rlabel metal3 s 88454 114450 88934 114570 6 mgmt_rdata_ro[11]
port 87 nsew default output
rlabel metal3 s 88454 115674 88934 115794 6 mgmt_rdata_ro[12]
port 88 nsew default output
rlabel metal3 s 88454 116898 88934 117018 6 mgmt_rdata_ro[13]
port 89 nsew default output
rlabel metal3 s 88454 118122 88934 118242 6 mgmt_rdata_ro[14]
port 90 nsew default output
rlabel metal3 s 88454 119346 88934 119466 6 mgmt_rdata_ro[15]
port 91 nsew default output
rlabel metal3 s 88454 120570 88934 120690 6 mgmt_rdata_ro[16]
port 92 nsew default output
rlabel metal3 s 88454 121794 88934 121914 6 mgmt_rdata_ro[17]
port 93 nsew default output
rlabel metal3 s 88454 122882 88934 123002 6 mgmt_rdata_ro[18]
port 94 nsew default output
rlabel metal3 s 88454 124106 88934 124226 6 mgmt_rdata_ro[19]
port 95 nsew default output
rlabel metal3 s 88454 102482 88934 102602 6 mgmt_rdata_ro[1]
port 96 nsew default output
rlabel metal3 s 88454 125330 88934 125450 6 mgmt_rdata_ro[20]
port 97 nsew default output
rlabel metal3 s 88454 126554 88934 126674 6 mgmt_rdata_ro[21]
port 98 nsew default output
rlabel metal3 s 88454 127778 88934 127898 6 mgmt_rdata_ro[22]
port 99 nsew default output
rlabel metal3 s 88454 129002 88934 129122 6 mgmt_rdata_ro[23]
port 100 nsew default output
rlabel metal3 s 88454 130090 88934 130210 6 mgmt_rdata_ro[24]
port 101 nsew default output
rlabel metal3 s 88454 131314 88934 131434 6 mgmt_rdata_ro[25]
port 102 nsew default output
rlabel metal3 s 88454 132538 88934 132658 6 mgmt_rdata_ro[26]
port 103 nsew default output
rlabel metal3 s 88454 133762 88934 133882 6 mgmt_rdata_ro[27]
port 104 nsew default output
rlabel metal3 s 88454 134986 88934 135106 6 mgmt_rdata_ro[28]
port 105 nsew default output
rlabel metal3 s 88454 136210 88934 136330 6 mgmt_rdata_ro[29]
port 106 nsew default output
rlabel metal3 s 88454 103706 88934 103826 6 mgmt_rdata_ro[2]
port 107 nsew default output
rlabel metal3 s 88454 137298 88934 137418 6 mgmt_rdata_ro[30]
port 108 nsew default output
rlabel metal3 s 88454 138522 88934 138642 6 mgmt_rdata_ro[31]
port 109 nsew default output
rlabel metal3 s 88454 104930 88934 105050 6 mgmt_rdata_ro[3]
port 110 nsew default output
rlabel metal3 s 88454 106154 88934 106274 6 mgmt_rdata_ro[4]
port 111 nsew default output
rlabel metal3 s 88454 107242 88934 107362 6 mgmt_rdata_ro[5]
port 112 nsew default output
rlabel metal3 s 88454 108466 88934 108586 6 mgmt_rdata_ro[6]
port 113 nsew default output
rlabel metal3 s 88454 109690 88934 109810 6 mgmt_rdata_ro[7]
port 114 nsew default output
rlabel metal3 s 88454 110914 88934 111034 6 mgmt_rdata_ro[8]
port 115 nsew default output
rlabel metal3 s 88454 112138 88934 112258 6 mgmt_rdata_ro[9]
port 116 nsew default output
rlabel metal3 s 88454 139746 88934 139866 6 mgmt_wdata[0]
port 117 nsew default input
rlabel metal3 s 88454 151850 88934 151970 6 mgmt_wdata[10]
port 118 nsew default input
rlabel metal3 s 88454 152938 88934 153058 6 mgmt_wdata[11]
port 119 nsew default input
rlabel metal3 s 88454 154162 88934 154282 6 mgmt_wdata[12]
port 120 nsew default input
rlabel metal3 s 88454 155386 88934 155506 6 mgmt_wdata[13]
port 121 nsew default input
rlabel metal3 s 88454 156610 88934 156730 6 mgmt_wdata[14]
port 122 nsew default input
rlabel metal3 s 88454 157834 88934 157954 6 mgmt_wdata[15]
port 123 nsew default input
rlabel metal3 s 88454 159058 88934 159178 6 mgmt_wdata[16]
port 124 nsew default input
rlabel metal3 s 88454 160146 88934 160266 6 mgmt_wdata[17]
port 125 nsew default input
rlabel metal3 s 88454 161370 88934 161490 6 mgmt_wdata[18]
port 126 nsew default input
rlabel metal3 s 88454 162594 88934 162714 6 mgmt_wdata[19]
port 127 nsew default input
rlabel metal3 s 88454 140970 88934 141090 6 mgmt_wdata[1]
port 128 nsew default input
rlabel metal3 s 88454 163818 88934 163938 6 mgmt_wdata[20]
port 129 nsew default input
rlabel metal3 s 88454 165042 88934 165162 6 mgmt_wdata[21]
port 130 nsew default input
rlabel metal3 s 88454 166266 88934 166386 6 mgmt_wdata[22]
port 131 nsew default input
rlabel metal3 s 88454 167490 88934 167610 6 mgmt_wdata[23]
port 132 nsew default input
rlabel metal3 s 88454 168578 88934 168698 6 mgmt_wdata[24]
port 133 nsew default input
rlabel metal3 s 88454 169802 88934 169922 6 mgmt_wdata[25]
port 134 nsew default input
rlabel metal3 s 88454 171026 88934 171146 6 mgmt_wdata[26]
port 135 nsew default input
rlabel metal3 s 88454 172250 88934 172370 6 mgmt_wdata[27]
port 136 nsew default input
rlabel metal3 s 88454 173474 88934 173594 6 mgmt_wdata[28]
port 137 nsew default input
rlabel metal3 s 88454 174698 88934 174818 6 mgmt_wdata[29]
port 138 nsew default input
rlabel metal3 s 88454 142194 88934 142314 6 mgmt_wdata[2]
port 139 nsew default input
rlabel metal3 s 88454 175786 88934 175906 6 mgmt_wdata[30]
port 140 nsew default input
rlabel metal3 s 88454 177010 88934 177130 6 mgmt_wdata[31]
port 141 nsew default input
rlabel metal3 s 88454 143418 88934 143538 6 mgmt_wdata[3]
port 142 nsew default input
rlabel metal3 s 88454 144642 88934 144762 6 mgmt_wdata[4]
port 143 nsew default input
rlabel metal3 s 88454 145730 88934 145850 6 mgmt_wdata[5]
port 144 nsew default input
rlabel metal3 s 88454 146954 88934 147074 6 mgmt_wdata[6]
port 145 nsew default input
rlabel metal3 s 88454 148178 88934 148298 6 mgmt_wdata[7]
port 146 nsew default input
rlabel metal3 s 88454 149402 88934 149522 6 mgmt_wdata[8]
port 147 nsew default input
rlabel metal3 s 88454 150626 88934 150746 6 mgmt_wdata[9]
port 148 nsew default input
rlabel metal3 s 88454 178234 88934 178354 6 mgmt_wen[0]
port 149 nsew default input
rlabel metal3 s 88454 179458 88934 179578 6 mgmt_wen[1]
port 150 nsew default input
rlabel metal3 s 88454 180682 88934 180802 6 mgmt_wen_mask[0]
port 151 nsew default input
rlabel metal3 s 88454 181906 88934 182026 6 mgmt_wen_mask[1]
port 152 nsew default input
rlabel metal3 s 88454 182994 88934 183114 6 mgmt_wen_mask[2]
port 153 nsew default input
rlabel metal3 s 88454 184218 88934 184338 6 mgmt_wen_mask[3]
port 154 nsew default input
rlabel metal3 s 88454 185442 88934 185562 6 mgmt_wen_mask[4]
port 155 nsew default input
rlabel metal3 s 88454 186666 88934 186786 6 mgmt_wen_mask[5]
port 156 nsew default input
rlabel metal3 s 88454 187890 88934 188010 6 mgmt_wen_mask[6]
port 157 nsew default input
rlabel metal3 s 88454 189114 88934 189234 6 mgmt_wen_mask[7]
port 158 nsew default input
rlabel metal5 s 38 5092 87806 5412 6 VPWR
port 159 nsew power input
rlabel metal5 s 38 10092 87806 10412 6 VGND
port 160 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 88934 189234
string LEFview TRUE
string GDS_FILE ../gds/storage.gds
string GDS_END 15067618
string GDS_START 13323184
<< end >>

