magic
tech sky130A
magscale 1 2
timestamp 1624446576
<< nwell >>
rect 1066 189029 5190 189350
rect 1066 187941 5190 188507
rect 1066 186853 5190 187419
rect 1066 185765 5190 186331
rect 1066 184677 5190 185243
rect 1066 183589 5190 184155
rect 1066 182501 5190 183067
rect 1066 181413 5190 181979
rect 1066 180325 5190 180891
rect 1066 179237 5190 179803
rect 1066 178149 5190 178715
rect 1066 177061 5190 177627
rect 1066 175973 5190 176539
rect 1066 174885 5190 175451
rect 1066 173797 5190 174363
rect 1066 172709 5190 173275
rect 1066 171621 5190 172187
rect 1066 170533 5190 171099
rect 1066 169445 5190 170011
rect 1066 168357 5190 168923
rect 1066 167269 5190 167835
rect 1066 166181 5190 166747
rect 1066 165093 5190 165659
rect 1066 164005 5190 164571
rect 1066 162917 5190 163483
rect 1066 161829 5190 162395
rect 1066 160741 5190 161307
rect 1066 159653 5190 160219
rect 1066 158565 5190 159131
rect 1066 157477 5190 158043
rect 1066 156389 5190 156955
rect 1066 155301 5190 155867
rect 1066 154213 5190 154779
rect 1066 153125 5190 153691
rect 1066 152037 5190 152603
rect 1066 150949 5190 151515
rect 1066 149861 5190 150427
rect 1066 148773 5190 149339
rect 1066 147685 5190 148251
rect 1066 146597 5190 147163
rect 1066 145509 5190 146075
rect 1066 144421 5190 144987
rect 1066 143333 5190 143899
rect 1066 142245 5190 142811
rect 1066 141157 5190 141723
rect 1066 140069 5190 140635
rect 1066 138981 5190 139547
rect 1066 137893 5190 138459
rect 1066 136805 5190 137371
rect 1066 135717 5190 136283
rect 1066 134629 5190 135195
rect 1066 133541 5190 134107
rect 1066 132453 5190 133019
rect 1066 131365 5190 131931
rect 1066 130277 5190 130843
rect 1066 129189 5190 129755
rect 1066 128101 5190 128667
rect 1066 127013 5190 127579
rect 1066 125925 5190 126491
rect 1066 124837 5190 125403
rect 1066 123749 5190 124315
rect 1066 122661 5190 123227
rect 1066 121573 5190 122139
rect 1066 120485 5190 121051
rect 1066 119397 5190 119963
rect 1066 118309 5190 118875
rect 1066 117221 5190 117787
rect 1066 116133 5190 116699
rect 1066 115045 5190 115611
rect 1066 113957 5190 114523
rect 1066 112869 5190 113435
rect 1066 111781 5190 112347
rect 1066 110693 5190 111259
rect 1066 109605 5190 110171
rect 1066 108517 5190 109083
rect 1066 107429 5190 107995
rect 1066 106341 5190 106907
rect 1066 105253 5190 105819
rect 1066 104165 5190 104731
rect 1066 103077 5190 103643
rect 1066 101989 5190 102555
rect 1066 100901 5190 101467
rect 1066 99813 5190 100379
rect 1066 98725 5190 99291
rect 1066 97637 5190 98203
rect 1066 96549 5190 97115
rect 1066 95461 5190 96027
rect 1066 94373 5190 94939
rect 1066 93285 5190 93851
rect 1066 92197 5190 92763
rect 1066 91109 5190 91675
rect 1066 90021 5190 90587
rect 1066 88933 5190 89499
rect 1066 87845 5190 88411
rect 1066 86757 5190 87323
rect 1066 85669 5190 86235
rect 1066 84581 5190 85147
rect 1066 83493 5190 84059
rect 1066 82405 5190 82971
rect 1066 81317 5190 81883
rect 1066 80229 5190 80795
rect 1066 79141 5190 79707
rect 1066 78053 5190 78619
rect 1066 76965 5190 77531
rect 1066 75877 5190 76443
rect 1066 74789 5190 75355
rect 1066 73701 5190 74267
rect 1066 72613 5190 73179
rect 1066 71525 5190 72091
rect 1066 70437 5190 71003
rect 1066 69349 5190 69915
rect 1066 68261 5190 68827
rect 1066 67173 5190 67739
rect 1066 66085 5190 66651
rect 1066 64997 5190 65563
rect 1066 63909 5190 64475
rect 1066 62821 5190 63387
rect 1066 61733 5190 62299
rect 1066 60645 5190 61211
rect 1066 59557 5190 60123
rect 1066 58469 5190 59035
rect 1066 57381 5190 57947
rect 1066 56293 5190 56859
rect 1066 55205 5190 55771
rect 1066 54117 5190 54683
rect 1066 53029 5190 53595
rect 1066 51941 5190 52507
rect 1066 50853 5190 51419
rect 1066 49765 5190 50331
rect 1066 48677 5190 49243
rect 1066 47589 5190 48155
rect 1066 46501 5190 47067
rect 1066 45413 5190 45979
rect 1066 44325 5190 44891
rect 1066 43237 5190 43803
rect 1066 42149 5190 42715
rect 1066 41061 5190 41627
rect 1066 39973 5190 40539
rect 1066 38885 5190 39451
rect 1066 37797 5190 38363
rect 1066 36709 5190 37275
rect 1066 35621 5190 36187
rect 1066 34533 5190 35099
rect 1066 33445 5190 34011
rect 1066 32357 5190 32923
rect 1066 31269 5190 31835
rect 1066 30181 5190 30747
rect 1066 29093 5190 29659
rect 1066 28005 5190 28571
rect 1066 26917 5190 27483
rect 1066 25829 5190 26395
rect 1066 24741 5190 25307
rect 1066 23653 5190 24219
rect 1066 22565 5190 23131
rect 1066 21477 5190 22043
rect 1066 20389 5190 20955
rect 1066 19301 5190 19867
rect 1066 18213 5190 18779
rect 1066 17125 5190 17691
rect 1066 16037 5190 16603
rect 1066 14949 5190 15515
rect 1066 13861 5190 14427
rect 1066 12773 5190 13339
rect 1066 11685 5190 12251
rect 1066 10597 5190 11163
rect 1066 9509 5190 10075
rect 1066 8421 5190 8987
rect 1066 7333 5190 7899
rect 1066 6245 5190 6811
rect 1066 5157 5190 5723
rect 1066 4069 5190 4635
rect 1066 2981 5190 3547
rect 1066 2138 5190 2459
<< obsli1 >>
rect 1104 1581 90896 189329
<< obsm1 >>
rect 1104 76 90896 189360
<< obsm2 >>
rect 1956 70 90418 189360
<< metal3 >>
rect 91200 191360 92000 191480
rect 91200 190136 92000 190256
rect 91200 188912 92000 189032
rect 91200 187688 92000 187808
rect 91200 186464 92000 186584
rect 91200 185240 92000 185360
rect 91200 184016 92000 184136
rect 91200 182792 92000 182912
rect 91200 181568 92000 181688
rect 91200 180344 92000 180464
rect 91200 179120 92000 179240
rect 91200 177896 92000 178016
rect 91200 176672 92000 176792
rect 91200 175448 92000 175568
rect 91200 174224 92000 174344
rect 91200 173136 92000 173256
rect 91200 171912 92000 172032
rect 91200 170688 92000 170808
rect 91200 169464 92000 169584
rect 91200 168240 92000 168360
rect 91200 167016 92000 167136
rect 91200 165792 92000 165912
rect 91200 164568 92000 164688
rect 91200 163344 92000 163464
rect 91200 162120 92000 162240
rect 91200 160896 92000 161016
rect 91200 159672 92000 159792
rect 91200 158448 92000 158568
rect 91200 157224 92000 157344
rect 91200 156000 92000 156120
rect 91200 154776 92000 154896
rect 91200 153688 92000 153808
rect 91200 152464 92000 152584
rect 91200 151240 92000 151360
rect 91200 150016 92000 150136
rect 91200 148792 92000 148912
rect 91200 147568 92000 147688
rect 91200 146344 92000 146464
rect 91200 145120 92000 145240
rect 91200 143896 92000 144016
rect 91200 142672 92000 142792
rect 91200 141448 92000 141568
rect 91200 140224 92000 140344
rect 91200 139000 92000 139120
rect 91200 137776 92000 137896
rect 91200 136552 92000 136672
rect 91200 135328 92000 135448
rect 91200 134240 92000 134360
rect 91200 133016 92000 133136
rect 91200 131792 92000 131912
rect 91200 130568 92000 130688
rect 91200 129344 92000 129464
rect 91200 128120 92000 128240
rect 91200 126896 92000 127016
rect 91200 125672 92000 125792
rect 91200 124448 92000 124568
rect 91200 123224 92000 123344
rect 91200 122000 92000 122120
rect 91200 120776 92000 120896
rect 91200 119552 92000 119672
rect 91200 118328 92000 118448
rect 91200 117104 92000 117224
rect 91200 115880 92000 116000
rect 91200 114792 92000 114912
rect 91200 113568 92000 113688
rect 91200 112344 92000 112464
rect 91200 111120 92000 111240
rect 91200 109896 92000 110016
rect 91200 108672 92000 108792
rect 91200 107448 92000 107568
rect 91200 106224 92000 106344
rect 91200 105000 92000 105120
rect 91200 103776 92000 103896
rect 91200 102552 92000 102672
rect 91200 101328 92000 101448
rect 91200 100104 92000 100224
rect 91200 98880 92000 99000
rect 91200 97656 92000 97776
rect 91200 96568 92000 96688
rect 91200 95344 92000 95464
rect 91200 94120 92000 94240
rect 91200 92896 92000 93016
rect 91200 91672 92000 91792
rect 91200 90448 92000 90568
rect 91200 89224 92000 89344
rect 91200 88000 92000 88120
rect 91200 86776 92000 86896
rect 91200 85552 92000 85672
rect 91200 84328 92000 84448
rect 91200 83104 92000 83224
rect 91200 81880 92000 82000
rect 91200 80656 92000 80776
rect 91200 79432 92000 79552
rect 91200 78208 92000 78328
rect 91200 77120 92000 77240
rect 91200 75896 92000 76016
rect 91200 74672 92000 74792
rect 91200 73448 92000 73568
rect 91200 72224 92000 72344
rect 91200 71000 92000 71120
rect 91200 69776 92000 69896
rect 91200 68552 92000 68672
rect 91200 67328 92000 67448
rect 91200 66104 92000 66224
rect 91200 64880 92000 65000
rect 91200 63656 92000 63776
rect 91200 62432 92000 62552
rect 91200 61208 92000 61328
rect 91200 59984 92000 60104
rect 91200 58760 92000 58880
rect 91200 57672 92000 57792
rect 91200 56448 92000 56568
rect 91200 55224 92000 55344
rect 91200 54000 92000 54120
rect 91200 52776 92000 52896
rect 91200 51552 92000 51672
rect 91200 50328 92000 50448
rect 91200 49104 92000 49224
rect 91200 47880 92000 48000
rect 91200 46656 92000 46776
rect 91200 45432 92000 45552
rect 91200 44208 92000 44328
rect 91200 42984 92000 43104
rect 91200 41760 92000 41880
rect 91200 40536 92000 40656
rect 91200 39312 92000 39432
rect 91200 38224 92000 38344
rect 91200 37000 92000 37120
rect 91200 35776 92000 35896
rect 91200 34552 92000 34672
rect 91200 33328 92000 33448
rect 91200 32104 92000 32224
rect 91200 30880 92000 31000
rect 91200 29656 92000 29776
rect 91200 28432 92000 28552
rect 91200 27208 92000 27328
rect 91200 25984 92000 26104
rect 91200 24760 92000 24880
rect 91200 23536 92000 23656
rect 91200 22312 92000 22432
rect 91200 21088 92000 21208
rect 91200 19864 92000 19984
rect 91200 18776 92000 18896
rect 91200 17552 92000 17672
rect 91200 16328 92000 16448
rect 91200 15104 92000 15224
rect 91200 13880 92000 14000
rect 91200 12656 92000 12776
rect 91200 11432 92000 11552
rect 91200 10208 92000 10328
rect 91200 8984 92000 9104
rect 91200 7760 92000 7880
rect 91200 6536 92000 6656
rect 91200 5312 92000 5432
rect 91200 4088 92000 4208
rect 91200 2864 92000 2984
rect 91200 1640 92000 1760
rect 91200 552 92000 672
<< obsm3 >>
rect 1944 191280 91120 191452
rect 1944 190336 91200 191280
rect 1944 190056 91120 190336
rect 1944 189112 91200 190056
rect 1944 188832 91120 189112
rect 1944 187888 91200 188832
rect 1944 187608 91120 187888
rect 1944 186664 91200 187608
rect 1944 186384 91120 186664
rect 1944 185440 91200 186384
rect 1944 185160 91120 185440
rect 1944 184216 91200 185160
rect 1944 183936 91120 184216
rect 1944 182992 91200 183936
rect 1944 182712 91120 182992
rect 1944 181768 91200 182712
rect 1944 181488 91120 181768
rect 1944 180544 91200 181488
rect 1944 180264 91120 180544
rect 1944 179320 91200 180264
rect 1944 179040 91120 179320
rect 1944 178096 91200 179040
rect 1944 177816 91120 178096
rect 1944 176872 91200 177816
rect 1944 176592 91120 176872
rect 1944 175648 91200 176592
rect 1944 175368 91120 175648
rect 1944 174424 91200 175368
rect 1944 174144 91120 174424
rect 1944 173336 91200 174144
rect 1944 173056 91120 173336
rect 1944 172112 91200 173056
rect 1944 171832 91120 172112
rect 1944 170888 91200 171832
rect 1944 170608 91120 170888
rect 1944 169664 91200 170608
rect 1944 169384 91120 169664
rect 1944 168440 91200 169384
rect 1944 168160 91120 168440
rect 1944 167216 91200 168160
rect 1944 166936 91120 167216
rect 1944 165992 91200 166936
rect 1944 165712 91120 165992
rect 1944 164768 91200 165712
rect 1944 164488 91120 164768
rect 1944 163544 91200 164488
rect 1944 163264 91120 163544
rect 1944 162320 91200 163264
rect 1944 162040 91120 162320
rect 1944 161096 91200 162040
rect 1944 160816 91120 161096
rect 1944 159872 91200 160816
rect 1944 159592 91120 159872
rect 1944 158648 91200 159592
rect 1944 158368 91120 158648
rect 1944 157424 91200 158368
rect 1944 157144 91120 157424
rect 1944 156200 91200 157144
rect 1944 155920 91120 156200
rect 1944 154976 91200 155920
rect 1944 154696 91120 154976
rect 1944 153888 91200 154696
rect 1944 153608 91120 153888
rect 1944 152664 91200 153608
rect 1944 152384 91120 152664
rect 1944 151440 91200 152384
rect 1944 151160 91120 151440
rect 1944 150216 91200 151160
rect 1944 149936 91120 150216
rect 1944 148992 91200 149936
rect 1944 148712 91120 148992
rect 1944 147768 91200 148712
rect 1944 147488 91120 147768
rect 1944 146544 91200 147488
rect 1944 146264 91120 146544
rect 1944 145320 91200 146264
rect 1944 145040 91120 145320
rect 1944 144096 91200 145040
rect 1944 143816 91120 144096
rect 1944 142872 91200 143816
rect 1944 142592 91120 142872
rect 1944 141648 91200 142592
rect 1944 141368 91120 141648
rect 1944 140424 91200 141368
rect 1944 140144 91120 140424
rect 1944 139200 91200 140144
rect 1944 138920 91120 139200
rect 1944 137976 91200 138920
rect 1944 137696 91120 137976
rect 1944 136752 91200 137696
rect 1944 136472 91120 136752
rect 1944 135528 91200 136472
rect 1944 135248 91120 135528
rect 1944 134440 91200 135248
rect 1944 134160 91120 134440
rect 1944 133216 91200 134160
rect 1944 132936 91120 133216
rect 1944 131992 91200 132936
rect 1944 131712 91120 131992
rect 1944 130768 91200 131712
rect 1944 130488 91120 130768
rect 1944 129544 91200 130488
rect 1944 129264 91120 129544
rect 1944 128320 91200 129264
rect 1944 128040 91120 128320
rect 1944 127096 91200 128040
rect 1944 126816 91120 127096
rect 1944 125872 91200 126816
rect 1944 125592 91120 125872
rect 1944 124648 91200 125592
rect 1944 124368 91120 124648
rect 1944 123424 91200 124368
rect 1944 123144 91120 123424
rect 1944 122200 91200 123144
rect 1944 121920 91120 122200
rect 1944 120976 91200 121920
rect 1944 120696 91120 120976
rect 1944 119752 91200 120696
rect 1944 119472 91120 119752
rect 1944 118528 91200 119472
rect 1944 118248 91120 118528
rect 1944 117304 91200 118248
rect 1944 117024 91120 117304
rect 1944 116080 91200 117024
rect 1944 115800 91120 116080
rect 1944 114992 91200 115800
rect 1944 114712 91120 114992
rect 1944 113768 91200 114712
rect 1944 113488 91120 113768
rect 1944 112544 91200 113488
rect 1944 112264 91120 112544
rect 1944 111320 91200 112264
rect 1944 111040 91120 111320
rect 1944 110096 91200 111040
rect 1944 109816 91120 110096
rect 1944 108872 91200 109816
rect 1944 108592 91120 108872
rect 1944 107648 91200 108592
rect 1944 107368 91120 107648
rect 1944 106424 91200 107368
rect 1944 106144 91120 106424
rect 1944 105200 91200 106144
rect 1944 104920 91120 105200
rect 1944 103976 91200 104920
rect 1944 103696 91120 103976
rect 1944 102752 91200 103696
rect 1944 102472 91120 102752
rect 1944 101528 91200 102472
rect 1944 101248 91120 101528
rect 1944 100304 91200 101248
rect 1944 100024 91120 100304
rect 1944 99080 91200 100024
rect 1944 98800 91120 99080
rect 1944 97856 91200 98800
rect 1944 97576 91120 97856
rect 1944 96768 91200 97576
rect 1944 96488 91120 96768
rect 1944 95544 91200 96488
rect 1944 95264 91120 95544
rect 1944 94320 91200 95264
rect 1944 94040 91120 94320
rect 1944 93096 91200 94040
rect 1944 92816 91120 93096
rect 1944 91872 91200 92816
rect 1944 91592 91120 91872
rect 1944 90648 91200 91592
rect 1944 90368 91120 90648
rect 1944 89424 91200 90368
rect 1944 89144 91120 89424
rect 1944 88200 91200 89144
rect 1944 87920 91120 88200
rect 1944 86976 91200 87920
rect 1944 86696 91120 86976
rect 1944 85752 91200 86696
rect 1944 85472 91120 85752
rect 1944 84528 91200 85472
rect 1944 84248 91120 84528
rect 1944 83304 91200 84248
rect 1944 83024 91120 83304
rect 1944 82080 91200 83024
rect 1944 81800 91120 82080
rect 1944 80856 91200 81800
rect 1944 80576 91120 80856
rect 1944 79632 91200 80576
rect 1944 79352 91120 79632
rect 1944 78408 91200 79352
rect 1944 78128 91120 78408
rect 1944 77320 91200 78128
rect 1944 77040 91120 77320
rect 1944 76096 91200 77040
rect 1944 75816 91120 76096
rect 1944 74872 91200 75816
rect 1944 74592 91120 74872
rect 1944 73648 91200 74592
rect 1944 73368 91120 73648
rect 1944 72424 91200 73368
rect 1944 72144 91120 72424
rect 1944 71200 91200 72144
rect 1944 70920 91120 71200
rect 1944 69976 91200 70920
rect 1944 69696 91120 69976
rect 1944 68752 91200 69696
rect 1944 68472 91120 68752
rect 1944 67528 91200 68472
rect 1944 67248 91120 67528
rect 1944 66304 91200 67248
rect 1944 66024 91120 66304
rect 1944 65080 91200 66024
rect 1944 64800 91120 65080
rect 1944 63856 91200 64800
rect 1944 63576 91120 63856
rect 1944 62632 91200 63576
rect 1944 62352 91120 62632
rect 1944 61408 91200 62352
rect 1944 61128 91120 61408
rect 1944 60184 91200 61128
rect 1944 59904 91120 60184
rect 1944 58960 91200 59904
rect 1944 58680 91120 58960
rect 1944 57872 91200 58680
rect 1944 57592 91120 57872
rect 1944 56648 91200 57592
rect 1944 56368 91120 56648
rect 1944 55424 91200 56368
rect 1944 55144 91120 55424
rect 1944 54200 91200 55144
rect 1944 53920 91120 54200
rect 1944 52976 91200 53920
rect 1944 52696 91120 52976
rect 1944 51752 91200 52696
rect 1944 51472 91120 51752
rect 1944 50528 91200 51472
rect 1944 50248 91120 50528
rect 1944 49304 91200 50248
rect 1944 49024 91120 49304
rect 1944 48080 91200 49024
rect 1944 47800 91120 48080
rect 1944 46856 91200 47800
rect 1944 46576 91120 46856
rect 1944 45632 91200 46576
rect 1944 45352 91120 45632
rect 1944 44408 91200 45352
rect 1944 44128 91120 44408
rect 1944 43184 91200 44128
rect 1944 42904 91120 43184
rect 1944 41960 91200 42904
rect 1944 41680 91120 41960
rect 1944 40736 91200 41680
rect 1944 40456 91120 40736
rect 1944 39512 91200 40456
rect 1944 39232 91120 39512
rect 1944 38424 91200 39232
rect 1944 38144 91120 38424
rect 1944 37200 91200 38144
rect 1944 36920 91120 37200
rect 1944 35976 91200 36920
rect 1944 35696 91120 35976
rect 1944 34752 91200 35696
rect 1944 34472 91120 34752
rect 1944 33528 91200 34472
rect 1944 33248 91120 33528
rect 1944 32304 91200 33248
rect 1944 32024 91120 32304
rect 1944 31080 91200 32024
rect 1944 30800 91120 31080
rect 1944 29856 91200 30800
rect 1944 29576 91120 29856
rect 1944 28632 91200 29576
rect 1944 28352 91120 28632
rect 1944 27408 91200 28352
rect 1944 27128 91120 27408
rect 1944 26184 91200 27128
rect 1944 25904 91120 26184
rect 1944 24960 91200 25904
rect 1944 24680 91120 24960
rect 1944 23736 91200 24680
rect 1944 23456 91120 23736
rect 1944 22512 91200 23456
rect 1944 22232 91120 22512
rect 1944 21288 91200 22232
rect 1944 21008 91120 21288
rect 1944 20064 91200 21008
rect 1944 19784 91120 20064
rect 1944 18976 91200 19784
rect 1944 18696 91120 18976
rect 1944 17752 91200 18696
rect 1944 17472 91120 17752
rect 1944 16528 91200 17472
rect 1944 16248 91120 16528
rect 1944 15304 91200 16248
rect 1944 15024 91120 15304
rect 1944 14080 91200 15024
rect 1944 13800 91120 14080
rect 1944 12856 91200 13800
rect 1944 12576 91120 12856
rect 1944 11632 91200 12576
rect 1944 11352 91120 11632
rect 1944 10408 91200 11352
rect 1944 10128 91120 10408
rect 1944 9184 91200 10128
rect 1944 8904 91120 9184
rect 1944 7960 91200 8904
rect 1944 7680 91120 7960
rect 1944 6736 91200 7680
rect 1944 6456 91120 6736
rect 1944 5512 91200 6456
rect 1944 5232 91120 5512
rect 1944 4288 91200 5232
rect 1944 4008 91120 4288
rect 1944 3064 91200 4008
rect 1944 2784 91120 3064
rect 1944 1840 91200 2784
rect 1944 1560 91120 1840
rect 1944 752 91200 1560
rect 1944 472 91120 752
rect 1944 171 91200 472
<< metal4 >>
rect 1944 2128 2264 189360
rect 3944 2128 4264 189360
rect 85944 2128 86264 189360
rect 87944 2128 88264 189360
rect 89944 2128 90264 189360
<< obsm4 >>
rect 4390 189440 90738 191453
rect 4390 2048 85864 189440
rect 86344 2048 87864 189440
rect 88344 2048 89864 189440
rect 90344 2048 90738 189440
rect 4390 171 90738 2048
<< metal5 >>
rect 1104 185298 90896 185618
rect 1104 180298 90896 180618
rect 1104 175298 90896 175618
rect 1104 170298 90896 170618
rect 1104 165298 90896 165618
rect 1104 160298 90896 160618
rect 1104 155298 90896 155618
rect 1104 150298 90896 150618
rect 1104 145298 90896 145618
rect 1104 140298 90896 140618
rect 1104 135298 90896 135618
rect 1104 130298 90896 130618
rect 1104 125298 90896 125618
rect 1104 120298 90896 120618
rect 1104 115298 90896 115618
rect 1104 110298 90896 110618
rect 1104 105298 90896 105618
rect 1104 100298 90896 100618
rect 1104 95298 90896 95618
rect 1104 90298 90896 90618
rect 1104 85298 90896 85618
rect 1104 80298 90896 80618
rect 1104 75298 90896 75618
rect 1104 70298 90896 70618
rect 1104 65298 90896 65618
rect 1104 60298 90896 60618
rect 1104 55298 90896 55618
rect 1104 50298 90896 50618
rect 1104 45298 90896 45618
rect 1104 40298 90896 40618
rect 1104 35298 90896 35618
rect 1104 30298 90896 30618
rect 1104 25298 90896 25618
rect 1104 20298 90896 20618
rect 1104 15298 90896 15618
rect 1104 10298 90896 10618
rect 1104 5298 90896 5618
<< obsm5 >>
rect 4348 125938 90780 126300
rect 4348 120938 90780 124978
rect 4348 115938 90780 119978
rect 4348 110938 90780 114978
rect 4348 105938 90780 109978
rect 4348 100938 90780 104978
rect 4348 95938 90780 99978
rect 4348 90938 90780 94978
rect 4348 85938 90780 89978
rect 4348 80938 90780 84978
rect 4348 75938 90780 79978
rect 4348 70938 90780 74978
rect 4348 65938 90780 69978
rect 4348 60938 90780 64978
rect 4348 55938 90780 59978
rect 4348 50938 90780 54978
rect 4348 45938 90780 49978
rect 4348 40938 90780 44978
rect 4348 35938 90780 39978
rect 4348 30938 90780 34978
rect 4348 25938 90780 29978
rect 4348 20938 90780 24978
rect 4348 15938 90780 19978
rect 4348 10938 90780 14978
rect 4348 5938 90780 9978
rect 4348 2220 90780 4978
<< labels >>
rlabel metal3 s 91200 88000 92000 88120 6 mgmt_addr[0]
port 1 nsew signal input
rlabel metal3 s 91200 89224 92000 89344 6 mgmt_addr[1]
port 2 nsew signal input
rlabel metal3 s 91200 90448 92000 90568 6 mgmt_addr[2]
port 3 nsew signal input
rlabel metal3 s 91200 91672 92000 91792 6 mgmt_addr[3]
port 4 nsew signal input
rlabel metal3 s 91200 92896 92000 93016 6 mgmt_addr[4]
port 5 nsew signal input
rlabel metal3 s 91200 94120 92000 94240 6 mgmt_addr[5]
port 6 nsew signal input
rlabel metal3 s 91200 95344 92000 95464 6 mgmt_addr[6]
port 7 nsew signal input
rlabel metal3 s 91200 96568 92000 96688 6 mgmt_addr[7]
port 8 nsew signal input
rlabel metal3 s 91200 97656 92000 97776 6 mgmt_addr_ro[0]
port 9 nsew signal input
rlabel metal3 s 91200 98880 92000 99000 6 mgmt_addr_ro[1]
port 10 nsew signal input
rlabel metal3 s 91200 100104 92000 100224 6 mgmt_addr_ro[2]
port 11 nsew signal input
rlabel metal3 s 91200 101328 92000 101448 6 mgmt_addr_ro[3]
port 12 nsew signal input
rlabel metal3 s 91200 102552 92000 102672 6 mgmt_addr_ro[4]
port 13 nsew signal input
rlabel metal3 s 91200 103776 92000 103896 6 mgmt_addr_ro[5]
port 14 nsew signal input
rlabel metal3 s 91200 105000 92000 105120 6 mgmt_addr_ro[6]
port 15 nsew signal input
rlabel metal3 s 91200 106224 92000 106344 6 mgmt_addr_ro[7]
port 16 nsew signal input
rlabel metal3 s 91200 86776 92000 86896 6 mgmt_clk
port 17 nsew signal input
rlabel metal3 s 91200 552 92000 672 6 mgmt_ena[0]
port 18 nsew signal input
rlabel metal3 s 91200 146344 92000 146464 6 mgmt_ena[1]
port 19 nsew signal input
rlabel metal3 s 91200 1640 92000 1760 6 mgmt_ena_ro
port 20 nsew signal input
rlabel metal3 s 91200 8984 92000 9104 6 mgmt_rdata[0]
port 21 nsew signal output
rlabel metal3 s 91200 21088 92000 21208 6 mgmt_rdata[10]
port 22 nsew signal output
rlabel metal3 s 91200 22312 92000 22432 6 mgmt_rdata[11]
port 23 nsew signal output
rlabel metal3 s 91200 23536 92000 23656 6 mgmt_rdata[12]
port 24 nsew signal output
rlabel metal3 s 91200 24760 92000 24880 6 mgmt_rdata[13]
port 25 nsew signal output
rlabel metal3 s 91200 25984 92000 26104 6 mgmt_rdata[14]
port 26 nsew signal output
rlabel metal3 s 91200 27208 92000 27328 6 mgmt_rdata[15]
port 27 nsew signal output
rlabel metal3 s 91200 28432 92000 28552 6 mgmt_rdata[16]
port 28 nsew signal output
rlabel metal3 s 91200 29656 92000 29776 6 mgmt_rdata[17]
port 29 nsew signal output
rlabel metal3 s 91200 30880 92000 31000 6 mgmt_rdata[18]
port 30 nsew signal output
rlabel metal3 s 91200 32104 92000 32224 6 mgmt_rdata[19]
port 31 nsew signal output
rlabel metal3 s 91200 10208 92000 10328 6 mgmt_rdata[1]
port 32 nsew signal output
rlabel metal3 s 91200 33328 92000 33448 6 mgmt_rdata[20]
port 33 nsew signal output
rlabel metal3 s 91200 34552 92000 34672 6 mgmt_rdata[21]
port 34 nsew signal output
rlabel metal3 s 91200 35776 92000 35896 6 mgmt_rdata[22]
port 35 nsew signal output
rlabel metal3 s 91200 37000 92000 37120 6 mgmt_rdata[23]
port 36 nsew signal output
rlabel metal3 s 91200 38224 92000 38344 6 mgmt_rdata[24]
port 37 nsew signal output
rlabel metal3 s 91200 39312 92000 39432 6 mgmt_rdata[25]
port 38 nsew signal output
rlabel metal3 s 91200 40536 92000 40656 6 mgmt_rdata[26]
port 39 nsew signal output
rlabel metal3 s 91200 41760 92000 41880 6 mgmt_rdata[27]
port 40 nsew signal output
rlabel metal3 s 91200 42984 92000 43104 6 mgmt_rdata[28]
port 41 nsew signal output
rlabel metal3 s 91200 44208 92000 44328 6 mgmt_rdata[29]
port 42 nsew signal output
rlabel metal3 s 91200 11432 92000 11552 6 mgmt_rdata[2]
port 43 nsew signal output
rlabel metal3 s 91200 45432 92000 45552 6 mgmt_rdata[30]
port 44 nsew signal output
rlabel metal3 s 91200 46656 92000 46776 6 mgmt_rdata[31]
port 45 nsew signal output
rlabel metal3 s 91200 153688 92000 153808 6 mgmt_rdata[32]
port 46 nsew signal output
rlabel metal3 s 91200 154776 92000 154896 6 mgmt_rdata[33]
port 47 nsew signal output
rlabel metal3 s 91200 156000 92000 156120 6 mgmt_rdata[34]
port 48 nsew signal output
rlabel metal3 s 91200 157224 92000 157344 6 mgmt_rdata[35]
port 49 nsew signal output
rlabel metal3 s 91200 158448 92000 158568 6 mgmt_rdata[36]
port 50 nsew signal output
rlabel metal3 s 91200 159672 92000 159792 6 mgmt_rdata[37]
port 51 nsew signal output
rlabel metal3 s 91200 160896 92000 161016 6 mgmt_rdata[38]
port 52 nsew signal output
rlabel metal3 s 91200 162120 92000 162240 6 mgmt_rdata[39]
port 53 nsew signal output
rlabel metal3 s 91200 12656 92000 12776 6 mgmt_rdata[3]
port 54 nsew signal output
rlabel metal3 s 91200 163344 92000 163464 6 mgmt_rdata[40]
port 55 nsew signal output
rlabel metal3 s 91200 164568 92000 164688 6 mgmt_rdata[41]
port 56 nsew signal output
rlabel metal3 s 91200 165792 92000 165912 6 mgmt_rdata[42]
port 57 nsew signal output
rlabel metal3 s 91200 167016 92000 167136 6 mgmt_rdata[43]
port 58 nsew signal output
rlabel metal3 s 91200 168240 92000 168360 6 mgmt_rdata[44]
port 59 nsew signal output
rlabel metal3 s 91200 169464 92000 169584 6 mgmt_rdata[45]
port 60 nsew signal output
rlabel metal3 s 91200 170688 92000 170808 6 mgmt_rdata[46]
port 61 nsew signal output
rlabel metal3 s 91200 171912 92000 172032 6 mgmt_rdata[47]
port 62 nsew signal output
rlabel metal3 s 91200 173136 92000 173256 6 mgmt_rdata[48]
port 63 nsew signal output
rlabel metal3 s 91200 174224 92000 174344 6 mgmt_rdata[49]
port 64 nsew signal output
rlabel metal3 s 91200 13880 92000 14000 6 mgmt_rdata[4]
port 65 nsew signal output
rlabel metal3 s 91200 175448 92000 175568 6 mgmt_rdata[50]
port 66 nsew signal output
rlabel metal3 s 91200 176672 92000 176792 6 mgmt_rdata[51]
port 67 nsew signal output
rlabel metal3 s 91200 177896 92000 178016 6 mgmt_rdata[52]
port 68 nsew signal output
rlabel metal3 s 91200 179120 92000 179240 6 mgmt_rdata[53]
port 69 nsew signal output
rlabel metal3 s 91200 180344 92000 180464 6 mgmt_rdata[54]
port 70 nsew signal output
rlabel metal3 s 91200 181568 92000 181688 6 mgmt_rdata[55]
port 71 nsew signal output
rlabel metal3 s 91200 182792 92000 182912 6 mgmt_rdata[56]
port 72 nsew signal output
rlabel metal3 s 91200 184016 92000 184136 6 mgmt_rdata[57]
port 73 nsew signal output
rlabel metal3 s 91200 185240 92000 185360 6 mgmt_rdata[58]
port 74 nsew signal output
rlabel metal3 s 91200 186464 92000 186584 6 mgmt_rdata[59]
port 75 nsew signal output
rlabel metal3 s 91200 15104 92000 15224 6 mgmt_rdata[5]
port 76 nsew signal output
rlabel metal3 s 91200 187688 92000 187808 6 mgmt_rdata[60]
port 77 nsew signal output
rlabel metal3 s 91200 188912 92000 189032 6 mgmt_rdata[61]
port 78 nsew signal output
rlabel metal3 s 91200 190136 92000 190256 6 mgmt_rdata[62]
port 79 nsew signal output
rlabel metal3 s 91200 191360 92000 191480 6 mgmt_rdata[63]
port 80 nsew signal output
rlabel metal3 s 91200 16328 92000 16448 6 mgmt_rdata[6]
port 81 nsew signal output
rlabel metal3 s 91200 17552 92000 17672 6 mgmt_rdata[7]
port 82 nsew signal output
rlabel metal3 s 91200 18776 92000 18896 6 mgmt_rdata[8]
port 83 nsew signal output
rlabel metal3 s 91200 19864 92000 19984 6 mgmt_rdata[9]
port 84 nsew signal output
rlabel metal3 s 91200 47880 92000 48000 6 mgmt_rdata_ro[0]
port 85 nsew signal output
rlabel metal3 s 91200 59984 92000 60104 6 mgmt_rdata_ro[10]
port 86 nsew signal output
rlabel metal3 s 91200 61208 92000 61328 6 mgmt_rdata_ro[11]
port 87 nsew signal output
rlabel metal3 s 91200 62432 92000 62552 6 mgmt_rdata_ro[12]
port 88 nsew signal output
rlabel metal3 s 91200 63656 92000 63776 6 mgmt_rdata_ro[13]
port 89 nsew signal output
rlabel metal3 s 91200 64880 92000 65000 6 mgmt_rdata_ro[14]
port 90 nsew signal output
rlabel metal3 s 91200 66104 92000 66224 6 mgmt_rdata_ro[15]
port 91 nsew signal output
rlabel metal3 s 91200 67328 92000 67448 6 mgmt_rdata_ro[16]
port 92 nsew signal output
rlabel metal3 s 91200 68552 92000 68672 6 mgmt_rdata_ro[17]
port 93 nsew signal output
rlabel metal3 s 91200 69776 92000 69896 6 mgmt_rdata_ro[18]
port 94 nsew signal output
rlabel metal3 s 91200 71000 92000 71120 6 mgmt_rdata_ro[19]
port 95 nsew signal output
rlabel metal3 s 91200 49104 92000 49224 6 mgmt_rdata_ro[1]
port 96 nsew signal output
rlabel metal3 s 91200 72224 92000 72344 6 mgmt_rdata_ro[20]
port 97 nsew signal output
rlabel metal3 s 91200 73448 92000 73568 6 mgmt_rdata_ro[21]
port 98 nsew signal output
rlabel metal3 s 91200 74672 92000 74792 6 mgmt_rdata_ro[22]
port 99 nsew signal output
rlabel metal3 s 91200 75896 92000 76016 6 mgmt_rdata_ro[23]
port 100 nsew signal output
rlabel metal3 s 91200 77120 92000 77240 6 mgmt_rdata_ro[24]
port 101 nsew signal output
rlabel metal3 s 91200 78208 92000 78328 6 mgmt_rdata_ro[25]
port 102 nsew signal output
rlabel metal3 s 91200 79432 92000 79552 6 mgmt_rdata_ro[26]
port 103 nsew signal output
rlabel metal3 s 91200 80656 92000 80776 6 mgmt_rdata_ro[27]
port 104 nsew signal output
rlabel metal3 s 91200 81880 92000 82000 6 mgmt_rdata_ro[28]
port 105 nsew signal output
rlabel metal3 s 91200 83104 92000 83224 6 mgmt_rdata_ro[29]
port 106 nsew signal output
rlabel metal3 s 91200 50328 92000 50448 6 mgmt_rdata_ro[2]
port 107 nsew signal output
rlabel metal3 s 91200 84328 92000 84448 6 mgmt_rdata_ro[30]
port 108 nsew signal output
rlabel metal3 s 91200 85552 92000 85672 6 mgmt_rdata_ro[31]
port 109 nsew signal output
rlabel metal3 s 91200 51552 92000 51672 6 mgmt_rdata_ro[3]
port 110 nsew signal output
rlabel metal3 s 91200 52776 92000 52896 6 mgmt_rdata_ro[4]
port 111 nsew signal output
rlabel metal3 s 91200 54000 92000 54120 6 mgmt_rdata_ro[5]
port 112 nsew signal output
rlabel metal3 s 91200 55224 92000 55344 6 mgmt_rdata_ro[6]
port 113 nsew signal output
rlabel metal3 s 91200 56448 92000 56568 6 mgmt_rdata_ro[7]
port 114 nsew signal output
rlabel metal3 s 91200 57672 92000 57792 6 mgmt_rdata_ro[8]
port 115 nsew signal output
rlabel metal3 s 91200 58760 92000 58880 6 mgmt_rdata_ro[9]
port 116 nsew signal output
rlabel metal3 s 91200 107448 92000 107568 6 mgmt_wdata[0]
port 117 nsew signal input
rlabel metal3 s 91200 119552 92000 119672 6 mgmt_wdata[10]
port 118 nsew signal input
rlabel metal3 s 91200 120776 92000 120896 6 mgmt_wdata[11]
port 119 nsew signal input
rlabel metal3 s 91200 122000 92000 122120 6 mgmt_wdata[12]
port 120 nsew signal input
rlabel metal3 s 91200 123224 92000 123344 6 mgmt_wdata[13]
port 121 nsew signal input
rlabel metal3 s 91200 124448 92000 124568 6 mgmt_wdata[14]
port 122 nsew signal input
rlabel metal3 s 91200 125672 92000 125792 6 mgmt_wdata[15]
port 123 nsew signal input
rlabel metal3 s 91200 126896 92000 127016 6 mgmt_wdata[16]
port 124 nsew signal input
rlabel metal3 s 91200 128120 92000 128240 6 mgmt_wdata[17]
port 125 nsew signal input
rlabel metal3 s 91200 129344 92000 129464 6 mgmt_wdata[18]
port 126 nsew signal input
rlabel metal3 s 91200 130568 92000 130688 6 mgmt_wdata[19]
port 127 nsew signal input
rlabel metal3 s 91200 108672 92000 108792 6 mgmt_wdata[1]
port 128 nsew signal input
rlabel metal3 s 91200 131792 92000 131912 6 mgmt_wdata[20]
port 129 nsew signal input
rlabel metal3 s 91200 133016 92000 133136 6 mgmt_wdata[21]
port 130 nsew signal input
rlabel metal3 s 91200 134240 92000 134360 6 mgmt_wdata[22]
port 131 nsew signal input
rlabel metal3 s 91200 135328 92000 135448 6 mgmt_wdata[23]
port 132 nsew signal input
rlabel metal3 s 91200 136552 92000 136672 6 mgmt_wdata[24]
port 133 nsew signal input
rlabel metal3 s 91200 137776 92000 137896 6 mgmt_wdata[25]
port 134 nsew signal input
rlabel metal3 s 91200 139000 92000 139120 6 mgmt_wdata[26]
port 135 nsew signal input
rlabel metal3 s 91200 140224 92000 140344 6 mgmt_wdata[27]
port 136 nsew signal input
rlabel metal3 s 91200 141448 92000 141568 6 mgmt_wdata[28]
port 137 nsew signal input
rlabel metal3 s 91200 142672 92000 142792 6 mgmt_wdata[29]
port 138 nsew signal input
rlabel metal3 s 91200 109896 92000 110016 6 mgmt_wdata[2]
port 139 nsew signal input
rlabel metal3 s 91200 143896 92000 144016 6 mgmt_wdata[30]
port 140 nsew signal input
rlabel metal3 s 91200 145120 92000 145240 6 mgmt_wdata[31]
port 141 nsew signal input
rlabel metal3 s 91200 111120 92000 111240 6 mgmt_wdata[3]
port 142 nsew signal input
rlabel metal3 s 91200 112344 92000 112464 6 mgmt_wdata[4]
port 143 nsew signal input
rlabel metal3 s 91200 113568 92000 113688 6 mgmt_wdata[5]
port 144 nsew signal input
rlabel metal3 s 91200 114792 92000 114912 6 mgmt_wdata[6]
port 145 nsew signal input
rlabel metal3 s 91200 115880 92000 116000 6 mgmt_wdata[7]
port 146 nsew signal input
rlabel metal3 s 91200 117104 92000 117224 6 mgmt_wdata[8]
port 147 nsew signal input
rlabel metal3 s 91200 118328 92000 118448 6 mgmt_wdata[9]
port 148 nsew signal input
rlabel metal3 s 91200 2864 92000 2984 6 mgmt_wen[0]
port 149 nsew signal input
rlabel metal3 s 91200 147568 92000 147688 6 mgmt_wen[1]
port 150 nsew signal input
rlabel metal3 s 91200 4088 92000 4208 6 mgmt_wen_mask[0]
port 151 nsew signal input
rlabel metal3 s 91200 5312 92000 5432 6 mgmt_wen_mask[1]
port 152 nsew signal input
rlabel metal3 s 91200 6536 92000 6656 6 mgmt_wen_mask[2]
port 153 nsew signal input
rlabel metal3 s 91200 7760 92000 7880 6 mgmt_wen_mask[3]
port 154 nsew signal input
rlabel metal3 s 91200 148792 92000 148912 6 mgmt_wen_mask[4]
port 155 nsew signal input
rlabel metal3 s 91200 150016 92000 150136 6 mgmt_wen_mask[5]
port 156 nsew signal input
rlabel metal3 s 91200 151240 92000 151360 6 mgmt_wen_mask[6]
port 157 nsew signal input
rlabel metal3 s 91200 152464 92000 152584 6 mgmt_wen_mask[7]
port 158 nsew signal input
rlabel metal4 s 89944 2128 90264 189360 6 VPWR
port 159 nsew power bidirectional
rlabel metal4 s 85944 2128 86264 189360 6 VPWR
port 160 nsew power bidirectional
rlabel metal4 s 1944 2128 2264 189360 6 VPWR
port 161 nsew power bidirectional
rlabel metal5 s 1104 185298 90896 185618 6 VPWR
port 162 nsew power bidirectional
rlabel metal5 s 1104 175298 90896 175618 6 VPWR
port 163 nsew power bidirectional
rlabel metal5 s 1104 165298 90896 165618 6 VPWR
port 164 nsew power bidirectional
rlabel metal5 s 1104 155298 90896 155618 6 VPWR
port 165 nsew power bidirectional
rlabel metal5 s 1104 145298 90896 145618 6 VPWR
port 166 nsew power bidirectional
rlabel metal5 s 1104 135298 90896 135618 6 VPWR
port 167 nsew power bidirectional
rlabel metal5 s 1104 125298 90896 125618 6 VPWR
port 168 nsew power bidirectional
rlabel metal5 s 1104 115298 90896 115618 6 VPWR
port 169 nsew power bidirectional
rlabel metal5 s 1104 105298 90896 105618 6 VPWR
port 170 nsew power bidirectional
rlabel metal5 s 1104 95298 90896 95618 6 VPWR
port 171 nsew power bidirectional
rlabel metal5 s 1104 85298 90896 85618 6 VPWR
port 172 nsew power bidirectional
rlabel metal5 s 1104 75298 90896 75618 6 VPWR
port 173 nsew power bidirectional
rlabel metal5 s 1104 65298 90896 65618 6 VPWR
port 174 nsew power bidirectional
rlabel metal5 s 1104 55298 90896 55618 6 VPWR
port 175 nsew power bidirectional
rlabel metal5 s 1104 45298 90896 45618 6 VPWR
port 176 nsew power bidirectional
rlabel metal5 s 1104 35298 90896 35618 6 VPWR
port 177 nsew power bidirectional
rlabel metal5 s 1104 25298 90896 25618 6 VPWR
port 178 nsew power bidirectional
rlabel metal5 s 1104 15298 90896 15618 6 VPWR
port 179 nsew power bidirectional
rlabel metal5 s 1104 5298 90896 5618 6 VPWR
port 180 nsew power bidirectional
rlabel metal4 s 87944 2128 88264 189360 6 VGND
port 181 nsew ground bidirectional
rlabel metal4 s 3944 2128 4264 189360 6 VGND
port 182 nsew ground bidirectional
rlabel metal5 s 1104 180298 90896 180618 6 VGND
port 183 nsew ground bidirectional
rlabel metal5 s 1104 170298 90896 170618 6 VGND
port 184 nsew ground bidirectional
rlabel metal5 s 1104 160298 90896 160618 6 VGND
port 185 nsew ground bidirectional
rlabel metal5 s 1104 150298 90896 150618 6 VGND
port 186 nsew ground bidirectional
rlabel metal5 s 1104 140298 90896 140618 6 VGND
port 187 nsew ground bidirectional
rlabel metal5 s 1104 130298 90896 130618 6 VGND
port 188 nsew ground bidirectional
rlabel metal5 s 1104 120298 90896 120618 6 VGND
port 189 nsew ground bidirectional
rlabel metal5 s 1104 110298 90896 110618 6 VGND
port 190 nsew ground bidirectional
rlabel metal5 s 1104 100298 90896 100618 6 VGND
port 191 nsew ground bidirectional
rlabel metal5 s 1104 90298 90896 90618 6 VGND
port 192 nsew ground bidirectional
rlabel metal5 s 1104 80298 90896 80618 6 VGND
port 193 nsew ground bidirectional
rlabel metal5 s 1104 70298 90896 70618 6 VGND
port 194 nsew ground bidirectional
rlabel metal5 s 1104 60298 90896 60618 6 VGND
port 195 nsew ground bidirectional
rlabel metal5 s 1104 50298 90896 50618 6 VGND
port 196 nsew ground bidirectional
rlabel metal5 s 1104 40298 90896 40618 6 VGND
port 197 nsew ground bidirectional
rlabel metal5 s 1104 30298 90896 30618 6 VGND
port 198 nsew ground bidirectional
rlabel metal5 s 1104 20298 90896 20618 6 VGND
port 199 nsew ground bidirectional
rlabel metal5 s 1104 10298 90896 10618 6 VGND
port 200 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 92000 192000
string LEFview TRUE
string GDS_FILE /project/openlane/storage/runs/storage/results/magic/storage.gds
string GDS_END 14864420
string GDS_START 12876356
<< end >>

