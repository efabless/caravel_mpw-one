* SPICE NETLIST
***************************************


***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808687 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 AD=0.98 AS=1.96 PD=7.28 PS=14.56 NRD=0 NRS=0 m=1 sa=90000.2 sb=90004.3 a=1.26 p=14.36
XM1 2 3 4 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=90000.7 sb=90003.9 a=1.26 p=14.36
XM2 4 3 2 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=90001.1 sb=90003.4 a=1.26 p=14.36
XM3 2 3 4 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=90001.6 sb=90002.9 a=1.26 p=14.36
XM4 4 3 2 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=90002 sb=90002.5 a=1.26 p=14.36
XM5 2 3 4 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=90002.5 sb=90002 a=1.26 p=14.36
XM6 4 3 2 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=90002.9 sb=90001.6 a=1.26 p=14.36
XM7 2 3 4 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=90003.4 sb=90001.1 a=1.26 p=14.36
XM8 4 3 2 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=90003.9 sb=90000.7 a=1.26 p=14.36
XM9 2 3 4 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 AD=1.96 AS=0.98 PD=14.56 PS=7.28 NRD=0 NRS=0 m=1 sa=90004.3 sb=90000.2 a=1.26 p=14.36
.ENDS
***************************************

***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808701 2
**
*.SEEDPROM
X0 2 2 sky130_fd_pr__diode_pw2nd_05v5 a=2.1 p=14.6 m=1
X1 2 2 sky130_fd_pr__diode_pw2nd_05v5 a=2.1 p=14.6 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808703 2
**
*.SEEDPROM
X0 2 2 sky130_fd_pr__diode_pw2nd_05v5 a=2.1 p=14.6 m=1
X1 2 2 sky130_fd_pr__diode_pw2nd_05v5 a=2.1 p=14.6 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808705 2
**
*.SEEDPROM
X0 2 2 sky130_fd_pr__diode_pw2nd_05v5 a=2.1 p=14.6 m=1
X1 2 2 sky130_fd_pr__diode_pw2nd_05v5 a=2.1 p=14.6 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808693 1
**
*.SEEDPROM
X0 1 1 sky130_fd_pr__diode_pw2nd_05v5 a=1.5 p=10.6 m=1
X1 1 1 sky130_fd_pr__diode_pw2nd_05v5 a=1.5 p=10.6 m=1
.ENDS
***************************************
.SUBCKT sky130_ef_io__vccd_lvc_clamped2_pad   VSSD VSSIO VCCD VDDIO VSSA VCCHIB VDDA VSWITCH AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
**
XM0 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90001.1 sb=90019.9 a=1.26 p=14.36
XM1 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90001.1 sb=90019.9 a=1.26 p=14.36
XM2 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90001.1 sb=90019.9 a=1.26 p=14.36
XM3 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90001.1 sb=90019.9 a=1.26 p=14.36
XM4 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90001.1 sb=90019.9 a=0.9 p=10.36
XM5 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90001.1 sb=90019.9 a=1.26 p=14.36
XM6 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90002.3 sb=90019.9 a=1.26 p=14.36
XM7 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90002.3 sb=90019.9 a=1.26 p=14.36
XM8 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90002.3 sb=90019.9 a=1.26 p=14.36
XM9 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90002.3 sb=90019.9 a=1.26 p=14.36
XM10 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90002.3 sb=90019.9 a=0.9 p=10.36
XM11 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90002.3 sb=90019.9 a=1.26 p=14.36
XM12 VSSD 9 VSSD VSSD sky130_fd_pr__nfet_01v8 L=4 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=2e+06 sb=2.00002e+06 a=20 p=18
XM13 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90003.9 sb=90019.9 a=1.26 p=14.36
XM14 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90003.9 sb=90019.9 a=1.26 p=14.36
XM15 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90003.9 sb=90019.9 a=1.26 p=14.36
XM16 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90003.9 sb=90019.9 a=1.26 p=14.36
XM17 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90003.9 sb=90019.9 a=0.9 p=10.36
XM18 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90001.1 sb=90019.9 a=1.26 p=14.36
XM19 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90003.9 sb=90019.9 a=1.26 p=14.36
XM20 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90001.7 sb=90019.9 a=1.26 p=14.36
XM21 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90001.7 sb=90019.9 a=1.26 p=14.36
XM22 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90001.7 sb=90019.9 a=1.26 p=14.36
XM23 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90005.1 sb=90019.9 a=1.26 p=14.36
XM24 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90005.1 sb=90019.9 a=1.26 p=14.36
XM25 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90005.1 sb=90019.9 a=1.26 p=14.36
XM26 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90005.1 sb=90019.9 a=1.26 p=14.36
XM27 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90005.1 sb=90019.9 a=0.9 p=10.36
XM28 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90002.3 sb=90019.9 a=1.26 p=14.36
XM29 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90005.1 sb=90019.9 a=1.26 p=14.36
XM30 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90003.1 sb=90019.9 a=1.26 p=14.36
XM31 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90003.1 sb=90019.9 a=1.26 p=14.36
XM32 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90003.1 sb=90019.9 a=1.26 p=14.36
XM33 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90006.6 sb=90019.9 a=1.26 p=14.36
XM34 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90006.6 sb=90019.9 a=1.26 p=14.36
XM35 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90006.6 sb=90019.9 a=1.26 p=14.36
XM36 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90006.6 sb=90019.9 a=1.26 p=14.36
XM37 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90006.6 sb=90019.9 a=0.9 p=10.36
XM38 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90003.9 sb=90019.9 a=1.26 p=14.36
XM39 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90006.6 sb=90019.9 a=1.26 p=14.36
XM40 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90007.8 sb=90019.9 a=1.26 p=14.36
XM41 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90007.8 sb=90019.9 a=1.26 p=14.36
XM42 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90007.8 sb=90019.9 a=1.26 p=14.36
XM43 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90007.8 sb=90019.9 a=1.26 p=14.36
XM44 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90007.8 sb=90019.9 a=0.9 p=10.36
XM45 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90005.1 sb=90019.9 a=1.26 p=14.36
XM46 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90007.8 sb=90019.9 a=1.26 p=14.36
XM47 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90005.9 sb=90019.9 a=1.26 p=14.36
XM48 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90005.9 sb=90019.9 a=1.26 p=14.36
XM49 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90005.9 sb=90019.9 a=1.26 p=14.36
XM50 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90009.4 sb=90019.9 a=1.26 p=14.36
XM51 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90009.4 sb=90019.9 a=1.26 p=14.36
XM52 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90009.4 sb=90019.9 a=1.26 p=14.36
XM53 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90009.4 sb=90019.9 a=1.26 p=14.36
XM54 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90009.4 sb=90019.9 a=0.9 p=10.36
XM55 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90006.6 sb=90019.9 a=1.26 p=14.36
XM56 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90009.4 sb=90019.9 a=1.26 p=14.36
XM57 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90007.3 sb=90019.9 a=1.26 p=14.36
XM58 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90007.3 sb=90019.9 a=1.26 p=14.36
XM59 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90007.3 sb=90019.9 a=1.26 p=14.36
XM60 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90010.6 sb=90019.9 a=1.26 p=14.36
XM61 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90010.6 sb=90019.9 a=1.26 p=14.36
XM62 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90010.6 sb=90019.9 a=1.26 p=14.36
XM63 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90010.6 sb=90019.9 a=1.26 p=14.36
XM64 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90010.6 sb=90019.9 a=0.9 p=10.36
XM65 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90007.8 sb=90019.9 a=1.26 p=14.36
XM66 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90010.6 sb=90019.9 a=1.26 p=14.36
XM67 VSSD 9 11 VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 sa=90000.6 sb=90019.9 a=1.26 p=14.36
XM68 VSSD 9 11 VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 sa=90000.6 sb=90019.9 a=1.26 p=14.36
XM69 VSSIO 5 7 VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 sa=90000.6 sb=90019.9 a=1.26 p=14.36
XM70 VSSIO 5 7 VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 sa=90000.6 sb=90019.9 a=1.26 p=14.36
XM71 VSSIO 5 7 VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 sa=90000.6 sb=90019.9 a=1.26 p=14.36
XM72 VSSD 9 VSSD VSSD sky130_fd_pr__nfet_01v8 L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=4e+06 sb=4.00002e+06 a=40 p=26
XM73 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90012.2 sb=90019.9 a=1.26 p=14.36
XM74 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90012.2 sb=90019.9 a=1.26 p=14.36
XM75 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90012.2 sb=90019.9 a=1.26 p=14.36
XM76 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90012.2 sb=90019.9 a=1.26 p=14.36
XM77 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90012.2 sb=90019.9 a=0.9 p=10.36
XM78 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90009.4 sb=90019.9 a=1.26 p=14.36
XM79 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90012.2 sb=90019.9 a=1.26 p=14.36
XM80 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90001.7 sb=90019.9 a=0.9 p=10.36
XM81 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90001.7 sb=90019.9 a=1.26 p=14.36
XM82 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90010.1 sb=90019.9 a=1.26 p=14.36
XM83 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90010.1 sb=90019.9 a=1.26 p=14.36
XM84 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90010.1 sb=90019.9 a=1.26 p=14.36
XM85 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90013.4 sb=90019.9 a=1.26 p=14.36
XM86 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90013.4 sb=90019.9 a=1.26 p=14.36
XM87 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90013.4 sb=90019.9 a=1.26 p=14.36
XM88 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90013.4 sb=90019.9 a=1.26 p=14.36
XM89 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90013.4 sb=90019.9 a=0.9 p=10.36
XM90 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90010.6 sb=90019.9 a=1.26 p=14.36
XM91 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90013.4 sb=90019.9 a=1.26 p=14.36
XM92 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90003.1 sb=90019.9 a=0.9 p=10.36
XM93 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90003.1 sb=90019.9 a=1.26 p=14.36
XM94 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90011.4 sb=90019.9 a=1.26 p=14.36
XM95 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90011.4 sb=90019.9 a=1.26 p=14.36
XM96 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90011.4 sb=90019.9 a=1.26 p=14.36
XM97 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90015 sb=90019.9 a=1.26 p=14.36
XM98 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90015 sb=90019.9 a=1.26 p=14.36
XM99 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90015 sb=90019.9 a=1.26 p=14.36
XM100 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90015 sb=90019.9 a=1.26 p=14.36
XM101 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90015 sb=90019.9 a=0.9 p=10.36
XM102 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90012.2 sb=90019.9 a=1.26 p=14.36
XM103 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90015 sb=90019.9 a=1.26 p=14.36
XM104 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90016.2 sb=90019.9 a=1.26 p=14.36
XM105 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90016.2 sb=90019.9 a=1.26 p=14.36
XM106 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90016.2 sb=90019.9 a=1.26 p=14.36
XM107 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90016.2 sb=90019.9 a=1.26 p=14.36
XM108 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90016.1 sb=90019.9 a=0.9 p=10.36
XM109 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90013.4 sb=90019.9 a=1.26 p=14.36
XM110 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90016.2 sb=90019.9 a=1.26 p=14.36
XM111 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90005.9 sb=90019.9 a=0.9 p=10.36
XM112 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90005.9 sb=90019.9 a=1.26 p=14.36
XM113 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90014.3 sb=90019.9 a=1.26 p=14.36
XM114 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90014.3 sb=90019.9 a=1.26 p=14.36
XM115 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90014.3 sb=90019.9 a=1.26 p=14.36
XM116 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90017.7 sb=90019.9 a=1.26 p=14.36
XM117 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90017.7 sb=90019.9 a=1.26 p=14.36
XM118 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90017.7 sb=90019.9 a=1.26 p=14.36
XM119 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90017.7 sb=90019.9 a=1.26 p=14.36
XM120 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90017.7 sb=90019.9 a=0.9 p=10.36
XM121 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90015 sb=90019.9 a=1.26 p=14.36
XM122 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90017.7 sb=90019.9 a=1.26 p=14.36
XM123 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90007.3 sb=90019.9 a=0.9 p=10.36
XM124 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90007.3 sb=90019.9 a=1.26 p=14.36
XM125 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90015.6 sb=90019.9 a=1.26 p=14.36
XM126 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90015.6 sb=90019.9 a=1.26 p=14.36
XM127 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90015.6 sb=90019.9 a=1.26 p=14.36
XM128 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90018.9 sb=90019.9 a=1.26 p=14.36
XM129 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90018.9 sb=90019.9 a=1.26 p=14.36
XM130 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90018.9 sb=90019.9 a=1.26 p=14.36
XM131 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90018.9 sb=90019.9 a=1.26 p=14.36
XM132 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90018.9 sb=90019.9 a=0.9 p=10.36
XM133 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90016.2 sb=90019.9 a=1.26 p=14.36
XM134 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90018.9 sb=90019.9 a=1.26 p=14.36
XM135 VSSD 9 VSSD VSSD sky130_fd_pr__nfet_01v8 L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00002e+06 a=40 p=26
XM136 VSSD 9 VSSD VSSD sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 sa=4e+06 sb=4.00002e+06 a=56 p=30
XM137 VSSD 9 VSSD VSSD sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 sa=4e+06 sb=4.00002e+06 a=56 p=30
XM138 VSSIO 5 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 sa=4e+06 sb=4.00002e+06 a=56 p=30
XM139 VSSIO 5 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 sa=4e+06 sb=4.00002e+06 a=56 p=30
XM140 VSSIO 5 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 sa=4e+06 sb=4.00002e+06 a=56 p=30
XM141 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM142 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM143 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM144 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM145 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM146 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90017.7 sb=90019.9 a=1.26 p=14.36
XM147 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM148 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90010.1 sb=90019.9 a=0.9 p=10.36
XM149 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90010.1 sb=90019.9 a=1.26 p=14.36
XM150 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90018.5 sb=90019.9 a=1.26 p=14.36
XM151 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90018.5 sb=90019.9 a=1.26 p=14.36
XM152 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90018.5 sb=90019.9 a=1.26 p=14.36
XM153 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM154 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM155 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM156 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM157 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM158 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90018.9 sb=90019.9 a=1.26 p=14.36
XM159 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM160 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90011.4 sb=90019.9 a=0.9 p=10.36
XM161 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90011.4 sb=90019.9 a=1.26 p=14.36
XM162 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.8 sb=90019.9 a=1.26 p=14.36
XM163 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.8 sb=90019.9 a=1.26 p=14.36
XM164 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.8 sb=90019.9 a=1.26 p=14.36
XM165 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM166 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM167 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM168 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM169 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM170 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM171 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM172 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM173 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM174 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM175 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM176 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM177 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM178 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM179 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90014.3 sb=90019.9 a=0.9 p=10.36
XM180 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90014.3 sb=90019.9 a=1.26 p=14.36
XM181 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM182 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM183 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM184 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM185 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM186 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM187 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM188 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM189 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM190 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM191 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90015.6 sb=90019.9 a=0.9 p=10.36
XM192 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90015.6 sb=90019.9 a=1.26 p=14.36
XM193 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM194 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM195 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM196 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM197 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM198 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM199 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM200 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM201 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM202 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM203 VSSD 9 VSSD VSSD sky130_fd_pr__nfet_01v8 L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4.00002e+06 a=40 p=26
XM204 VSSD 9 VSSD VSSD sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30
XM205 VSSD 9 VSSD VSSD sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30
XM206 VSSIO 5 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30
XM207 VSSIO 5 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30
XM208 VSSIO 5 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30
XM209 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM210 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM211 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM212 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM213 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM214 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM215 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM216 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90018.5 sb=90019.9 a=0.9 p=10.36
XM217 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90018.5 sb=90019.9 a=1.26 p=14.36
XM218 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM219 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM220 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM221 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM222 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM223 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM224 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM225 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM226 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM227 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM228 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90019.8 sb=90019.9 a=0.9 p=10.36
XM229 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.8 sb=90019.9 a=1.26 p=14.36
XM230 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM231 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM232 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM233 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM234 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM235 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM236 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM237 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM238 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM239 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM240 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM241 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM242 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM243 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM244 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM245 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM246 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM247 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90019.9 sb=90019.8 a=0.9 p=10.36
XM248 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.8 a=1.26 p=14.36
XM249 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.8 a=1.26 p=14.36
XM250 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.8 a=1.26 p=14.36
XM251 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.8 a=1.26 p=14.36
XM252 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90018.9 a=1.26 p=14.36
XM253 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90018.9 a=1.26 p=14.36
XM254 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90018.9 a=1.26 p=14.36
XM255 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90018.9 a=1.26 p=14.36
XM256 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90018.9 a=0.9 p=10.36
XM257 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90018.9 a=1.26 p=14.36
XM258 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90018.9 a=1.26 p=14.36
XM259 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90019.9 sb=90018.5 a=0.9 p=10.36
XM260 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90018.5 a=1.26 p=14.36
XM261 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90018.5 a=1.26 p=14.36
XM262 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90018.5 a=1.26 p=14.36
XM263 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90018.5 a=1.26 p=14.36
XM264 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90017.7 a=1.26 p=14.36
XM265 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90017.7 a=1.26 p=14.36
XM266 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90017.7 a=1.26 p=14.36
XM267 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90017.7 a=1.26 p=14.36
XM268 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90017.7 a=0.9 p=10.36
XM269 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90017.7 a=1.26 p=14.36
XM270 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90017.7 a=1.26 p=14.36
XM271 VSSD 9 VSSD VSSD sky130_fd_pr__nfet_01v8 L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4.00001e+06 a=40 p=26
XM272 VSSD 9 VSSD VSSD sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30
XM273 VSSD 9 VSSD VSSD sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30
XM274 VSSIO 5 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30
XM275 VSSIO 5 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30
XM276 VSSIO 5 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30
XM277 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90016.2 a=1.26 p=14.36
XM278 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90016.2 a=1.26 p=14.36
XM279 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90016.2 a=1.26 p=14.36
XM280 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90016.2 a=1.26 p=14.36
XM281 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90016.1 a=0.9 p=10.36
XM282 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90016.2 a=1.26 p=14.36
XM283 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90016.2 a=1.26 p=14.36
XM284 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90019.9 sb=90015.6 a=0.9 p=10.36
XM285 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90015.6 a=1.26 p=14.36
XM286 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90015.6 a=1.26 p=14.36
XM287 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90015.6 a=1.26 p=14.36
XM288 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90015.6 a=1.26 p=14.36
XM289 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90015 a=1.26 p=14.36
XM290 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90015 a=1.26 p=14.36
XM291 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90015 a=1.26 p=14.36
XM292 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90015 a=1.26 p=14.36
XM293 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90015 a=0.9 p=10.36
XM294 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90015 a=1.26 p=14.36
XM295 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90015 a=1.26 p=14.36
XM296 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90019.9 sb=90014.3 a=0.9 p=10.36
XM297 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90014.3 a=1.26 p=14.36
XM298 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90014.3 a=1.26 p=14.36
XM299 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90014.3 a=1.26 p=14.36
XM300 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90014.3 a=1.26 p=14.36
XM301 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90013.4 a=1.26 p=14.36
XM302 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90013.4 a=1.26 p=14.36
XM303 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90013.4 a=1.26 p=14.36
XM304 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90013.4 a=1.26 p=14.36
XM305 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90013.4 a=0.9 p=10.36
XM306 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90013.4 a=1.26 p=14.36
XM307 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90013.4 a=1.26 p=14.36
XM308 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90012.2 a=1.26 p=14.36
XM309 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90012.2 a=1.26 p=14.36
XM310 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90012.2 a=1.26 p=14.36
XM311 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90012.2 a=1.26 p=14.36
XM312 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90012.2 a=0.9 p=10.36
XM313 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90012.2 a=1.26 p=14.36
XM314 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90012.2 a=1.26 p=14.36
XM315 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90019.9 sb=90011.4 a=0.9 p=10.36
XM316 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90011.4 a=1.26 p=14.36
XM317 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90011.4 a=1.26 p=14.36
XM318 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90011.4 a=1.26 p=14.36
XM319 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90011.4 a=1.26 p=14.36
XM320 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90010.6 a=1.26 p=14.36
XM321 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90010.6 a=1.26 p=14.36
XM322 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90010.6 a=1.26 p=14.36
XM323 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90010.6 a=1.26 p=14.36
XM324 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90010.6 a=0.9 p=10.36
XM325 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90010.6 a=1.26 p=14.36
XM326 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90010.6 a=1.26 p=14.36
XM327 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90019.9 sb=90010.1 a=0.9 p=10.36
XM328 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90010.1 a=1.26 p=14.36
XM329 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90010.1 a=1.26 p=14.36
XM330 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90010.1 a=1.26 p=14.36
XM331 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90010.1 a=1.26 p=14.36
XM332 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90009.4 a=1.26 p=14.36
XM333 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90009.4 a=1.26 p=14.36
XM334 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90009.4 a=1.26 p=14.36
XM335 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90009.4 a=1.26 p=14.36
XM336 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90009.4 a=0.9 p=10.36
XM337 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90009.4 a=1.26 p=14.36
XM338 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90009.4 a=1.26 p=14.36
XM339 VSSD 9 VSSD VSSD sky130_fd_pr__nfet_01v8 L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=40 p=26
XM340 VSSD 9 VSSD VSSD sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM341 VSSD 9 VSSD VSSD sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM342 VSSIO 5 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM343 VSSIO 5 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM344 VSSIO 5 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM345 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90007.8 a=1.26 p=14.36
XM346 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90007.8 a=1.26 p=14.36
XM347 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90007.8 a=1.26 p=14.36
XM348 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90007.8 a=1.26 p=14.36
XM349 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90007.8 a=0.9 p=10.36
XM350 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90007.8 a=1.26 p=14.36
XM351 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90007.8 a=1.26 p=14.36
XM352 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90019.9 sb=90007.3 a=0.9 p=10.36
XM353 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90007.3 a=1.26 p=14.36
XM354 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90007.3 a=1.26 p=14.36
XM355 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90007.3 a=1.26 p=14.36
XM356 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90007.3 a=1.26 p=14.36
XM357 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90006.6 a=1.26 p=14.36
XM358 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90006.6 a=1.26 p=14.36
XM359 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90006.6 a=1.26 p=14.36
XM360 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90006.6 a=1.26 p=14.36
XM361 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90006.6 a=0.9 p=10.36
XM362 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90006.6 a=1.26 p=14.36
XM363 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90006.6 a=1.26 p=14.36
XM364 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90019.9 sb=90005.9 a=0.9 p=10.36
XM365 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90005.9 a=1.26 p=14.36
XM366 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90005.9 a=1.26 p=14.36
XM367 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90005.9 a=1.26 p=14.36
XM368 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90005.9 a=1.26 p=14.36
XM369 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90005.1 a=1.26 p=14.36
XM370 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90005.1 a=1.26 p=14.36
XM371 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90005.1 a=1.26 p=14.36
XM372 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90005.1 a=1.26 p=14.36
XM373 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90005.1 a=0.9 p=10.36
XM374 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90005.1 a=1.26 p=14.36
XM375 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90005.1 a=1.26 p=14.36
XM376 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90003.9 a=1.26 p=14.36
XM377 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90003.9 a=1.26 p=14.36
XM378 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90003.9 a=1.26 p=14.36
XM379 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90003.9 a=1.26 p=14.36
XM380 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90003.9 a=0.9 p=10.36
XM381 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90003.9 a=1.26 p=14.36
XM382 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90003.9 a=1.26 p=14.36
XM383 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90019.9 sb=90003.1 a=0.9 p=10.36
XM384 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90003.1 a=1.26 p=14.36
XM385 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90003.1 a=1.26 p=14.36
XM386 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90003.1 a=1.26 p=14.36
XM387 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90003.1 a=1.26 p=14.36
XM388 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90002.3 a=1.26 p=14.36
XM389 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90002.3 a=1.26 p=14.36
XM390 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90002.3 a=1.26 p=14.36
XM391 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90002.3 a=1.26 p=14.36
XM392 VCCD 11 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90002.3 a=0.9 p=10.36
XM393 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90002.3 a=1.26 p=14.36
XM394 VCCD 7 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90002.3 a=1.26 p=14.36
XM395 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90019.9 sb=90001.7 a=0.9 p=10.36
XM396 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90001.7 a=1.26 p=14.36
XM397 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90001.7 a=1.26 p=14.36
XM398 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90001.7 a=1.26 p=14.36
XM399 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90001.7 a=1.26 p=14.36
XM400 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90001.1 a=1.26 p=14.36
XM401 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90001.1 a=1.26 p=14.36
XM402 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90001.1 a=1.26 p=14.36
XM403 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90001.1 a=1.26 p=14.36
XM404 VSSD 11 VCCD VSSD sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90001.1 a=0.9 p=10.36
XM405 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90001.1 a=1.26 p=14.36
XM406 VSSIO 7 VCCD VSSIO sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90001.1 a=1.26 p=14.36
XM407 VSSD 9 VSSD VSSD sky130_fd_pr__nfet_01v8 L=8 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=40 p=26
XM408 VSSD 9 VSSD VSSD sky130_fd_pr__nfet_01v8 L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM409 VSSD 9 VSSD VSSD sky130_fd_pr__nfet_01v8 L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM410 VSSIO 5 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM411 VSSIO 5 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM412 VSSIO 5 VSSIO VSSIO sky130_fd_pr__nfet_01v8 L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
X413 VSSIO VDDIO condiode a=1e-06 p=0.004 m=1
X414 VSSD VDDIO condiode a=1e-06 p=0.004 m=1
X415 VSSIO VDDIO condiode a=1e-06 p=0.004 m=1
XD416 VSSIO VSSA sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
XD417 VSSIO VSSA sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
XD418 VSSIO VSSA sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
XD419 VSSIO VSSA sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
XD420 VSSA VSSIO sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
XD421 VSSA VSSIO sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
XD422 VSSA VSSIO sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
XD423 VSSA VSSIO sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
X424 VSSIO VSSIO sky130_fd_pr__diode_pw2nd_05v5 a=1.5 p=10.6 m=1
X425 VSSIO VSSIO sky130_fd_pr__diode_pw2nd_05v5 a=2.1 p=14.6 m=1
X426 VSSIO VSSIO sky130_fd_pr__diode_pw2nd_05v5 a=1.5 p=10.6 m=1
X427 VSSIO VSSIO sky130_fd_pr__diode_pw2nd_05v5 a=2.1 p=14.6 m=1
X428 VSSD VCCD sky130_fd_pr__model__parasitic__diode_ps2nw a=108.41 p=46.58 m=1
X429 VSSD VCCD sky130_fd_pr__model__parasitic__diode_ps2nw a=108.41 p=46.58 m=1
X430 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2dn a=10516.3 p=468.87 m=1
X431 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn a=4115.42 p=264.63 m=1
X432 VSSIO VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn a=5703.29 p=340.89 m=1
R433 VCCD 5 sky130_fd_pr__res_generic_po L=1950 W=0.33 m=1
R434 8 6 sky130_fd_pr__res_generic_po L=720 W=0.33 m=1
R435 8 9 sky130_fd_pr__res_generic_po L=200 W=0.33 m=1
R436 10 6 sky130_fd_pr__res_generic_po L=300 W=0.33 m=1
R437 10 VCCD sky130_fd_pr__res_generic_po L=900 W=0.33 m=1
R438 VCCD VCCD 0.01 short m=1
X439 VCCD 5 7 sky130_fd_pr__pfet_01v8__example_55959141808687
X440 VCCD 5 7 sky130_fd_pr__pfet_01v8__example_55959141808687
X441 VCCD 9 11 sky130_fd_pr__pfet_01v8__example_55959141808687
X442 VCCD 9 11 sky130_fd_pr__pfet_01v8__example_55959141808687
X662 VSSD VSSA sky130_fd_io__gnd2gnd_sub_dnwl
X663 VSSD VSSIO sky130_fd_io__gnd2gnd_sub_dnwl
X674 VSSIO sky130_fd_pr__nfet_01v8__example_55959141808701
X675 VSSIO sky130_fd_pr__nfet_01v8__example_55959141808703
X676 VSSIO sky130_fd_pr__nfet_01v8__example_55959141808703
X677 VSSIO sky130_fd_pr__nfet_01v8__example_55959141808703
X678 VSSD sky130_fd_pr__nfet_01v8__example_55959141808705
X679 VSSD sky130_fd_pr__nfet_01v8__example_55959141808705
X680 VSSD sky130_fd_pr__nfet_01v8__example_55959141808705
X681 VSSD sky130_fd_pr__nfet_01v8__example_55959141808705
X682 VSSIO sky130_fd_pr__nfet_01v8__example_55959141808705
X683 VSSD sky130_fd_pr__nfet_01v8__example_55959141808693
.ENDS
***************************************
