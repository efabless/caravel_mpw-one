magic
tech sky130A
timestamp 1606942031
<< metal2 >>
rect 4043 351760 4099 352480
rect 12139 351760 12195 352480
rect 20235 351760 20291 352480
rect 28377 351760 28433 352480
rect 36473 351760 36529 352480
rect 44569 351760 44625 352480
rect 52711 351760 52767 352480
rect 60807 351760 60863 352480
rect 68903 351760 68959 352480
rect 77045 351760 77101 352480
rect 85141 351760 85197 352480
rect 93237 351760 93293 352480
rect 101379 351760 101435 352480
rect 109475 351760 109531 352480
rect 117571 351760 117627 352480
rect 125713 351760 125769 352480
rect 133809 351760 133865 352480
rect 141905 351760 141961 352480
rect 150047 351760 150103 352480
rect 158143 351760 158199 352480
rect 166239 351760 166295 352480
rect 174381 351760 174437 352480
rect 182477 351760 182533 352480
rect 190573 351760 190629 352480
rect 198715 351760 198771 352480
rect 206811 351760 206867 352480
rect 214907 351760 214963 352480
rect 223049 351760 223105 352480
rect 231145 351760 231201 352480
rect 239241 351760 239297 352480
rect 247383 351760 247439 352480
rect 255479 351760 255535 352480
rect 263575 351760 263631 352480
rect 271717 351760 271773 352480
rect 279813 351760 279869 352480
rect 287909 351760 287965 352480
rect 271 -480 327 240
rect 823 -480 879 240
rect 1421 -480 1477 240
rect 2019 -480 2075 240
rect 2617 -480 2673 240
rect 3215 -480 3271 240
rect 3813 -480 3869 240
rect 4411 -480 4467 240
rect 5009 -480 5065 240
rect 5607 -480 5663 240
rect 6205 -480 6261 240
rect 6803 -480 6859 240
rect 7401 -480 7457 240
rect 7999 -480 8055 240
rect 8597 -480 8653 240
rect 9149 -480 9205 240
rect 9747 -480 9803 240
rect 10345 -480 10401 240
rect 10943 -480 10999 240
rect 11541 -480 11597 240
rect 12139 -480 12195 240
rect 12737 -480 12793 240
rect 13335 -480 13391 240
rect 13933 -480 13989 240
rect 14531 -480 14587 240
rect 15129 -480 15185 240
rect 15727 -480 15783 240
rect 16325 -480 16381 240
rect 16923 -480 16979 240
rect 17475 -480 17531 240
rect 18073 -480 18129 240
rect 18671 -480 18727 240
rect 19269 -480 19325 240
rect 19867 -480 19923 240
rect 20465 -480 20521 240
rect 21063 -480 21119 240
rect 21661 -480 21717 240
rect 22259 -480 22315 240
rect 22857 -480 22913 240
rect 23455 -480 23511 240
rect 24053 -480 24109 240
rect 24651 -480 24707 240
rect 25249 -480 25305 240
rect 25801 -480 25857 240
rect 26399 -480 26455 240
rect 26997 -480 27053 240
rect 27595 -480 27651 240
rect 28193 -480 28249 240
rect 28791 -480 28847 240
rect 29389 -480 29445 240
rect 29987 -480 30043 240
rect 30585 -480 30641 240
rect 31183 -480 31239 240
rect 31781 -480 31837 240
rect 32379 -480 32435 240
rect 32977 -480 33033 240
rect 33575 -480 33631 240
rect 34127 -480 34183 240
rect 34725 -480 34781 240
rect 35323 -480 35379 240
rect 35921 -480 35977 240
rect 36519 -480 36575 240
rect 37117 -480 37173 240
rect 37715 -480 37771 240
rect 38313 -480 38369 240
rect 38911 -480 38967 240
rect 39509 -480 39565 240
rect 40107 -480 40163 240
rect 40705 -480 40761 240
rect 41303 -480 41359 240
rect 41901 -480 41957 240
rect 42453 -480 42509 240
rect 43051 -480 43107 240
rect 43649 -480 43705 240
rect 44247 -480 44303 240
rect 44845 -480 44901 240
rect 45443 -480 45499 240
rect 46041 -480 46097 240
rect 46639 -480 46695 240
rect 47237 -480 47293 240
rect 47835 -480 47891 240
rect 48433 -480 48489 240
rect 49031 -480 49087 240
rect 49629 -480 49685 240
rect 50227 -480 50283 240
rect 50779 -480 50835 240
rect 51377 -480 51433 240
rect 51975 -480 52031 240
rect 52573 -480 52629 240
rect 53171 -480 53227 240
rect 53769 -480 53825 240
rect 54367 -480 54423 240
rect 54965 -480 55021 240
rect 55563 -480 55619 240
rect 56161 -480 56217 240
rect 56759 -480 56815 240
rect 57357 -480 57413 240
rect 57955 -480 58011 240
rect 58553 -480 58609 240
rect 59105 -480 59161 240
rect 59703 -480 59759 240
rect 60301 -480 60357 240
rect 60899 -480 60955 240
rect 61497 -480 61553 240
rect 62095 -480 62151 240
rect 62693 -480 62749 240
rect 63291 -480 63347 240
rect 63889 -480 63945 240
rect 64487 -480 64543 240
rect 65085 -480 65141 240
rect 65683 -480 65739 240
rect 66281 -480 66337 240
rect 66879 -480 66935 240
rect 67431 -480 67487 240
rect 68029 -480 68085 240
rect 68627 -480 68683 240
rect 69225 -480 69281 240
rect 69823 -480 69879 240
rect 70421 -480 70477 240
rect 71019 -480 71075 240
rect 71617 -480 71673 240
rect 72215 -480 72271 240
rect 72813 -480 72869 240
rect 73411 -480 73467 240
rect 74009 -480 74065 240
rect 74607 -480 74663 240
rect 75205 -480 75261 240
rect 75757 -480 75813 240
rect 76355 -480 76411 240
rect 76953 -480 77009 240
rect 77551 -480 77607 240
rect 78149 -480 78205 240
rect 78747 -480 78803 240
rect 79345 -480 79401 240
rect 79943 -480 79999 240
rect 80541 -480 80597 240
rect 81139 -480 81195 240
rect 81737 -480 81793 240
rect 82335 -480 82391 240
rect 82933 -480 82989 240
rect 83531 -480 83587 240
rect 84083 -480 84139 240
rect 84681 -480 84737 240
rect 85279 -480 85335 240
rect 85877 -480 85933 240
rect 86475 -480 86531 240
rect 87073 -480 87129 240
rect 87671 -480 87727 240
rect 88269 -480 88325 240
rect 88867 -480 88923 240
rect 89465 -480 89521 240
rect 90063 -480 90119 240
rect 90661 -480 90717 240
rect 91259 -480 91315 240
rect 91857 -480 91913 240
rect 92409 -480 92465 240
rect 93007 -480 93063 240
rect 93605 -480 93661 240
rect 94203 -480 94259 240
rect 94801 -480 94857 240
rect 95399 -480 95455 240
rect 95997 -480 96053 240
rect 96595 -480 96651 240
rect 97193 -480 97249 240
rect 97791 -480 97847 240
rect 98389 -480 98445 240
rect 98987 -480 99043 240
rect 99585 -480 99641 240
rect 100183 -480 100239 240
rect 100735 -480 100791 240
rect 101333 -480 101389 240
rect 101931 -480 101987 240
rect 102529 -480 102585 240
rect 103127 -480 103183 240
rect 103725 -480 103781 240
rect 104323 -480 104379 240
rect 104921 -480 104977 240
rect 105519 -480 105575 240
rect 106117 -480 106173 240
rect 106715 -480 106771 240
rect 107313 -480 107369 240
rect 107911 -480 107967 240
rect 108509 -480 108565 240
rect 109061 -480 109117 240
rect 109659 -480 109715 240
rect 110257 -480 110313 240
rect 110855 -480 110911 240
rect 111453 -480 111509 240
rect 112051 -480 112107 240
rect 112649 -480 112705 240
rect 113247 -480 113303 240
rect 113845 -480 113901 240
rect 114443 -480 114499 240
rect 115041 -480 115097 240
rect 115639 -480 115695 240
rect 116237 -480 116293 240
rect 116835 -480 116891 240
rect 117387 -480 117443 240
rect 117985 -480 118041 240
rect 118583 -480 118639 240
rect 119181 -480 119237 240
rect 119779 -480 119835 240
rect 120377 -480 120433 240
rect 120975 -480 121031 240
rect 121573 -480 121629 240
rect 122171 -480 122227 240
rect 122769 -480 122825 240
rect 123367 -480 123423 240
rect 123965 -480 124021 240
rect 124563 -480 124619 240
rect 125161 -480 125217 240
rect 125713 -480 125769 240
rect 126311 -480 126367 240
rect 126909 -480 126965 240
rect 127507 -480 127563 240
rect 128105 -480 128161 240
rect 128703 -480 128759 240
rect 129301 -480 129357 240
rect 129899 -480 129955 240
rect 130497 -480 130553 240
rect 131095 -480 131151 240
rect 131693 -480 131749 240
rect 132291 -480 132347 240
rect 132889 -480 132945 240
rect 133487 -480 133543 240
rect 134039 -480 134095 240
rect 134637 -480 134693 240
rect 135235 -480 135291 240
rect 135833 -480 135889 240
rect 136431 -480 136487 240
rect 137029 -480 137085 240
rect 137627 -480 137683 240
rect 138225 -480 138281 240
rect 138823 -480 138879 240
rect 139421 -480 139477 240
rect 140019 -480 140075 240
rect 140617 -480 140673 240
rect 141215 -480 141271 240
rect 141813 -480 141869 240
rect 142365 -480 142421 240
rect 142963 -480 143019 240
rect 143561 -480 143617 240
rect 144159 -480 144215 240
rect 144757 -480 144813 240
rect 145355 -480 145411 240
rect 145953 -480 146009 240
rect 146551 -480 146607 240
rect 147149 -480 147205 240
rect 147747 -480 147803 240
rect 148345 -480 148401 240
rect 148943 -480 148999 240
rect 149541 -480 149597 240
rect 150139 -480 150195 240
rect 150691 -480 150747 240
rect 151289 -480 151345 240
rect 151887 -480 151943 240
rect 152485 -480 152541 240
rect 153083 -480 153139 240
rect 153681 -480 153737 240
rect 154279 -480 154335 240
rect 154877 -480 154933 240
rect 155475 -480 155531 240
rect 156073 -480 156129 240
rect 156671 -480 156727 240
rect 157269 -480 157325 240
rect 157867 -480 157923 240
rect 158465 -480 158521 240
rect 159017 -480 159073 240
rect 159615 -480 159671 240
rect 160213 -480 160269 240
rect 160811 -480 160867 240
rect 161409 -480 161465 240
rect 162007 -480 162063 240
rect 162605 -480 162661 240
rect 163203 -480 163259 240
rect 163801 -480 163857 240
rect 164399 -480 164455 240
rect 164997 -480 165053 240
rect 165595 -480 165651 240
rect 166193 -480 166249 240
rect 166791 -480 166847 240
rect 167343 -480 167399 240
rect 167941 -480 167997 240
rect 168539 -480 168595 240
rect 169137 -480 169193 240
rect 169735 -480 169791 240
rect 170333 -480 170389 240
rect 170931 -480 170987 240
rect 171529 -480 171585 240
rect 172127 -480 172183 240
rect 172725 -480 172781 240
rect 173323 -480 173379 240
rect 173921 -480 173977 240
rect 174519 -480 174575 240
rect 175117 -480 175173 240
rect 175669 -480 175725 240
rect 176267 -480 176323 240
rect 176865 -480 176921 240
rect 177463 -480 177519 240
rect 178061 -480 178117 240
rect 178659 -480 178715 240
rect 179257 -480 179313 240
rect 179855 -480 179911 240
rect 180453 -480 180509 240
rect 181051 -480 181107 240
rect 181649 -480 181705 240
rect 182247 -480 182303 240
rect 182845 -480 182901 240
rect 183443 -480 183499 240
rect 183995 -480 184051 240
rect 184593 -480 184649 240
rect 185191 -480 185247 240
rect 185789 -480 185845 240
rect 186387 -480 186443 240
rect 186985 -480 187041 240
rect 187583 -480 187639 240
rect 188181 -480 188237 240
rect 188779 -480 188835 240
rect 189377 -480 189433 240
rect 189975 -480 190031 240
rect 190573 -480 190629 240
rect 191171 -480 191227 240
rect 191769 -480 191825 240
rect 192321 -480 192377 240
rect 192919 -480 192975 240
rect 193517 -480 193573 240
rect 194115 -480 194171 240
rect 194713 -480 194769 240
rect 195311 -480 195367 240
rect 195909 -480 195965 240
rect 196507 -480 196563 240
rect 197105 -480 197161 240
rect 197703 -480 197759 240
rect 198301 -480 198357 240
rect 198899 -480 198955 240
rect 199497 -480 199553 240
rect 200095 -480 200151 240
rect 200647 -480 200703 240
rect 201245 -480 201301 240
rect 201843 -480 201899 240
rect 202441 -480 202497 240
rect 203039 -480 203095 240
rect 203637 -480 203693 240
rect 204235 -480 204291 240
rect 204833 -480 204889 240
rect 205431 -480 205487 240
rect 206029 -480 206085 240
rect 206627 -480 206683 240
rect 207225 -480 207281 240
rect 207823 -480 207879 240
rect 208421 -480 208477 240
rect 208973 -480 209029 240
rect 209571 -480 209627 240
rect 210169 -480 210225 240
rect 210767 -480 210823 240
rect 211365 -480 211421 240
rect 211963 -480 212019 240
rect 212561 -480 212617 240
rect 213159 -480 213215 240
rect 213757 -480 213813 240
rect 214355 -480 214411 240
rect 214953 -480 215009 240
rect 215551 -480 215607 240
rect 216149 -480 216205 240
rect 216747 -480 216803 240
rect 217299 -480 217355 240
rect 217897 -480 217953 240
rect 218495 -480 218551 240
rect 219093 -480 219149 240
rect 219691 -480 219747 240
rect 220289 -480 220345 240
rect 220887 -480 220943 240
rect 221485 -480 221541 240
rect 222083 -480 222139 240
rect 222681 -480 222737 240
rect 223279 -480 223335 240
rect 223877 -480 223933 240
rect 224475 -480 224531 240
rect 225073 -480 225129 240
rect 225625 -480 225681 240
rect 226223 -480 226279 240
rect 226821 -480 226877 240
rect 227419 -480 227475 240
rect 228017 -480 228073 240
rect 228615 -480 228671 240
rect 229213 -480 229269 240
rect 229811 -480 229867 240
rect 230409 -480 230465 240
rect 231007 -480 231063 240
rect 231605 -480 231661 240
rect 232203 -480 232259 240
rect 232801 -480 232857 240
rect 233399 -480 233455 240
rect 233951 -480 234007 240
rect 234549 -480 234605 240
rect 235147 -480 235203 240
rect 235745 -480 235801 240
rect 236343 -480 236399 240
rect 236941 -480 236997 240
rect 237539 -480 237595 240
rect 238137 -480 238193 240
rect 238735 -480 238791 240
rect 239333 -480 239389 240
rect 239931 -480 239987 240
rect 240529 -480 240585 240
rect 241127 -480 241183 240
rect 241725 -480 241781 240
rect 242277 -480 242333 240
rect 242875 -480 242931 240
rect 243473 -480 243529 240
rect 244071 -480 244127 240
rect 244669 -480 244725 240
rect 245267 -480 245323 240
rect 245865 -480 245921 240
rect 246463 -480 246519 240
rect 247061 -480 247117 240
rect 247659 -480 247715 240
rect 248257 -480 248313 240
rect 248855 -480 248911 240
rect 249453 -480 249509 240
rect 250051 -480 250107 240
rect 250603 -480 250659 240
rect 251201 -480 251257 240
rect 251799 -480 251855 240
rect 252397 -480 252453 240
rect 252995 -480 253051 240
rect 253593 -480 253649 240
rect 254191 -480 254247 240
rect 254789 -480 254845 240
rect 255387 -480 255443 240
rect 255985 -480 256041 240
rect 256583 -480 256639 240
rect 257181 -480 257237 240
rect 257779 -480 257835 240
rect 258377 -480 258433 240
rect 258929 -480 258985 240
rect 259527 -480 259583 240
rect 260125 -480 260181 240
rect 260723 -480 260779 240
rect 261321 -480 261377 240
rect 261919 -480 261975 240
rect 262517 -480 262573 240
rect 263115 -480 263171 240
rect 263713 -480 263769 240
rect 264311 -480 264367 240
rect 264909 -480 264965 240
rect 265507 -480 265563 240
rect 266105 -480 266161 240
rect 266703 -480 266759 240
rect 267255 -480 267311 240
rect 267853 -480 267909 240
rect 268451 -480 268507 240
rect 269049 -480 269105 240
rect 269647 -480 269703 240
rect 270245 -480 270301 240
rect 270843 -480 270899 240
rect 271441 -480 271497 240
rect 272039 -480 272095 240
rect 272637 -480 272693 240
rect 273235 -480 273291 240
rect 273833 -480 273889 240
rect 274431 -480 274487 240
rect 275029 -480 275085 240
rect 275581 -480 275637 240
rect 276179 -480 276235 240
rect 276777 -480 276833 240
rect 277375 -480 277431 240
rect 277973 -480 278029 240
rect 278571 -480 278627 240
rect 279169 -480 279225 240
rect 279767 -480 279823 240
rect 280365 -480 280421 240
rect 280963 -480 281019 240
rect 281561 -480 281617 240
rect 282159 -480 282215 240
rect 282757 -480 282813 240
rect 283355 -480 283411 240
rect 283907 -480 283963 240
rect 284505 -480 284561 240
rect 285103 -480 285159 240
rect 285701 -480 285757 240
rect 286299 -480 286355 240
rect 286897 -480 286953 240
rect 287495 -480 287551 240
rect 288093 -480 288149 240
rect 288691 -480 288747 240
rect 289289 -480 289345 240
rect 289887 -480 289943 240
rect 290485 -480 290541 240
rect 291083 -480 291139 240
rect 291681 -480 291737 240
<< metal3 >>
rect 291760 348950 292480 349070
rect -480 348270 240 348390
rect 291760 343102 292480 343222
rect -480 341062 240 341182
rect 291760 337254 292480 337374
rect -480 333922 240 334042
rect 291760 331338 292480 331458
rect -480 326714 240 326834
rect 291760 325490 292480 325610
rect 291760 319642 292480 319762
rect -480 319506 240 319626
rect 291760 313794 292480 313914
rect -480 312366 240 312486
rect 291760 307878 292480 307998
rect -480 305158 240 305278
rect 291760 302030 292480 302150
rect -480 297950 240 298070
rect 291760 296182 292480 296302
rect -480 290810 240 290930
rect 291760 290334 292480 290454
rect 291760 284418 292480 284538
rect -480 283602 240 283722
rect 291760 278570 292480 278690
rect -480 276462 240 276582
rect 291760 272722 292480 272842
rect -480 269254 240 269374
rect 291760 266874 292480 266994
rect -480 262046 240 262166
rect 291760 260958 292480 261078
rect 291760 255110 292480 255230
rect -480 254906 240 255026
rect 291760 249262 292480 249382
rect -480 247698 240 247818
rect 291760 243346 292480 243466
rect -480 240490 240 240610
rect 291760 237498 292480 237618
rect -480 233350 240 233470
rect 291760 231650 292480 231770
rect -480 226142 240 226262
rect 291760 225802 292480 225922
rect 291760 219886 292480 220006
rect -480 218934 240 219054
rect 291760 214038 292480 214158
rect -480 211794 240 211914
rect 291760 208190 292480 208310
rect -480 204586 240 204706
rect 291760 202342 292480 202462
rect -480 197446 240 197566
rect 291760 196426 292480 196546
rect 291760 190578 292480 190698
rect -480 190238 240 190358
rect 291760 184730 292480 184850
rect -480 183030 240 183150
rect 291760 178882 292480 179002
rect -480 175890 240 176010
rect 291760 172966 292480 173086
rect -480 168682 240 168802
rect 291760 167118 292480 167238
rect -480 161474 240 161594
rect 291760 161270 292480 161390
rect 291760 155354 292480 155474
rect -480 154334 240 154454
rect 291760 149506 292480 149626
rect -480 147126 240 147246
rect 291760 143658 292480 143778
rect -480 139986 240 140106
rect 291760 137810 292480 137930
rect -480 132778 240 132898
rect 291760 131894 292480 132014
rect 291760 126046 292480 126166
rect -480 125570 240 125690
rect 291760 120198 292480 120318
rect -480 118430 240 118550
rect 291760 114350 292480 114470
rect -480 111222 240 111342
rect 291760 108434 292480 108554
rect -480 104014 240 104134
rect 291760 102586 292480 102706
rect -480 96874 240 96994
rect 291760 96738 292480 96858
rect 291760 90890 292480 91010
rect -480 89666 240 89786
rect 291760 84974 292480 85094
rect -480 82458 240 82578
rect 291760 79126 292480 79246
rect -480 75318 240 75438
rect 291760 73278 292480 73398
rect -480 68110 240 68230
rect 291760 67362 292480 67482
rect 291760 61514 292480 61634
rect -480 60970 240 61090
rect 291760 55666 292480 55786
rect -480 53762 240 53882
rect 291760 49818 292480 49938
rect -480 46554 240 46674
rect 291760 43902 292480 44022
rect -480 39414 240 39534
rect 291760 38054 292480 38174
rect -480 32206 240 32326
rect 291760 32206 292480 32326
rect 291760 26358 292480 26478
rect -480 24998 240 25118
rect 291760 20442 292480 20562
rect -480 17858 240 17978
rect 291760 14594 292480 14714
rect -480 10650 240 10770
rect 291760 8746 292480 8866
rect -480 3510 240 3630
rect 291760 2898 292480 3018
<< metal4 >>
rect -4288 355709 -3988 355720
rect -4288 355591 -4197 355709
rect -4079 355591 -3988 355709
rect -4288 355549 -3988 355591
rect -4288 355431 -4197 355549
rect -4079 355431 -3988 355549
rect -4288 339627 -3988 355431
rect -4288 339509 -4197 339627
rect -4079 339509 -3988 339627
rect -4288 339467 -3988 339509
rect -4288 339349 -4197 339467
rect -4079 339349 -3988 339467
rect -4288 321627 -3988 339349
rect -4288 321509 -4197 321627
rect -4079 321509 -3988 321627
rect -4288 321467 -3988 321509
rect -4288 321349 -4197 321467
rect -4079 321349 -3988 321467
rect -4288 303627 -3988 321349
rect -4288 303509 -4197 303627
rect -4079 303509 -3988 303627
rect -4288 303467 -3988 303509
rect -4288 303349 -4197 303467
rect -4079 303349 -3988 303467
rect -4288 285627 -3988 303349
rect -4288 285509 -4197 285627
rect -4079 285509 -3988 285627
rect -4288 285467 -3988 285509
rect -4288 285349 -4197 285467
rect -4079 285349 -3988 285467
rect -4288 267627 -3988 285349
rect -4288 267509 -4197 267627
rect -4079 267509 -3988 267627
rect -4288 267467 -3988 267509
rect -4288 267349 -4197 267467
rect -4079 267349 -3988 267467
rect -4288 249627 -3988 267349
rect -4288 249509 -4197 249627
rect -4079 249509 -3988 249627
rect -4288 249467 -3988 249509
rect -4288 249349 -4197 249467
rect -4079 249349 -3988 249467
rect -4288 231627 -3988 249349
rect -4288 231509 -4197 231627
rect -4079 231509 -3988 231627
rect -4288 231467 -3988 231509
rect -4288 231349 -4197 231467
rect -4079 231349 -3988 231467
rect -4288 213627 -3988 231349
rect -4288 213509 -4197 213627
rect -4079 213509 -3988 213627
rect -4288 213467 -3988 213509
rect -4288 213349 -4197 213467
rect -4079 213349 -3988 213467
rect -4288 195627 -3988 213349
rect -4288 195509 -4197 195627
rect -4079 195509 -3988 195627
rect -4288 195467 -3988 195509
rect -4288 195349 -4197 195467
rect -4079 195349 -3988 195467
rect -4288 177627 -3988 195349
rect -4288 177509 -4197 177627
rect -4079 177509 -3988 177627
rect -4288 177467 -3988 177509
rect -4288 177349 -4197 177467
rect -4079 177349 -3988 177467
rect -4288 159627 -3988 177349
rect -4288 159509 -4197 159627
rect -4079 159509 -3988 159627
rect -4288 159467 -3988 159509
rect -4288 159349 -4197 159467
rect -4079 159349 -3988 159467
rect -4288 141627 -3988 159349
rect -4288 141509 -4197 141627
rect -4079 141509 -3988 141627
rect -4288 141467 -3988 141509
rect -4288 141349 -4197 141467
rect -4079 141349 -3988 141467
rect -4288 123627 -3988 141349
rect -4288 123509 -4197 123627
rect -4079 123509 -3988 123627
rect -4288 123467 -3988 123509
rect -4288 123349 -4197 123467
rect -4079 123349 -3988 123467
rect -4288 105627 -3988 123349
rect -4288 105509 -4197 105627
rect -4079 105509 -3988 105627
rect -4288 105467 -3988 105509
rect -4288 105349 -4197 105467
rect -4079 105349 -3988 105467
rect -4288 87627 -3988 105349
rect -4288 87509 -4197 87627
rect -4079 87509 -3988 87627
rect -4288 87467 -3988 87509
rect -4288 87349 -4197 87467
rect -4079 87349 -3988 87467
rect -4288 69627 -3988 87349
rect -4288 69509 -4197 69627
rect -4079 69509 -3988 69627
rect -4288 69467 -3988 69509
rect -4288 69349 -4197 69467
rect -4079 69349 -3988 69467
rect -4288 51627 -3988 69349
rect -4288 51509 -4197 51627
rect -4079 51509 -3988 51627
rect -4288 51467 -3988 51509
rect -4288 51349 -4197 51467
rect -4079 51349 -3988 51467
rect -4288 33627 -3988 51349
rect -4288 33509 -4197 33627
rect -4079 33509 -3988 33627
rect -4288 33467 -3988 33509
rect -4288 33349 -4197 33467
rect -4079 33349 -3988 33467
rect -4288 15627 -3988 33349
rect -4288 15509 -4197 15627
rect -4079 15509 -3988 15627
rect -4288 15467 -3988 15509
rect -4288 15349 -4197 15467
rect -4079 15349 -3988 15467
rect -4288 -3463 -3988 15349
rect -3818 355239 -3518 355250
rect -3818 355121 -3727 355239
rect -3609 355121 -3518 355239
rect -3818 355079 -3518 355121
rect -3818 354961 -3727 355079
rect -3609 354961 -3518 355079
rect -3818 348627 -3518 354961
rect 5802 355239 6102 355720
rect 5802 355121 5893 355239
rect 6011 355121 6102 355239
rect 5802 355079 6102 355121
rect 5802 354961 5893 355079
rect 6011 354961 6102 355079
rect -3818 348509 -3727 348627
rect -3609 348509 -3518 348627
rect -3818 348467 -3518 348509
rect -3818 348349 -3727 348467
rect -3609 348349 -3518 348467
rect -3818 330627 -3518 348349
rect -3818 330509 -3727 330627
rect -3609 330509 -3518 330627
rect -3818 330467 -3518 330509
rect -3818 330349 -3727 330467
rect -3609 330349 -3518 330467
rect -3818 312627 -3518 330349
rect -3818 312509 -3727 312627
rect -3609 312509 -3518 312627
rect -3818 312467 -3518 312509
rect -3818 312349 -3727 312467
rect -3609 312349 -3518 312467
rect -3818 294627 -3518 312349
rect -3818 294509 -3727 294627
rect -3609 294509 -3518 294627
rect -3818 294467 -3518 294509
rect -3818 294349 -3727 294467
rect -3609 294349 -3518 294467
rect -3818 276627 -3518 294349
rect -3818 276509 -3727 276627
rect -3609 276509 -3518 276627
rect -3818 276467 -3518 276509
rect -3818 276349 -3727 276467
rect -3609 276349 -3518 276467
rect -3818 258627 -3518 276349
rect -3818 258509 -3727 258627
rect -3609 258509 -3518 258627
rect -3818 258467 -3518 258509
rect -3818 258349 -3727 258467
rect -3609 258349 -3518 258467
rect -3818 240627 -3518 258349
rect -3818 240509 -3727 240627
rect -3609 240509 -3518 240627
rect -3818 240467 -3518 240509
rect -3818 240349 -3727 240467
rect -3609 240349 -3518 240467
rect -3818 222627 -3518 240349
rect -3818 222509 -3727 222627
rect -3609 222509 -3518 222627
rect -3818 222467 -3518 222509
rect -3818 222349 -3727 222467
rect -3609 222349 -3518 222467
rect -3818 204627 -3518 222349
rect -3818 204509 -3727 204627
rect -3609 204509 -3518 204627
rect -3818 204467 -3518 204509
rect -3818 204349 -3727 204467
rect -3609 204349 -3518 204467
rect -3818 186627 -3518 204349
rect -3818 186509 -3727 186627
rect -3609 186509 -3518 186627
rect -3818 186467 -3518 186509
rect -3818 186349 -3727 186467
rect -3609 186349 -3518 186467
rect -3818 168627 -3518 186349
rect -3818 168509 -3727 168627
rect -3609 168509 -3518 168627
rect -3818 168467 -3518 168509
rect -3818 168349 -3727 168467
rect -3609 168349 -3518 168467
rect -3818 150627 -3518 168349
rect -3818 150509 -3727 150627
rect -3609 150509 -3518 150627
rect -3818 150467 -3518 150509
rect -3818 150349 -3727 150467
rect -3609 150349 -3518 150467
rect -3818 132627 -3518 150349
rect -3818 132509 -3727 132627
rect -3609 132509 -3518 132627
rect -3818 132467 -3518 132509
rect -3818 132349 -3727 132467
rect -3609 132349 -3518 132467
rect -3818 114627 -3518 132349
rect -3818 114509 -3727 114627
rect -3609 114509 -3518 114627
rect -3818 114467 -3518 114509
rect -3818 114349 -3727 114467
rect -3609 114349 -3518 114467
rect -3818 96627 -3518 114349
rect -3818 96509 -3727 96627
rect -3609 96509 -3518 96627
rect -3818 96467 -3518 96509
rect -3818 96349 -3727 96467
rect -3609 96349 -3518 96467
rect -3818 78627 -3518 96349
rect -3818 78509 -3727 78627
rect -3609 78509 -3518 78627
rect -3818 78467 -3518 78509
rect -3818 78349 -3727 78467
rect -3609 78349 -3518 78467
rect -3818 60627 -3518 78349
rect -3818 60509 -3727 60627
rect -3609 60509 -3518 60627
rect -3818 60467 -3518 60509
rect -3818 60349 -3727 60467
rect -3609 60349 -3518 60467
rect -3818 42627 -3518 60349
rect -3818 42509 -3727 42627
rect -3609 42509 -3518 42627
rect -3818 42467 -3518 42509
rect -3818 42349 -3727 42467
rect -3609 42349 -3518 42467
rect -3818 24627 -3518 42349
rect -3818 24509 -3727 24627
rect -3609 24509 -3518 24627
rect -3818 24467 -3518 24509
rect -3818 24349 -3727 24467
rect -3609 24349 -3518 24467
rect -3818 6627 -3518 24349
rect -3818 6509 -3727 6627
rect -3609 6509 -3518 6627
rect -3818 6467 -3518 6509
rect -3818 6349 -3727 6467
rect -3609 6349 -3518 6467
rect -3818 -2993 -3518 6349
rect -3348 354769 -3048 354780
rect -3348 354651 -3257 354769
rect -3139 354651 -3048 354769
rect -3348 354609 -3048 354651
rect -3348 354491 -3257 354609
rect -3139 354491 -3048 354609
rect -3348 337827 -3048 354491
rect -3348 337709 -3257 337827
rect -3139 337709 -3048 337827
rect -3348 337667 -3048 337709
rect -3348 337549 -3257 337667
rect -3139 337549 -3048 337667
rect -3348 319827 -3048 337549
rect -3348 319709 -3257 319827
rect -3139 319709 -3048 319827
rect -3348 319667 -3048 319709
rect -3348 319549 -3257 319667
rect -3139 319549 -3048 319667
rect -3348 301827 -3048 319549
rect -3348 301709 -3257 301827
rect -3139 301709 -3048 301827
rect -3348 301667 -3048 301709
rect -3348 301549 -3257 301667
rect -3139 301549 -3048 301667
rect -3348 283827 -3048 301549
rect -3348 283709 -3257 283827
rect -3139 283709 -3048 283827
rect -3348 283667 -3048 283709
rect -3348 283549 -3257 283667
rect -3139 283549 -3048 283667
rect -3348 265827 -3048 283549
rect -3348 265709 -3257 265827
rect -3139 265709 -3048 265827
rect -3348 265667 -3048 265709
rect -3348 265549 -3257 265667
rect -3139 265549 -3048 265667
rect -3348 247827 -3048 265549
rect -3348 247709 -3257 247827
rect -3139 247709 -3048 247827
rect -3348 247667 -3048 247709
rect -3348 247549 -3257 247667
rect -3139 247549 -3048 247667
rect -3348 229827 -3048 247549
rect -3348 229709 -3257 229827
rect -3139 229709 -3048 229827
rect -3348 229667 -3048 229709
rect -3348 229549 -3257 229667
rect -3139 229549 -3048 229667
rect -3348 211827 -3048 229549
rect -3348 211709 -3257 211827
rect -3139 211709 -3048 211827
rect -3348 211667 -3048 211709
rect -3348 211549 -3257 211667
rect -3139 211549 -3048 211667
rect -3348 193827 -3048 211549
rect -3348 193709 -3257 193827
rect -3139 193709 -3048 193827
rect -3348 193667 -3048 193709
rect -3348 193549 -3257 193667
rect -3139 193549 -3048 193667
rect -3348 175827 -3048 193549
rect -3348 175709 -3257 175827
rect -3139 175709 -3048 175827
rect -3348 175667 -3048 175709
rect -3348 175549 -3257 175667
rect -3139 175549 -3048 175667
rect -3348 157827 -3048 175549
rect -3348 157709 -3257 157827
rect -3139 157709 -3048 157827
rect -3348 157667 -3048 157709
rect -3348 157549 -3257 157667
rect -3139 157549 -3048 157667
rect -3348 139827 -3048 157549
rect -3348 139709 -3257 139827
rect -3139 139709 -3048 139827
rect -3348 139667 -3048 139709
rect -3348 139549 -3257 139667
rect -3139 139549 -3048 139667
rect -3348 121827 -3048 139549
rect -3348 121709 -3257 121827
rect -3139 121709 -3048 121827
rect -3348 121667 -3048 121709
rect -3348 121549 -3257 121667
rect -3139 121549 -3048 121667
rect -3348 103827 -3048 121549
rect -3348 103709 -3257 103827
rect -3139 103709 -3048 103827
rect -3348 103667 -3048 103709
rect -3348 103549 -3257 103667
rect -3139 103549 -3048 103667
rect -3348 85827 -3048 103549
rect -3348 85709 -3257 85827
rect -3139 85709 -3048 85827
rect -3348 85667 -3048 85709
rect -3348 85549 -3257 85667
rect -3139 85549 -3048 85667
rect -3348 67827 -3048 85549
rect -3348 67709 -3257 67827
rect -3139 67709 -3048 67827
rect -3348 67667 -3048 67709
rect -3348 67549 -3257 67667
rect -3139 67549 -3048 67667
rect -3348 49827 -3048 67549
rect -3348 49709 -3257 49827
rect -3139 49709 -3048 49827
rect -3348 49667 -3048 49709
rect -3348 49549 -3257 49667
rect -3139 49549 -3048 49667
rect -3348 31827 -3048 49549
rect -3348 31709 -3257 31827
rect -3139 31709 -3048 31827
rect -3348 31667 -3048 31709
rect -3348 31549 -3257 31667
rect -3139 31549 -3048 31667
rect -3348 13827 -3048 31549
rect -3348 13709 -3257 13827
rect -3139 13709 -3048 13827
rect -3348 13667 -3048 13709
rect -3348 13549 -3257 13667
rect -3139 13549 -3048 13667
rect -3348 -2523 -3048 13549
rect -2878 354299 -2578 354310
rect -2878 354181 -2787 354299
rect -2669 354181 -2578 354299
rect -2878 354139 -2578 354181
rect -2878 354021 -2787 354139
rect -2669 354021 -2578 354139
rect -2878 346827 -2578 354021
rect 4002 354299 4302 354780
rect 4002 354181 4093 354299
rect 4211 354181 4302 354299
rect 4002 354139 4302 354181
rect 4002 354021 4093 354139
rect 4211 354021 4302 354139
rect -2878 346709 -2787 346827
rect -2669 346709 -2578 346827
rect -2878 346667 -2578 346709
rect -2878 346549 -2787 346667
rect -2669 346549 -2578 346667
rect -2878 328827 -2578 346549
rect -2878 328709 -2787 328827
rect -2669 328709 -2578 328827
rect -2878 328667 -2578 328709
rect -2878 328549 -2787 328667
rect -2669 328549 -2578 328667
rect -2878 310827 -2578 328549
rect -2878 310709 -2787 310827
rect -2669 310709 -2578 310827
rect -2878 310667 -2578 310709
rect -2878 310549 -2787 310667
rect -2669 310549 -2578 310667
rect -2878 292827 -2578 310549
rect -2878 292709 -2787 292827
rect -2669 292709 -2578 292827
rect -2878 292667 -2578 292709
rect -2878 292549 -2787 292667
rect -2669 292549 -2578 292667
rect -2878 274827 -2578 292549
rect -2878 274709 -2787 274827
rect -2669 274709 -2578 274827
rect -2878 274667 -2578 274709
rect -2878 274549 -2787 274667
rect -2669 274549 -2578 274667
rect -2878 256827 -2578 274549
rect -2878 256709 -2787 256827
rect -2669 256709 -2578 256827
rect -2878 256667 -2578 256709
rect -2878 256549 -2787 256667
rect -2669 256549 -2578 256667
rect -2878 238827 -2578 256549
rect -2878 238709 -2787 238827
rect -2669 238709 -2578 238827
rect -2878 238667 -2578 238709
rect -2878 238549 -2787 238667
rect -2669 238549 -2578 238667
rect -2878 220827 -2578 238549
rect -2878 220709 -2787 220827
rect -2669 220709 -2578 220827
rect -2878 220667 -2578 220709
rect -2878 220549 -2787 220667
rect -2669 220549 -2578 220667
rect -2878 202827 -2578 220549
rect -2878 202709 -2787 202827
rect -2669 202709 -2578 202827
rect -2878 202667 -2578 202709
rect -2878 202549 -2787 202667
rect -2669 202549 -2578 202667
rect -2878 184827 -2578 202549
rect -2878 184709 -2787 184827
rect -2669 184709 -2578 184827
rect -2878 184667 -2578 184709
rect -2878 184549 -2787 184667
rect -2669 184549 -2578 184667
rect -2878 166827 -2578 184549
rect -2878 166709 -2787 166827
rect -2669 166709 -2578 166827
rect -2878 166667 -2578 166709
rect -2878 166549 -2787 166667
rect -2669 166549 -2578 166667
rect -2878 148827 -2578 166549
rect -2878 148709 -2787 148827
rect -2669 148709 -2578 148827
rect -2878 148667 -2578 148709
rect -2878 148549 -2787 148667
rect -2669 148549 -2578 148667
rect -2878 130827 -2578 148549
rect -2878 130709 -2787 130827
rect -2669 130709 -2578 130827
rect -2878 130667 -2578 130709
rect -2878 130549 -2787 130667
rect -2669 130549 -2578 130667
rect -2878 112827 -2578 130549
rect -2878 112709 -2787 112827
rect -2669 112709 -2578 112827
rect -2878 112667 -2578 112709
rect -2878 112549 -2787 112667
rect -2669 112549 -2578 112667
rect -2878 94827 -2578 112549
rect -2878 94709 -2787 94827
rect -2669 94709 -2578 94827
rect -2878 94667 -2578 94709
rect -2878 94549 -2787 94667
rect -2669 94549 -2578 94667
rect -2878 76827 -2578 94549
rect -2878 76709 -2787 76827
rect -2669 76709 -2578 76827
rect -2878 76667 -2578 76709
rect -2878 76549 -2787 76667
rect -2669 76549 -2578 76667
rect -2878 58827 -2578 76549
rect -2878 58709 -2787 58827
rect -2669 58709 -2578 58827
rect -2878 58667 -2578 58709
rect -2878 58549 -2787 58667
rect -2669 58549 -2578 58667
rect -2878 40827 -2578 58549
rect -2878 40709 -2787 40827
rect -2669 40709 -2578 40827
rect -2878 40667 -2578 40709
rect -2878 40549 -2787 40667
rect -2669 40549 -2578 40667
rect -2878 22827 -2578 40549
rect -2878 22709 -2787 22827
rect -2669 22709 -2578 22827
rect -2878 22667 -2578 22709
rect -2878 22549 -2787 22667
rect -2669 22549 -2578 22667
rect -2878 4827 -2578 22549
rect -2878 4709 -2787 4827
rect -2669 4709 -2578 4827
rect -2878 4667 -2578 4709
rect -2878 4549 -2787 4667
rect -2669 4549 -2578 4667
rect -2878 -2053 -2578 4549
rect -2408 353829 -2108 353840
rect -2408 353711 -2317 353829
rect -2199 353711 -2108 353829
rect -2408 353669 -2108 353711
rect -2408 353551 -2317 353669
rect -2199 353551 -2108 353669
rect -2408 336027 -2108 353551
rect -2408 335909 -2317 336027
rect -2199 335909 -2108 336027
rect -2408 335867 -2108 335909
rect -2408 335749 -2317 335867
rect -2199 335749 -2108 335867
rect -2408 318027 -2108 335749
rect -2408 317909 -2317 318027
rect -2199 317909 -2108 318027
rect -2408 317867 -2108 317909
rect -2408 317749 -2317 317867
rect -2199 317749 -2108 317867
rect -2408 300027 -2108 317749
rect -2408 299909 -2317 300027
rect -2199 299909 -2108 300027
rect -2408 299867 -2108 299909
rect -2408 299749 -2317 299867
rect -2199 299749 -2108 299867
rect -2408 282027 -2108 299749
rect -2408 281909 -2317 282027
rect -2199 281909 -2108 282027
rect -2408 281867 -2108 281909
rect -2408 281749 -2317 281867
rect -2199 281749 -2108 281867
rect -2408 264027 -2108 281749
rect -2408 263909 -2317 264027
rect -2199 263909 -2108 264027
rect -2408 263867 -2108 263909
rect -2408 263749 -2317 263867
rect -2199 263749 -2108 263867
rect -2408 246027 -2108 263749
rect -2408 245909 -2317 246027
rect -2199 245909 -2108 246027
rect -2408 245867 -2108 245909
rect -2408 245749 -2317 245867
rect -2199 245749 -2108 245867
rect -2408 228027 -2108 245749
rect -2408 227909 -2317 228027
rect -2199 227909 -2108 228027
rect -2408 227867 -2108 227909
rect -2408 227749 -2317 227867
rect -2199 227749 -2108 227867
rect -2408 210027 -2108 227749
rect -2408 209909 -2317 210027
rect -2199 209909 -2108 210027
rect -2408 209867 -2108 209909
rect -2408 209749 -2317 209867
rect -2199 209749 -2108 209867
rect -2408 192027 -2108 209749
rect -2408 191909 -2317 192027
rect -2199 191909 -2108 192027
rect -2408 191867 -2108 191909
rect -2408 191749 -2317 191867
rect -2199 191749 -2108 191867
rect -2408 174027 -2108 191749
rect -2408 173909 -2317 174027
rect -2199 173909 -2108 174027
rect -2408 173867 -2108 173909
rect -2408 173749 -2317 173867
rect -2199 173749 -2108 173867
rect -2408 156027 -2108 173749
rect -2408 155909 -2317 156027
rect -2199 155909 -2108 156027
rect -2408 155867 -2108 155909
rect -2408 155749 -2317 155867
rect -2199 155749 -2108 155867
rect -2408 138027 -2108 155749
rect -2408 137909 -2317 138027
rect -2199 137909 -2108 138027
rect -2408 137867 -2108 137909
rect -2408 137749 -2317 137867
rect -2199 137749 -2108 137867
rect -2408 120027 -2108 137749
rect -2408 119909 -2317 120027
rect -2199 119909 -2108 120027
rect -2408 119867 -2108 119909
rect -2408 119749 -2317 119867
rect -2199 119749 -2108 119867
rect -2408 102027 -2108 119749
rect -2408 101909 -2317 102027
rect -2199 101909 -2108 102027
rect -2408 101867 -2108 101909
rect -2408 101749 -2317 101867
rect -2199 101749 -2108 101867
rect -2408 84027 -2108 101749
rect -2408 83909 -2317 84027
rect -2199 83909 -2108 84027
rect -2408 83867 -2108 83909
rect -2408 83749 -2317 83867
rect -2199 83749 -2108 83867
rect -2408 66027 -2108 83749
rect -2408 65909 -2317 66027
rect -2199 65909 -2108 66027
rect -2408 65867 -2108 65909
rect -2408 65749 -2317 65867
rect -2199 65749 -2108 65867
rect -2408 48027 -2108 65749
rect -2408 47909 -2317 48027
rect -2199 47909 -2108 48027
rect -2408 47867 -2108 47909
rect -2408 47749 -2317 47867
rect -2199 47749 -2108 47867
rect -2408 30027 -2108 47749
rect -2408 29909 -2317 30027
rect -2199 29909 -2108 30027
rect -2408 29867 -2108 29909
rect -2408 29749 -2317 29867
rect -2199 29749 -2108 29867
rect -2408 12027 -2108 29749
rect -2408 11909 -2317 12027
rect -2199 11909 -2108 12027
rect -2408 11867 -2108 11909
rect -2408 11749 -2317 11867
rect -2199 11749 -2108 11867
rect -2408 -1583 -2108 11749
rect -1938 353359 -1638 353370
rect -1938 353241 -1847 353359
rect -1729 353241 -1638 353359
rect -1938 353199 -1638 353241
rect -1938 353081 -1847 353199
rect -1729 353081 -1638 353199
rect -1938 345027 -1638 353081
rect 2202 353359 2502 353840
rect 2202 353241 2293 353359
rect 2411 353241 2502 353359
rect 2202 353199 2502 353241
rect 2202 353081 2293 353199
rect 2411 353081 2502 353199
rect -1938 344909 -1847 345027
rect -1729 344909 -1638 345027
rect -1938 344867 -1638 344909
rect -1938 344749 -1847 344867
rect -1729 344749 -1638 344867
rect -1938 327027 -1638 344749
rect -1938 326909 -1847 327027
rect -1729 326909 -1638 327027
rect -1938 326867 -1638 326909
rect -1938 326749 -1847 326867
rect -1729 326749 -1638 326867
rect -1938 309027 -1638 326749
rect -1938 308909 -1847 309027
rect -1729 308909 -1638 309027
rect -1938 308867 -1638 308909
rect -1938 308749 -1847 308867
rect -1729 308749 -1638 308867
rect -1938 291027 -1638 308749
rect -1938 290909 -1847 291027
rect -1729 290909 -1638 291027
rect -1938 290867 -1638 290909
rect -1938 290749 -1847 290867
rect -1729 290749 -1638 290867
rect -1938 273027 -1638 290749
rect -1938 272909 -1847 273027
rect -1729 272909 -1638 273027
rect -1938 272867 -1638 272909
rect -1938 272749 -1847 272867
rect -1729 272749 -1638 272867
rect -1938 255027 -1638 272749
rect -1938 254909 -1847 255027
rect -1729 254909 -1638 255027
rect -1938 254867 -1638 254909
rect -1938 254749 -1847 254867
rect -1729 254749 -1638 254867
rect -1938 237027 -1638 254749
rect -1938 236909 -1847 237027
rect -1729 236909 -1638 237027
rect -1938 236867 -1638 236909
rect -1938 236749 -1847 236867
rect -1729 236749 -1638 236867
rect -1938 219027 -1638 236749
rect -1938 218909 -1847 219027
rect -1729 218909 -1638 219027
rect -1938 218867 -1638 218909
rect -1938 218749 -1847 218867
rect -1729 218749 -1638 218867
rect -1938 201027 -1638 218749
rect -1938 200909 -1847 201027
rect -1729 200909 -1638 201027
rect -1938 200867 -1638 200909
rect -1938 200749 -1847 200867
rect -1729 200749 -1638 200867
rect -1938 183027 -1638 200749
rect -1938 182909 -1847 183027
rect -1729 182909 -1638 183027
rect -1938 182867 -1638 182909
rect -1938 182749 -1847 182867
rect -1729 182749 -1638 182867
rect -1938 165027 -1638 182749
rect -1938 164909 -1847 165027
rect -1729 164909 -1638 165027
rect -1938 164867 -1638 164909
rect -1938 164749 -1847 164867
rect -1729 164749 -1638 164867
rect -1938 147027 -1638 164749
rect -1938 146909 -1847 147027
rect -1729 146909 -1638 147027
rect -1938 146867 -1638 146909
rect -1938 146749 -1847 146867
rect -1729 146749 -1638 146867
rect -1938 129027 -1638 146749
rect -1938 128909 -1847 129027
rect -1729 128909 -1638 129027
rect -1938 128867 -1638 128909
rect -1938 128749 -1847 128867
rect -1729 128749 -1638 128867
rect -1938 111027 -1638 128749
rect -1938 110909 -1847 111027
rect -1729 110909 -1638 111027
rect -1938 110867 -1638 110909
rect -1938 110749 -1847 110867
rect -1729 110749 -1638 110867
rect -1938 93027 -1638 110749
rect -1938 92909 -1847 93027
rect -1729 92909 -1638 93027
rect -1938 92867 -1638 92909
rect -1938 92749 -1847 92867
rect -1729 92749 -1638 92867
rect -1938 75027 -1638 92749
rect -1938 74909 -1847 75027
rect -1729 74909 -1638 75027
rect -1938 74867 -1638 74909
rect -1938 74749 -1847 74867
rect -1729 74749 -1638 74867
rect -1938 57027 -1638 74749
rect -1938 56909 -1847 57027
rect -1729 56909 -1638 57027
rect -1938 56867 -1638 56909
rect -1938 56749 -1847 56867
rect -1729 56749 -1638 56867
rect -1938 39027 -1638 56749
rect -1938 38909 -1847 39027
rect -1729 38909 -1638 39027
rect -1938 38867 -1638 38909
rect -1938 38749 -1847 38867
rect -1729 38749 -1638 38867
rect -1938 21027 -1638 38749
rect -1938 20909 -1847 21027
rect -1729 20909 -1638 21027
rect -1938 20867 -1638 20909
rect -1938 20749 -1847 20867
rect -1729 20749 -1638 20867
rect -1938 3027 -1638 20749
rect -1938 2909 -1847 3027
rect -1729 2909 -1638 3027
rect -1938 2867 -1638 2909
rect -1938 2749 -1847 2867
rect -1729 2749 -1638 2867
rect -1938 -1113 -1638 2749
rect -1468 352889 -1168 352900
rect -1468 352771 -1377 352889
rect -1259 352771 -1168 352889
rect -1468 352729 -1168 352771
rect -1468 352611 -1377 352729
rect -1259 352611 -1168 352729
rect -1468 334227 -1168 352611
rect -1468 334109 -1377 334227
rect -1259 334109 -1168 334227
rect -1468 334067 -1168 334109
rect -1468 333949 -1377 334067
rect -1259 333949 -1168 334067
rect -1468 316227 -1168 333949
rect -1468 316109 -1377 316227
rect -1259 316109 -1168 316227
rect -1468 316067 -1168 316109
rect -1468 315949 -1377 316067
rect -1259 315949 -1168 316067
rect -1468 298227 -1168 315949
rect -1468 298109 -1377 298227
rect -1259 298109 -1168 298227
rect -1468 298067 -1168 298109
rect -1468 297949 -1377 298067
rect -1259 297949 -1168 298067
rect -1468 280227 -1168 297949
rect -1468 280109 -1377 280227
rect -1259 280109 -1168 280227
rect -1468 280067 -1168 280109
rect -1468 279949 -1377 280067
rect -1259 279949 -1168 280067
rect -1468 262227 -1168 279949
rect -1468 262109 -1377 262227
rect -1259 262109 -1168 262227
rect -1468 262067 -1168 262109
rect -1468 261949 -1377 262067
rect -1259 261949 -1168 262067
rect -1468 244227 -1168 261949
rect -1468 244109 -1377 244227
rect -1259 244109 -1168 244227
rect -1468 244067 -1168 244109
rect -1468 243949 -1377 244067
rect -1259 243949 -1168 244067
rect -1468 226227 -1168 243949
rect -1468 226109 -1377 226227
rect -1259 226109 -1168 226227
rect -1468 226067 -1168 226109
rect -1468 225949 -1377 226067
rect -1259 225949 -1168 226067
rect -1468 208227 -1168 225949
rect -1468 208109 -1377 208227
rect -1259 208109 -1168 208227
rect -1468 208067 -1168 208109
rect -1468 207949 -1377 208067
rect -1259 207949 -1168 208067
rect -1468 190227 -1168 207949
rect -1468 190109 -1377 190227
rect -1259 190109 -1168 190227
rect -1468 190067 -1168 190109
rect -1468 189949 -1377 190067
rect -1259 189949 -1168 190067
rect -1468 172227 -1168 189949
rect -1468 172109 -1377 172227
rect -1259 172109 -1168 172227
rect -1468 172067 -1168 172109
rect -1468 171949 -1377 172067
rect -1259 171949 -1168 172067
rect -1468 154227 -1168 171949
rect -1468 154109 -1377 154227
rect -1259 154109 -1168 154227
rect -1468 154067 -1168 154109
rect -1468 153949 -1377 154067
rect -1259 153949 -1168 154067
rect -1468 136227 -1168 153949
rect -1468 136109 -1377 136227
rect -1259 136109 -1168 136227
rect -1468 136067 -1168 136109
rect -1468 135949 -1377 136067
rect -1259 135949 -1168 136067
rect -1468 118227 -1168 135949
rect -1468 118109 -1377 118227
rect -1259 118109 -1168 118227
rect -1468 118067 -1168 118109
rect -1468 117949 -1377 118067
rect -1259 117949 -1168 118067
rect -1468 100227 -1168 117949
rect -1468 100109 -1377 100227
rect -1259 100109 -1168 100227
rect -1468 100067 -1168 100109
rect -1468 99949 -1377 100067
rect -1259 99949 -1168 100067
rect -1468 82227 -1168 99949
rect -1468 82109 -1377 82227
rect -1259 82109 -1168 82227
rect -1468 82067 -1168 82109
rect -1468 81949 -1377 82067
rect -1259 81949 -1168 82067
rect -1468 64227 -1168 81949
rect -1468 64109 -1377 64227
rect -1259 64109 -1168 64227
rect -1468 64067 -1168 64109
rect -1468 63949 -1377 64067
rect -1259 63949 -1168 64067
rect -1468 46227 -1168 63949
rect -1468 46109 -1377 46227
rect -1259 46109 -1168 46227
rect -1468 46067 -1168 46109
rect -1468 45949 -1377 46067
rect -1259 45949 -1168 46067
rect -1468 28227 -1168 45949
rect -1468 28109 -1377 28227
rect -1259 28109 -1168 28227
rect -1468 28067 -1168 28109
rect -1468 27949 -1377 28067
rect -1259 27949 -1168 28067
rect -1468 10227 -1168 27949
rect -1468 10109 -1377 10227
rect -1259 10109 -1168 10227
rect -1468 10067 -1168 10109
rect -1468 9949 -1377 10067
rect -1259 9949 -1168 10067
rect -1468 -643 -1168 9949
rect -998 352419 -698 352430
rect -998 352301 -907 352419
rect -789 352301 -698 352419
rect -998 352259 -698 352301
rect -998 352141 -907 352259
rect -789 352141 -698 352259
rect -998 343227 -698 352141
rect 402 352419 702 352900
rect 402 352301 493 352419
rect 611 352301 702 352419
rect 402 352259 702 352301
rect 402 352141 493 352259
rect 611 352141 702 352259
rect 402 351760 702 352141
rect 2202 351760 2502 353081
rect 4002 351760 4302 354021
rect 5802 351760 6102 354961
rect 14802 355709 15102 355720
rect 14802 355591 14893 355709
rect 15011 355591 15102 355709
rect 14802 355549 15102 355591
rect 14802 355431 14893 355549
rect 15011 355431 15102 355549
rect 13002 354769 13302 354780
rect 13002 354651 13093 354769
rect 13211 354651 13302 354769
rect 13002 354609 13302 354651
rect 13002 354491 13093 354609
rect 13211 354491 13302 354609
rect 11202 353829 11502 353840
rect 11202 353711 11293 353829
rect 11411 353711 11502 353829
rect 11202 353669 11502 353711
rect 11202 353551 11293 353669
rect 11411 353551 11502 353669
rect 9402 352889 9702 352900
rect 9402 352771 9493 352889
rect 9611 352771 9702 352889
rect 9402 352729 9702 352771
rect 9402 352611 9493 352729
rect 9611 352611 9702 352729
rect 9402 351760 9702 352611
rect 11202 351760 11502 353551
rect 13002 351760 13302 354491
rect 14802 351760 15102 355431
rect 23802 355239 24102 355720
rect 23802 355121 23893 355239
rect 24011 355121 24102 355239
rect 23802 355079 24102 355121
rect 23802 354961 23893 355079
rect 24011 354961 24102 355079
rect 22002 354299 22302 354780
rect 22002 354181 22093 354299
rect 22211 354181 22302 354299
rect 22002 354139 22302 354181
rect 22002 354021 22093 354139
rect 22211 354021 22302 354139
rect 20202 353359 20502 353840
rect 20202 353241 20293 353359
rect 20411 353241 20502 353359
rect 20202 353199 20502 353241
rect 20202 353081 20293 353199
rect 20411 353081 20502 353199
rect 18402 352419 18702 352900
rect 18402 352301 18493 352419
rect 18611 352301 18702 352419
rect 18402 352259 18702 352301
rect 18402 352141 18493 352259
rect 18611 352141 18702 352259
rect 18402 351760 18702 352141
rect 20202 351760 20502 353081
rect 22002 351760 22302 354021
rect 23802 351760 24102 354961
rect 32802 355709 33102 355720
rect 32802 355591 32893 355709
rect 33011 355591 33102 355709
rect 32802 355549 33102 355591
rect 32802 355431 32893 355549
rect 33011 355431 33102 355549
rect 31002 354769 31302 354780
rect 31002 354651 31093 354769
rect 31211 354651 31302 354769
rect 31002 354609 31302 354651
rect 31002 354491 31093 354609
rect 31211 354491 31302 354609
rect 29202 353829 29502 353840
rect 29202 353711 29293 353829
rect 29411 353711 29502 353829
rect 29202 353669 29502 353711
rect 29202 353551 29293 353669
rect 29411 353551 29502 353669
rect 27402 352889 27702 352900
rect 27402 352771 27493 352889
rect 27611 352771 27702 352889
rect 27402 352729 27702 352771
rect 27402 352611 27493 352729
rect 27611 352611 27702 352729
rect 27402 351760 27702 352611
rect 29202 351760 29502 353551
rect 31002 351760 31302 354491
rect 32802 351760 33102 355431
rect 41802 355239 42102 355720
rect 41802 355121 41893 355239
rect 42011 355121 42102 355239
rect 41802 355079 42102 355121
rect 41802 354961 41893 355079
rect 42011 354961 42102 355079
rect 40002 354299 40302 354780
rect 40002 354181 40093 354299
rect 40211 354181 40302 354299
rect 40002 354139 40302 354181
rect 40002 354021 40093 354139
rect 40211 354021 40302 354139
rect 38202 353359 38502 353840
rect 38202 353241 38293 353359
rect 38411 353241 38502 353359
rect 38202 353199 38502 353241
rect 38202 353081 38293 353199
rect 38411 353081 38502 353199
rect 36402 352419 36702 352900
rect 36402 352301 36493 352419
rect 36611 352301 36702 352419
rect 36402 352259 36702 352301
rect 36402 352141 36493 352259
rect 36611 352141 36702 352259
rect 36402 351760 36702 352141
rect 38202 351760 38502 353081
rect 40002 351760 40302 354021
rect 41802 351760 42102 354961
rect 50802 355709 51102 355720
rect 50802 355591 50893 355709
rect 51011 355591 51102 355709
rect 50802 355549 51102 355591
rect 50802 355431 50893 355549
rect 51011 355431 51102 355549
rect 49002 354769 49302 354780
rect 49002 354651 49093 354769
rect 49211 354651 49302 354769
rect 49002 354609 49302 354651
rect 49002 354491 49093 354609
rect 49211 354491 49302 354609
rect 47202 353829 47502 353840
rect 47202 353711 47293 353829
rect 47411 353711 47502 353829
rect 47202 353669 47502 353711
rect 47202 353551 47293 353669
rect 47411 353551 47502 353669
rect 45402 352889 45702 352900
rect 45402 352771 45493 352889
rect 45611 352771 45702 352889
rect 45402 352729 45702 352771
rect 45402 352611 45493 352729
rect 45611 352611 45702 352729
rect 45402 351760 45702 352611
rect 47202 351760 47502 353551
rect 49002 351760 49302 354491
rect 50802 351760 51102 355431
rect 59802 355239 60102 355720
rect 59802 355121 59893 355239
rect 60011 355121 60102 355239
rect 59802 355079 60102 355121
rect 59802 354961 59893 355079
rect 60011 354961 60102 355079
rect 58002 354299 58302 354780
rect 58002 354181 58093 354299
rect 58211 354181 58302 354299
rect 58002 354139 58302 354181
rect 58002 354021 58093 354139
rect 58211 354021 58302 354139
rect 56202 353359 56502 353840
rect 56202 353241 56293 353359
rect 56411 353241 56502 353359
rect 56202 353199 56502 353241
rect 56202 353081 56293 353199
rect 56411 353081 56502 353199
rect 54402 352419 54702 352900
rect 54402 352301 54493 352419
rect 54611 352301 54702 352419
rect 54402 352259 54702 352301
rect 54402 352141 54493 352259
rect 54611 352141 54702 352259
rect 54402 351760 54702 352141
rect 56202 351760 56502 353081
rect 58002 351760 58302 354021
rect 59802 351760 60102 354961
rect 68802 355709 69102 355720
rect 68802 355591 68893 355709
rect 69011 355591 69102 355709
rect 68802 355549 69102 355591
rect 68802 355431 68893 355549
rect 69011 355431 69102 355549
rect 67002 354769 67302 354780
rect 67002 354651 67093 354769
rect 67211 354651 67302 354769
rect 67002 354609 67302 354651
rect 67002 354491 67093 354609
rect 67211 354491 67302 354609
rect 65202 353829 65502 353840
rect 65202 353711 65293 353829
rect 65411 353711 65502 353829
rect 65202 353669 65502 353711
rect 65202 353551 65293 353669
rect 65411 353551 65502 353669
rect 63402 352889 63702 352900
rect 63402 352771 63493 352889
rect 63611 352771 63702 352889
rect 63402 352729 63702 352771
rect 63402 352611 63493 352729
rect 63611 352611 63702 352729
rect 63402 351760 63702 352611
rect 65202 351760 65502 353551
rect 67002 351760 67302 354491
rect 68802 351760 69102 355431
rect 77802 355239 78102 355720
rect 77802 355121 77893 355239
rect 78011 355121 78102 355239
rect 77802 355079 78102 355121
rect 77802 354961 77893 355079
rect 78011 354961 78102 355079
rect 76002 354299 76302 354780
rect 76002 354181 76093 354299
rect 76211 354181 76302 354299
rect 76002 354139 76302 354181
rect 76002 354021 76093 354139
rect 76211 354021 76302 354139
rect 74202 353359 74502 353840
rect 74202 353241 74293 353359
rect 74411 353241 74502 353359
rect 74202 353199 74502 353241
rect 74202 353081 74293 353199
rect 74411 353081 74502 353199
rect 72402 352419 72702 352900
rect 72402 352301 72493 352419
rect 72611 352301 72702 352419
rect 72402 352259 72702 352301
rect 72402 352141 72493 352259
rect 72611 352141 72702 352259
rect 72402 351760 72702 352141
rect 74202 351760 74502 353081
rect 76002 351760 76302 354021
rect 77802 351760 78102 354961
rect 86802 355709 87102 355720
rect 86802 355591 86893 355709
rect 87011 355591 87102 355709
rect 86802 355549 87102 355591
rect 86802 355431 86893 355549
rect 87011 355431 87102 355549
rect 85002 354769 85302 354780
rect 85002 354651 85093 354769
rect 85211 354651 85302 354769
rect 85002 354609 85302 354651
rect 85002 354491 85093 354609
rect 85211 354491 85302 354609
rect 83202 353829 83502 353840
rect 83202 353711 83293 353829
rect 83411 353711 83502 353829
rect 83202 353669 83502 353711
rect 83202 353551 83293 353669
rect 83411 353551 83502 353669
rect 81402 352889 81702 352900
rect 81402 352771 81493 352889
rect 81611 352771 81702 352889
rect 81402 352729 81702 352771
rect 81402 352611 81493 352729
rect 81611 352611 81702 352729
rect 81402 351760 81702 352611
rect 83202 351760 83502 353551
rect 85002 351760 85302 354491
rect 86802 351760 87102 355431
rect 95802 355239 96102 355720
rect 95802 355121 95893 355239
rect 96011 355121 96102 355239
rect 95802 355079 96102 355121
rect 95802 354961 95893 355079
rect 96011 354961 96102 355079
rect 94002 354299 94302 354780
rect 94002 354181 94093 354299
rect 94211 354181 94302 354299
rect 94002 354139 94302 354181
rect 94002 354021 94093 354139
rect 94211 354021 94302 354139
rect 92202 353359 92502 353840
rect 92202 353241 92293 353359
rect 92411 353241 92502 353359
rect 92202 353199 92502 353241
rect 92202 353081 92293 353199
rect 92411 353081 92502 353199
rect 90402 352419 90702 352900
rect 90402 352301 90493 352419
rect 90611 352301 90702 352419
rect 90402 352259 90702 352301
rect 90402 352141 90493 352259
rect 90611 352141 90702 352259
rect 90402 351760 90702 352141
rect 92202 351760 92502 353081
rect 94002 351760 94302 354021
rect 95802 351760 96102 354961
rect 104802 355709 105102 355720
rect 104802 355591 104893 355709
rect 105011 355591 105102 355709
rect 104802 355549 105102 355591
rect 104802 355431 104893 355549
rect 105011 355431 105102 355549
rect 103002 354769 103302 354780
rect 103002 354651 103093 354769
rect 103211 354651 103302 354769
rect 103002 354609 103302 354651
rect 103002 354491 103093 354609
rect 103211 354491 103302 354609
rect 101202 353829 101502 353840
rect 101202 353711 101293 353829
rect 101411 353711 101502 353829
rect 101202 353669 101502 353711
rect 101202 353551 101293 353669
rect 101411 353551 101502 353669
rect 99402 352889 99702 352900
rect 99402 352771 99493 352889
rect 99611 352771 99702 352889
rect 99402 352729 99702 352771
rect 99402 352611 99493 352729
rect 99611 352611 99702 352729
rect 99402 351760 99702 352611
rect 101202 351760 101502 353551
rect 103002 351760 103302 354491
rect 104802 351760 105102 355431
rect 113802 355239 114102 355720
rect 113802 355121 113893 355239
rect 114011 355121 114102 355239
rect 113802 355079 114102 355121
rect 113802 354961 113893 355079
rect 114011 354961 114102 355079
rect 112002 354299 112302 354780
rect 112002 354181 112093 354299
rect 112211 354181 112302 354299
rect 112002 354139 112302 354181
rect 112002 354021 112093 354139
rect 112211 354021 112302 354139
rect 110202 353359 110502 353840
rect 110202 353241 110293 353359
rect 110411 353241 110502 353359
rect 110202 353199 110502 353241
rect 110202 353081 110293 353199
rect 110411 353081 110502 353199
rect 108402 352419 108702 352900
rect 108402 352301 108493 352419
rect 108611 352301 108702 352419
rect 108402 352259 108702 352301
rect 108402 352141 108493 352259
rect 108611 352141 108702 352259
rect 108402 351760 108702 352141
rect 110202 351760 110502 353081
rect 112002 351760 112302 354021
rect 113802 351760 114102 354961
rect 122802 355709 123102 355720
rect 122802 355591 122893 355709
rect 123011 355591 123102 355709
rect 122802 355549 123102 355591
rect 122802 355431 122893 355549
rect 123011 355431 123102 355549
rect 121002 354769 121302 354780
rect 121002 354651 121093 354769
rect 121211 354651 121302 354769
rect 121002 354609 121302 354651
rect 121002 354491 121093 354609
rect 121211 354491 121302 354609
rect 119202 353829 119502 353840
rect 119202 353711 119293 353829
rect 119411 353711 119502 353829
rect 119202 353669 119502 353711
rect 119202 353551 119293 353669
rect 119411 353551 119502 353669
rect 117402 352889 117702 352900
rect 117402 352771 117493 352889
rect 117611 352771 117702 352889
rect 117402 352729 117702 352771
rect 117402 352611 117493 352729
rect 117611 352611 117702 352729
rect 117402 351760 117702 352611
rect 119202 351760 119502 353551
rect 121002 351760 121302 354491
rect 122802 351760 123102 355431
rect 131802 355239 132102 355720
rect 131802 355121 131893 355239
rect 132011 355121 132102 355239
rect 131802 355079 132102 355121
rect 131802 354961 131893 355079
rect 132011 354961 132102 355079
rect 130002 354299 130302 354780
rect 130002 354181 130093 354299
rect 130211 354181 130302 354299
rect 130002 354139 130302 354181
rect 130002 354021 130093 354139
rect 130211 354021 130302 354139
rect 128202 353359 128502 353840
rect 128202 353241 128293 353359
rect 128411 353241 128502 353359
rect 128202 353199 128502 353241
rect 128202 353081 128293 353199
rect 128411 353081 128502 353199
rect 126402 352419 126702 352900
rect 126402 352301 126493 352419
rect 126611 352301 126702 352419
rect 126402 352259 126702 352301
rect 126402 352141 126493 352259
rect 126611 352141 126702 352259
rect 126402 351760 126702 352141
rect 128202 351760 128502 353081
rect 130002 351760 130302 354021
rect 131802 351760 132102 354961
rect 140802 355709 141102 355720
rect 140802 355591 140893 355709
rect 141011 355591 141102 355709
rect 140802 355549 141102 355591
rect 140802 355431 140893 355549
rect 141011 355431 141102 355549
rect 139002 354769 139302 354780
rect 139002 354651 139093 354769
rect 139211 354651 139302 354769
rect 139002 354609 139302 354651
rect 139002 354491 139093 354609
rect 139211 354491 139302 354609
rect 137202 353829 137502 353840
rect 137202 353711 137293 353829
rect 137411 353711 137502 353829
rect 137202 353669 137502 353711
rect 137202 353551 137293 353669
rect 137411 353551 137502 353669
rect 135402 352889 135702 352900
rect 135402 352771 135493 352889
rect 135611 352771 135702 352889
rect 135402 352729 135702 352771
rect 135402 352611 135493 352729
rect 135611 352611 135702 352729
rect 135402 351760 135702 352611
rect 137202 351760 137502 353551
rect 139002 351760 139302 354491
rect 140802 351760 141102 355431
rect 149802 355239 150102 355720
rect 149802 355121 149893 355239
rect 150011 355121 150102 355239
rect 149802 355079 150102 355121
rect 149802 354961 149893 355079
rect 150011 354961 150102 355079
rect 148002 354299 148302 354780
rect 148002 354181 148093 354299
rect 148211 354181 148302 354299
rect 148002 354139 148302 354181
rect 148002 354021 148093 354139
rect 148211 354021 148302 354139
rect 146202 353359 146502 353840
rect 146202 353241 146293 353359
rect 146411 353241 146502 353359
rect 146202 353199 146502 353241
rect 146202 353081 146293 353199
rect 146411 353081 146502 353199
rect 144402 352419 144702 352900
rect 144402 352301 144493 352419
rect 144611 352301 144702 352419
rect 144402 352259 144702 352301
rect 144402 352141 144493 352259
rect 144611 352141 144702 352259
rect 144402 351760 144702 352141
rect 146202 351760 146502 353081
rect 148002 351760 148302 354021
rect 149802 351760 150102 354961
rect 158802 355709 159102 355720
rect 158802 355591 158893 355709
rect 159011 355591 159102 355709
rect 158802 355549 159102 355591
rect 158802 355431 158893 355549
rect 159011 355431 159102 355549
rect 157002 354769 157302 354780
rect 157002 354651 157093 354769
rect 157211 354651 157302 354769
rect 157002 354609 157302 354651
rect 157002 354491 157093 354609
rect 157211 354491 157302 354609
rect 155202 353829 155502 353840
rect 155202 353711 155293 353829
rect 155411 353711 155502 353829
rect 155202 353669 155502 353711
rect 155202 353551 155293 353669
rect 155411 353551 155502 353669
rect 153402 352889 153702 352900
rect 153402 352771 153493 352889
rect 153611 352771 153702 352889
rect 153402 352729 153702 352771
rect 153402 352611 153493 352729
rect 153611 352611 153702 352729
rect 153402 351760 153702 352611
rect 155202 351760 155502 353551
rect 157002 351760 157302 354491
rect 158802 351760 159102 355431
rect 167802 355239 168102 355720
rect 167802 355121 167893 355239
rect 168011 355121 168102 355239
rect 167802 355079 168102 355121
rect 167802 354961 167893 355079
rect 168011 354961 168102 355079
rect 166002 354299 166302 354780
rect 166002 354181 166093 354299
rect 166211 354181 166302 354299
rect 166002 354139 166302 354181
rect 166002 354021 166093 354139
rect 166211 354021 166302 354139
rect 164202 353359 164502 353840
rect 164202 353241 164293 353359
rect 164411 353241 164502 353359
rect 164202 353199 164502 353241
rect 164202 353081 164293 353199
rect 164411 353081 164502 353199
rect 162402 352419 162702 352900
rect 162402 352301 162493 352419
rect 162611 352301 162702 352419
rect 162402 352259 162702 352301
rect 162402 352141 162493 352259
rect 162611 352141 162702 352259
rect 162402 351760 162702 352141
rect 164202 351760 164502 353081
rect 166002 351760 166302 354021
rect 167802 351760 168102 354961
rect 176802 355709 177102 355720
rect 176802 355591 176893 355709
rect 177011 355591 177102 355709
rect 176802 355549 177102 355591
rect 176802 355431 176893 355549
rect 177011 355431 177102 355549
rect 175002 354769 175302 354780
rect 175002 354651 175093 354769
rect 175211 354651 175302 354769
rect 175002 354609 175302 354651
rect 175002 354491 175093 354609
rect 175211 354491 175302 354609
rect 173202 353829 173502 353840
rect 173202 353711 173293 353829
rect 173411 353711 173502 353829
rect 173202 353669 173502 353711
rect 173202 353551 173293 353669
rect 173411 353551 173502 353669
rect 171402 352889 171702 352900
rect 171402 352771 171493 352889
rect 171611 352771 171702 352889
rect 171402 352729 171702 352771
rect 171402 352611 171493 352729
rect 171611 352611 171702 352729
rect 171402 351760 171702 352611
rect 173202 351760 173502 353551
rect 175002 351760 175302 354491
rect 176802 351760 177102 355431
rect 185802 355239 186102 355720
rect 185802 355121 185893 355239
rect 186011 355121 186102 355239
rect 185802 355079 186102 355121
rect 185802 354961 185893 355079
rect 186011 354961 186102 355079
rect 184002 354299 184302 354780
rect 184002 354181 184093 354299
rect 184211 354181 184302 354299
rect 184002 354139 184302 354181
rect 184002 354021 184093 354139
rect 184211 354021 184302 354139
rect 182202 353359 182502 353840
rect 182202 353241 182293 353359
rect 182411 353241 182502 353359
rect 182202 353199 182502 353241
rect 182202 353081 182293 353199
rect 182411 353081 182502 353199
rect 180402 352419 180702 352900
rect 180402 352301 180493 352419
rect 180611 352301 180702 352419
rect 180402 352259 180702 352301
rect 180402 352141 180493 352259
rect 180611 352141 180702 352259
rect 180402 351760 180702 352141
rect 182202 351760 182502 353081
rect 184002 351760 184302 354021
rect 185802 351760 186102 354961
rect 194802 355709 195102 355720
rect 194802 355591 194893 355709
rect 195011 355591 195102 355709
rect 194802 355549 195102 355591
rect 194802 355431 194893 355549
rect 195011 355431 195102 355549
rect 193002 354769 193302 354780
rect 193002 354651 193093 354769
rect 193211 354651 193302 354769
rect 193002 354609 193302 354651
rect 193002 354491 193093 354609
rect 193211 354491 193302 354609
rect 191202 353829 191502 353840
rect 191202 353711 191293 353829
rect 191411 353711 191502 353829
rect 191202 353669 191502 353711
rect 191202 353551 191293 353669
rect 191411 353551 191502 353669
rect 189402 352889 189702 352900
rect 189402 352771 189493 352889
rect 189611 352771 189702 352889
rect 189402 352729 189702 352771
rect 189402 352611 189493 352729
rect 189611 352611 189702 352729
rect 189402 351760 189702 352611
rect 191202 351760 191502 353551
rect 193002 351760 193302 354491
rect 194802 351760 195102 355431
rect 203802 355239 204102 355720
rect 203802 355121 203893 355239
rect 204011 355121 204102 355239
rect 203802 355079 204102 355121
rect 203802 354961 203893 355079
rect 204011 354961 204102 355079
rect 202002 354299 202302 354780
rect 202002 354181 202093 354299
rect 202211 354181 202302 354299
rect 202002 354139 202302 354181
rect 202002 354021 202093 354139
rect 202211 354021 202302 354139
rect 200202 353359 200502 353840
rect 200202 353241 200293 353359
rect 200411 353241 200502 353359
rect 200202 353199 200502 353241
rect 200202 353081 200293 353199
rect 200411 353081 200502 353199
rect 198402 352419 198702 352900
rect 198402 352301 198493 352419
rect 198611 352301 198702 352419
rect 198402 352259 198702 352301
rect 198402 352141 198493 352259
rect 198611 352141 198702 352259
rect 198402 351760 198702 352141
rect 200202 351760 200502 353081
rect 202002 351760 202302 354021
rect 203802 351760 204102 354961
rect 212802 355709 213102 355720
rect 212802 355591 212893 355709
rect 213011 355591 213102 355709
rect 212802 355549 213102 355591
rect 212802 355431 212893 355549
rect 213011 355431 213102 355549
rect 211002 354769 211302 354780
rect 211002 354651 211093 354769
rect 211211 354651 211302 354769
rect 211002 354609 211302 354651
rect 211002 354491 211093 354609
rect 211211 354491 211302 354609
rect 209202 353829 209502 353840
rect 209202 353711 209293 353829
rect 209411 353711 209502 353829
rect 209202 353669 209502 353711
rect 209202 353551 209293 353669
rect 209411 353551 209502 353669
rect 207402 352889 207702 352900
rect 207402 352771 207493 352889
rect 207611 352771 207702 352889
rect 207402 352729 207702 352771
rect 207402 352611 207493 352729
rect 207611 352611 207702 352729
rect 207402 351760 207702 352611
rect 209202 351760 209502 353551
rect 211002 351760 211302 354491
rect 212802 351760 213102 355431
rect 221802 355239 222102 355720
rect 221802 355121 221893 355239
rect 222011 355121 222102 355239
rect 221802 355079 222102 355121
rect 221802 354961 221893 355079
rect 222011 354961 222102 355079
rect 220002 354299 220302 354780
rect 220002 354181 220093 354299
rect 220211 354181 220302 354299
rect 220002 354139 220302 354181
rect 220002 354021 220093 354139
rect 220211 354021 220302 354139
rect 218202 353359 218502 353840
rect 218202 353241 218293 353359
rect 218411 353241 218502 353359
rect 218202 353199 218502 353241
rect 218202 353081 218293 353199
rect 218411 353081 218502 353199
rect 216402 352419 216702 352900
rect 216402 352301 216493 352419
rect 216611 352301 216702 352419
rect 216402 352259 216702 352301
rect 216402 352141 216493 352259
rect 216611 352141 216702 352259
rect 216402 351760 216702 352141
rect 218202 351760 218502 353081
rect 220002 351760 220302 354021
rect 221802 351760 222102 354961
rect 230802 355709 231102 355720
rect 230802 355591 230893 355709
rect 231011 355591 231102 355709
rect 230802 355549 231102 355591
rect 230802 355431 230893 355549
rect 231011 355431 231102 355549
rect 229002 354769 229302 354780
rect 229002 354651 229093 354769
rect 229211 354651 229302 354769
rect 229002 354609 229302 354651
rect 229002 354491 229093 354609
rect 229211 354491 229302 354609
rect 227202 353829 227502 353840
rect 227202 353711 227293 353829
rect 227411 353711 227502 353829
rect 227202 353669 227502 353711
rect 227202 353551 227293 353669
rect 227411 353551 227502 353669
rect 225402 352889 225702 352900
rect 225402 352771 225493 352889
rect 225611 352771 225702 352889
rect 225402 352729 225702 352771
rect 225402 352611 225493 352729
rect 225611 352611 225702 352729
rect 225402 351760 225702 352611
rect 227202 351760 227502 353551
rect 229002 351760 229302 354491
rect 230802 351760 231102 355431
rect 239802 355239 240102 355720
rect 239802 355121 239893 355239
rect 240011 355121 240102 355239
rect 239802 355079 240102 355121
rect 239802 354961 239893 355079
rect 240011 354961 240102 355079
rect 238002 354299 238302 354780
rect 238002 354181 238093 354299
rect 238211 354181 238302 354299
rect 238002 354139 238302 354181
rect 238002 354021 238093 354139
rect 238211 354021 238302 354139
rect 236202 353359 236502 353840
rect 236202 353241 236293 353359
rect 236411 353241 236502 353359
rect 236202 353199 236502 353241
rect 236202 353081 236293 353199
rect 236411 353081 236502 353199
rect 234402 352419 234702 352900
rect 234402 352301 234493 352419
rect 234611 352301 234702 352419
rect 234402 352259 234702 352301
rect 234402 352141 234493 352259
rect 234611 352141 234702 352259
rect 234402 351760 234702 352141
rect 236202 351760 236502 353081
rect 238002 351760 238302 354021
rect 239802 351760 240102 354961
rect 248802 355709 249102 355720
rect 248802 355591 248893 355709
rect 249011 355591 249102 355709
rect 248802 355549 249102 355591
rect 248802 355431 248893 355549
rect 249011 355431 249102 355549
rect 247002 354769 247302 354780
rect 247002 354651 247093 354769
rect 247211 354651 247302 354769
rect 247002 354609 247302 354651
rect 247002 354491 247093 354609
rect 247211 354491 247302 354609
rect 245202 353829 245502 353840
rect 245202 353711 245293 353829
rect 245411 353711 245502 353829
rect 245202 353669 245502 353711
rect 245202 353551 245293 353669
rect 245411 353551 245502 353669
rect 243402 352889 243702 352900
rect 243402 352771 243493 352889
rect 243611 352771 243702 352889
rect 243402 352729 243702 352771
rect 243402 352611 243493 352729
rect 243611 352611 243702 352729
rect 243402 351760 243702 352611
rect 245202 351760 245502 353551
rect 247002 351760 247302 354491
rect 248802 351760 249102 355431
rect 257802 355239 258102 355720
rect 257802 355121 257893 355239
rect 258011 355121 258102 355239
rect 257802 355079 258102 355121
rect 257802 354961 257893 355079
rect 258011 354961 258102 355079
rect 256002 354299 256302 354780
rect 256002 354181 256093 354299
rect 256211 354181 256302 354299
rect 256002 354139 256302 354181
rect 256002 354021 256093 354139
rect 256211 354021 256302 354139
rect 254202 353359 254502 353840
rect 254202 353241 254293 353359
rect 254411 353241 254502 353359
rect 254202 353199 254502 353241
rect 254202 353081 254293 353199
rect 254411 353081 254502 353199
rect 252402 352419 252702 352900
rect 252402 352301 252493 352419
rect 252611 352301 252702 352419
rect 252402 352259 252702 352301
rect 252402 352141 252493 352259
rect 252611 352141 252702 352259
rect 252402 351760 252702 352141
rect 254202 351760 254502 353081
rect 256002 351760 256302 354021
rect 257802 351760 258102 354961
rect 266802 355709 267102 355720
rect 266802 355591 266893 355709
rect 267011 355591 267102 355709
rect 266802 355549 267102 355591
rect 266802 355431 266893 355549
rect 267011 355431 267102 355549
rect 265002 354769 265302 354780
rect 265002 354651 265093 354769
rect 265211 354651 265302 354769
rect 265002 354609 265302 354651
rect 265002 354491 265093 354609
rect 265211 354491 265302 354609
rect 263202 353829 263502 353840
rect 263202 353711 263293 353829
rect 263411 353711 263502 353829
rect 263202 353669 263502 353711
rect 263202 353551 263293 353669
rect 263411 353551 263502 353669
rect 261402 352889 261702 352900
rect 261402 352771 261493 352889
rect 261611 352771 261702 352889
rect 261402 352729 261702 352771
rect 261402 352611 261493 352729
rect 261611 352611 261702 352729
rect 261402 351760 261702 352611
rect 263202 351760 263502 353551
rect 265002 351760 265302 354491
rect 266802 351760 267102 355431
rect 275802 355239 276102 355720
rect 275802 355121 275893 355239
rect 276011 355121 276102 355239
rect 275802 355079 276102 355121
rect 275802 354961 275893 355079
rect 276011 354961 276102 355079
rect 274002 354299 274302 354780
rect 274002 354181 274093 354299
rect 274211 354181 274302 354299
rect 274002 354139 274302 354181
rect 274002 354021 274093 354139
rect 274211 354021 274302 354139
rect 272202 353359 272502 353840
rect 272202 353241 272293 353359
rect 272411 353241 272502 353359
rect 272202 353199 272502 353241
rect 272202 353081 272293 353199
rect 272411 353081 272502 353199
rect 270402 352419 270702 352900
rect 270402 352301 270493 352419
rect 270611 352301 270702 352419
rect 270402 352259 270702 352301
rect 270402 352141 270493 352259
rect 270611 352141 270702 352259
rect 270402 351760 270702 352141
rect 272202 351760 272502 353081
rect 274002 351760 274302 354021
rect 275802 351760 276102 354961
rect 284802 355709 285102 355720
rect 284802 355591 284893 355709
rect 285011 355591 285102 355709
rect 284802 355549 285102 355591
rect 284802 355431 284893 355549
rect 285011 355431 285102 355549
rect 283002 354769 283302 354780
rect 283002 354651 283093 354769
rect 283211 354651 283302 354769
rect 283002 354609 283302 354651
rect 283002 354491 283093 354609
rect 283211 354491 283302 354609
rect 281202 353829 281502 353840
rect 281202 353711 281293 353829
rect 281411 353711 281502 353829
rect 281202 353669 281502 353711
rect 281202 353551 281293 353669
rect 281411 353551 281502 353669
rect 279402 352889 279702 352900
rect 279402 352771 279493 352889
rect 279611 352771 279702 352889
rect 279402 352729 279702 352771
rect 279402 352611 279493 352729
rect 279611 352611 279702 352729
rect 279402 351760 279702 352611
rect 281202 351760 281502 353551
rect 283002 351760 283302 354491
rect 284802 351760 285102 355431
rect 295950 355709 296250 355720
rect 295950 355591 296041 355709
rect 296159 355591 296250 355709
rect 295950 355549 296250 355591
rect 295950 355431 296041 355549
rect 296159 355431 296250 355549
rect 295480 355239 295780 355250
rect 295480 355121 295571 355239
rect 295689 355121 295780 355239
rect 295480 355079 295780 355121
rect 295480 354961 295571 355079
rect 295689 354961 295780 355079
rect 295010 354769 295310 354780
rect 295010 354651 295101 354769
rect 295219 354651 295310 354769
rect 295010 354609 295310 354651
rect 295010 354491 295101 354609
rect 295219 354491 295310 354609
rect 294540 354299 294840 354310
rect 294540 354181 294631 354299
rect 294749 354181 294840 354299
rect 294540 354139 294840 354181
rect 294540 354021 294631 354139
rect 294749 354021 294840 354139
rect 290202 353359 290502 353840
rect 294070 353829 294370 353840
rect 294070 353711 294161 353829
rect 294279 353711 294370 353829
rect 294070 353669 294370 353711
rect 294070 353551 294161 353669
rect 294279 353551 294370 353669
rect 290202 353241 290293 353359
rect 290411 353241 290502 353359
rect 290202 353199 290502 353241
rect 290202 353081 290293 353199
rect 290411 353081 290502 353199
rect 288402 352419 288702 352900
rect 288402 352301 288493 352419
rect 288611 352301 288702 352419
rect 288402 352259 288702 352301
rect 288402 352141 288493 352259
rect 288611 352141 288702 352259
rect 288402 351760 288702 352141
rect 290202 351760 290502 353081
rect 293600 353359 293900 353370
rect 293600 353241 293691 353359
rect 293809 353241 293900 353359
rect 293600 353199 293900 353241
rect 293600 353081 293691 353199
rect 293809 353081 293900 353199
rect 293130 352889 293430 352900
rect 293130 352771 293221 352889
rect 293339 352771 293430 352889
rect 293130 352729 293430 352771
rect 293130 352611 293221 352729
rect 293339 352611 293430 352729
rect 292660 352419 292960 352430
rect 292660 352301 292751 352419
rect 292869 352301 292960 352419
rect 292660 352259 292960 352301
rect 292660 352141 292751 352259
rect 292869 352141 292960 352259
rect -998 343109 -907 343227
rect -789 343109 -698 343227
rect -998 343067 -698 343109
rect -998 342949 -907 343067
rect -789 342949 -698 343067
rect -998 325227 -698 342949
rect -998 325109 -907 325227
rect -789 325109 -698 325227
rect -998 325067 -698 325109
rect -998 324949 -907 325067
rect -789 324949 -698 325067
rect -998 307227 -698 324949
rect -998 307109 -907 307227
rect -789 307109 -698 307227
rect -998 307067 -698 307109
rect -998 306949 -907 307067
rect -789 306949 -698 307067
rect -998 289227 -698 306949
rect -998 289109 -907 289227
rect -789 289109 -698 289227
rect -998 289067 -698 289109
rect -998 288949 -907 289067
rect -789 288949 -698 289067
rect -998 271227 -698 288949
rect -998 271109 -907 271227
rect -789 271109 -698 271227
rect -998 271067 -698 271109
rect -998 270949 -907 271067
rect -789 270949 -698 271067
rect -998 253227 -698 270949
rect -998 253109 -907 253227
rect -789 253109 -698 253227
rect -998 253067 -698 253109
rect -998 252949 -907 253067
rect -789 252949 -698 253067
rect -998 235227 -698 252949
rect -998 235109 -907 235227
rect -789 235109 -698 235227
rect -998 235067 -698 235109
rect -998 234949 -907 235067
rect -789 234949 -698 235067
rect -998 217227 -698 234949
rect -998 217109 -907 217227
rect -789 217109 -698 217227
rect -998 217067 -698 217109
rect -998 216949 -907 217067
rect -789 216949 -698 217067
rect -998 199227 -698 216949
rect -998 199109 -907 199227
rect -789 199109 -698 199227
rect -998 199067 -698 199109
rect -998 198949 -907 199067
rect -789 198949 -698 199067
rect -998 181227 -698 198949
rect -998 181109 -907 181227
rect -789 181109 -698 181227
rect -998 181067 -698 181109
rect -998 180949 -907 181067
rect -789 180949 -698 181067
rect -998 163227 -698 180949
rect -998 163109 -907 163227
rect -789 163109 -698 163227
rect -998 163067 -698 163109
rect -998 162949 -907 163067
rect -789 162949 -698 163067
rect -998 145227 -698 162949
rect -998 145109 -907 145227
rect -789 145109 -698 145227
rect -998 145067 -698 145109
rect -998 144949 -907 145067
rect -789 144949 -698 145067
rect -998 127227 -698 144949
rect -998 127109 -907 127227
rect -789 127109 -698 127227
rect -998 127067 -698 127109
rect -998 126949 -907 127067
rect -789 126949 -698 127067
rect -998 109227 -698 126949
rect -998 109109 -907 109227
rect -789 109109 -698 109227
rect -998 109067 -698 109109
rect -998 108949 -907 109067
rect -789 108949 -698 109067
rect -998 91227 -698 108949
rect -998 91109 -907 91227
rect -789 91109 -698 91227
rect -998 91067 -698 91109
rect -998 90949 -907 91067
rect -789 90949 -698 91067
rect -998 73227 -698 90949
rect -998 73109 -907 73227
rect -789 73109 -698 73227
rect -998 73067 -698 73109
rect -998 72949 -907 73067
rect -789 72949 -698 73067
rect -998 55227 -698 72949
rect -998 55109 -907 55227
rect -789 55109 -698 55227
rect -998 55067 -698 55109
rect -998 54949 -907 55067
rect -789 54949 -698 55067
rect -998 37227 -698 54949
rect -998 37109 -907 37227
rect -789 37109 -698 37227
rect -998 37067 -698 37109
rect -998 36949 -907 37067
rect -789 36949 -698 37067
rect -998 19227 -698 36949
rect -998 19109 -907 19227
rect -789 19109 -698 19227
rect -998 19067 -698 19109
rect -998 18949 -907 19067
rect -789 18949 -698 19067
rect -998 1227 -698 18949
rect -998 1109 -907 1227
rect -789 1109 -698 1227
rect -998 1067 -698 1109
rect -998 949 -907 1067
rect -789 949 -698 1067
rect -998 -173 -698 949
rect 292660 343227 292960 352141
rect 292660 343109 292751 343227
rect 292869 343109 292960 343227
rect 292660 343067 292960 343109
rect 292660 342949 292751 343067
rect 292869 342949 292960 343067
rect 292660 325227 292960 342949
rect 292660 325109 292751 325227
rect 292869 325109 292960 325227
rect 292660 325067 292960 325109
rect 292660 324949 292751 325067
rect 292869 324949 292960 325067
rect 292660 307227 292960 324949
rect 292660 307109 292751 307227
rect 292869 307109 292960 307227
rect 292660 307067 292960 307109
rect 292660 306949 292751 307067
rect 292869 306949 292960 307067
rect 292660 289227 292960 306949
rect 292660 289109 292751 289227
rect 292869 289109 292960 289227
rect 292660 289067 292960 289109
rect 292660 288949 292751 289067
rect 292869 288949 292960 289067
rect 292660 271227 292960 288949
rect 292660 271109 292751 271227
rect 292869 271109 292960 271227
rect 292660 271067 292960 271109
rect 292660 270949 292751 271067
rect 292869 270949 292960 271067
rect 292660 253227 292960 270949
rect 292660 253109 292751 253227
rect 292869 253109 292960 253227
rect 292660 253067 292960 253109
rect 292660 252949 292751 253067
rect 292869 252949 292960 253067
rect 292660 235227 292960 252949
rect 292660 235109 292751 235227
rect 292869 235109 292960 235227
rect 292660 235067 292960 235109
rect 292660 234949 292751 235067
rect 292869 234949 292960 235067
rect 292660 217227 292960 234949
rect 292660 217109 292751 217227
rect 292869 217109 292960 217227
rect 292660 217067 292960 217109
rect 292660 216949 292751 217067
rect 292869 216949 292960 217067
rect 292660 199227 292960 216949
rect 292660 199109 292751 199227
rect 292869 199109 292960 199227
rect 292660 199067 292960 199109
rect 292660 198949 292751 199067
rect 292869 198949 292960 199067
rect 292660 181227 292960 198949
rect 292660 181109 292751 181227
rect 292869 181109 292960 181227
rect 292660 181067 292960 181109
rect 292660 180949 292751 181067
rect 292869 180949 292960 181067
rect 292660 163227 292960 180949
rect 292660 163109 292751 163227
rect 292869 163109 292960 163227
rect 292660 163067 292960 163109
rect 292660 162949 292751 163067
rect 292869 162949 292960 163067
rect 292660 145227 292960 162949
rect 292660 145109 292751 145227
rect 292869 145109 292960 145227
rect 292660 145067 292960 145109
rect 292660 144949 292751 145067
rect 292869 144949 292960 145067
rect 292660 127227 292960 144949
rect 292660 127109 292751 127227
rect 292869 127109 292960 127227
rect 292660 127067 292960 127109
rect 292660 126949 292751 127067
rect 292869 126949 292960 127067
rect 292660 109227 292960 126949
rect 292660 109109 292751 109227
rect 292869 109109 292960 109227
rect 292660 109067 292960 109109
rect 292660 108949 292751 109067
rect 292869 108949 292960 109067
rect 292660 91227 292960 108949
rect 292660 91109 292751 91227
rect 292869 91109 292960 91227
rect 292660 91067 292960 91109
rect 292660 90949 292751 91067
rect 292869 90949 292960 91067
rect 292660 73227 292960 90949
rect 292660 73109 292751 73227
rect 292869 73109 292960 73227
rect 292660 73067 292960 73109
rect 292660 72949 292751 73067
rect 292869 72949 292960 73067
rect 292660 55227 292960 72949
rect 292660 55109 292751 55227
rect 292869 55109 292960 55227
rect 292660 55067 292960 55109
rect 292660 54949 292751 55067
rect 292869 54949 292960 55067
rect 292660 37227 292960 54949
rect 292660 37109 292751 37227
rect 292869 37109 292960 37227
rect 292660 37067 292960 37109
rect 292660 36949 292751 37067
rect 292869 36949 292960 37067
rect 292660 19227 292960 36949
rect 292660 19109 292751 19227
rect 292869 19109 292960 19227
rect 292660 19067 292960 19109
rect 292660 18949 292751 19067
rect 292869 18949 292960 19067
rect 292660 1227 292960 18949
rect 292660 1109 292751 1227
rect 292869 1109 292960 1227
rect 292660 1067 292960 1109
rect 292660 949 292751 1067
rect 292869 949 292960 1067
rect -998 -291 -907 -173
rect -789 -291 -698 -173
rect -998 -333 -698 -291
rect -998 -451 -907 -333
rect -789 -451 -698 -333
rect -998 -462 -698 -451
rect 402 -173 702 240
rect 402 -291 493 -173
rect 611 -291 702 -173
rect 402 -333 702 -291
rect 402 -451 493 -333
rect 611 -451 702 -333
rect -1468 -761 -1377 -643
rect -1259 -761 -1168 -643
rect -1468 -803 -1168 -761
rect -1468 -921 -1377 -803
rect -1259 -921 -1168 -803
rect -1468 -932 -1168 -921
rect 402 -932 702 -451
rect -1938 -1231 -1847 -1113
rect -1729 -1231 -1638 -1113
rect -1938 -1273 -1638 -1231
rect -1938 -1391 -1847 -1273
rect -1729 -1391 -1638 -1273
rect -1938 -1402 -1638 -1391
rect 2202 -1113 2502 240
rect 2202 -1231 2293 -1113
rect 2411 -1231 2502 -1113
rect 2202 -1273 2502 -1231
rect 2202 -1391 2293 -1273
rect 2411 -1391 2502 -1273
rect -2408 -1701 -2317 -1583
rect -2199 -1701 -2108 -1583
rect -2408 -1743 -2108 -1701
rect -2408 -1861 -2317 -1743
rect -2199 -1861 -2108 -1743
rect -2408 -1872 -2108 -1861
rect 2202 -1872 2502 -1391
rect -2878 -2171 -2787 -2053
rect -2669 -2171 -2578 -2053
rect -2878 -2213 -2578 -2171
rect -2878 -2331 -2787 -2213
rect -2669 -2331 -2578 -2213
rect -2878 -2342 -2578 -2331
rect 4002 -2053 4302 240
rect 4002 -2171 4093 -2053
rect 4211 -2171 4302 -2053
rect 4002 -2213 4302 -2171
rect 4002 -2331 4093 -2213
rect 4211 -2331 4302 -2213
rect -3348 -2641 -3257 -2523
rect -3139 -2641 -3048 -2523
rect -3348 -2683 -3048 -2641
rect -3348 -2801 -3257 -2683
rect -3139 -2801 -3048 -2683
rect -3348 -2812 -3048 -2801
rect 4002 -2812 4302 -2331
rect -3818 -3111 -3727 -2993
rect -3609 -3111 -3518 -2993
rect -3818 -3153 -3518 -3111
rect -3818 -3271 -3727 -3153
rect -3609 -3271 -3518 -3153
rect -3818 -3282 -3518 -3271
rect 5802 -2993 6102 240
rect 9402 -643 9702 240
rect 9402 -761 9493 -643
rect 9611 -761 9702 -643
rect 9402 -803 9702 -761
rect 9402 -921 9493 -803
rect 9611 -921 9702 -803
rect 9402 -932 9702 -921
rect 11202 -1583 11502 240
rect 11202 -1701 11293 -1583
rect 11411 -1701 11502 -1583
rect 11202 -1743 11502 -1701
rect 11202 -1861 11293 -1743
rect 11411 -1861 11502 -1743
rect 11202 -1872 11502 -1861
rect 13002 -2523 13302 240
rect 13002 -2641 13093 -2523
rect 13211 -2641 13302 -2523
rect 13002 -2683 13302 -2641
rect 13002 -2801 13093 -2683
rect 13211 -2801 13302 -2683
rect 13002 -2812 13302 -2801
rect 5802 -3111 5893 -2993
rect 6011 -3111 6102 -2993
rect 5802 -3153 6102 -3111
rect 5802 -3271 5893 -3153
rect 6011 -3271 6102 -3153
rect -4288 -3581 -4197 -3463
rect -4079 -3581 -3988 -3463
rect -4288 -3623 -3988 -3581
rect -4288 -3741 -4197 -3623
rect -4079 -3741 -3988 -3623
rect -4288 -3752 -3988 -3741
rect 5802 -3752 6102 -3271
rect 14802 -3463 15102 240
rect 18402 -173 18702 240
rect 18402 -291 18493 -173
rect 18611 -291 18702 -173
rect 18402 -333 18702 -291
rect 18402 -451 18493 -333
rect 18611 -451 18702 -333
rect 18402 -932 18702 -451
rect 20202 -1113 20502 240
rect 20202 -1231 20293 -1113
rect 20411 -1231 20502 -1113
rect 20202 -1273 20502 -1231
rect 20202 -1391 20293 -1273
rect 20411 -1391 20502 -1273
rect 20202 -1872 20502 -1391
rect 22002 -2053 22302 240
rect 22002 -2171 22093 -2053
rect 22211 -2171 22302 -2053
rect 22002 -2213 22302 -2171
rect 22002 -2331 22093 -2213
rect 22211 -2331 22302 -2213
rect 22002 -2812 22302 -2331
rect 14802 -3581 14893 -3463
rect 15011 -3581 15102 -3463
rect 14802 -3623 15102 -3581
rect 14802 -3741 14893 -3623
rect 15011 -3741 15102 -3623
rect 14802 -3752 15102 -3741
rect 23802 -2993 24102 240
rect 27402 -643 27702 240
rect 27402 -761 27493 -643
rect 27611 -761 27702 -643
rect 27402 -803 27702 -761
rect 27402 -921 27493 -803
rect 27611 -921 27702 -803
rect 27402 -932 27702 -921
rect 29202 -1583 29502 240
rect 29202 -1701 29293 -1583
rect 29411 -1701 29502 -1583
rect 29202 -1743 29502 -1701
rect 29202 -1861 29293 -1743
rect 29411 -1861 29502 -1743
rect 29202 -1872 29502 -1861
rect 31002 -2523 31302 240
rect 31002 -2641 31093 -2523
rect 31211 -2641 31302 -2523
rect 31002 -2683 31302 -2641
rect 31002 -2801 31093 -2683
rect 31211 -2801 31302 -2683
rect 31002 -2812 31302 -2801
rect 23802 -3111 23893 -2993
rect 24011 -3111 24102 -2993
rect 23802 -3153 24102 -3111
rect 23802 -3271 23893 -3153
rect 24011 -3271 24102 -3153
rect 23802 -3752 24102 -3271
rect 32802 -3463 33102 240
rect 36402 -173 36702 240
rect 36402 -291 36493 -173
rect 36611 -291 36702 -173
rect 36402 -333 36702 -291
rect 36402 -451 36493 -333
rect 36611 -451 36702 -333
rect 36402 -932 36702 -451
rect 38202 -1113 38502 240
rect 38202 -1231 38293 -1113
rect 38411 -1231 38502 -1113
rect 38202 -1273 38502 -1231
rect 38202 -1391 38293 -1273
rect 38411 -1391 38502 -1273
rect 38202 -1872 38502 -1391
rect 40002 -2053 40302 240
rect 40002 -2171 40093 -2053
rect 40211 -2171 40302 -2053
rect 40002 -2213 40302 -2171
rect 40002 -2331 40093 -2213
rect 40211 -2331 40302 -2213
rect 40002 -2812 40302 -2331
rect 32802 -3581 32893 -3463
rect 33011 -3581 33102 -3463
rect 32802 -3623 33102 -3581
rect 32802 -3741 32893 -3623
rect 33011 -3741 33102 -3623
rect 32802 -3752 33102 -3741
rect 41802 -2993 42102 240
rect 45402 -643 45702 240
rect 45402 -761 45493 -643
rect 45611 -761 45702 -643
rect 45402 -803 45702 -761
rect 45402 -921 45493 -803
rect 45611 -921 45702 -803
rect 45402 -932 45702 -921
rect 47202 -1583 47502 240
rect 47202 -1701 47293 -1583
rect 47411 -1701 47502 -1583
rect 47202 -1743 47502 -1701
rect 47202 -1861 47293 -1743
rect 47411 -1861 47502 -1743
rect 47202 -1872 47502 -1861
rect 49002 -2523 49302 240
rect 49002 -2641 49093 -2523
rect 49211 -2641 49302 -2523
rect 49002 -2683 49302 -2641
rect 49002 -2801 49093 -2683
rect 49211 -2801 49302 -2683
rect 49002 -2812 49302 -2801
rect 41802 -3111 41893 -2993
rect 42011 -3111 42102 -2993
rect 41802 -3153 42102 -3111
rect 41802 -3271 41893 -3153
rect 42011 -3271 42102 -3153
rect 41802 -3752 42102 -3271
rect 50802 -3463 51102 240
rect 54402 -173 54702 240
rect 54402 -291 54493 -173
rect 54611 -291 54702 -173
rect 54402 -333 54702 -291
rect 54402 -451 54493 -333
rect 54611 -451 54702 -333
rect 54402 -932 54702 -451
rect 56202 -1113 56502 240
rect 56202 -1231 56293 -1113
rect 56411 -1231 56502 -1113
rect 56202 -1273 56502 -1231
rect 56202 -1391 56293 -1273
rect 56411 -1391 56502 -1273
rect 56202 -1872 56502 -1391
rect 58002 -2053 58302 240
rect 58002 -2171 58093 -2053
rect 58211 -2171 58302 -2053
rect 58002 -2213 58302 -2171
rect 58002 -2331 58093 -2213
rect 58211 -2331 58302 -2213
rect 58002 -2812 58302 -2331
rect 50802 -3581 50893 -3463
rect 51011 -3581 51102 -3463
rect 50802 -3623 51102 -3581
rect 50802 -3741 50893 -3623
rect 51011 -3741 51102 -3623
rect 50802 -3752 51102 -3741
rect 59802 -2993 60102 240
rect 63402 -643 63702 240
rect 63402 -761 63493 -643
rect 63611 -761 63702 -643
rect 63402 -803 63702 -761
rect 63402 -921 63493 -803
rect 63611 -921 63702 -803
rect 63402 -932 63702 -921
rect 65202 -1583 65502 240
rect 65202 -1701 65293 -1583
rect 65411 -1701 65502 -1583
rect 65202 -1743 65502 -1701
rect 65202 -1861 65293 -1743
rect 65411 -1861 65502 -1743
rect 65202 -1872 65502 -1861
rect 67002 -2523 67302 240
rect 67002 -2641 67093 -2523
rect 67211 -2641 67302 -2523
rect 67002 -2683 67302 -2641
rect 67002 -2801 67093 -2683
rect 67211 -2801 67302 -2683
rect 67002 -2812 67302 -2801
rect 59802 -3111 59893 -2993
rect 60011 -3111 60102 -2993
rect 59802 -3153 60102 -3111
rect 59802 -3271 59893 -3153
rect 60011 -3271 60102 -3153
rect 59802 -3752 60102 -3271
rect 68802 -3463 69102 240
rect 72402 -173 72702 240
rect 72402 -291 72493 -173
rect 72611 -291 72702 -173
rect 72402 -333 72702 -291
rect 72402 -451 72493 -333
rect 72611 -451 72702 -333
rect 72402 -932 72702 -451
rect 74202 -1113 74502 240
rect 74202 -1231 74293 -1113
rect 74411 -1231 74502 -1113
rect 74202 -1273 74502 -1231
rect 74202 -1391 74293 -1273
rect 74411 -1391 74502 -1273
rect 74202 -1872 74502 -1391
rect 76002 -2053 76302 240
rect 76002 -2171 76093 -2053
rect 76211 -2171 76302 -2053
rect 76002 -2213 76302 -2171
rect 76002 -2331 76093 -2213
rect 76211 -2331 76302 -2213
rect 76002 -2812 76302 -2331
rect 68802 -3581 68893 -3463
rect 69011 -3581 69102 -3463
rect 68802 -3623 69102 -3581
rect 68802 -3741 68893 -3623
rect 69011 -3741 69102 -3623
rect 68802 -3752 69102 -3741
rect 77802 -2993 78102 240
rect 81402 -643 81702 240
rect 81402 -761 81493 -643
rect 81611 -761 81702 -643
rect 81402 -803 81702 -761
rect 81402 -921 81493 -803
rect 81611 -921 81702 -803
rect 81402 -932 81702 -921
rect 83202 -1583 83502 240
rect 83202 -1701 83293 -1583
rect 83411 -1701 83502 -1583
rect 83202 -1743 83502 -1701
rect 83202 -1861 83293 -1743
rect 83411 -1861 83502 -1743
rect 83202 -1872 83502 -1861
rect 85002 -2523 85302 240
rect 85002 -2641 85093 -2523
rect 85211 -2641 85302 -2523
rect 85002 -2683 85302 -2641
rect 85002 -2801 85093 -2683
rect 85211 -2801 85302 -2683
rect 85002 -2812 85302 -2801
rect 77802 -3111 77893 -2993
rect 78011 -3111 78102 -2993
rect 77802 -3153 78102 -3111
rect 77802 -3271 77893 -3153
rect 78011 -3271 78102 -3153
rect 77802 -3752 78102 -3271
rect 86802 -3463 87102 240
rect 90402 -173 90702 240
rect 90402 -291 90493 -173
rect 90611 -291 90702 -173
rect 90402 -333 90702 -291
rect 90402 -451 90493 -333
rect 90611 -451 90702 -333
rect 90402 -932 90702 -451
rect 92202 -1113 92502 240
rect 92202 -1231 92293 -1113
rect 92411 -1231 92502 -1113
rect 92202 -1273 92502 -1231
rect 92202 -1391 92293 -1273
rect 92411 -1391 92502 -1273
rect 92202 -1872 92502 -1391
rect 94002 -2053 94302 240
rect 94002 -2171 94093 -2053
rect 94211 -2171 94302 -2053
rect 94002 -2213 94302 -2171
rect 94002 -2331 94093 -2213
rect 94211 -2331 94302 -2213
rect 94002 -2812 94302 -2331
rect 86802 -3581 86893 -3463
rect 87011 -3581 87102 -3463
rect 86802 -3623 87102 -3581
rect 86802 -3741 86893 -3623
rect 87011 -3741 87102 -3623
rect 86802 -3752 87102 -3741
rect 95802 -2993 96102 240
rect 99402 -643 99702 240
rect 99402 -761 99493 -643
rect 99611 -761 99702 -643
rect 99402 -803 99702 -761
rect 99402 -921 99493 -803
rect 99611 -921 99702 -803
rect 99402 -932 99702 -921
rect 101202 -1583 101502 240
rect 101202 -1701 101293 -1583
rect 101411 -1701 101502 -1583
rect 101202 -1743 101502 -1701
rect 101202 -1861 101293 -1743
rect 101411 -1861 101502 -1743
rect 101202 -1872 101502 -1861
rect 103002 -2523 103302 240
rect 103002 -2641 103093 -2523
rect 103211 -2641 103302 -2523
rect 103002 -2683 103302 -2641
rect 103002 -2801 103093 -2683
rect 103211 -2801 103302 -2683
rect 103002 -2812 103302 -2801
rect 95802 -3111 95893 -2993
rect 96011 -3111 96102 -2993
rect 95802 -3153 96102 -3111
rect 95802 -3271 95893 -3153
rect 96011 -3271 96102 -3153
rect 95802 -3752 96102 -3271
rect 104802 -3463 105102 240
rect 108402 -173 108702 240
rect 108402 -291 108493 -173
rect 108611 -291 108702 -173
rect 108402 -333 108702 -291
rect 108402 -451 108493 -333
rect 108611 -451 108702 -333
rect 108402 -932 108702 -451
rect 110202 -1113 110502 240
rect 110202 -1231 110293 -1113
rect 110411 -1231 110502 -1113
rect 110202 -1273 110502 -1231
rect 110202 -1391 110293 -1273
rect 110411 -1391 110502 -1273
rect 110202 -1872 110502 -1391
rect 112002 -2053 112302 240
rect 112002 -2171 112093 -2053
rect 112211 -2171 112302 -2053
rect 112002 -2213 112302 -2171
rect 112002 -2331 112093 -2213
rect 112211 -2331 112302 -2213
rect 112002 -2812 112302 -2331
rect 104802 -3581 104893 -3463
rect 105011 -3581 105102 -3463
rect 104802 -3623 105102 -3581
rect 104802 -3741 104893 -3623
rect 105011 -3741 105102 -3623
rect 104802 -3752 105102 -3741
rect 113802 -2993 114102 240
rect 117402 -643 117702 240
rect 117402 -761 117493 -643
rect 117611 -761 117702 -643
rect 117402 -803 117702 -761
rect 117402 -921 117493 -803
rect 117611 -921 117702 -803
rect 117402 -932 117702 -921
rect 119202 -1583 119502 240
rect 119202 -1701 119293 -1583
rect 119411 -1701 119502 -1583
rect 119202 -1743 119502 -1701
rect 119202 -1861 119293 -1743
rect 119411 -1861 119502 -1743
rect 119202 -1872 119502 -1861
rect 121002 -2523 121302 240
rect 121002 -2641 121093 -2523
rect 121211 -2641 121302 -2523
rect 121002 -2683 121302 -2641
rect 121002 -2801 121093 -2683
rect 121211 -2801 121302 -2683
rect 121002 -2812 121302 -2801
rect 113802 -3111 113893 -2993
rect 114011 -3111 114102 -2993
rect 113802 -3153 114102 -3111
rect 113802 -3271 113893 -3153
rect 114011 -3271 114102 -3153
rect 113802 -3752 114102 -3271
rect 122802 -3463 123102 240
rect 126402 -173 126702 240
rect 126402 -291 126493 -173
rect 126611 -291 126702 -173
rect 126402 -333 126702 -291
rect 126402 -451 126493 -333
rect 126611 -451 126702 -333
rect 126402 -932 126702 -451
rect 128202 -1113 128502 240
rect 128202 -1231 128293 -1113
rect 128411 -1231 128502 -1113
rect 128202 -1273 128502 -1231
rect 128202 -1391 128293 -1273
rect 128411 -1391 128502 -1273
rect 128202 -1872 128502 -1391
rect 130002 -2053 130302 240
rect 130002 -2171 130093 -2053
rect 130211 -2171 130302 -2053
rect 130002 -2213 130302 -2171
rect 130002 -2331 130093 -2213
rect 130211 -2331 130302 -2213
rect 130002 -2812 130302 -2331
rect 122802 -3581 122893 -3463
rect 123011 -3581 123102 -3463
rect 122802 -3623 123102 -3581
rect 122802 -3741 122893 -3623
rect 123011 -3741 123102 -3623
rect 122802 -3752 123102 -3741
rect 131802 -2993 132102 240
rect 135402 -643 135702 240
rect 135402 -761 135493 -643
rect 135611 -761 135702 -643
rect 135402 -803 135702 -761
rect 135402 -921 135493 -803
rect 135611 -921 135702 -803
rect 135402 -932 135702 -921
rect 137202 -1583 137502 240
rect 137202 -1701 137293 -1583
rect 137411 -1701 137502 -1583
rect 137202 -1743 137502 -1701
rect 137202 -1861 137293 -1743
rect 137411 -1861 137502 -1743
rect 137202 -1872 137502 -1861
rect 139002 -2523 139302 240
rect 139002 -2641 139093 -2523
rect 139211 -2641 139302 -2523
rect 139002 -2683 139302 -2641
rect 139002 -2801 139093 -2683
rect 139211 -2801 139302 -2683
rect 139002 -2812 139302 -2801
rect 131802 -3111 131893 -2993
rect 132011 -3111 132102 -2993
rect 131802 -3153 132102 -3111
rect 131802 -3271 131893 -3153
rect 132011 -3271 132102 -3153
rect 131802 -3752 132102 -3271
rect 140802 -3463 141102 240
rect 144402 -173 144702 240
rect 144402 -291 144493 -173
rect 144611 -291 144702 -173
rect 144402 -333 144702 -291
rect 144402 -451 144493 -333
rect 144611 -451 144702 -333
rect 144402 -932 144702 -451
rect 146202 -1113 146502 240
rect 146202 -1231 146293 -1113
rect 146411 -1231 146502 -1113
rect 146202 -1273 146502 -1231
rect 146202 -1391 146293 -1273
rect 146411 -1391 146502 -1273
rect 146202 -1872 146502 -1391
rect 148002 -2053 148302 240
rect 148002 -2171 148093 -2053
rect 148211 -2171 148302 -2053
rect 148002 -2213 148302 -2171
rect 148002 -2331 148093 -2213
rect 148211 -2331 148302 -2213
rect 148002 -2812 148302 -2331
rect 140802 -3581 140893 -3463
rect 141011 -3581 141102 -3463
rect 140802 -3623 141102 -3581
rect 140802 -3741 140893 -3623
rect 141011 -3741 141102 -3623
rect 140802 -3752 141102 -3741
rect 149802 -2993 150102 240
rect 153402 -643 153702 240
rect 153402 -761 153493 -643
rect 153611 -761 153702 -643
rect 153402 -803 153702 -761
rect 153402 -921 153493 -803
rect 153611 -921 153702 -803
rect 153402 -932 153702 -921
rect 155202 -1583 155502 240
rect 155202 -1701 155293 -1583
rect 155411 -1701 155502 -1583
rect 155202 -1743 155502 -1701
rect 155202 -1861 155293 -1743
rect 155411 -1861 155502 -1743
rect 155202 -1872 155502 -1861
rect 157002 -2523 157302 240
rect 157002 -2641 157093 -2523
rect 157211 -2641 157302 -2523
rect 157002 -2683 157302 -2641
rect 157002 -2801 157093 -2683
rect 157211 -2801 157302 -2683
rect 157002 -2812 157302 -2801
rect 149802 -3111 149893 -2993
rect 150011 -3111 150102 -2993
rect 149802 -3153 150102 -3111
rect 149802 -3271 149893 -3153
rect 150011 -3271 150102 -3153
rect 149802 -3752 150102 -3271
rect 158802 -3463 159102 240
rect 162402 -173 162702 240
rect 162402 -291 162493 -173
rect 162611 -291 162702 -173
rect 162402 -333 162702 -291
rect 162402 -451 162493 -333
rect 162611 -451 162702 -333
rect 162402 -932 162702 -451
rect 164202 -1113 164502 240
rect 164202 -1231 164293 -1113
rect 164411 -1231 164502 -1113
rect 164202 -1273 164502 -1231
rect 164202 -1391 164293 -1273
rect 164411 -1391 164502 -1273
rect 164202 -1872 164502 -1391
rect 166002 -2053 166302 240
rect 166002 -2171 166093 -2053
rect 166211 -2171 166302 -2053
rect 166002 -2213 166302 -2171
rect 166002 -2331 166093 -2213
rect 166211 -2331 166302 -2213
rect 166002 -2812 166302 -2331
rect 158802 -3581 158893 -3463
rect 159011 -3581 159102 -3463
rect 158802 -3623 159102 -3581
rect 158802 -3741 158893 -3623
rect 159011 -3741 159102 -3623
rect 158802 -3752 159102 -3741
rect 167802 -2993 168102 240
rect 171402 -643 171702 240
rect 171402 -761 171493 -643
rect 171611 -761 171702 -643
rect 171402 -803 171702 -761
rect 171402 -921 171493 -803
rect 171611 -921 171702 -803
rect 171402 -932 171702 -921
rect 173202 -1583 173502 240
rect 173202 -1701 173293 -1583
rect 173411 -1701 173502 -1583
rect 173202 -1743 173502 -1701
rect 173202 -1861 173293 -1743
rect 173411 -1861 173502 -1743
rect 173202 -1872 173502 -1861
rect 175002 -2523 175302 240
rect 175002 -2641 175093 -2523
rect 175211 -2641 175302 -2523
rect 175002 -2683 175302 -2641
rect 175002 -2801 175093 -2683
rect 175211 -2801 175302 -2683
rect 175002 -2812 175302 -2801
rect 167802 -3111 167893 -2993
rect 168011 -3111 168102 -2993
rect 167802 -3153 168102 -3111
rect 167802 -3271 167893 -3153
rect 168011 -3271 168102 -3153
rect 167802 -3752 168102 -3271
rect 176802 -3463 177102 240
rect 180402 -173 180702 240
rect 180402 -291 180493 -173
rect 180611 -291 180702 -173
rect 180402 -333 180702 -291
rect 180402 -451 180493 -333
rect 180611 -451 180702 -333
rect 180402 -932 180702 -451
rect 182202 -1113 182502 240
rect 182202 -1231 182293 -1113
rect 182411 -1231 182502 -1113
rect 182202 -1273 182502 -1231
rect 182202 -1391 182293 -1273
rect 182411 -1391 182502 -1273
rect 182202 -1872 182502 -1391
rect 184002 -2053 184302 240
rect 184002 -2171 184093 -2053
rect 184211 -2171 184302 -2053
rect 184002 -2213 184302 -2171
rect 184002 -2331 184093 -2213
rect 184211 -2331 184302 -2213
rect 184002 -2812 184302 -2331
rect 176802 -3581 176893 -3463
rect 177011 -3581 177102 -3463
rect 176802 -3623 177102 -3581
rect 176802 -3741 176893 -3623
rect 177011 -3741 177102 -3623
rect 176802 -3752 177102 -3741
rect 185802 -2993 186102 240
rect 189402 -643 189702 240
rect 189402 -761 189493 -643
rect 189611 -761 189702 -643
rect 189402 -803 189702 -761
rect 189402 -921 189493 -803
rect 189611 -921 189702 -803
rect 189402 -932 189702 -921
rect 191202 -1583 191502 240
rect 191202 -1701 191293 -1583
rect 191411 -1701 191502 -1583
rect 191202 -1743 191502 -1701
rect 191202 -1861 191293 -1743
rect 191411 -1861 191502 -1743
rect 191202 -1872 191502 -1861
rect 193002 -2523 193302 240
rect 193002 -2641 193093 -2523
rect 193211 -2641 193302 -2523
rect 193002 -2683 193302 -2641
rect 193002 -2801 193093 -2683
rect 193211 -2801 193302 -2683
rect 193002 -2812 193302 -2801
rect 185802 -3111 185893 -2993
rect 186011 -3111 186102 -2993
rect 185802 -3153 186102 -3111
rect 185802 -3271 185893 -3153
rect 186011 -3271 186102 -3153
rect 185802 -3752 186102 -3271
rect 194802 -3463 195102 240
rect 198402 -173 198702 240
rect 198402 -291 198493 -173
rect 198611 -291 198702 -173
rect 198402 -333 198702 -291
rect 198402 -451 198493 -333
rect 198611 -451 198702 -333
rect 198402 -932 198702 -451
rect 200202 -1113 200502 240
rect 200202 -1231 200293 -1113
rect 200411 -1231 200502 -1113
rect 200202 -1273 200502 -1231
rect 200202 -1391 200293 -1273
rect 200411 -1391 200502 -1273
rect 200202 -1872 200502 -1391
rect 202002 -2053 202302 240
rect 202002 -2171 202093 -2053
rect 202211 -2171 202302 -2053
rect 202002 -2213 202302 -2171
rect 202002 -2331 202093 -2213
rect 202211 -2331 202302 -2213
rect 202002 -2812 202302 -2331
rect 194802 -3581 194893 -3463
rect 195011 -3581 195102 -3463
rect 194802 -3623 195102 -3581
rect 194802 -3741 194893 -3623
rect 195011 -3741 195102 -3623
rect 194802 -3752 195102 -3741
rect 203802 -2993 204102 240
rect 207402 -643 207702 240
rect 207402 -761 207493 -643
rect 207611 -761 207702 -643
rect 207402 -803 207702 -761
rect 207402 -921 207493 -803
rect 207611 -921 207702 -803
rect 207402 -932 207702 -921
rect 209202 -1583 209502 240
rect 209202 -1701 209293 -1583
rect 209411 -1701 209502 -1583
rect 209202 -1743 209502 -1701
rect 209202 -1861 209293 -1743
rect 209411 -1861 209502 -1743
rect 209202 -1872 209502 -1861
rect 211002 -2523 211302 240
rect 211002 -2641 211093 -2523
rect 211211 -2641 211302 -2523
rect 211002 -2683 211302 -2641
rect 211002 -2801 211093 -2683
rect 211211 -2801 211302 -2683
rect 211002 -2812 211302 -2801
rect 203802 -3111 203893 -2993
rect 204011 -3111 204102 -2993
rect 203802 -3153 204102 -3111
rect 203802 -3271 203893 -3153
rect 204011 -3271 204102 -3153
rect 203802 -3752 204102 -3271
rect 212802 -3463 213102 240
rect 216402 -173 216702 240
rect 216402 -291 216493 -173
rect 216611 -291 216702 -173
rect 216402 -333 216702 -291
rect 216402 -451 216493 -333
rect 216611 -451 216702 -333
rect 216402 -932 216702 -451
rect 218202 -1113 218502 240
rect 218202 -1231 218293 -1113
rect 218411 -1231 218502 -1113
rect 218202 -1273 218502 -1231
rect 218202 -1391 218293 -1273
rect 218411 -1391 218502 -1273
rect 218202 -1872 218502 -1391
rect 220002 -2053 220302 240
rect 220002 -2171 220093 -2053
rect 220211 -2171 220302 -2053
rect 220002 -2213 220302 -2171
rect 220002 -2331 220093 -2213
rect 220211 -2331 220302 -2213
rect 220002 -2812 220302 -2331
rect 212802 -3581 212893 -3463
rect 213011 -3581 213102 -3463
rect 212802 -3623 213102 -3581
rect 212802 -3741 212893 -3623
rect 213011 -3741 213102 -3623
rect 212802 -3752 213102 -3741
rect 221802 -2993 222102 240
rect 225402 -643 225702 240
rect 225402 -761 225493 -643
rect 225611 -761 225702 -643
rect 225402 -803 225702 -761
rect 225402 -921 225493 -803
rect 225611 -921 225702 -803
rect 225402 -932 225702 -921
rect 227202 -1583 227502 240
rect 227202 -1701 227293 -1583
rect 227411 -1701 227502 -1583
rect 227202 -1743 227502 -1701
rect 227202 -1861 227293 -1743
rect 227411 -1861 227502 -1743
rect 227202 -1872 227502 -1861
rect 229002 -2523 229302 240
rect 229002 -2641 229093 -2523
rect 229211 -2641 229302 -2523
rect 229002 -2683 229302 -2641
rect 229002 -2801 229093 -2683
rect 229211 -2801 229302 -2683
rect 229002 -2812 229302 -2801
rect 221802 -3111 221893 -2993
rect 222011 -3111 222102 -2993
rect 221802 -3153 222102 -3111
rect 221802 -3271 221893 -3153
rect 222011 -3271 222102 -3153
rect 221802 -3752 222102 -3271
rect 230802 -3463 231102 240
rect 234402 -173 234702 240
rect 234402 -291 234493 -173
rect 234611 -291 234702 -173
rect 234402 -333 234702 -291
rect 234402 -451 234493 -333
rect 234611 -451 234702 -333
rect 234402 -932 234702 -451
rect 236202 -1113 236502 240
rect 236202 -1231 236293 -1113
rect 236411 -1231 236502 -1113
rect 236202 -1273 236502 -1231
rect 236202 -1391 236293 -1273
rect 236411 -1391 236502 -1273
rect 236202 -1872 236502 -1391
rect 238002 -2053 238302 240
rect 238002 -2171 238093 -2053
rect 238211 -2171 238302 -2053
rect 238002 -2213 238302 -2171
rect 238002 -2331 238093 -2213
rect 238211 -2331 238302 -2213
rect 238002 -2812 238302 -2331
rect 230802 -3581 230893 -3463
rect 231011 -3581 231102 -3463
rect 230802 -3623 231102 -3581
rect 230802 -3741 230893 -3623
rect 231011 -3741 231102 -3623
rect 230802 -3752 231102 -3741
rect 239802 -2993 240102 240
rect 243402 -643 243702 240
rect 243402 -761 243493 -643
rect 243611 -761 243702 -643
rect 243402 -803 243702 -761
rect 243402 -921 243493 -803
rect 243611 -921 243702 -803
rect 243402 -932 243702 -921
rect 245202 -1583 245502 240
rect 245202 -1701 245293 -1583
rect 245411 -1701 245502 -1583
rect 245202 -1743 245502 -1701
rect 245202 -1861 245293 -1743
rect 245411 -1861 245502 -1743
rect 245202 -1872 245502 -1861
rect 247002 -2523 247302 240
rect 247002 -2641 247093 -2523
rect 247211 -2641 247302 -2523
rect 247002 -2683 247302 -2641
rect 247002 -2801 247093 -2683
rect 247211 -2801 247302 -2683
rect 247002 -2812 247302 -2801
rect 239802 -3111 239893 -2993
rect 240011 -3111 240102 -2993
rect 239802 -3153 240102 -3111
rect 239802 -3271 239893 -3153
rect 240011 -3271 240102 -3153
rect 239802 -3752 240102 -3271
rect 248802 -3463 249102 240
rect 252402 -173 252702 240
rect 252402 -291 252493 -173
rect 252611 -291 252702 -173
rect 252402 -333 252702 -291
rect 252402 -451 252493 -333
rect 252611 -451 252702 -333
rect 252402 -932 252702 -451
rect 254202 -1113 254502 240
rect 254202 -1231 254293 -1113
rect 254411 -1231 254502 -1113
rect 254202 -1273 254502 -1231
rect 254202 -1391 254293 -1273
rect 254411 -1391 254502 -1273
rect 254202 -1872 254502 -1391
rect 256002 -2053 256302 240
rect 256002 -2171 256093 -2053
rect 256211 -2171 256302 -2053
rect 256002 -2213 256302 -2171
rect 256002 -2331 256093 -2213
rect 256211 -2331 256302 -2213
rect 256002 -2812 256302 -2331
rect 248802 -3581 248893 -3463
rect 249011 -3581 249102 -3463
rect 248802 -3623 249102 -3581
rect 248802 -3741 248893 -3623
rect 249011 -3741 249102 -3623
rect 248802 -3752 249102 -3741
rect 257802 -2993 258102 240
rect 261402 -643 261702 240
rect 261402 -761 261493 -643
rect 261611 -761 261702 -643
rect 261402 -803 261702 -761
rect 261402 -921 261493 -803
rect 261611 -921 261702 -803
rect 261402 -932 261702 -921
rect 263202 -1583 263502 240
rect 263202 -1701 263293 -1583
rect 263411 -1701 263502 -1583
rect 263202 -1743 263502 -1701
rect 263202 -1861 263293 -1743
rect 263411 -1861 263502 -1743
rect 263202 -1872 263502 -1861
rect 265002 -2523 265302 240
rect 265002 -2641 265093 -2523
rect 265211 -2641 265302 -2523
rect 265002 -2683 265302 -2641
rect 265002 -2801 265093 -2683
rect 265211 -2801 265302 -2683
rect 265002 -2812 265302 -2801
rect 257802 -3111 257893 -2993
rect 258011 -3111 258102 -2993
rect 257802 -3153 258102 -3111
rect 257802 -3271 257893 -3153
rect 258011 -3271 258102 -3153
rect 257802 -3752 258102 -3271
rect 266802 -3463 267102 240
rect 270402 -173 270702 240
rect 270402 -291 270493 -173
rect 270611 -291 270702 -173
rect 270402 -333 270702 -291
rect 270402 -451 270493 -333
rect 270611 -451 270702 -333
rect 270402 -932 270702 -451
rect 272202 -1113 272502 240
rect 272202 -1231 272293 -1113
rect 272411 -1231 272502 -1113
rect 272202 -1273 272502 -1231
rect 272202 -1391 272293 -1273
rect 272411 -1391 272502 -1273
rect 272202 -1872 272502 -1391
rect 274002 -2053 274302 240
rect 274002 -2171 274093 -2053
rect 274211 -2171 274302 -2053
rect 274002 -2213 274302 -2171
rect 274002 -2331 274093 -2213
rect 274211 -2331 274302 -2213
rect 274002 -2812 274302 -2331
rect 266802 -3581 266893 -3463
rect 267011 -3581 267102 -3463
rect 266802 -3623 267102 -3581
rect 266802 -3741 266893 -3623
rect 267011 -3741 267102 -3623
rect 266802 -3752 267102 -3741
rect 275802 -2993 276102 240
rect 279402 -643 279702 240
rect 279402 -761 279493 -643
rect 279611 -761 279702 -643
rect 279402 -803 279702 -761
rect 279402 -921 279493 -803
rect 279611 -921 279702 -803
rect 279402 -932 279702 -921
rect 281202 -1583 281502 240
rect 281202 -1701 281293 -1583
rect 281411 -1701 281502 -1583
rect 281202 -1743 281502 -1701
rect 281202 -1861 281293 -1743
rect 281411 -1861 281502 -1743
rect 281202 -1872 281502 -1861
rect 283002 -2523 283302 240
rect 283002 -2641 283093 -2523
rect 283211 -2641 283302 -2523
rect 283002 -2683 283302 -2641
rect 283002 -2801 283093 -2683
rect 283211 -2801 283302 -2683
rect 283002 -2812 283302 -2801
rect 275802 -3111 275893 -2993
rect 276011 -3111 276102 -2993
rect 275802 -3153 276102 -3111
rect 275802 -3271 275893 -3153
rect 276011 -3271 276102 -3153
rect 275802 -3752 276102 -3271
rect 284802 -3463 285102 240
rect 288402 -173 288702 240
rect 288402 -291 288493 -173
rect 288611 -291 288702 -173
rect 288402 -333 288702 -291
rect 288402 -451 288493 -333
rect 288611 -451 288702 -333
rect 288402 -932 288702 -451
rect 290202 -1113 290502 240
rect 292660 -173 292960 949
rect 292660 -291 292751 -173
rect 292869 -291 292960 -173
rect 292660 -333 292960 -291
rect 292660 -451 292751 -333
rect 292869 -451 292960 -333
rect 292660 -462 292960 -451
rect 293130 334227 293430 352611
rect 293130 334109 293221 334227
rect 293339 334109 293430 334227
rect 293130 334067 293430 334109
rect 293130 333949 293221 334067
rect 293339 333949 293430 334067
rect 293130 316227 293430 333949
rect 293130 316109 293221 316227
rect 293339 316109 293430 316227
rect 293130 316067 293430 316109
rect 293130 315949 293221 316067
rect 293339 315949 293430 316067
rect 293130 298227 293430 315949
rect 293130 298109 293221 298227
rect 293339 298109 293430 298227
rect 293130 298067 293430 298109
rect 293130 297949 293221 298067
rect 293339 297949 293430 298067
rect 293130 280227 293430 297949
rect 293130 280109 293221 280227
rect 293339 280109 293430 280227
rect 293130 280067 293430 280109
rect 293130 279949 293221 280067
rect 293339 279949 293430 280067
rect 293130 262227 293430 279949
rect 293130 262109 293221 262227
rect 293339 262109 293430 262227
rect 293130 262067 293430 262109
rect 293130 261949 293221 262067
rect 293339 261949 293430 262067
rect 293130 244227 293430 261949
rect 293130 244109 293221 244227
rect 293339 244109 293430 244227
rect 293130 244067 293430 244109
rect 293130 243949 293221 244067
rect 293339 243949 293430 244067
rect 293130 226227 293430 243949
rect 293130 226109 293221 226227
rect 293339 226109 293430 226227
rect 293130 226067 293430 226109
rect 293130 225949 293221 226067
rect 293339 225949 293430 226067
rect 293130 208227 293430 225949
rect 293130 208109 293221 208227
rect 293339 208109 293430 208227
rect 293130 208067 293430 208109
rect 293130 207949 293221 208067
rect 293339 207949 293430 208067
rect 293130 190227 293430 207949
rect 293130 190109 293221 190227
rect 293339 190109 293430 190227
rect 293130 190067 293430 190109
rect 293130 189949 293221 190067
rect 293339 189949 293430 190067
rect 293130 172227 293430 189949
rect 293130 172109 293221 172227
rect 293339 172109 293430 172227
rect 293130 172067 293430 172109
rect 293130 171949 293221 172067
rect 293339 171949 293430 172067
rect 293130 154227 293430 171949
rect 293130 154109 293221 154227
rect 293339 154109 293430 154227
rect 293130 154067 293430 154109
rect 293130 153949 293221 154067
rect 293339 153949 293430 154067
rect 293130 136227 293430 153949
rect 293130 136109 293221 136227
rect 293339 136109 293430 136227
rect 293130 136067 293430 136109
rect 293130 135949 293221 136067
rect 293339 135949 293430 136067
rect 293130 118227 293430 135949
rect 293130 118109 293221 118227
rect 293339 118109 293430 118227
rect 293130 118067 293430 118109
rect 293130 117949 293221 118067
rect 293339 117949 293430 118067
rect 293130 100227 293430 117949
rect 293130 100109 293221 100227
rect 293339 100109 293430 100227
rect 293130 100067 293430 100109
rect 293130 99949 293221 100067
rect 293339 99949 293430 100067
rect 293130 82227 293430 99949
rect 293130 82109 293221 82227
rect 293339 82109 293430 82227
rect 293130 82067 293430 82109
rect 293130 81949 293221 82067
rect 293339 81949 293430 82067
rect 293130 64227 293430 81949
rect 293130 64109 293221 64227
rect 293339 64109 293430 64227
rect 293130 64067 293430 64109
rect 293130 63949 293221 64067
rect 293339 63949 293430 64067
rect 293130 46227 293430 63949
rect 293130 46109 293221 46227
rect 293339 46109 293430 46227
rect 293130 46067 293430 46109
rect 293130 45949 293221 46067
rect 293339 45949 293430 46067
rect 293130 28227 293430 45949
rect 293130 28109 293221 28227
rect 293339 28109 293430 28227
rect 293130 28067 293430 28109
rect 293130 27949 293221 28067
rect 293339 27949 293430 28067
rect 293130 10227 293430 27949
rect 293130 10109 293221 10227
rect 293339 10109 293430 10227
rect 293130 10067 293430 10109
rect 293130 9949 293221 10067
rect 293339 9949 293430 10067
rect 293130 -643 293430 9949
rect 293130 -761 293221 -643
rect 293339 -761 293430 -643
rect 293130 -803 293430 -761
rect 293130 -921 293221 -803
rect 293339 -921 293430 -803
rect 293130 -932 293430 -921
rect 293600 345027 293900 353081
rect 293600 344909 293691 345027
rect 293809 344909 293900 345027
rect 293600 344867 293900 344909
rect 293600 344749 293691 344867
rect 293809 344749 293900 344867
rect 293600 327027 293900 344749
rect 293600 326909 293691 327027
rect 293809 326909 293900 327027
rect 293600 326867 293900 326909
rect 293600 326749 293691 326867
rect 293809 326749 293900 326867
rect 293600 309027 293900 326749
rect 293600 308909 293691 309027
rect 293809 308909 293900 309027
rect 293600 308867 293900 308909
rect 293600 308749 293691 308867
rect 293809 308749 293900 308867
rect 293600 291027 293900 308749
rect 293600 290909 293691 291027
rect 293809 290909 293900 291027
rect 293600 290867 293900 290909
rect 293600 290749 293691 290867
rect 293809 290749 293900 290867
rect 293600 273027 293900 290749
rect 293600 272909 293691 273027
rect 293809 272909 293900 273027
rect 293600 272867 293900 272909
rect 293600 272749 293691 272867
rect 293809 272749 293900 272867
rect 293600 255027 293900 272749
rect 293600 254909 293691 255027
rect 293809 254909 293900 255027
rect 293600 254867 293900 254909
rect 293600 254749 293691 254867
rect 293809 254749 293900 254867
rect 293600 237027 293900 254749
rect 293600 236909 293691 237027
rect 293809 236909 293900 237027
rect 293600 236867 293900 236909
rect 293600 236749 293691 236867
rect 293809 236749 293900 236867
rect 293600 219027 293900 236749
rect 293600 218909 293691 219027
rect 293809 218909 293900 219027
rect 293600 218867 293900 218909
rect 293600 218749 293691 218867
rect 293809 218749 293900 218867
rect 293600 201027 293900 218749
rect 293600 200909 293691 201027
rect 293809 200909 293900 201027
rect 293600 200867 293900 200909
rect 293600 200749 293691 200867
rect 293809 200749 293900 200867
rect 293600 183027 293900 200749
rect 293600 182909 293691 183027
rect 293809 182909 293900 183027
rect 293600 182867 293900 182909
rect 293600 182749 293691 182867
rect 293809 182749 293900 182867
rect 293600 165027 293900 182749
rect 293600 164909 293691 165027
rect 293809 164909 293900 165027
rect 293600 164867 293900 164909
rect 293600 164749 293691 164867
rect 293809 164749 293900 164867
rect 293600 147027 293900 164749
rect 293600 146909 293691 147027
rect 293809 146909 293900 147027
rect 293600 146867 293900 146909
rect 293600 146749 293691 146867
rect 293809 146749 293900 146867
rect 293600 129027 293900 146749
rect 293600 128909 293691 129027
rect 293809 128909 293900 129027
rect 293600 128867 293900 128909
rect 293600 128749 293691 128867
rect 293809 128749 293900 128867
rect 293600 111027 293900 128749
rect 293600 110909 293691 111027
rect 293809 110909 293900 111027
rect 293600 110867 293900 110909
rect 293600 110749 293691 110867
rect 293809 110749 293900 110867
rect 293600 93027 293900 110749
rect 293600 92909 293691 93027
rect 293809 92909 293900 93027
rect 293600 92867 293900 92909
rect 293600 92749 293691 92867
rect 293809 92749 293900 92867
rect 293600 75027 293900 92749
rect 293600 74909 293691 75027
rect 293809 74909 293900 75027
rect 293600 74867 293900 74909
rect 293600 74749 293691 74867
rect 293809 74749 293900 74867
rect 293600 57027 293900 74749
rect 293600 56909 293691 57027
rect 293809 56909 293900 57027
rect 293600 56867 293900 56909
rect 293600 56749 293691 56867
rect 293809 56749 293900 56867
rect 293600 39027 293900 56749
rect 293600 38909 293691 39027
rect 293809 38909 293900 39027
rect 293600 38867 293900 38909
rect 293600 38749 293691 38867
rect 293809 38749 293900 38867
rect 293600 21027 293900 38749
rect 293600 20909 293691 21027
rect 293809 20909 293900 21027
rect 293600 20867 293900 20909
rect 293600 20749 293691 20867
rect 293809 20749 293900 20867
rect 293600 3027 293900 20749
rect 293600 2909 293691 3027
rect 293809 2909 293900 3027
rect 293600 2867 293900 2909
rect 293600 2749 293691 2867
rect 293809 2749 293900 2867
rect 290202 -1231 290293 -1113
rect 290411 -1231 290502 -1113
rect 290202 -1273 290502 -1231
rect 290202 -1391 290293 -1273
rect 290411 -1391 290502 -1273
rect 290202 -1872 290502 -1391
rect 293600 -1113 293900 2749
rect 293600 -1231 293691 -1113
rect 293809 -1231 293900 -1113
rect 293600 -1273 293900 -1231
rect 293600 -1391 293691 -1273
rect 293809 -1391 293900 -1273
rect 293600 -1402 293900 -1391
rect 294070 336027 294370 353551
rect 294070 335909 294161 336027
rect 294279 335909 294370 336027
rect 294070 335867 294370 335909
rect 294070 335749 294161 335867
rect 294279 335749 294370 335867
rect 294070 318027 294370 335749
rect 294070 317909 294161 318027
rect 294279 317909 294370 318027
rect 294070 317867 294370 317909
rect 294070 317749 294161 317867
rect 294279 317749 294370 317867
rect 294070 300027 294370 317749
rect 294070 299909 294161 300027
rect 294279 299909 294370 300027
rect 294070 299867 294370 299909
rect 294070 299749 294161 299867
rect 294279 299749 294370 299867
rect 294070 282027 294370 299749
rect 294070 281909 294161 282027
rect 294279 281909 294370 282027
rect 294070 281867 294370 281909
rect 294070 281749 294161 281867
rect 294279 281749 294370 281867
rect 294070 264027 294370 281749
rect 294070 263909 294161 264027
rect 294279 263909 294370 264027
rect 294070 263867 294370 263909
rect 294070 263749 294161 263867
rect 294279 263749 294370 263867
rect 294070 246027 294370 263749
rect 294070 245909 294161 246027
rect 294279 245909 294370 246027
rect 294070 245867 294370 245909
rect 294070 245749 294161 245867
rect 294279 245749 294370 245867
rect 294070 228027 294370 245749
rect 294070 227909 294161 228027
rect 294279 227909 294370 228027
rect 294070 227867 294370 227909
rect 294070 227749 294161 227867
rect 294279 227749 294370 227867
rect 294070 210027 294370 227749
rect 294070 209909 294161 210027
rect 294279 209909 294370 210027
rect 294070 209867 294370 209909
rect 294070 209749 294161 209867
rect 294279 209749 294370 209867
rect 294070 192027 294370 209749
rect 294070 191909 294161 192027
rect 294279 191909 294370 192027
rect 294070 191867 294370 191909
rect 294070 191749 294161 191867
rect 294279 191749 294370 191867
rect 294070 174027 294370 191749
rect 294070 173909 294161 174027
rect 294279 173909 294370 174027
rect 294070 173867 294370 173909
rect 294070 173749 294161 173867
rect 294279 173749 294370 173867
rect 294070 156027 294370 173749
rect 294070 155909 294161 156027
rect 294279 155909 294370 156027
rect 294070 155867 294370 155909
rect 294070 155749 294161 155867
rect 294279 155749 294370 155867
rect 294070 138027 294370 155749
rect 294070 137909 294161 138027
rect 294279 137909 294370 138027
rect 294070 137867 294370 137909
rect 294070 137749 294161 137867
rect 294279 137749 294370 137867
rect 294070 120027 294370 137749
rect 294070 119909 294161 120027
rect 294279 119909 294370 120027
rect 294070 119867 294370 119909
rect 294070 119749 294161 119867
rect 294279 119749 294370 119867
rect 294070 102027 294370 119749
rect 294070 101909 294161 102027
rect 294279 101909 294370 102027
rect 294070 101867 294370 101909
rect 294070 101749 294161 101867
rect 294279 101749 294370 101867
rect 294070 84027 294370 101749
rect 294070 83909 294161 84027
rect 294279 83909 294370 84027
rect 294070 83867 294370 83909
rect 294070 83749 294161 83867
rect 294279 83749 294370 83867
rect 294070 66027 294370 83749
rect 294070 65909 294161 66027
rect 294279 65909 294370 66027
rect 294070 65867 294370 65909
rect 294070 65749 294161 65867
rect 294279 65749 294370 65867
rect 294070 48027 294370 65749
rect 294070 47909 294161 48027
rect 294279 47909 294370 48027
rect 294070 47867 294370 47909
rect 294070 47749 294161 47867
rect 294279 47749 294370 47867
rect 294070 30027 294370 47749
rect 294070 29909 294161 30027
rect 294279 29909 294370 30027
rect 294070 29867 294370 29909
rect 294070 29749 294161 29867
rect 294279 29749 294370 29867
rect 294070 12027 294370 29749
rect 294070 11909 294161 12027
rect 294279 11909 294370 12027
rect 294070 11867 294370 11909
rect 294070 11749 294161 11867
rect 294279 11749 294370 11867
rect 294070 -1583 294370 11749
rect 294070 -1701 294161 -1583
rect 294279 -1701 294370 -1583
rect 294070 -1743 294370 -1701
rect 294070 -1861 294161 -1743
rect 294279 -1861 294370 -1743
rect 294070 -1872 294370 -1861
rect 294540 346827 294840 354021
rect 294540 346709 294631 346827
rect 294749 346709 294840 346827
rect 294540 346667 294840 346709
rect 294540 346549 294631 346667
rect 294749 346549 294840 346667
rect 294540 328827 294840 346549
rect 294540 328709 294631 328827
rect 294749 328709 294840 328827
rect 294540 328667 294840 328709
rect 294540 328549 294631 328667
rect 294749 328549 294840 328667
rect 294540 310827 294840 328549
rect 294540 310709 294631 310827
rect 294749 310709 294840 310827
rect 294540 310667 294840 310709
rect 294540 310549 294631 310667
rect 294749 310549 294840 310667
rect 294540 292827 294840 310549
rect 294540 292709 294631 292827
rect 294749 292709 294840 292827
rect 294540 292667 294840 292709
rect 294540 292549 294631 292667
rect 294749 292549 294840 292667
rect 294540 274827 294840 292549
rect 294540 274709 294631 274827
rect 294749 274709 294840 274827
rect 294540 274667 294840 274709
rect 294540 274549 294631 274667
rect 294749 274549 294840 274667
rect 294540 256827 294840 274549
rect 294540 256709 294631 256827
rect 294749 256709 294840 256827
rect 294540 256667 294840 256709
rect 294540 256549 294631 256667
rect 294749 256549 294840 256667
rect 294540 238827 294840 256549
rect 294540 238709 294631 238827
rect 294749 238709 294840 238827
rect 294540 238667 294840 238709
rect 294540 238549 294631 238667
rect 294749 238549 294840 238667
rect 294540 220827 294840 238549
rect 294540 220709 294631 220827
rect 294749 220709 294840 220827
rect 294540 220667 294840 220709
rect 294540 220549 294631 220667
rect 294749 220549 294840 220667
rect 294540 202827 294840 220549
rect 294540 202709 294631 202827
rect 294749 202709 294840 202827
rect 294540 202667 294840 202709
rect 294540 202549 294631 202667
rect 294749 202549 294840 202667
rect 294540 184827 294840 202549
rect 294540 184709 294631 184827
rect 294749 184709 294840 184827
rect 294540 184667 294840 184709
rect 294540 184549 294631 184667
rect 294749 184549 294840 184667
rect 294540 166827 294840 184549
rect 294540 166709 294631 166827
rect 294749 166709 294840 166827
rect 294540 166667 294840 166709
rect 294540 166549 294631 166667
rect 294749 166549 294840 166667
rect 294540 148827 294840 166549
rect 294540 148709 294631 148827
rect 294749 148709 294840 148827
rect 294540 148667 294840 148709
rect 294540 148549 294631 148667
rect 294749 148549 294840 148667
rect 294540 130827 294840 148549
rect 294540 130709 294631 130827
rect 294749 130709 294840 130827
rect 294540 130667 294840 130709
rect 294540 130549 294631 130667
rect 294749 130549 294840 130667
rect 294540 112827 294840 130549
rect 294540 112709 294631 112827
rect 294749 112709 294840 112827
rect 294540 112667 294840 112709
rect 294540 112549 294631 112667
rect 294749 112549 294840 112667
rect 294540 94827 294840 112549
rect 294540 94709 294631 94827
rect 294749 94709 294840 94827
rect 294540 94667 294840 94709
rect 294540 94549 294631 94667
rect 294749 94549 294840 94667
rect 294540 76827 294840 94549
rect 294540 76709 294631 76827
rect 294749 76709 294840 76827
rect 294540 76667 294840 76709
rect 294540 76549 294631 76667
rect 294749 76549 294840 76667
rect 294540 58827 294840 76549
rect 294540 58709 294631 58827
rect 294749 58709 294840 58827
rect 294540 58667 294840 58709
rect 294540 58549 294631 58667
rect 294749 58549 294840 58667
rect 294540 40827 294840 58549
rect 294540 40709 294631 40827
rect 294749 40709 294840 40827
rect 294540 40667 294840 40709
rect 294540 40549 294631 40667
rect 294749 40549 294840 40667
rect 294540 22827 294840 40549
rect 294540 22709 294631 22827
rect 294749 22709 294840 22827
rect 294540 22667 294840 22709
rect 294540 22549 294631 22667
rect 294749 22549 294840 22667
rect 294540 4827 294840 22549
rect 294540 4709 294631 4827
rect 294749 4709 294840 4827
rect 294540 4667 294840 4709
rect 294540 4549 294631 4667
rect 294749 4549 294840 4667
rect 294540 -2053 294840 4549
rect 294540 -2171 294631 -2053
rect 294749 -2171 294840 -2053
rect 294540 -2213 294840 -2171
rect 294540 -2331 294631 -2213
rect 294749 -2331 294840 -2213
rect 294540 -2342 294840 -2331
rect 295010 337827 295310 354491
rect 295010 337709 295101 337827
rect 295219 337709 295310 337827
rect 295010 337667 295310 337709
rect 295010 337549 295101 337667
rect 295219 337549 295310 337667
rect 295010 319827 295310 337549
rect 295010 319709 295101 319827
rect 295219 319709 295310 319827
rect 295010 319667 295310 319709
rect 295010 319549 295101 319667
rect 295219 319549 295310 319667
rect 295010 301827 295310 319549
rect 295010 301709 295101 301827
rect 295219 301709 295310 301827
rect 295010 301667 295310 301709
rect 295010 301549 295101 301667
rect 295219 301549 295310 301667
rect 295010 283827 295310 301549
rect 295010 283709 295101 283827
rect 295219 283709 295310 283827
rect 295010 283667 295310 283709
rect 295010 283549 295101 283667
rect 295219 283549 295310 283667
rect 295010 265827 295310 283549
rect 295010 265709 295101 265827
rect 295219 265709 295310 265827
rect 295010 265667 295310 265709
rect 295010 265549 295101 265667
rect 295219 265549 295310 265667
rect 295010 247827 295310 265549
rect 295010 247709 295101 247827
rect 295219 247709 295310 247827
rect 295010 247667 295310 247709
rect 295010 247549 295101 247667
rect 295219 247549 295310 247667
rect 295010 229827 295310 247549
rect 295010 229709 295101 229827
rect 295219 229709 295310 229827
rect 295010 229667 295310 229709
rect 295010 229549 295101 229667
rect 295219 229549 295310 229667
rect 295010 211827 295310 229549
rect 295010 211709 295101 211827
rect 295219 211709 295310 211827
rect 295010 211667 295310 211709
rect 295010 211549 295101 211667
rect 295219 211549 295310 211667
rect 295010 193827 295310 211549
rect 295010 193709 295101 193827
rect 295219 193709 295310 193827
rect 295010 193667 295310 193709
rect 295010 193549 295101 193667
rect 295219 193549 295310 193667
rect 295010 175827 295310 193549
rect 295010 175709 295101 175827
rect 295219 175709 295310 175827
rect 295010 175667 295310 175709
rect 295010 175549 295101 175667
rect 295219 175549 295310 175667
rect 295010 157827 295310 175549
rect 295010 157709 295101 157827
rect 295219 157709 295310 157827
rect 295010 157667 295310 157709
rect 295010 157549 295101 157667
rect 295219 157549 295310 157667
rect 295010 139827 295310 157549
rect 295010 139709 295101 139827
rect 295219 139709 295310 139827
rect 295010 139667 295310 139709
rect 295010 139549 295101 139667
rect 295219 139549 295310 139667
rect 295010 121827 295310 139549
rect 295010 121709 295101 121827
rect 295219 121709 295310 121827
rect 295010 121667 295310 121709
rect 295010 121549 295101 121667
rect 295219 121549 295310 121667
rect 295010 103827 295310 121549
rect 295010 103709 295101 103827
rect 295219 103709 295310 103827
rect 295010 103667 295310 103709
rect 295010 103549 295101 103667
rect 295219 103549 295310 103667
rect 295010 85827 295310 103549
rect 295010 85709 295101 85827
rect 295219 85709 295310 85827
rect 295010 85667 295310 85709
rect 295010 85549 295101 85667
rect 295219 85549 295310 85667
rect 295010 67827 295310 85549
rect 295010 67709 295101 67827
rect 295219 67709 295310 67827
rect 295010 67667 295310 67709
rect 295010 67549 295101 67667
rect 295219 67549 295310 67667
rect 295010 49827 295310 67549
rect 295010 49709 295101 49827
rect 295219 49709 295310 49827
rect 295010 49667 295310 49709
rect 295010 49549 295101 49667
rect 295219 49549 295310 49667
rect 295010 31827 295310 49549
rect 295010 31709 295101 31827
rect 295219 31709 295310 31827
rect 295010 31667 295310 31709
rect 295010 31549 295101 31667
rect 295219 31549 295310 31667
rect 295010 13827 295310 31549
rect 295010 13709 295101 13827
rect 295219 13709 295310 13827
rect 295010 13667 295310 13709
rect 295010 13549 295101 13667
rect 295219 13549 295310 13667
rect 295010 -2523 295310 13549
rect 295010 -2641 295101 -2523
rect 295219 -2641 295310 -2523
rect 295010 -2683 295310 -2641
rect 295010 -2801 295101 -2683
rect 295219 -2801 295310 -2683
rect 295010 -2812 295310 -2801
rect 295480 348627 295780 354961
rect 295480 348509 295571 348627
rect 295689 348509 295780 348627
rect 295480 348467 295780 348509
rect 295480 348349 295571 348467
rect 295689 348349 295780 348467
rect 295480 330627 295780 348349
rect 295480 330509 295571 330627
rect 295689 330509 295780 330627
rect 295480 330467 295780 330509
rect 295480 330349 295571 330467
rect 295689 330349 295780 330467
rect 295480 312627 295780 330349
rect 295480 312509 295571 312627
rect 295689 312509 295780 312627
rect 295480 312467 295780 312509
rect 295480 312349 295571 312467
rect 295689 312349 295780 312467
rect 295480 294627 295780 312349
rect 295480 294509 295571 294627
rect 295689 294509 295780 294627
rect 295480 294467 295780 294509
rect 295480 294349 295571 294467
rect 295689 294349 295780 294467
rect 295480 276627 295780 294349
rect 295480 276509 295571 276627
rect 295689 276509 295780 276627
rect 295480 276467 295780 276509
rect 295480 276349 295571 276467
rect 295689 276349 295780 276467
rect 295480 258627 295780 276349
rect 295480 258509 295571 258627
rect 295689 258509 295780 258627
rect 295480 258467 295780 258509
rect 295480 258349 295571 258467
rect 295689 258349 295780 258467
rect 295480 240627 295780 258349
rect 295480 240509 295571 240627
rect 295689 240509 295780 240627
rect 295480 240467 295780 240509
rect 295480 240349 295571 240467
rect 295689 240349 295780 240467
rect 295480 222627 295780 240349
rect 295480 222509 295571 222627
rect 295689 222509 295780 222627
rect 295480 222467 295780 222509
rect 295480 222349 295571 222467
rect 295689 222349 295780 222467
rect 295480 204627 295780 222349
rect 295480 204509 295571 204627
rect 295689 204509 295780 204627
rect 295480 204467 295780 204509
rect 295480 204349 295571 204467
rect 295689 204349 295780 204467
rect 295480 186627 295780 204349
rect 295480 186509 295571 186627
rect 295689 186509 295780 186627
rect 295480 186467 295780 186509
rect 295480 186349 295571 186467
rect 295689 186349 295780 186467
rect 295480 168627 295780 186349
rect 295480 168509 295571 168627
rect 295689 168509 295780 168627
rect 295480 168467 295780 168509
rect 295480 168349 295571 168467
rect 295689 168349 295780 168467
rect 295480 150627 295780 168349
rect 295480 150509 295571 150627
rect 295689 150509 295780 150627
rect 295480 150467 295780 150509
rect 295480 150349 295571 150467
rect 295689 150349 295780 150467
rect 295480 132627 295780 150349
rect 295480 132509 295571 132627
rect 295689 132509 295780 132627
rect 295480 132467 295780 132509
rect 295480 132349 295571 132467
rect 295689 132349 295780 132467
rect 295480 114627 295780 132349
rect 295480 114509 295571 114627
rect 295689 114509 295780 114627
rect 295480 114467 295780 114509
rect 295480 114349 295571 114467
rect 295689 114349 295780 114467
rect 295480 96627 295780 114349
rect 295480 96509 295571 96627
rect 295689 96509 295780 96627
rect 295480 96467 295780 96509
rect 295480 96349 295571 96467
rect 295689 96349 295780 96467
rect 295480 78627 295780 96349
rect 295480 78509 295571 78627
rect 295689 78509 295780 78627
rect 295480 78467 295780 78509
rect 295480 78349 295571 78467
rect 295689 78349 295780 78467
rect 295480 60627 295780 78349
rect 295480 60509 295571 60627
rect 295689 60509 295780 60627
rect 295480 60467 295780 60509
rect 295480 60349 295571 60467
rect 295689 60349 295780 60467
rect 295480 42627 295780 60349
rect 295480 42509 295571 42627
rect 295689 42509 295780 42627
rect 295480 42467 295780 42509
rect 295480 42349 295571 42467
rect 295689 42349 295780 42467
rect 295480 24627 295780 42349
rect 295480 24509 295571 24627
rect 295689 24509 295780 24627
rect 295480 24467 295780 24509
rect 295480 24349 295571 24467
rect 295689 24349 295780 24467
rect 295480 6627 295780 24349
rect 295480 6509 295571 6627
rect 295689 6509 295780 6627
rect 295480 6467 295780 6509
rect 295480 6349 295571 6467
rect 295689 6349 295780 6467
rect 295480 -2993 295780 6349
rect 295480 -3111 295571 -2993
rect 295689 -3111 295780 -2993
rect 295480 -3153 295780 -3111
rect 295480 -3271 295571 -3153
rect 295689 -3271 295780 -3153
rect 295480 -3282 295780 -3271
rect 295950 339627 296250 355431
rect 295950 339509 296041 339627
rect 296159 339509 296250 339627
rect 295950 339467 296250 339509
rect 295950 339349 296041 339467
rect 296159 339349 296250 339467
rect 295950 321627 296250 339349
rect 295950 321509 296041 321627
rect 296159 321509 296250 321627
rect 295950 321467 296250 321509
rect 295950 321349 296041 321467
rect 296159 321349 296250 321467
rect 295950 303627 296250 321349
rect 295950 303509 296041 303627
rect 296159 303509 296250 303627
rect 295950 303467 296250 303509
rect 295950 303349 296041 303467
rect 296159 303349 296250 303467
rect 295950 285627 296250 303349
rect 295950 285509 296041 285627
rect 296159 285509 296250 285627
rect 295950 285467 296250 285509
rect 295950 285349 296041 285467
rect 296159 285349 296250 285467
rect 295950 267627 296250 285349
rect 295950 267509 296041 267627
rect 296159 267509 296250 267627
rect 295950 267467 296250 267509
rect 295950 267349 296041 267467
rect 296159 267349 296250 267467
rect 295950 249627 296250 267349
rect 295950 249509 296041 249627
rect 296159 249509 296250 249627
rect 295950 249467 296250 249509
rect 295950 249349 296041 249467
rect 296159 249349 296250 249467
rect 295950 231627 296250 249349
rect 295950 231509 296041 231627
rect 296159 231509 296250 231627
rect 295950 231467 296250 231509
rect 295950 231349 296041 231467
rect 296159 231349 296250 231467
rect 295950 213627 296250 231349
rect 295950 213509 296041 213627
rect 296159 213509 296250 213627
rect 295950 213467 296250 213509
rect 295950 213349 296041 213467
rect 296159 213349 296250 213467
rect 295950 195627 296250 213349
rect 295950 195509 296041 195627
rect 296159 195509 296250 195627
rect 295950 195467 296250 195509
rect 295950 195349 296041 195467
rect 296159 195349 296250 195467
rect 295950 177627 296250 195349
rect 295950 177509 296041 177627
rect 296159 177509 296250 177627
rect 295950 177467 296250 177509
rect 295950 177349 296041 177467
rect 296159 177349 296250 177467
rect 295950 159627 296250 177349
rect 295950 159509 296041 159627
rect 296159 159509 296250 159627
rect 295950 159467 296250 159509
rect 295950 159349 296041 159467
rect 296159 159349 296250 159467
rect 295950 141627 296250 159349
rect 295950 141509 296041 141627
rect 296159 141509 296250 141627
rect 295950 141467 296250 141509
rect 295950 141349 296041 141467
rect 296159 141349 296250 141467
rect 295950 123627 296250 141349
rect 295950 123509 296041 123627
rect 296159 123509 296250 123627
rect 295950 123467 296250 123509
rect 295950 123349 296041 123467
rect 296159 123349 296250 123467
rect 295950 105627 296250 123349
rect 295950 105509 296041 105627
rect 296159 105509 296250 105627
rect 295950 105467 296250 105509
rect 295950 105349 296041 105467
rect 296159 105349 296250 105467
rect 295950 87627 296250 105349
rect 295950 87509 296041 87627
rect 296159 87509 296250 87627
rect 295950 87467 296250 87509
rect 295950 87349 296041 87467
rect 296159 87349 296250 87467
rect 295950 69627 296250 87349
rect 295950 69509 296041 69627
rect 296159 69509 296250 69627
rect 295950 69467 296250 69509
rect 295950 69349 296041 69467
rect 296159 69349 296250 69467
rect 295950 51627 296250 69349
rect 295950 51509 296041 51627
rect 296159 51509 296250 51627
rect 295950 51467 296250 51509
rect 295950 51349 296041 51467
rect 296159 51349 296250 51467
rect 295950 33627 296250 51349
rect 295950 33509 296041 33627
rect 296159 33509 296250 33627
rect 295950 33467 296250 33509
rect 295950 33349 296041 33467
rect 296159 33349 296250 33467
rect 295950 15627 296250 33349
rect 295950 15509 296041 15627
rect 296159 15509 296250 15627
rect 295950 15467 296250 15509
rect 295950 15349 296041 15467
rect 296159 15349 296250 15467
rect 284802 -3581 284893 -3463
rect 285011 -3581 285102 -3463
rect 284802 -3623 285102 -3581
rect 284802 -3741 284893 -3623
rect 285011 -3741 285102 -3623
rect 284802 -3752 285102 -3741
rect 295950 -3463 296250 15349
rect 295950 -3581 296041 -3463
rect 296159 -3581 296250 -3463
rect 295950 -3623 296250 -3581
rect 295950 -3741 296041 -3623
rect 296159 -3741 296250 -3623
rect 295950 -3752 296250 -3741
<< via4 >>
rect -4197 355591 -4079 355709
rect -4197 355431 -4079 355549
rect -4197 339509 -4079 339627
rect -4197 339349 -4079 339467
rect -4197 321509 -4079 321627
rect -4197 321349 -4079 321467
rect -4197 303509 -4079 303627
rect -4197 303349 -4079 303467
rect -4197 285509 -4079 285627
rect -4197 285349 -4079 285467
rect -4197 267509 -4079 267627
rect -4197 267349 -4079 267467
rect -4197 249509 -4079 249627
rect -4197 249349 -4079 249467
rect -4197 231509 -4079 231627
rect -4197 231349 -4079 231467
rect -4197 213509 -4079 213627
rect -4197 213349 -4079 213467
rect -4197 195509 -4079 195627
rect -4197 195349 -4079 195467
rect -4197 177509 -4079 177627
rect -4197 177349 -4079 177467
rect -4197 159509 -4079 159627
rect -4197 159349 -4079 159467
rect -4197 141509 -4079 141627
rect -4197 141349 -4079 141467
rect -4197 123509 -4079 123627
rect -4197 123349 -4079 123467
rect -4197 105509 -4079 105627
rect -4197 105349 -4079 105467
rect -4197 87509 -4079 87627
rect -4197 87349 -4079 87467
rect -4197 69509 -4079 69627
rect -4197 69349 -4079 69467
rect -4197 51509 -4079 51627
rect -4197 51349 -4079 51467
rect -4197 33509 -4079 33627
rect -4197 33349 -4079 33467
rect -4197 15509 -4079 15627
rect -4197 15349 -4079 15467
rect -3727 355121 -3609 355239
rect -3727 354961 -3609 355079
rect 5893 355121 6011 355239
rect 5893 354961 6011 355079
rect -3727 348509 -3609 348627
rect -3727 348349 -3609 348467
rect -3727 330509 -3609 330627
rect -3727 330349 -3609 330467
rect -3727 312509 -3609 312627
rect -3727 312349 -3609 312467
rect -3727 294509 -3609 294627
rect -3727 294349 -3609 294467
rect -3727 276509 -3609 276627
rect -3727 276349 -3609 276467
rect -3727 258509 -3609 258627
rect -3727 258349 -3609 258467
rect -3727 240509 -3609 240627
rect -3727 240349 -3609 240467
rect -3727 222509 -3609 222627
rect -3727 222349 -3609 222467
rect -3727 204509 -3609 204627
rect -3727 204349 -3609 204467
rect -3727 186509 -3609 186627
rect -3727 186349 -3609 186467
rect -3727 168509 -3609 168627
rect -3727 168349 -3609 168467
rect -3727 150509 -3609 150627
rect -3727 150349 -3609 150467
rect -3727 132509 -3609 132627
rect -3727 132349 -3609 132467
rect -3727 114509 -3609 114627
rect -3727 114349 -3609 114467
rect -3727 96509 -3609 96627
rect -3727 96349 -3609 96467
rect -3727 78509 -3609 78627
rect -3727 78349 -3609 78467
rect -3727 60509 -3609 60627
rect -3727 60349 -3609 60467
rect -3727 42509 -3609 42627
rect -3727 42349 -3609 42467
rect -3727 24509 -3609 24627
rect -3727 24349 -3609 24467
rect -3727 6509 -3609 6627
rect -3727 6349 -3609 6467
rect -3257 354651 -3139 354769
rect -3257 354491 -3139 354609
rect -3257 337709 -3139 337827
rect -3257 337549 -3139 337667
rect -3257 319709 -3139 319827
rect -3257 319549 -3139 319667
rect -3257 301709 -3139 301827
rect -3257 301549 -3139 301667
rect -3257 283709 -3139 283827
rect -3257 283549 -3139 283667
rect -3257 265709 -3139 265827
rect -3257 265549 -3139 265667
rect -3257 247709 -3139 247827
rect -3257 247549 -3139 247667
rect -3257 229709 -3139 229827
rect -3257 229549 -3139 229667
rect -3257 211709 -3139 211827
rect -3257 211549 -3139 211667
rect -3257 193709 -3139 193827
rect -3257 193549 -3139 193667
rect -3257 175709 -3139 175827
rect -3257 175549 -3139 175667
rect -3257 157709 -3139 157827
rect -3257 157549 -3139 157667
rect -3257 139709 -3139 139827
rect -3257 139549 -3139 139667
rect -3257 121709 -3139 121827
rect -3257 121549 -3139 121667
rect -3257 103709 -3139 103827
rect -3257 103549 -3139 103667
rect -3257 85709 -3139 85827
rect -3257 85549 -3139 85667
rect -3257 67709 -3139 67827
rect -3257 67549 -3139 67667
rect -3257 49709 -3139 49827
rect -3257 49549 -3139 49667
rect -3257 31709 -3139 31827
rect -3257 31549 -3139 31667
rect -3257 13709 -3139 13827
rect -3257 13549 -3139 13667
rect -2787 354181 -2669 354299
rect -2787 354021 -2669 354139
rect 4093 354181 4211 354299
rect 4093 354021 4211 354139
rect -2787 346709 -2669 346827
rect -2787 346549 -2669 346667
rect -2787 328709 -2669 328827
rect -2787 328549 -2669 328667
rect -2787 310709 -2669 310827
rect -2787 310549 -2669 310667
rect -2787 292709 -2669 292827
rect -2787 292549 -2669 292667
rect -2787 274709 -2669 274827
rect -2787 274549 -2669 274667
rect -2787 256709 -2669 256827
rect -2787 256549 -2669 256667
rect -2787 238709 -2669 238827
rect -2787 238549 -2669 238667
rect -2787 220709 -2669 220827
rect -2787 220549 -2669 220667
rect -2787 202709 -2669 202827
rect -2787 202549 -2669 202667
rect -2787 184709 -2669 184827
rect -2787 184549 -2669 184667
rect -2787 166709 -2669 166827
rect -2787 166549 -2669 166667
rect -2787 148709 -2669 148827
rect -2787 148549 -2669 148667
rect -2787 130709 -2669 130827
rect -2787 130549 -2669 130667
rect -2787 112709 -2669 112827
rect -2787 112549 -2669 112667
rect -2787 94709 -2669 94827
rect -2787 94549 -2669 94667
rect -2787 76709 -2669 76827
rect -2787 76549 -2669 76667
rect -2787 58709 -2669 58827
rect -2787 58549 -2669 58667
rect -2787 40709 -2669 40827
rect -2787 40549 -2669 40667
rect -2787 22709 -2669 22827
rect -2787 22549 -2669 22667
rect -2787 4709 -2669 4827
rect -2787 4549 -2669 4667
rect -2317 353711 -2199 353829
rect -2317 353551 -2199 353669
rect -2317 335909 -2199 336027
rect -2317 335749 -2199 335867
rect -2317 317909 -2199 318027
rect -2317 317749 -2199 317867
rect -2317 299909 -2199 300027
rect -2317 299749 -2199 299867
rect -2317 281909 -2199 282027
rect -2317 281749 -2199 281867
rect -2317 263909 -2199 264027
rect -2317 263749 -2199 263867
rect -2317 245909 -2199 246027
rect -2317 245749 -2199 245867
rect -2317 227909 -2199 228027
rect -2317 227749 -2199 227867
rect -2317 209909 -2199 210027
rect -2317 209749 -2199 209867
rect -2317 191909 -2199 192027
rect -2317 191749 -2199 191867
rect -2317 173909 -2199 174027
rect -2317 173749 -2199 173867
rect -2317 155909 -2199 156027
rect -2317 155749 -2199 155867
rect -2317 137909 -2199 138027
rect -2317 137749 -2199 137867
rect -2317 119909 -2199 120027
rect -2317 119749 -2199 119867
rect -2317 101909 -2199 102027
rect -2317 101749 -2199 101867
rect -2317 83909 -2199 84027
rect -2317 83749 -2199 83867
rect -2317 65909 -2199 66027
rect -2317 65749 -2199 65867
rect -2317 47909 -2199 48027
rect -2317 47749 -2199 47867
rect -2317 29909 -2199 30027
rect -2317 29749 -2199 29867
rect -2317 11909 -2199 12027
rect -2317 11749 -2199 11867
rect -1847 353241 -1729 353359
rect -1847 353081 -1729 353199
rect 2293 353241 2411 353359
rect 2293 353081 2411 353199
rect -1847 344909 -1729 345027
rect -1847 344749 -1729 344867
rect -1847 326909 -1729 327027
rect -1847 326749 -1729 326867
rect -1847 308909 -1729 309027
rect -1847 308749 -1729 308867
rect -1847 290909 -1729 291027
rect -1847 290749 -1729 290867
rect -1847 272909 -1729 273027
rect -1847 272749 -1729 272867
rect -1847 254909 -1729 255027
rect -1847 254749 -1729 254867
rect -1847 236909 -1729 237027
rect -1847 236749 -1729 236867
rect -1847 218909 -1729 219027
rect -1847 218749 -1729 218867
rect -1847 200909 -1729 201027
rect -1847 200749 -1729 200867
rect -1847 182909 -1729 183027
rect -1847 182749 -1729 182867
rect -1847 164909 -1729 165027
rect -1847 164749 -1729 164867
rect -1847 146909 -1729 147027
rect -1847 146749 -1729 146867
rect -1847 128909 -1729 129027
rect -1847 128749 -1729 128867
rect -1847 110909 -1729 111027
rect -1847 110749 -1729 110867
rect -1847 92909 -1729 93027
rect -1847 92749 -1729 92867
rect -1847 74909 -1729 75027
rect -1847 74749 -1729 74867
rect -1847 56909 -1729 57027
rect -1847 56749 -1729 56867
rect -1847 38909 -1729 39027
rect -1847 38749 -1729 38867
rect -1847 20909 -1729 21027
rect -1847 20749 -1729 20867
rect -1847 2909 -1729 3027
rect -1847 2749 -1729 2867
rect -1377 352771 -1259 352889
rect -1377 352611 -1259 352729
rect -1377 334109 -1259 334227
rect -1377 333949 -1259 334067
rect -1377 316109 -1259 316227
rect -1377 315949 -1259 316067
rect -1377 298109 -1259 298227
rect -1377 297949 -1259 298067
rect -1377 280109 -1259 280227
rect -1377 279949 -1259 280067
rect -1377 262109 -1259 262227
rect -1377 261949 -1259 262067
rect -1377 244109 -1259 244227
rect -1377 243949 -1259 244067
rect -1377 226109 -1259 226227
rect -1377 225949 -1259 226067
rect -1377 208109 -1259 208227
rect -1377 207949 -1259 208067
rect -1377 190109 -1259 190227
rect -1377 189949 -1259 190067
rect -1377 172109 -1259 172227
rect -1377 171949 -1259 172067
rect -1377 154109 -1259 154227
rect -1377 153949 -1259 154067
rect -1377 136109 -1259 136227
rect -1377 135949 -1259 136067
rect -1377 118109 -1259 118227
rect -1377 117949 -1259 118067
rect -1377 100109 -1259 100227
rect -1377 99949 -1259 100067
rect -1377 82109 -1259 82227
rect -1377 81949 -1259 82067
rect -1377 64109 -1259 64227
rect -1377 63949 -1259 64067
rect -1377 46109 -1259 46227
rect -1377 45949 -1259 46067
rect -1377 28109 -1259 28227
rect -1377 27949 -1259 28067
rect -1377 10109 -1259 10227
rect -1377 9949 -1259 10067
rect -907 352301 -789 352419
rect -907 352141 -789 352259
rect 493 352301 611 352419
rect 493 352141 611 352259
rect 14893 355591 15011 355709
rect 14893 355431 15011 355549
rect 13093 354651 13211 354769
rect 13093 354491 13211 354609
rect 11293 353711 11411 353829
rect 11293 353551 11411 353669
rect 9493 352771 9611 352889
rect 9493 352611 9611 352729
rect 23893 355121 24011 355239
rect 23893 354961 24011 355079
rect 22093 354181 22211 354299
rect 22093 354021 22211 354139
rect 20293 353241 20411 353359
rect 20293 353081 20411 353199
rect 18493 352301 18611 352419
rect 18493 352141 18611 352259
rect 32893 355591 33011 355709
rect 32893 355431 33011 355549
rect 31093 354651 31211 354769
rect 31093 354491 31211 354609
rect 29293 353711 29411 353829
rect 29293 353551 29411 353669
rect 27493 352771 27611 352889
rect 27493 352611 27611 352729
rect 41893 355121 42011 355239
rect 41893 354961 42011 355079
rect 40093 354181 40211 354299
rect 40093 354021 40211 354139
rect 38293 353241 38411 353359
rect 38293 353081 38411 353199
rect 36493 352301 36611 352419
rect 36493 352141 36611 352259
rect 50893 355591 51011 355709
rect 50893 355431 51011 355549
rect 49093 354651 49211 354769
rect 49093 354491 49211 354609
rect 47293 353711 47411 353829
rect 47293 353551 47411 353669
rect 45493 352771 45611 352889
rect 45493 352611 45611 352729
rect 59893 355121 60011 355239
rect 59893 354961 60011 355079
rect 58093 354181 58211 354299
rect 58093 354021 58211 354139
rect 56293 353241 56411 353359
rect 56293 353081 56411 353199
rect 54493 352301 54611 352419
rect 54493 352141 54611 352259
rect 68893 355591 69011 355709
rect 68893 355431 69011 355549
rect 67093 354651 67211 354769
rect 67093 354491 67211 354609
rect 65293 353711 65411 353829
rect 65293 353551 65411 353669
rect 63493 352771 63611 352889
rect 63493 352611 63611 352729
rect 77893 355121 78011 355239
rect 77893 354961 78011 355079
rect 76093 354181 76211 354299
rect 76093 354021 76211 354139
rect 74293 353241 74411 353359
rect 74293 353081 74411 353199
rect 72493 352301 72611 352419
rect 72493 352141 72611 352259
rect 86893 355591 87011 355709
rect 86893 355431 87011 355549
rect 85093 354651 85211 354769
rect 85093 354491 85211 354609
rect 83293 353711 83411 353829
rect 83293 353551 83411 353669
rect 81493 352771 81611 352889
rect 81493 352611 81611 352729
rect 95893 355121 96011 355239
rect 95893 354961 96011 355079
rect 94093 354181 94211 354299
rect 94093 354021 94211 354139
rect 92293 353241 92411 353359
rect 92293 353081 92411 353199
rect 90493 352301 90611 352419
rect 90493 352141 90611 352259
rect 104893 355591 105011 355709
rect 104893 355431 105011 355549
rect 103093 354651 103211 354769
rect 103093 354491 103211 354609
rect 101293 353711 101411 353829
rect 101293 353551 101411 353669
rect 99493 352771 99611 352889
rect 99493 352611 99611 352729
rect 113893 355121 114011 355239
rect 113893 354961 114011 355079
rect 112093 354181 112211 354299
rect 112093 354021 112211 354139
rect 110293 353241 110411 353359
rect 110293 353081 110411 353199
rect 108493 352301 108611 352419
rect 108493 352141 108611 352259
rect 122893 355591 123011 355709
rect 122893 355431 123011 355549
rect 121093 354651 121211 354769
rect 121093 354491 121211 354609
rect 119293 353711 119411 353829
rect 119293 353551 119411 353669
rect 117493 352771 117611 352889
rect 117493 352611 117611 352729
rect 131893 355121 132011 355239
rect 131893 354961 132011 355079
rect 130093 354181 130211 354299
rect 130093 354021 130211 354139
rect 128293 353241 128411 353359
rect 128293 353081 128411 353199
rect 126493 352301 126611 352419
rect 126493 352141 126611 352259
rect 140893 355591 141011 355709
rect 140893 355431 141011 355549
rect 139093 354651 139211 354769
rect 139093 354491 139211 354609
rect 137293 353711 137411 353829
rect 137293 353551 137411 353669
rect 135493 352771 135611 352889
rect 135493 352611 135611 352729
rect 149893 355121 150011 355239
rect 149893 354961 150011 355079
rect 148093 354181 148211 354299
rect 148093 354021 148211 354139
rect 146293 353241 146411 353359
rect 146293 353081 146411 353199
rect 144493 352301 144611 352419
rect 144493 352141 144611 352259
rect 158893 355591 159011 355709
rect 158893 355431 159011 355549
rect 157093 354651 157211 354769
rect 157093 354491 157211 354609
rect 155293 353711 155411 353829
rect 155293 353551 155411 353669
rect 153493 352771 153611 352889
rect 153493 352611 153611 352729
rect 167893 355121 168011 355239
rect 167893 354961 168011 355079
rect 166093 354181 166211 354299
rect 166093 354021 166211 354139
rect 164293 353241 164411 353359
rect 164293 353081 164411 353199
rect 162493 352301 162611 352419
rect 162493 352141 162611 352259
rect 176893 355591 177011 355709
rect 176893 355431 177011 355549
rect 175093 354651 175211 354769
rect 175093 354491 175211 354609
rect 173293 353711 173411 353829
rect 173293 353551 173411 353669
rect 171493 352771 171611 352889
rect 171493 352611 171611 352729
rect 185893 355121 186011 355239
rect 185893 354961 186011 355079
rect 184093 354181 184211 354299
rect 184093 354021 184211 354139
rect 182293 353241 182411 353359
rect 182293 353081 182411 353199
rect 180493 352301 180611 352419
rect 180493 352141 180611 352259
rect 194893 355591 195011 355709
rect 194893 355431 195011 355549
rect 193093 354651 193211 354769
rect 193093 354491 193211 354609
rect 191293 353711 191411 353829
rect 191293 353551 191411 353669
rect 189493 352771 189611 352889
rect 189493 352611 189611 352729
rect 203893 355121 204011 355239
rect 203893 354961 204011 355079
rect 202093 354181 202211 354299
rect 202093 354021 202211 354139
rect 200293 353241 200411 353359
rect 200293 353081 200411 353199
rect 198493 352301 198611 352419
rect 198493 352141 198611 352259
rect 212893 355591 213011 355709
rect 212893 355431 213011 355549
rect 211093 354651 211211 354769
rect 211093 354491 211211 354609
rect 209293 353711 209411 353829
rect 209293 353551 209411 353669
rect 207493 352771 207611 352889
rect 207493 352611 207611 352729
rect 221893 355121 222011 355239
rect 221893 354961 222011 355079
rect 220093 354181 220211 354299
rect 220093 354021 220211 354139
rect 218293 353241 218411 353359
rect 218293 353081 218411 353199
rect 216493 352301 216611 352419
rect 216493 352141 216611 352259
rect 230893 355591 231011 355709
rect 230893 355431 231011 355549
rect 229093 354651 229211 354769
rect 229093 354491 229211 354609
rect 227293 353711 227411 353829
rect 227293 353551 227411 353669
rect 225493 352771 225611 352889
rect 225493 352611 225611 352729
rect 239893 355121 240011 355239
rect 239893 354961 240011 355079
rect 238093 354181 238211 354299
rect 238093 354021 238211 354139
rect 236293 353241 236411 353359
rect 236293 353081 236411 353199
rect 234493 352301 234611 352419
rect 234493 352141 234611 352259
rect 248893 355591 249011 355709
rect 248893 355431 249011 355549
rect 247093 354651 247211 354769
rect 247093 354491 247211 354609
rect 245293 353711 245411 353829
rect 245293 353551 245411 353669
rect 243493 352771 243611 352889
rect 243493 352611 243611 352729
rect 257893 355121 258011 355239
rect 257893 354961 258011 355079
rect 256093 354181 256211 354299
rect 256093 354021 256211 354139
rect 254293 353241 254411 353359
rect 254293 353081 254411 353199
rect 252493 352301 252611 352419
rect 252493 352141 252611 352259
rect 266893 355591 267011 355709
rect 266893 355431 267011 355549
rect 265093 354651 265211 354769
rect 265093 354491 265211 354609
rect 263293 353711 263411 353829
rect 263293 353551 263411 353669
rect 261493 352771 261611 352889
rect 261493 352611 261611 352729
rect 275893 355121 276011 355239
rect 275893 354961 276011 355079
rect 274093 354181 274211 354299
rect 274093 354021 274211 354139
rect 272293 353241 272411 353359
rect 272293 353081 272411 353199
rect 270493 352301 270611 352419
rect 270493 352141 270611 352259
rect 284893 355591 285011 355709
rect 284893 355431 285011 355549
rect 283093 354651 283211 354769
rect 283093 354491 283211 354609
rect 281293 353711 281411 353829
rect 281293 353551 281411 353669
rect 279493 352771 279611 352889
rect 279493 352611 279611 352729
rect 296041 355591 296159 355709
rect 296041 355431 296159 355549
rect 295571 355121 295689 355239
rect 295571 354961 295689 355079
rect 295101 354651 295219 354769
rect 295101 354491 295219 354609
rect 294631 354181 294749 354299
rect 294631 354021 294749 354139
rect 294161 353711 294279 353829
rect 294161 353551 294279 353669
rect 290293 353241 290411 353359
rect 290293 353081 290411 353199
rect 288493 352301 288611 352419
rect 288493 352141 288611 352259
rect 293691 353241 293809 353359
rect 293691 353081 293809 353199
rect 293221 352771 293339 352889
rect 293221 352611 293339 352729
rect 292751 352301 292869 352419
rect 292751 352141 292869 352259
rect -907 343109 -789 343227
rect -907 342949 -789 343067
rect -907 325109 -789 325227
rect -907 324949 -789 325067
rect -907 307109 -789 307227
rect -907 306949 -789 307067
rect -907 289109 -789 289227
rect -907 288949 -789 289067
rect -907 271109 -789 271227
rect -907 270949 -789 271067
rect -907 253109 -789 253227
rect -907 252949 -789 253067
rect -907 235109 -789 235227
rect -907 234949 -789 235067
rect -907 217109 -789 217227
rect -907 216949 -789 217067
rect -907 199109 -789 199227
rect -907 198949 -789 199067
rect -907 181109 -789 181227
rect -907 180949 -789 181067
rect -907 163109 -789 163227
rect -907 162949 -789 163067
rect -907 145109 -789 145227
rect -907 144949 -789 145067
rect -907 127109 -789 127227
rect -907 126949 -789 127067
rect -907 109109 -789 109227
rect -907 108949 -789 109067
rect -907 91109 -789 91227
rect -907 90949 -789 91067
rect -907 73109 -789 73227
rect -907 72949 -789 73067
rect -907 55109 -789 55227
rect -907 54949 -789 55067
rect -907 37109 -789 37227
rect -907 36949 -789 37067
rect -907 19109 -789 19227
rect -907 18949 -789 19067
rect -907 1109 -789 1227
rect -907 949 -789 1067
rect 292751 343109 292869 343227
rect 292751 342949 292869 343067
rect 292751 325109 292869 325227
rect 292751 324949 292869 325067
rect 292751 307109 292869 307227
rect 292751 306949 292869 307067
rect 292751 289109 292869 289227
rect 292751 288949 292869 289067
rect 292751 271109 292869 271227
rect 292751 270949 292869 271067
rect 292751 253109 292869 253227
rect 292751 252949 292869 253067
rect 292751 235109 292869 235227
rect 292751 234949 292869 235067
rect 292751 217109 292869 217227
rect 292751 216949 292869 217067
rect 292751 199109 292869 199227
rect 292751 198949 292869 199067
rect 292751 181109 292869 181227
rect 292751 180949 292869 181067
rect 292751 163109 292869 163227
rect 292751 162949 292869 163067
rect 292751 145109 292869 145227
rect 292751 144949 292869 145067
rect 292751 127109 292869 127227
rect 292751 126949 292869 127067
rect 292751 109109 292869 109227
rect 292751 108949 292869 109067
rect 292751 91109 292869 91227
rect 292751 90949 292869 91067
rect 292751 73109 292869 73227
rect 292751 72949 292869 73067
rect 292751 55109 292869 55227
rect 292751 54949 292869 55067
rect 292751 37109 292869 37227
rect 292751 36949 292869 37067
rect 292751 19109 292869 19227
rect 292751 18949 292869 19067
rect 292751 1109 292869 1227
rect 292751 949 292869 1067
rect -907 -291 -789 -173
rect -907 -451 -789 -333
rect 493 -291 611 -173
rect 493 -451 611 -333
rect -1377 -761 -1259 -643
rect -1377 -921 -1259 -803
rect -1847 -1231 -1729 -1113
rect -1847 -1391 -1729 -1273
rect 2293 -1231 2411 -1113
rect 2293 -1391 2411 -1273
rect -2317 -1701 -2199 -1583
rect -2317 -1861 -2199 -1743
rect -2787 -2171 -2669 -2053
rect -2787 -2331 -2669 -2213
rect 4093 -2171 4211 -2053
rect 4093 -2331 4211 -2213
rect -3257 -2641 -3139 -2523
rect -3257 -2801 -3139 -2683
rect -3727 -3111 -3609 -2993
rect -3727 -3271 -3609 -3153
rect 9493 -761 9611 -643
rect 9493 -921 9611 -803
rect 11293 -1701 11411 -1583
rect 11293 -1861 11411 -1743
rect 13093 -2641 13211 -2523
rect 13093 -2801 13211 -2683
rect 5893 -3111 6011 -2993
rect 5893 -3271 6011 -3153
rect -4197 -3581 -4079 -3463
rect -4197 -3741 -4079 -3623
rect 18493 -291 18611 -173
rect 18493 -451 18611 -333
rect 20293 -1231 20411 -1113
rect 20293 -1391 20411 -1273
rect 22093 -2171 22211 -2053
rect 22093 -2331 22211 -2213
rect 14893 -3581 15011 -3463
rect 14893 -3741 15011 -3623
rect 27493 -761 27611 -643
rect 27493 -921 27611 -803
rect 29293 -1701 29411 -1583
rect 29293 -1861 29411 -1743
rect 31093 -2641 31211 -2523
rect 31093 -2801 31211 -2683
rect 23893 -3111 24011 -2993
rect 23893 -3271 24011 -3153
rect 36493 -291 36611 -173
rect 36493 -451 36611 -333
rect 38293 -1231 38411 -1113
rect 38293 -1391 38411 -1273
rect 40093 -2171 40211 -2053
rect 40093 -2331 40211 -2213
rect 32893 -3581 33011 -3463
rect 32893 -3741 33011 -3623
rect 45493 -761 45611 -643
rect 45493 -921 45611 -803
rect 47293 -1701 47411 -1583
rect 47293 -1861 47411 -1743
rect 49093 -2641 49211 -2523
rect 49093 -2801 49211 -2683
rect 41893 -3111 42011 -2993
rect 41893 -3271 42011 -3153
rect 54493 -291 54611 -173
rect 54493 -451 54611 -333
rect 56293 -1231 56411 -1113
rect 56293 -1391 56411 -1273
rect 58093 -2171 58211 -2053
rect 58093 -2331 58211 -2213
rect 50893 -3581 51011 -3463
rect 50893 -3741 51011 -3623
rect 63493 -761 63611 -643
rect 63493 -921 63611 -803
rect 65293 -1701 65411 -1583
rect 65293 -1861 65411 -1743
rect 67093 -2641 67211 -2523
rect 67093 -2801 67211 -2683
rect 59893 -3111 60011 -2993
rect 59893 -3271 60011 -3153
rect 72493 -291 72611 -173
rect 72493 -451 72611 -333
rect 74293 -1231 74411 -1113
rect 74293 -1391 74411 -1273
rect 76093 -2171 76211 -2053
rect 76093 -2331 76211 -2213
rect 68893 -3581 69011 -3463
rect 68893 -3741 69011 -3623
rect 81493 -761 81611 -643
rect 81493 -921 81611 -803
rect 83293 -1701 83411 -1583
rect 83293 -1861 83411 -1743
rect 85093 -2641 85211 -2523
rect 85093 -2801 85211 -2683
rect 77893 -3111 78011 -2993
rect 77893 -3271 78011 -3153
rect 90493 -291 90611 -173
rect 90493 -451 90611 -333
rect 92293 -1231 92411 -1113
rect 92293 -1391 92411 -1273
rect 94093 -2171 94211 -2053
rect 94093 -2331 94211 -2213
rect 86893 -3581 87011 -3463
rect 86893 -3741 87011 -3623
rect 99493 -761 99611 -643
rect 99493 -921 99611 -803
rect 101293 -1701 101411 -1583
rect 101293 -1861 101411 -1743
rect 103093 -2641 103211 -2523
rect 103093 -2801 103211 -2683
rect 95893 -3111 96011 -2993
rect 95893 -3271 96011 -3153
rect 108493 -291 108611 -173
rect 108493 -451 108611 -333
rect 110293 -1231 110411 -1113
rect 110293 -1391 110411 -1273
rect 112093 -2171 112211 -2053
rect 112093 -2331 112211 -2213
rect 104893 -3581 105011 -3463
rect 104893 -3741 105011 -3623
rect 117493 -761 117611 -643
rect 117493 -921 117611 -803
rect 119293 -1701 119411 -1583
rect 119293 -1861 119411 -1743
rect 121093 -2641 121211 -2523
rect 121093 -2801 121211 -2683
rect 113893 -3111 114011 -2993
rect 113893 -3271 114011 -3153
rect 126493 -291 126611 -173
rect 126493 -451 126611 -333
rect 128293 -1231 128411 -1113
rect 128293 -1391 128411 -1273
rect 130093 -2171 130211 -2053
rect 130093 -2331 130211 -2213
rect 122893 -3581 123011 -3463
rect 122893 -3741 123011 -3623
rect 135493 -761 135611 -643
rect 135493 -921 135611 -803
rect 137293 -1701 137411 -1583
rect 137293 -1861 137411 -1743
rect 139093 -2641 139211 -2523
rect 139093 -2801 139211 -2683
rect 131893 -3111 132011 -2993
rect 131893 -3271 132011 -3153
rect 144493 -291 144611 -173
rect 144493 -451 144611 -333
rect 146293 -1231 146411 -1113
rect 146293 -1391 146411 -1273
rect 148093 -2171 148211 -2053
rect 148093 -2331 148211 -2213
rect 140893 -3581 141011 -3463
rect 140893 -3741 141011 -3623
rect 153493 -761 153611 -643
rect 153493 -921 153611 -803
rect 155293 -1701 155411 -1583
rect 155293 -1861 155411 -1743
rect 157093 -2641 157211 -2523
rect 157093 -2801 157211 -2683
rect 149893 -3111 150011 -2993
rect 149893 -3271 150011 -3153
rect 162493 -291 162611 -173
rect 162493 -451 162611 -333
rect 164293 -1231 164411 -1113
rect 164293 -1391 164411 -1273
rect 166093 -2171 166211 -2053
rect 166093 -2331 166211 -2213
rect 158893 -3581 159011 -3463
rect 158893 -3741 159011 -3623
rect 171493 -761 171611 -643
rect 171493 -921 171611 -803
rect 173293 -1701 173411 -1583
rect 173293 -1861 173411 -1743
rect 175093 -2641 175211 -2523
rect 175093 -2801 175211 -2683
rect 167893 -3111 168011 -2993
rect 167893 -3271 168011 -3153
rect 180493 -291 180611 -173
rect 180493 -451 180611 -333
rect 182293 -1231 182411 -1113
rect 182293 -1391 182411 -1273
rect 184093 -2171 184211 -2053
rect 184093 -2331 184211 -2213
rect 176893 -3581 177011 -3463
rect 176893 -3741 177011 -3623
rect 189493 -761 189611 -643
rect 189493 -921 189611 -803
rect 191293 -1701 191411 -1583
rect 191293 -1861 191411 -1743
rect 193093 -2641 193211 -2523
rect 193093 -2801 193211 -2683
rect 185893 -3111 186011 -2993
rect 185893 -3271 186011 -3153
rect 198493 -291 198611 -173
rect 198493 -451 198611 -333
rect 200293 -1231 200411 -1113
rect 200293 -1391 200411 -1273
rect 202093 -2171 202211 -2053
rect 202093 -2331 202211 -2213
rect 194893 -3581 195011 -3463
rect 194893 -3741 195011 -3623
rect 207493 -761 207611 -643
rect 207493 -921 207611 -803
rect 209293 -1701 209411 -1583
rect 209293 -1861 209411 -1743
rect 211093 -2641 211211 -2523
rect 211093 -2801 211211 -2683
rect 203893 -3111 204011 -2993
rect 203893 -3271 204011 -3153
rect 216493 -291 216611 -173
rect 216493 -451 216611 -333
rect 218293 -1231 218411 -1113
rect 218293 -1391 218411 -1273
rect 220093 -2171 220211 -2053
rect 220093 -2331 220211 -2213
rect 212893 -3581 213011 -3463
rect 212893 -3741 213011 -3623
rect 225493 -761 225611 -643
rect 225493 -921 225611 -803
rect 227293 -1701 227411 -1583
rect 227293 -1861 227411 -1743
rect 229093 -2641 229211 -2523
rect 229093 -2801 229211 -2683
rect 221893 -3111 222011 -2993
rect 221893 -3271 222011 -3153
rect 234493 -291 234611 -173
rect 234493 -451 234611 -333
rect 236293 -1231 236411 -1113
rect 236293 -1391 236411 -1273
rect 238093 -2171 238211 -2053
rect 238093 -2331 238211 -2213
rect 230893 -3581 231011 -3463
rect 230893 -3741 231011 -3623
rect 243493 -761 243611 -643
rect 243493 -921 243611 -803
rect 245293 -1701 245411 -1583
rect 245293 -1861 245411 -1743
rect 247093 -2641 247211 -2523
rect 247093 -2801 247211 -2683
rect 239893 -3111 240011 -2993
rect 239893 -3271 240011 -3153
rect 252493 -291 252611 -173
rect 252493 -451 252611 -333
rect 254293 -1231 254411 -1113
rect 254293 -1391 254411 -1273
rect 256093 -2171 256211 -2053
rect 256093 -2331 256211 -2213
rect 248893 -3581 249011 -3463
rect 248893 -3741 249011 -3623
rect 261493 -761 261611 -643
rect 261493 -921 261611 -803
rect 263293 -1701 263411 -1583
rect 263293 -1861 263411 -1743
rect 265093 -2641 265211 -2523
rect 265093 -2801 265211 -2683
rect 257893 -3111 258011 -2993
rect 257893 -3271 258011 -3153
rect 270493 -291 270611 -173
rect 270493 -451 270611 -333
rect 272293 -1231 272411 -1113
rect 272293 -1391 272411 -1273
rect 274093 -2171 274211 -2053
rect 274093 -2331 274211 -2213
rect 266893 -3581 267011 -3463
rect 266893 -3741 267011 -3623
rect 279493 -761 279611 -643
rect 279493 -921 279611 -803
rect 281293 -1701 281411 -1583
rect 281293 -1861 281411 -1743
rect 283093 -2641 283211 -2523
rect 283093 -2801 283211 -2683
rect 275893 -3111 276011 -2993
rect 275893 -3271 276011 -3153
rect 288493 -291 288611 -173
rect 288493 -451 288611 -333
rect 292751 -291 292869 -173
rect 292751 -451 292869 -333
rect 293221 334109 293339 334227
rect 293221 333949 293339 334067
rect 293221 316109 293339 316227
rect 293221 315949 293339 316067
rect 293221 298109 293339 298227
rect 293221 297949 293339 298067
rect 293221 280109 293339 280227
rect 293221 279949 293339 280067
rect 293221 262109 293339 262227
rect 293221 261949 293339 262067
rect 293221 244109 293339 244227
rect 293221 243949 293339 244067
rect 293221 226109 293339 226227
rect 293221 225949 293339 226067
rect 293221 208109 293339 208227
rect 293221 207949 293339 208067
rect 293221 190109 293339 190227
rect 293221 189949 293339 190067
rect 293221 172109 293339 172227
rect 293221 171949 293339 172067
rect 293221 154109 293339 154227
rect 293221 153949 293339 154067
rect 293221 136109 293339 136227
rect 293221 135949 293339 136067
rect 293221 118109 293339 118227
rect 293221 117949 293339 118067
rect 293221 100109 293339 100227
rect 293221 99949 293339 100067
rect 293221 82109 293339 82227
rect 293221 81949 293339 82067
rect 293221 64109 293339 64227
rect 293221 63949 293339 64067
rect 293221 46109 293339 46227
rect 293221 45949 293339 46067
rect 293221 28109 293339 28227
rect 293221 27949 293339 28067
rect 293221 10109 293339 10227
rect 293221 9949 293339 10067
rect 293221 -761 293339 -643
rect 293221 -921 293339 -803
rect 293691 344909 293809 345027
rect 293691 344749 293809 344867
rect 293691 326909 293809 327027
rect 293691 326749 293809 326867
rect 293691 308909 293809 309027
rect 293691 308749 293809 308867
rect 293691 290909 293809 291027
rect 293691 290749 293809 290867
rect 293691 272909 293809 273027
rect 293691 272749 293809 272867
rect 293691 254909 293809 255027
rect 293691 254749 293809 254867
rect 293691 236909 293809 237027
rect 293691 236749 293809 236867
rect 293691 218909 293809 219027
rect 293691 218749 293809 218867
rect 293691 200909 293809 201027
rect 293691 200749 293809 200867
rect 293691 182909 293809 183027
rect 293691 182749 293809 182867
rect 293691 164909 293809 165027
rect 293691 164749 293809 164867
rect 293691 146909 293809 147027
rect 293691 146749 293809 146867
rect 293691 128909 293809 129027
rect 293691 128749 293809 128867
rect 293691 110909 293809 111027
rect 293691 110749 293809 110867
rect 293691 92909 293809 93027
rect 293691 92749 293809 92867
rect 293691 74909 293809 75027
rect 293691 74749 293809 74867
rect 293691 56909 293809 57027
rect 293691 56749 293809 56867
rect 293691 38909 293809 39027
rect 293691 38749 293809 38867
rect 293691 20909 293809 21027
rect 293691 20749 293809 20867
rect 293691 2909 293809 3027
rect 293691 2749 293809 2867
rect 290293 -1231 290411 -1113
rect 290293 -1391 290411 -1273
rect 293691 -1231 293809 -1113
rect 293691 -1391 293809 -1273
rect 294161 335909 294279 336027
rect 294161 335749 294279 335867
rect 294161 317909 294279 318027
rect 294161 317749 294279 317867
rect 294161 299909 294279 300027
rect 294161 299749 294279 299867
rect 294161 281909 294279 282027
rect 294161 281749 294279 281867
rect 294161 263909 294279 264027
rect 294161 263749 294279 263867
rect 294161 245909 294279 246027
rect 294161 245749 294279 245867
rect 294161 227909 294279 228027
rect 294161 227749 294279 227867
rect 294161 209909 294279 210027
rect 294161 209749 294279 209867
rect 294161 191909 294279 192027
rect 294161 191749 294279 191867
rect 294161 173909 294279 174027
rect 294161 173749 294279 173867
rect 294161 155909 294279 156027
rect 294161 155749 294279 155867
rect 294161 137909 294279 138027
rect 294161 137749 294279 137867
rect 294161 119909 294279 120027
rect 294161 119749 294279 119867
rect 294161 101909 294279 102027
rect 294161 101749 294279 101867
rect 294161 83909 294279 84027
rect 294161 83749 294279 83867
rect 294161 65909 294279 66027
rect 294161 65749 294279 65867
rect 294161 47909 294279 48027
rect 294161 47749 294279 47867
rect 294161 29909 294279 30027
rect 294161 29749 294279 29867
rect 294161 11909 294279 12027
rect 294161 11749 294279 11867
rect 294161 -1701 294279 -1583
rect 294161 -1861 294279 -1743
rect 294631 346709 294749 346827
rect 294631 346549 294749 346667
rect 294631 328709 294749 328827
rect 294631 328549 294749 328667
rect 294631 310709 294749 310827
rect 294631 310549 294749 310667
rect 294631 292709 294749 292827
rect 294631 292549 294749 292667
rect 294631 274709 294749 274827
rect 294631 274549 294749 274667
rect 294631 256709 294749 256827
rect 294631 256549 294749 256667
rect 294631 238709 294749 238827
rect 294631 238549 294749 238667
rect 294631 220709 294749 220827
rect 294631 220549 294749 220667
rect 294631 202709 294749 202827
rect 294631 202549 294749 202667
rect 294631 184709 294749 184827
rect 294631 184549 294749 184667
rect 294631 166709 294749 166827
rect 294631 166549 294749 166667
rect 294631 148709 294749 148827
rect 294631 148549 294749 148667
rect 294631 130709 294749 130827
rect 294631 130549 294749 130667
rect 294631 112709 294749 112827
rect 294631 112549 294749 112667
rect 294631 94709 294749 94827
rect 294631 94549 294749 94667
rect 294631 76709 294749 76827
rect 294631 76549 294749 76667
rect 294631 58709 294749 58827
rect 294631 58549 294749 58667
rect 294631 40709 294749 40827
rect 294631 40549 294749 40667
rect 294631 22709 294749 22827
rect 294631 22549 294749 22667
rect 294631 4709 294749 4827
rect 294631 4549 294749 4667
rect 294631 -2171 294749 -2053
rect 294631 -2331 294749 -2213
rect 295101 337709 295219 337827
rect 295101 337549 295219 337667
rect 295101 319709 295219 319827
rect 295101 319549 295219 319667
rect 295101 301709 295219 301827
rect 295101 301549 295219 301667
rect 295101 283709 295219 283827
rect 295101 283549 295219 283667
rect 295101 265709 295219 265827
rect 295101 265549 295219 265667
rect 295101 247709 295219 247827
rect 295101 247549 295219 247667
rect 295101 229709 295219 229827
rect 295101 229549 295219 229667
rect 295101 211709 295219 211827
rect 295101 211549 295219 211667
rect 295101 193709 295219 193827
rect 295101 193549 295219 193667
rect 295101 175709 295219 175827
rect 295101 175549 295219 175667
rect 295101 157709 295219 157827
rect 295101 157549 295219 157667
rect 295101 139709 295219 139827
rect 295101 139549 295219 139667
rect 295101 121709 295219 121827
rect 295101 121549 295219 121667
rect 295101 103709 295219 103827
rect 295101 103549 295219 103667
rect 295101 85709 295219 85827
rect 295101 85549 295219 85667
rect 295101 67709 295219 67827
rect 295101 67549 295219 67667
rect 295101 49709 295219 49827
rect 295101 49549 295219 49667
rect 295101 31709 295219 31827
rect 295101 31549 295219 31667
rect 295101 13709 295219 13827
rect 295101 13549 295219 13667
rect 295101 -2641 295219 -2523
rect 295101 -2801 295219 -2683
rect 295571 348509 295689 348627
rect 295571 348349 295689 348467
rect 295571 330509 295689 330627
rect 295571 330349 295689 330467
rect 295571 312509 295689 312627
rect 295571 312349 295689 312467
rect 295571 294509 295689 294627
rect 295571 294349 295689 294467
rect 295571 276509 295689 276627
rect 295571 276349 295689 276467
rect 295571 258509 295689 258627
rect 295571 258349 295689 258467
rect 295571 240509 295689 240627
rect 295571 240349 295689 240467
rect 295571 222509 295689 222627
rect 295571 222349 295689 222467
rect 295571 204509 295689 204627
rect 295571 204349 295689 204467
rect 295571 186509 295689 186627
rect 295571 186349 295689 186467
rect 295571 168509 295689 168627
rect 295571 168349 295689 168467
rect 295571 150509 295689 150627
rect 295571 150349 295689 150467
rect 295571 132509 295689 132627
rect 295571 132349 295689 132467
rect 295571 114509 295689 114627
rect 295571 114349 295689 114467
rect 295571 96509 295689 96627
rect 295571 96349 295689 96467
rect 295571 78509 295689 78627
rect 295571 78349 295689 78467
rect 295571 60509 295689 60627
rect 295571 60349 295689 60467
rect 295571 42509 295689 42627
rect 295571 42349 295689 42467
rect 295571 24509 295689 24627
rect 295571 24349 295689 24467
rect 295571 6509 295689 6627
rect 295571 6349 295689 6467
rect 295571 -3111 295689 -2993
rect 295571 -3271 295689 -3153
rect 296041 339509 296159 339627
rect 296041 339349 296159 339467
rect 296041 321509 296159 321627
rect 296041 321349 296159 321467
rect 296041 303509 296159 303627
rect 296041 303349 296159 303467
rect 296041 285509 296159 285627
rect 296041 285349 296159 285467
rect 296041 267509 296159 267627
rect 296041 267349 296159 267467
rect 296041 249509 296159 249627
rect 296041 249349 296159 249467
rect 296041 231509 296159 231627
rect 296041 231349 296159 231467
rect 296041 213509 296159 213627
rect 296041 213349 296159 213467
rect 296041 195509 296159 195627
rect 296041 195349 296159 195467
rect 296041 177509 296159 177627
rect 296041 177349 296159 177467
rect 296041 159509 296159 159627
rect 296041 159349 296159 159467
rect 296041 141509 296159 141627
rect 296041 141349 296159 141467
rect 296041 123509 296159 123627
rect 296041 123349 296159 123467
rect 296041 105509 296159 105627
rect 296041 105349 296159 105467
rect 296041 87509 296159 87627
rect 296041 87349 296159 87467
rect 296041 69509 296159 69627
rect 296041 69349 296159 69467
rect 296041 51509 296159 51627
rect 296041 51349 296159 51467
rect 296041 33509 296159 33627
rect 296041 33349 296159 33467
rect 296041 15509 296159 15627
rect 296041 15349 296159 15467
rect 284893 -3581 285011 -3463
rect 284893 -3741 285011 -3623
rect 296041 -3581 296159 -3463
rect 296041 -3741 296159 -3623
<< metal5 >>
rect -4288 355720 -3988 355721
rect 14802 355720 15102 355721
rect 32802 355720 33102 355721
rect 50802 355720 51102 355721
rect 68802 355720 69102 355721
rect 86802 355720 87102 355721
rect 104802 355720 105102 355721
rect 122802 355720 123102 355721
rect 140802 355720 141102 355721
rect 158802 355720 159102 355721
rect 176802 355720 177102 355721
rect 194802 355720 195102 355721
rect 212802 355720 213102 355721
rect 230802 355720 231102 355721
rect 248802 355720 249102 355721
rect 266802 355720 267102 355721
rect 284802 355720 285102 355721
rect 295950 355720 296250 355721
rect -4288 355709 296250 355720
rect -4288 355591 -4197 355709
rect -4079 355591 14893 355709
rect 15011 355591 32893 355709
rect 33011 355591 50893 355709
rect 51011 355591 68893 355709
rect 69011 355591 86893 355709
rect 87011 355591 104893 355709
rect 105011 355591 122893 355709
rect 123011 355591 140893 355709
rect 141011 355591 158893 355709
rect 159011 355591 176893 355709
rect 177011 355591 194893 355709
rect 195011 355591 212893 355709
rect 213011 355591 230893 355709
rect 231011 355591 248893 355709
rect 249011 355591 266893 355709
rect 267011 355591 284893 355709
rect 285011 355591 296041 355709
rect 296159 355591 296250 355709
rect -4288 355549 296250 355591
rect -4288 355431 -4197 355549
rect -4079 355431 14893 355549
rect 15011 355431 32893 355549
rect 33011 355431 50893 355549
rect 51011 355431 68893 355549
rect 69011 355431 86893 355549
rect 87011 355431 104893 355549
rect 105011 355431 122893 355549
rect 123011 355431 140893 355549
rect 141011 355431 158893 355549
rect 159011 355431 176893 355549
rect 177011 355431 194893 355549
rect 195011 355431 212893 355549
rect 213011 355431 230893 355549
rect 231011 355431 248893 355549
rect 249011 355431 266893 355549
rect 267011 355431 284893 355549
rect 285011 355431 296041 355549
rect 296159 355431 296250 355549
rect -4288 355420 296250 355431
rect -4288 355419 -3988 355420
rect 14802 355419 15102 355420
rect 32802 355419 33102 355420
rect 50802 355419 51102 355420
rect 68802 355419 69102 355420
rect 86802 355419 87102 355420
rect 104802 355419 105102 355420
rect 122802 355419 123102 355420
rect 140802 355419 141102 355420
rect 158802 355419 159102 355420
rect 176802 355419 177102 355420
rect 194802 355419 195102 355420
rect 212802 355419 213102 355420
rect 230802 355419 231102 355420
rect 248802 355419 249102 355420
rect 266802 355419 267102 355420
rect 284802 355419 285102 355420
rect 295950 355419 296250 355420
rect -3818 355250 -3518 355251
rect 5802 355250 6102 355251
rect 23802 355250 24102 355251
rect 41802 355250 42102 355251
rect 59802 355250 60102 355251
rect 77802 355250 78102 355251
rect 95802 355250 96102 355251
rect 113802 355250 114102 355251
rect 131802 355250 132102 355251
rect 149802 355250 150102 355251
rect 167802 355250 168102 355251
rect 185802 355250 186102 355251
rect 203802 355250 204102 355251
rect 221802 355250 222102 355251
rect 239802 355250 240102 355251
rect 257802 355250 258102 355251
rect 275802 355250 276102 355251
rect 295480 355250 295780 355251
rect -3818 355239 295780 355250
rect -3818 355121 -3727 355239
rect -3609 355121 5893 355239
rect 6011 355121 23893 355239
rect 24011 355121 41893 355239
rect 42011 355121 59893 355239
rect 60011 355121 77893 355239
rect 78011 355121 95893 355239
rect 96011 355121 113893 355239
rect 114011 355121 131893 355239
rect 132011 355121 149893 355239
rect 150011 355121 167893 355239
rect 168011 355121 185893 355239
rect 186011 355121 203893 355239
rect 204011 355121 221893 355239
rect 222011 355121 239893 355239
rect 240011 355121 257893 355239
rect 258011 355121 275893 355239
rect 276011 355121 295571 355239
rect 295689 355121 295780 355239
rect -3818 355079 295780 355121
rect -3818 354961 -3727 355079
rect -3609 354961 5893 355079
rect 6011 354961 23893 355079
rect 24011 354961 41893 355079
rect 42011 354961 59893 355079
rect 60011 354961 77893 355079
rect 78011 354961 95893 355079
rect 96011 354961 113893 355079
rect 114011 354961 131893 355079
rect 132011 354961 149893 355079
rect 150011 354961 167893 355079
rect 168011 354961 185893 355079
rect 186011 354961 203893 355079
rect 204011 354961 221893 355079
rect 222011 354961 239893 355079
rect 240011 354961 257893 355079
rect 258011 354961 275893 355079
rect 276011 354961 295571 355079
rect 295689 354961 295780 355079
rect -3818 354950 295780 354961
rect -3818 354949 -3518 354950
rect 5802 354949 6102 354950
rect 23802 354949 24102 354950
rect 41802 354949 42102 354950
rect 59802 354949 60102 354950
rect 77802 354949 78102 354950
rect 95802 354949 96102 354950
rect 113802 354949 114102 354950
rect 131802 354949 132102 354950
rect 149802 354949 150102 354950
rect 167802 354949 168102 354950
rect 185802 354949 186102 354950
rect 203802 354949 204102 354950
rect 221802 354949 222102 354950
rect 239802 354949 240102 354950
rect 257802 354949 258102 354950
rect 275802 354949 276102 354950
rect 295480 354949 295780 354950
rect -3348 354780 -3048 354781
rect 13002 354780 13302 354781
rect 31002 354780 31302 354781
rect 49002 354780 49302 354781
rect 67002 354780 67302 354781
rect 85002 354780 85302 354781
rect 103002 354780 103302 354781
rect 121002 354780 121302 354781
rect 139002 354780 139302 354781
rect 157002 354780 157302 354781
rect 175002 354780 175302 354781
rect 193002 354780 193302 354781
rect 211002 354780 211302 354781
rect 229002 354780 229302 354781
rect 247002 354780 247302 354781
rect 265002 354780 265302 354781
rect 283002 354780 283302 354781
rect 295010 354780 295310 354781
rect -3348 354769 295310 354780
rect -3348 354651 -3257 354769
rect -3139 354651 13093 354769
rect 13211 354651 31093 354769
rect 31211 354651 49093 354769
rect 49211 354651 67093 354769
rect 67211 354651 85093 354769
rect 85211 354651 103093 354769
rect 103211 354651 121093 354769
rect 121211 354651 139093 354769
rect 139211 354651 157093 354769
rect 157211 354651 175093 354769
rect 175211 354651 193093 354769
rect 193211 354651 211093 354769
rect 211211 354651 229093 354769
rect 229211 354651 247093 354769
rect 247211 354651 265093 354769
rect 265211 354651 283093 354769
rect 283211 354651 295101 354769
rect 295219 354651 295310 354769
rect -3348 354609 295310 354651
rect -3348 354491 -3257 354609
rect -3139 354491 13093 354609
rect 13211 354491 31093 354609
rect 31211 354491 49093 354609
rect 49211 354491 67093 354609
rect 67211 354491 85093 354609
rect 85211 354491 103093 354609
rect 103211 354491 121093 354609
rect 121211 354491 139093 354609
rect 139211 354491 157093 354609
rect 157211 354491 175093 354609
rect 175211 354491 193093 354609
rect 193211 354491 211093 354609
rect 211211 354491 229093 354609
rect 229211 354491 247093 354609
rect 247211 354491 265093 354609
rect 265211 354491 283093 354609
rect 283211 354491 295101 354609
rect 295219 354491 295310 354609
rect -3348 354480 295310 354491
rect -3348 354479 -3048 354480
rect 13002 354479 13302 354480
rect 31002 354479 31302 354480
rect 49002 354479 49302 354480
rect 67002 354479 67302 354480
rect 85002 354479 85302 354480
rect 103002 354479 103302 354480
rect 121002 354479 121302 354480
rect 139002 354479 139302 354480
rect 157002 354479 157302 354480
rect 175002 354479 175302 354480
rect 193002 354479 193302 354480
rect 211002 354479 211302 354480
rect 229002 354479 229302 354480
rect 247002 354479 247302 354480
rect 265002 354479 265302 354480
rect 283002 354479 283302 354480
rect 295010 354479 295310 354480
rect -2878 354310 -2578 354311
rect 4002 354310 4302 354311
rect 22002 354310 22302 354311
rect 40002 354310 40302 354311
rect 58002 354310 58302 354311
rect 76002 354310 76302 354311
rect 94002 354310 94302 354311
rect 112002 354310 112302 354311
rect 130002 354310 130302 354311
rect 148002 354310 148302 354311
rect 166002 354310 166302 354311
rect 184002 354310 184302 354311
rect 202002 354310 202302 354311
rect 220002 354310 220302 354311
rect 238002 354310 238302 354311
rect 256002 354310 256302 354311
rect 274002 354310 274302 354311
rect 294540 354310 294840 354311
rect -2878 354299 294840 354310
rect -2878 354181 -2787 354299
rect -2669 354181 4093 354299
rect 4211 354181 22093 354299
rect 22211 354181 40093 354299
rect 40211 354181 58093 354299
rect 58211 354181 76093 354299
rect 76211 354181 94093 354299
rect 94211 354181 112093 354299
rect 112211 354181 130093 354299
rect 130211 354181 148093 354299
rect 148211 354181 166093 354299
rect 166211 354181 184093 354299
rect 184211 354181 202093 354299
rect 202211 354181 220093 354299
rect 220211 354181 238093 354299
rect 238211 354181 256093 354299
rect 256211 354181 274093 354299
rect 274211 354181 294631 354299
rect 294749 354181 294840 354299
rect -2878 354139 294840 354181
rect -2878 354021 -2787 354139
rect -2669 354021 4093 354139
rect 4211 354021 22093 354139
rect 22211 354021 40093 354139
rect 40211 354021 58093 354139
rect 58211 354021 76093 354139
rect 76211 354021 94093 354139
rect 94211 354021 112093 354139
rect 112211 354021 130093 354139
rect 130211 354021 148093 354139
rect 148211 354021 166093 354139
rect 166211 354021 184093 354139
rect 184211 354021 202093 354139
rect 202211 354021 220093 354139
rect 220211 354021 238093 354139
rect 238211 354021 256093 354139
rect 256211 354021 274093 354139
rect 274211 354021 294631 354139
rect 294749 354021 294840 354139
rect -2878 354010 294840 354021
rect -2878 354009 -2578 354010
rect 4002 354009 4302 354010
rect 22002 354009 22302 354010
rect 40002 354009 40302 354010
rect 58002 354009 58302 354010
rect 76002 354009 76302 354010
rect 94002 354009 94302 354010
rect 112002 354009 112302 354010
rect 130002 354009 130302 354010
rect 148002 354009 148302 354010
rect 166002 354009 166302 354010
rect 184002 354009 184302 354010
rect 202002 354009 202302 354010
rect 220002 354009 220302 354010
rect 238002 354009 238302 354010
rect 256002 354009 256302 354010
rect 274002 354009 274302 354010
rect 294540 354009 294840 354010
rect -2408 353840 -2108 353841
rect 11202 353840 11502 353841
rect 29202 353840 29502 353841
rect 47202 353840 47502 353841
rect 65202 353840 65502 353841
rect 83202 353840 83502 353841
rect 101202 353840 101502 353841
rect 119202 353840 119502 353841
rect 137202 353840 137502 353841
rect 155202 353840 155502 353841
rect 173202 353840 173502 353841
rect 191202 353840 191502 353841
rect 209202 353840 209502 353841
rect 227202 353840 227502 353841
rect 245202 353840 245502 353841
rect 263202 353840 263502 353841
rect 281202 353840 281502 353841
rect 294070 353840 294370 353841
rect -2408 353829 294370 353840
rect -2408 353711 -2317 353829
rect -2199 353711 11293 353829
rect 11411 353711 29293 353829
rect 29411 353711 47293 353829
rect 47411 353711 65293 353829
rect 65411 353711 83293 353829
rect 83411 353711 101293 353829
rect 101411 353711 119293 353829
rect 119411 353711 137293 353829
rect 137411 353711 155293 353829
rect 155411 353711 173293 353829
rect 173411 353711 191293 353829
rect 191411 353711 209293 353829
rect 209411 353711 227293 353829
rect 227411 353711 245293 353829
rect 245411 353711 263293 353829
rect 263411 353711 281293 353829
rect 281411 353711 294161 353829
rect 294279 353711 294370 353829
rect -2408 353669 294370 353711
rect -2408 353551 -2317 353669
rect -2199 353551 11293 353669
rect 11411 353551 29293 353669
rect 29411 353551 47293 353669
rect 47411 353551 65293 353669
rect 65411 353551 83293 353669
rect 83411 353551 101293 353669
rect 101411 353551 119293 353669
rect 119411 353551 137293 353669
rect 137411 353551 155293 353669
rect 155411 353551 173293 353669
rect 173411 353551 191293 353669
rect 191411 353551 209293 353669
rect 209411 353551 227293 353669
rect 227411 353551 245293 353669
rect 245411 353551 263293 353669
rect 263411 353551 281293 353669
rect 281411 353551 294161 353669
rect 294279 353551 294370 353669
rect -2408 353540 294370 353551
rect -2408 353539 -2108 353540
rect 11202 353539 11502 353540
rect 29202 353539 29502 353540
rect 47202 353539 47502 353540
rect 65202 353539 65502 353540
rect 83202 353539 83502 353540
rect 101202 353539 101502 353540
rect 119202 353539 119502 353540
rect 137202 353539 137502 353540
rect 155202 353539 155502 353540
rect 173202 353539 173502 353540
rect 191202 353539 191502 353540
rect 209202 353539 209502 353540
rect 227202 353539 227502 353540
rect 245202 353539 245502 353540
rect 263202 353539 263502 353540
rect 281202 353539 281502 353540
rect 294070 353539 294370 353540
rect -1938 353370 -1638 353371
rect 2202 353370 2502 353371
rect 20202 353370 20502 353371
rect 38202 353370 38502 353371
rect 56202 353370 56502 353371
rect 74202 353370 74502 353371
rect 92202 353370 92502 353371
rect 110202 353370 110502 353371
rect 128202 353370 128502 353371
rect 146202 353370 146502 353371
rect 164202 353370 164502 353371
rect 182202 353370 182502 353371
rect 200202 353370 200502 353371
rect 218202 353370 218502 353371
rect 236202 353370 236502 353371
rect 254202 353370 254502 353371
rect 272202 353370 272502 353371
rect 290202 353370 290502 353371
rect 293600 353370 293900 353371
rect -1938 353359 293900 353370
rect -1938 353241 -1847 353359
rect -1729 353241 2293 353359
rect 2411 353241 20293 353359
rect 20411 353241 38293 353359
rect 38411 353241 56293 353359
rect 56411 353241 74293 353359
rect 74411 353241 92293 353359
rect 92411 353241 110293 353359
rect 110411 353241 128293 353359
rect 128411 353241 146293 353359
rect 146411 353241 164293 353359
rect 164411 353241 182293 353359
rect 182411 353241 200293 353359
rect 200411 353241 218293 353359
rect 218411 353241 236293 353359
rect 236411 353241 254293 353359
rect 254411 353241 272293 353359
rect 272411 353241 290293 353359
rect 290411 353241 293691 353359
rect 293809 353241 293900 353359
rect -1938 353199 293900 353241
rect -1938 353081 -1847 353199
rect -1729 353081 2293 353199
rect 2411 353081 20293 353199
rect 20411 353081 38293 353199
rect 38411 353081 56293 353199
rect 56411 353081 74293 353199
rect 74411 353081 92293 353199
rect 92411 353081 110293 353199
rect 110411 353081 128293 353199
rect 128411 353081 146293 353199
rect 146411 353081 164293 353199
rect 164411 353081 182293 353199
rect 182411 353081 200293 353199
rect 200411 353081 218293 353199
rect 218411 353081 236293 353199
rect 236411 353081 254293 353199
rect 254411 353081 272293 353199
rect 272411 353081 290293 353199
rect 290411 353081 293691 353199
rect 293809 353081 293900 353199
rect -1938 353070 293900 353081
rect -1938 353069 -1638 353070
rect 2202 353069 2502 353070
rect 20202 353069 20502 353070
rect 38202 353069 38502 353070
rect 56202 353069 56502 353070
rect 74202 353069 74502 353070
rect 92202 353069 92502 353070
rect 110202 353069 110502 353070
rect 128202 353069 128502 353070
rect 146202 353069 146502 353070
rect 164202 353069 164502 353070
rect 182202 353069 182502 353070
rect 200202 353069 200502 353070
rect 218202 353069 218502 353070
rect 236202 353069 236502 353070
rect 254202 353069 254502 353070
rect 272202 353069 272502 353070
rect 290202 353069 290502 353070
rect 293600 353069 293900 353070
rect -1468 352900 -1168 352901
rect 9402 352900 9702 352901
rect 27402 352900 27702 352901
rect 45402 352900 45702 352901
rect 63402 352900 63702 352901
rect 81402 352900 81702 352901
rect 99402 352900 99702 352901
rect 117402 352900 117702 352901
rect 135402 352900 135702 352901
rect 153402 352900 153702 352901
rect 171402 352900 171702 352901
rect 189402 352900 189702 352901
rect 207402 352900 207702 352901
rect 225402 352900 225702 352901
rect 243402 352900 243702 352901
rect 261402 352900 261702 352901
rect 279402 352900 279702 352901
rect 293130 352900 293430 352901
rect -1468 352889 293430 352900
rect -1468 352771 -1377 352889
rect -1259 352771 9493 352889
rect 9611 352771 27493 352889
rect 27611 352771 45493 352889
rect 45611 352771 63493 352889
rect 63611 352771 81493 352889
rect 81611 352771 99493 352889
rect 99611 352771 117493 352889
rect 117611 352771 135493 352889
rect 135611 352771 153493 352889
rect 153611 352771 171493 352889
rect 171611 352771 189493 352889
rect 189611 352771 207493 352889
rect 207611 352771 225493 352889
rect 225611 352771 243493 352889
rect 243611 352771 261493 352889
rect 261611 352771 279493 352889
rect 279611 352771 293221 352889
rect 293339 352771 293430 352889
rect -1468 352729 293430 352771
rect -1468 352611 -1377 352729
rect -1259 352611 9493 352729
rect 9611 352611 27493 352729
rect 27611 352611 45493 352729
rect 45611 352611 63493 352729
rect 63611 352611 81493 352729
rect 81611 352611 99493 352729
rect 99611 352611 117493 352729
rect 117611 352611 135493 352729
rect 135611 352611 153493 352729
rect 153611 352611 171493 352729
rect 171611 352611 189493 352729
rect 189611 352611 207493 352729
rect 207611 352611 225493 352729
rect 225611 352611 243493 352729
rect 243611 352611 261493 352729
rect 261611 352611 279493 352729
rect 279611 352611 293221 352729
rect 293339 352611 293430 352729
rect -1468 352600 293430 352611
rect -1468 352599 -1168 352600
rect 9402 352599 9702 352600
rect 27402 352599 27702 352600
rect 45402 352599 45702 352600
rect 63402 352599 63702 352600
rect 81402 352599 81702 352600
rect 99402 352599 99702 352600
rect 117402 352599 117702 352600
rect 135402 352599 135702 352600
rect 153402 352599 153702 352600
rect 171402 352599 171702 352600
rect 189402 352599 189702 352600
rect 207402 352599 207702 352600
rect 225402 352599 225702 352600
rect 243402 352599 243702 352600
rect 261402 352599 261702 352600
rect 279402 352599 279702 352600
rect 293130 352599 293430 352600
rect -998 352430 -698 352431
rect 402 352430 702 352431
rect 18402 352430 18702 352431
rect 36402 352430 36702 352431
rect 54402 352430 54702 352431
rect 72402 352430 72702 352431
rect 90402 352430 90702 352431
rect 108402 352430 108702 352431
rect 126402 352430 126702 352431
rect 144402 352430 144702 352431
rect 162402 352430 162702 352431
rect 180402 352430 180702 352431
rect 198402 352430 198702 352431
rect 216402 352430 216702 352431
rect 234402 352430 234702 352431
rect 252402 352430 252702 352431
rect 270402 352430 270702 352431
rect 288402 352430 288702 352431
rect 292660 352430 292960 352431
rect -998 352419 292960 352430
rect -998 352301 -907 352419
rect -789 352301 493 352419
rect 611 352301 18493 352419
rect 18611 352301 36493 352419
rect 36611 352301 54493 352419
rect 54611 352301 72493 352419
rect 72611 352301 90493 352419
rect 90611 352301 108493 352419
rect 108611 352301 126493 352419
rect 126611 352301 144493 352419
rect 144611 352301 162493 352419
rect 162611 352301 180493 352419
rect 180611 352301 198493 352419
rect 198611 352301 216493 352419
rect 216611 352301 234493 352419
rect 234611 352301 252493 352419
rect 252611 352301 270493 352419
rect 270611 352301 288493 352419
rect 288611 352301 292751 352419
rect 292869 352301 292960 352419
rect -998 352259 292960 352301
rect -998 352141 -907 352259
rect -789 352141 493 352259
rect 611 352141 18493 352259
rect 18611 352141 36493 352259
rect 36611 352141 54493 352259
rect 54611 352141 72493 352259
rect 72611 352141 90493 352259
rect 90611 352141 108493 352259
rect 108611 352141 126493 352259
rect 126611 352141 144493 352259
rect 144611 352141 162493 352259
rect 162611 352141 180493 352259
rect 180611 352141 198493 352259
rect 198611 352141 216493 352259
rect 216611 352141 234493 352259
rect 234611 352141 252493 352259
rect 252611 352141 270493 352259
rect 270611 352141 288493 352259
rect 288611 352141 292751 352259
rect 292869 352141 292960 352259
rect -998 352130 292960 352141
rect -998 352129 -698 352130
rect 402 352129 702 352130
rect 18402 352129 18702 352130
rect 36402 352129 36702 352130
rect 54402 352129 54702 352130
rect 72402 352129 72702 352130
rect 90402 352129 90702 352130
rect 108402 352129 108702 352130
rect 126402 352129 126702 352130
rect 144402 352129 144702 352130
rect 162402 352129 162702 352130
rect 180402 352129 180702 352130
rect 198402 352129 198702 352130
rect 216402 352129 216702 352130
rect 234402 352129 234702 352130
rect 252402 352129 252702 352130
rect 270402 352129 270702 352130
rect 288402 352129 288702 352130
rect 292660 352129 292960 352130
rect -3818 348638 -3518 348639
rect 295480 348638 295780 348639
rect -4288 348627 240 348638
rect -4288 348509 -3727 348627
rect -3609 348509 240 348627
rect -4288 348467 240 348509
rect -4288 348349 -3727 348467
rect -3609 348349 240 348467
rect -4288 348338 240 348349
rect 291760 348627 296250 348638
rect 291760 348509 295571 348627
rect 295689 348509 296250 348627
rect 291760 348467 296250 348509
rect 291760 348349 295571 348467
rect 295689 348349 296250 348467
rect 291760 348338 296250 348349
rect -3818 348337 -3518 348338
rect 295480 348337 295780 348338
rect -2878 346838 -2578 346839
rect 294540 346838 294840 346839
rect -3348 346827 240 346838
rect -3348 346709 -2787 346827
rect -2669 346709 240 346827
rect -3348 346667 240 346709
rect -3348 346549 -2787 346667
rect -2669 346549 240 346667
rect -3348 346538 240 346549
rect 291760 346827 295310 346838
rect 291760 346709 294631 346827
rect 294749 346709 295310 346827
rect 291760 346667 295310 346709
rect 291760 346549 294631 346667
rect 294749 346549 295310 346667
rect 291760 346538 295310 346549
rect -2878 346537 -2578 346538
rect 294540 346537 294840 346538
rect -1938 345038 -1638 345039
rect 293600 345038 293900 345039
rect -2408 345027 240 345038
rect -2408 344909 -1847 345027
rect -1729 344909 240 345027
rect -2408 344867 240 344909
rect -2408 344749 -1847 344867
rect -1729 344749 240 344867
rect -2408 344738 240 344749
rect 291760 345027 294370 345038
rect 291760 344909 293691 345027
rect 293809 344909 294370 345027
rect 291760 344867 294370 344909
rect 291760 344749 293691 344867
rect 293809 344749 294370 344867
rect 291760 344738 294370 344749
rect -1938 344737 -1638 344738
rect 293600 344737 293900 344738
rect -998 343238 -698 343239
rect 292660 343238 292960 343239
rect -1468 343227 240 343238
rect -1468 343109 -907 343227
rect -789 343109 240 343227
rect -1468 343067 240 343109
rect -1468 342949 -907 343067
rect -789 342949 240 343067
rect -1468 342938 240 342949
rect 291760 343227 293430 343238
rect 291760 343109 292751 343227
rect 292869 343109 293430 343227
rect 291760 343067 293430 343109
rect 291760 342949 292751 343067
rect 292869 342949 293430 343067
rect 291760 342938 293430 342949
rect -998 342937 -698 342938
rect 292660 342937 292960 342938
rect -4288 339638 -3988 339639
rect 295950 339638 296250 339639
rect -4288 339627 240 339638
rect -4288 339509 -4197 339627
rect -4079 339509 240 339627
rect -4288 339467 240 339509
rect -4288 339349 -4197 339467
rect -4079 339349 240 339467
rect -4288 339338 240 339349
rect 291760 339627 296250 339638
rect 291760 339509 296041 339627
rect 296159 339509 296250 339627
rect 291760 339467 296250 339509
rect 291760 339349 296041 339467
rect 296159 339349 296250 339467
rect 291760 339338 296250 339349
rect -4288 339337 -3988 339338
rect 295950 339337 296250 339338
rect -3348 337838 -3048 337839
rect 295010 337838 295310 337839
rect -3348 337827 240 337838
rect -3348 337709 -3257 337827
rect -3139 337709 240 337827
rect -3348 337667 240 337709
rect -3348 337549 -3257 337667
rect -3139 337549 240 337667
rect -3348 337538 240 337549
rect 291760 337827 295310 337838
rect 291760 337709 295101 337827
rect 295219 337709 295310 337827
rect 291760 337667 295310 337709
rect 291760 337549 295101 337667
rect 295219 337549 295310 337667
rect 291760 337538 295310 337549
rect -3348 337537 -3048 337538
rect 295010 337537 295310 337538
rect -2408 336038 -2108 336039
rect 294070 336038 294370 336039
rect -2408 336027 240 336038
rect -2408 335909 -2317 336027
rect -2199 335909 240 336027
rect -2408 335867 240 335909
rect -2408 335749 -2317 335867
rect -2199 335749 240 335867
rect -2408 335738 240 335749
rect 291760 336027 294370 336038
rect 291760 335909 294161 336027
rect 294279 335909 294370 336027
rect 291760 335867 294370 335909
rect 291760 335749 294161 335867
rect 294279 335749 294370 335867
rect 291760 335738 294370 335749
rect -2408 335737 -2108 335738
rect 294070 335737 294370 335738
rect -1468 334238 -1168 334239
rect 293130 334238 293430 334239
rect -1468 334227 240 334238
rect -1468 334109 -1377 334227
rect -1259 334109 240 334227
rect -1468 334067 240 334109
rect -1468 333949 -1377 334067
rect -1259 333949 240 334067
rect -1468 333938 240 333949
rect 291760 334227 293430 334238
rect 291760 334109 293221 334227
rect 293339 334109 293430 334227
rect 291760 334067 293430 334109
rect 291760 333949 293221 334067
rect 293339 333949 293430 334067
rect 291760 333938 293430 333949
rect -1468 333937 -1168 333938
rect 293130 333937 293430 333938
rect -3818 330638 -3518 330639
rect 295480 330638 295780 330639
rect -4288 330627 240 330638
rect -4288 330509 -3727 330627
rect -3609 330509 240 330627
rect -4288 330467 240 330509
rect -4288 330349 -3727 330467
rect -3609 330349 240 330467
rect -4288 330338 240 330349
rect 291760 330627 296250 330638
rect 291760 330509 295571 330627
rect 295689 330509 296250 330627
rect 291760 330467 296250 330509
rect 291760 330349 295571 330467
rect 295689 330349 296250 330467
rect 291760 330338 296250 330349
rect -3818 330337 -3518 330338
rect 295480 330337 295780 330338
rect -2878 328838 -2578 328839
rect 294540 328838 294840 328839
rect -3348 328827 240 328838
rect -3348 328709 -2787 328827
rect -2669 328709 240 328827
rect -3348 328667 240 328709
rect -3348 328549 -2787 328667
rect -2669 328549 240 328667
rect -3348 328538 240 328549
rect 291760 328827 295310 328838
rect 291760 328709 294631 328827
rect 294749 328709 295310 328827
rect 291760 328667 295310 328709
rect 291760 328549 294631 328667
rect 294749 328549 295310 328667
rect 291760 328538 295310 328549
rect -2878 328537 -2578 328538
rect 294540 328537 294840 328538
rect -1938 327038 -1638 327039
rect 293600 327038 293900 327039
rect -2408 327027 240 327038
rect -2408 326909 -1847 327027
rect -1729 326909 240 327027
rect -2408 326867 240 326909
rect -2408 326749 -1847 326867
rect -1729 326749 240 326867
rect -2408 326738 240 326749
rect 291760 327027 294370 327038
rect 291760 326909 293691 327027
rect 293809 326909 294370 327027
rect 291760 326867 294370 326909
rect 291760 326749 293691 326867
rect 293809 326749 294370 326867
rect 291760 326738 294370 326749
rect -1938 326737 -1638 326738
rect 293600 326737 293900 326738
rect -998 325238 -698 325239
rect 292660 325238 292960 325239
rect -1468 325227 240 325238
rect -1468 325109 -907 325227
rect -789 325109 240 325227
rect -1468 325067 240 325109
rect -1468 324949 -907 325067
rect -789 324949 240 325067
rect -1468 324938 240 324949
rect 291760 325227 293430 325238
rect 291760 325109 292751 325227
rect 292869 325109 293430 325227
rect 291760 325067 293430 325109
rect 291760 324949 292751 325067
rect 292869 324949 293430 325067
rect 291760 324938 293430 324949
rect -998 324937 -698 324938
rect 292660 324937 292960 324938
rect -4288 321638 -3988 321639
rect 295950 321638 296250 321639
rect -4288 321627 240 321638
rect -4288 321509 -4197 321627
rect -4079 321509 240 321627
rect -4288 321467 240 321509
rect -4288 321349 -4197 321467
rect -4079 321349 240 321467
rect -4288 321338 240 321349
rect 291760 321627 296250 321638
rect 291760 321509 296041 321627
rect 296159 321509 296250 321627
rect 291760 321467 296250 321509
rect 291760 321349 296041 321467
rect 296159 321349 296250 321467
rect 291760 321338 296250 321349
rect -4288 321337 -3988 321338
rect 295950 321337 296250 321338
rect -3348 319838 -3048 319839
rect 295010 319838 295310 319839
rect -3348 319827 240 319838
rect -3348 319709 -3257 319827
rect -3139 319709 240 319827
rect -3348 319667 240 319709
rect -3348 319549 -3257 319667
rect -3139 319549 240 319667
rect -3348 319538 240 319549
rect 291760 319827 295310 319838
rect 291760 319709 295101 319827
rect 295219 319709 295310 319827
rect 291760 319667 295310 319709
rect 291760 319549 295101 319667
rect 295219 319549 295310 319667
rect 291760 319538 295310 319549
rect -3348 319537 -3048 319538
rect 295010 319537 295310 319538
rect -2408 318038 -2108 318039
rect 294070 318038 294370 318039
rect -2408 318027 240 318038
rect -2408 317909 -2317 318027
rect -2199 317909 240 318027
rect -2408 317867 240 317909
rect -2408 317749 -2317 317867
rect -2199 317749 240 317867
rect -2408 317738 240 317749
rect 291760 318027 294370 318038
rect 291760 317909 294161 318027
rect 294279 317909 294370 318027
rect 291760 317867 294370 317909
rect 291760 317749 294161 317867
rect 294279 317749 294370 317867
rect 291760 317738 294370 317749
rect -2408 317737 -2108 317738
rect 294070 317737 294370 317738
rect -1468 316238 -1168 316239
rect 293130 316238 293430 316239
rect -1468 316227 240 316238
rect -1468 316109 -1377 316227
rect -1259 316109 240 316227
rect -1468 316067 240 316109
rect -1468 315949 -1377 316067
rect -1259 315949 240 316067
rect -1468 315938 240 315949
rect 291760 316227 293430 316238
rect 291760 316109 293221 316227
rect 293339 316109 293430 316227
rect 291760 316067 293430 316109
rect 291760 315949 293221 316067
rect 293339 315949 293430 316067
rect 291760 315938 293430 315949
rect -1468 315937 -1168 315938
rect 293130 315937 293430 315938
rect -3818 312638 -3518 312639
rect 295480 312638 295780 312639
rect -4288 312627 240 312638
rect -4288 312509 -3727 312627
rect -3609 312509 240 312627
rect -4288 312467 240 312509
rect -4288 312349 -3727 312467
rect -3609 312349 240 312467
rect -4288 312338 240 312349
rect 291760 312627 296250 312638
rect 291760 312509 295571 312627
rect 295689 312509 296250 312627
rect 291760 312467 296250 312509
rect 291760 312349 295571 312467
rect 295689 312349 296250 312467
rect 291760 312338 296250 312349
rect -3818 312337 -3518 312338
rect 295480 312337 295780 312338
rect -2878 310838 -2578 310839
rect 294540 310838 294840 310839
rect -3348 310827 240 310838
rect -3348 310709 -2787 310827
rect -2669 310709 240 310827
rect -3348 310667 240 310709
rect -3348 310549 -2787 310667
rect -2669 310549 240 310667
rect -3348 310538 240 310549
rect 291760 310827 295310 310838
rect 291760 310709 294631 310827
rect 294749 310709 295310 310827
rect 291760 310667 295310 310709
rect 291760 310549 294631 310667
rect 294749 310549 295310 310667
rect 291760 310538 295310 310549
rect -2878 310537 -2578 310538
rect 294540 310537 294840 310538
rect -1938 309038 -1638 309039
rect 293600 309038 293900 309039
rect -2408 309027 240 309038
rect -2408 308909 -1847 309027
rect -1729 308909 240 309027
rect -2408 308867 240 308909
rect -2408 308749 -1847 308867
rect -1729 308749 240 308867
rect -2408 308738 240 308749
rect 291760 309027 294370 309038
rect 291760 308909 293691 309027
rect 293809 308909 294370 309027
rect 291760 308867 294370 308909
rect 291760 308749 293691 308867
rect 293809 308749 294370 308867
rect 291760 308738 294370 308749
rect -1938 308737 -1638 308738
rect 293600 308737 293900 308738
rect -998 307238 -698 307239
rect 292660 307238 292960 307239
rect -1468 307227 240 307238
rect -1468 307109 -907 307227
rect -789 307109 240 307227
rect -1468 307067 240 307109
rect -1468 306949 -907 307067
rect -789 306949 240 307067
rect -1468 306938 240 306949
rect 291760 307227 293430 307238
rect 291760 307109 292751 307227
rect 292869 307109 293430 307227
rect 291760 307067 293430 307109
rect 291760 306949 292751 307067
rect 292869 306949 293430 307067
rect 291760 306938 293430 306949
rect -998 306937 -698 306938
rect 292660 306937 292960 306938
rect -4288 303638 -3988 303639
rect 295950 303638 296250 303639
rect -4288 303627 240 303638
rect -4288 303509 -4197 303627
rect -4079 303509 240 303627
rect -4288 303467 240 303509
rect -4288 303349 -4197 303467
rect -4079 303349 240 303467
rect -4288 303338 240 303349
rect 291760 303627 296250 303638
rect 291760 303509 296041 303627
rect 296159 303509 296250 303627
rect 291760 303467 296250 303509
rect 291760 303349 296041 303467
rect 296159 303349 296250 303467
rect 291760 303338 296250 303349
rect -4288 303337 -3988 303338
rect 295950 303337 296250 303338
rect -3348 301838 -3048 301839
rect 295010 301838 295310 301839
rect -3348 301827 240 301838
rect -3348 301709 -3257 301827
rect -3139 301709 240 301827
rect -3348 301667 240 301709
rect -3348 301549 -3257 301667
rect -3139 301549 240 301667
rect -3348 301538 240 301549
rect 291760 301827 295310 301838
rect 291760 301709 295101 301827
rect 295219 301709 295310 301827
rect 291760 301667 295310 301709
rect 291760 301549 295101 301667
rect 295219 301549 295310 301667
rect 291760 301538 295310 301549
rect -3348 301537 -3048 301538
rect 295010 301537 295310 301538
rect -2408 300038 -2108 300039
rect 294070 300038 294370 300039
rect -2408 300027 240 300038
rect -2408 299909 -2317 300027
rect -2199 299909 240 300027
rect -2408 299867 240 299909
rect -2408 299749 -2317 299867
rect -2199 299749 240 299867
rect -2408 299738 240 299749
rect 291760 300027 294370 300038
rect 291760 299909 294161 300027
rect 294279 299909 294370 300027
rect 291760 299867 294370 299909
rect 291760 299749 294161 299867
rect 294279 299749 294370 299867
rect 291760 299738 294370 299749
rect -2408 299737 -2108 299738
rect 294070 299737 294370 299738
rect -1468 298238 -1168 298239
rect 293130 298238 293430 298239
rect -1468 298227 240 298238
rect -1468 298109 -1377 298227
rect -1259 298109 240 298227
rect -1468 298067 240 298109
rect -1468 297949 -1377 298067
rect -1259 297949 240 298067
rect -1468 297938 240 297949
rect 291760 298227 293430 298238
rect 291760 298109 293221 298227
rect 293339 298109 293430 298227
rect 291760 298067 293430 298109
rect 291760 297949 293221 298067
rect 293339 297949 293430 298067
rect 291760 297938 293430 297949
rect -1468 297937 -1168 297938
rect 293130 297937 293430 297938
rect -3818 294638 -3518 294639
rect 295480 294638 295780 294639
rect -4288 294627 240 294638
rect -4288 294509 -3727 294627
rect -3609 294509 240 294627
rect -4288 294467 240 294509
rect -4288 294349 -3727 294467
rect -3609 294349 240 294467
rect -4288 294338 240 294349
rect 291760 294627 296250 294638
rect 291760 294509 295571 294627
rect 295689 294509 296250 294627
rect 291760 294467 296250 294509
rect 291760 294349 295571 294467
rect 295689 294349 296250 294467
rect 291760 294338 296250 294349
rect -3818 294337 -3518 294338
rect 295480 294337 295780 294338
rect -2878 292838 -2578 292839
rect 294540 292838 294840 292839
rect -3348 292827 240 292838
rect -3348 292709 -2787 292827
rect -2669 292709 240 292827
rect -3348 292667 240 292709
rect -3348 292549 -2787 292667
rect -2669 292549 240 292667
rect -3348 292538 240 292549
rect 291760 292827 295310 292838
rect 291760 292709 294631 292827
rect 294749 292709 295310 292827
rect 291760 292667 295310 292709
rect 291760 292549 294631 292667
rect 294749 292549 295310 292667
rect 291760 292538 295310 292549
rect -2878 292537 -2578 292538
rect 294540 292537 294840 292538
rect -1938 291038 -1638 291039
rect 293600 291038 293900 291039
rect -2408 291027 240 291038
rect -2408 290909 -1847 291027
rect -1729 290909 240 291027
rect -2408 290867 240 290909
rect -2408 290749 -1847 290867
rect -1729 290749 240 290867
rect -2408 290738 240 290749
rect 291760 291027 294370 291038
rect 291760 290909 293691 291027
rect 293809 290909 294370 291027
rect 291760 290867 294370 290909
rect 291760 290749 293691 290867
rect 293809 290749 294370 290867
rect 291760 290738 294370 290749
rect -1938 290737 -1638 290738
rect 293600 290737 293900 290738
rect -998 289238 -698 289239
rect 292660 289238 292960 289239
rect -1468 289227 240 289238
rect -1468 289109 -907 289227
rect -789 289109 240 289227
rect -1468 289067 240 289109
rect -1468 288949 -907 289067
rect -789 288949 240 289067
rect -1468 288938 240 288949
rect 291760 289227 293430 289238
rect 291760 289109 292751 289227
rect 292869 289109 293430 289227
rect 291760 289067 293430 289109
rect 291760 288949 292751 289067
rect 292869 288949 293430 289067
rect 291760 288938 293430 288949
rect -998 288937 -698 288938
rect 292660 288937 292960 288938
rect -4288 285638 -3988 285639
rect 295950 285638 296250 285639
rect -4288 285627 240 285638
rect -4288 285509 -4197 285627
rect -4079 285509 240 285627
rect -4288 285467 240 285509
rect -4288 285349 -4197 285467
rect -4079 285349 240 285467
rect -4288 285338 240 285349
rect 291760 285627 296250 285638
rect 291760 285509 296041 285627
rect 296159 285509 296250 285627
rect 291760 285467 296250 285509
rect 291760 285349 296041 285467
rect 296159 285349 296250 285467
rect 291760 285338 296250 285349
rect -4288 285337 -3988 285338
rect 295950 285337 296250 285338
rect -3348 283838 -3048 283839
rect 295010 283838 295310 283839
rect -3348 283827 240 283838
rect -3348 283709 -3257 283827
rect -3139 283709 240 283827
rect -3348 283667 240 283709
rect -3348 283549 -3257 283667
rect -3139 283549 240 283667
rect -3348 283538 240 283549
rect 291760 283827 295310 283838
rect 291760 283709 295101 283827
rect 295219 283709 295310 283827
rect 291760 283667 295310 283709
rect 291760 283549 295101 283667
rect 295219 283549 295310 283667
rect 291760 283538 295310 283549
rect -3348 283537 -3048 283538
rect 295010 283537 295310 283538
rect -2408 282038 -2108 282039
rect 294070 282038 294370 282039
rect -2408 282027 240 282038
rect -2408 281909 -2317 282027
rect -2199 281909 240 282027
rect -2408 281867 240 281909
rect -2408 281749 -2317 281867
rect -2199 281749 240 281867
rect -2408 281738 240 281749
rect 291760 282027 294370 282038
rect 291760 281909 294161 282027
rect 294279 281909 294370 282027
rect 291760 281867 294370 281909
rect 291760 281749 294161 281867
rect 294279 281749 294370 281867
rect 291760 281738 294370 281749
rect -2408 281737 -2108 281738
rect 294070 281737 294370 281738
rect -1468 280238 -1168 280239
rect 293130 280238 293430 280239
rect -1468 280227 240 280238
rect -1468 280109 -1377 280227
rect -1259 280109 240 280227
rect -1468 280067 240 280109
rect -1468 279949 -1377 280067
rect -1259 279949 240 280067
rect -1468 279938 240 279949
rect 291760 280227 293430 280238
rect 291760 280109 293221 280227
rect 293339 280109 293430 280227
rect 291760 280067 293430 280109
rect 291760 279949 293221 280067
rect 293339 279949 293430 280067
rect 291760 279938 293430 279949
rect -1468 279937 -1168 279938
rect 293130 279937 293430 279938
rect -3818 276638 -3518 276639
rect 295480 276638 295780 276639
rect -4288 276627 240 276638
rect -4288 276509 -3727 276627
rect -3609 276509 240 276627
rect -4288 276467 240 276509
rect -4288 276349 -3727 276467
rect -3609 276349 240 276467
rect -4288 276338 240 276349
rect 291760 276627 296250 276638
rect 291760 276509 295571 276627
rect 295689 276509 296250 276627
rect 291760 276467 296250 276509
rect 291760 276349 295571 276467
rect 295689 276349 296250 276467
rect 291760 276338 296250 276349
rect -3818 276337 -3518 276338
rect 295480 276337 295780 276338
rect -2878 274838 -2578 274839
rect 294540 274838 294840 274839
rect -3348 274827 240 274838
rect -3348 274709 -2787 274827
rect -2669 274709 240 274827
rect -3348 274667 240 274709
rect -3348 274549 -2787 274667
rect -2669 274549 240 274667
rect -3348 274538 240 274549
rect 291760 274827 295310 274838
rect 291760 274709 294631 274827
rect 294749 274709 295310 274827
rect 291760 274667 295310 274709
rect 291760 274549 294631 274667
rect 294749 274549 295310 274667
rect 291760 274538 295310 274549
rect -2878 274537 -2578 274538
rect 294540 274537 294840 274538
rect -1938 273038 -1638 273039
rect 293600 273038 293900 273039
rect -2408 273027 240 273038
rect -2408 272909 -1847 273027
rect -1729 272909 240 273027
rect -2408 272867 240 272909
rect -2408 272749 -1847 272867
rect -1729 272749 240 272867
rect -2408 272738 240 272749
rect 291760 273027 294370 273038
rect 291760 272909 293691 273027
rect 293809 272909 294370 273027
rect 291760 272867 294370 272909
rect 291760 272749 293691 272867
rect 293809 272749 294370 272867
rect 291760 272738 294370 272749
rect -1938 272737 -1638 272738
rect 293600 272737 293900 272738
rect -998 271238 -698 271239
rect 292660 271238 292960 271239
rect -1468 271227 240 271238
rect -1468 271109 -907 271227
rect -789 271109 240 271227
rect -1468 271067 240 271109
rect -1468 270949 -907 271067
rect -789 270949 240 271067
rect -1468 270938 240 270949
rect 291760 271227 293430 271238
rect 291760 271109 292751 271227
rect 292869 271109 293430 271227
rect 291760 271067 293430 271109
rect 291760 270949 292751 271067
rect 292869 270949 293430 271067
rect 291760 270938 293430 270949
rect -998 270937 -698 270938
rect 292660 270937 292960 270938
rect -4288 267638 -3988 267639
rect 295950 267638 296250 267639
rect -4288 267627 240 267638
rect -4288 267509 -4197 267627
rect -4079 267509 240 267627
rect -4288 267467 240 267509
rect -4288 267349 -4197 267467
rect -4079 267349 240 267467
rect -4288 267338 240 267349
rect 291760 267627 296250 267638
rect 291760 267509 296041 267627
rect 296159 267509 296250 267627
rect 291760 267467 296250 267509
rect 291760 267349 296041 267467
rect 296159 267349 296250 267467
rect 291760 267338 296250 267349
rect -4288 267337 -3988 267338
rect 295950 267337 296250 267338
rect -3348 265838 -3048 265839
rect 295010 265838 295310 265839
rect -3348 265827 240 265838
rect -3348 265709 -3257 265827
rect -3139 265709 240 265827
rect -3348 265667 240 265709
rect -3348 265549 -3257 265667
rect -3139 265549 240 265667
rect -3348 265538 240 265549
rect 291760 265827 295310 265838
rect 291760 265709 295101 265827
rect 295219 265709 295310 265827
rect 291760 265667 295310 265709
rect 291760 265549 295101 265667
rect 295219 265549 295310 265667
rect 291760 265538 295310 265549
rect -3348 265537 -3048 265538
rect 295010 265537 295310 265538
rect -2408 264038 -2108 264039
rect 294070 264038 294370 264039
rect -2408 264027 240 264038
rect -2408 263909 -2317 264027
rect -2199 263909 240 264027
rect -2408 263867 240 263909
rect -2408 263749 -2317 263867
rect -2199 263749 240 263867
rect -2408 263738 240 263749
rect 291760 264027 294370 264038
rect 291760 263909 294161 264027
rect 294279 263909 294370 264027
rect 291760 263867 294370 263909
rect 291760 263749 294161 263867
rect 294279 263749 294370 263867
rect 291760 263738 294370 263749
rect -2408 263737 -2108 263738
rect 294070 263737 294370 263738
rect -1468 262238 -1168 262239
rect 293130 262238 293430 262239
rect -1468 262227 240 262238
rect -1468 262109 -1377 262227
rect -1259 262109 240 262227
rect -1468 262067 240 262109
rect -1468 261949 -1377 262067
rect -1259 261949 240 262067
rect -1468 261938 240 261949
rect 291760 262227 293430 262238
rect 291760 262109 293221 262227
rect 293339 262109 293430 262227
rect 291760 262067 293430 262109
rect 291760 261949 293221 262067
rect 293339 261949 293430 262067
rect 291760 261938 293430 261949
rect -1468 261937 -1168 261938
rect 293130 261937 293430 261938
rect -3818 258638 -3518 258639
rect 295480 258638 295780 258639
rect -4288 258627 240 258638
rect -4288 258509 -3727 258627
rect -3609 258509 240 258627
rect -4288 258467 240 258509
rect -4288 258349 -3727 258467
rect -3609 258349 240 258467
rect -4288 258338 240 258349
rect 291760 258627 296250 258638
rect 291760 258509 295571 258627
rect 295689 258509 296250 258627
rect 291760 258467 296250 258509
rect 291760 258349 295571 258467
rect 295689 258349 296250 258467
rect 291760 258338 296250 258349
rect -3818 258337 -3518 258338
rect 295480 258337 295780 258338
rect -2878 256838 -2578 256839
rect 294540 256838 294840 256839
rect -3348 256827 240 256838
rect -3348 256709 -2787 256827
rect -2669 256709 240 256827
rect -3348 256667 240 256709
rect -3348 256549 -2787 256667
rect -2669 256549 240 256667
rect -3348 256538 240 256549
rect 291760 256827 295310 256838
rect 291760 256709 294631 256827
rect 294749 256709 295310 256827
rect 291760 256667 295310 256709
rect 291760 256549 294631 256667
rect 294749 256549 295310 256667
rect 291760 256538 295310 256549
rect -2878 256537 -2578 256538
rect 294540 256537 294840 256538
rect -1938 255038 -1638 255039
rect 293600 255038 293900 255039
rect -2408 255027 240 255038
rect -2408 254909 -1847 255027
rect -1729 254909 240 255027
rect -2408 254867 240 254909
rect -2408 254749 -1847 254867
rect -1729 254749 240 254867
rect -2408 254738 240 254749
rect 291760 255027 294370 255038
rect 291760 254909 293691 255027
rect 293809 254909 294370 255027
rect 291760 254867 294370 254909
rect 291760 254749 293691 254867
rect 293809 254749 294370 254867
rect 291760 254738 294370 254749
rect -1938 254737 -1638 254738
rect 293600 254737 293900 254738
rect -998 253238 -698 253239
rect 292660 253238 292960 253239
rect -1468 253227 240 253238
rect -1468 253109 -907 253227
rect -789 253109 240 253227
rect -1468 253067 240 253109
rect -1468 252949 -907 253067
rect -789 252949 240 253067
rect -1468 252938 240 252949
rect 291760 253227 293430 253238
rect 291760 253109 292751 253227
rect 292869 253109 293430 253227
rect 291760 253067 293430 253109
rect 291760 252949 292751 253067
rect 292869 252949 293430 253067
rect 291760 252938 293430 252949
rect -998 252937 -698 252938
rect 292660 252937 292960 252938
rect -4288 249638 -3988 249639
rect 295950 249638 296250 249639
rect -4288 249627 240 249638
rect -4288 249509 -4197 249627
rect -4079 249509 240 249627
rect -4288 249467 240 249509
rect -4288 249349 -4197 249467
rect -4079 249349 240 249467
rect -4288 249338 240 249349
rect 291760 249627 296250 249638
rect 291760 249509 296041 249627
rect 296159 249509 296250 249627
rect 291760 249467 296250 249509
rect 291760 249349 296041 249467
rect 296159 249349 296250 249467
rect 291760 249338 296250 249349
rect -4288 249337 -3988 249338
rect 295950 249337 296250 249338
rect -3348 247838 -3048 247839
rect 295010 247838 295310 247839
rect -3348 247827 240 247838
rect -3348 247709 -3257 247827
rect -3139 247709 240 247827
rect -3348 247667 240 247709
rect -3348 247549 -3257 247667
rect -3139 247549 240 247667
rect -3348 247538 240 247549
rect 291760 247827 295310 247838
rect 291760 247709 295101 247827
rect 295219 247709 295310 247827
rect 291760 247667 295310 247709
rect 291760 247549 295101 247667
rect 295219 247549 295310 247667
rect 291760 247538 295310 247549
rect -3348 247537 -3048 247538
rect 295010 247537 295310 247538
rect -2408 246038 -2108 246039
rect 294070 246038 294370 246039
rect -2408 246027 240 246038
rect -2408 245909 -2317 246027
rect -2199 245909 240 246027
rect -2408 245867 240 245909
rect -2408 245749 -2317 245867
rect -2199 245749 240 245867
rect -2408 245738 240 245749
rect 291760 246027 294370 246038
rect 291760 245909 294161 246027
rect 294279 245909 294370 246027
rect 291760 245867 294370 245909
rect 291760 245749 294161 245867
rect 294279 245749 294370 245867
rect 291760 245738 294370 245749
rect -2408 245737 -2108 245738
rect 294070 245737 294370 245738
rect -1468 244238 -1168 244239
rect 293130 244238 293430 244239
rect -1468 244227 240 244238
rect -1468 244109 -1377 244227
rect -1259 244109 240 244227
rect -1468 244067 240 244109
rect -1468 243949 -1377 244067
rect -1259 243949 240 244067
rect -1468 243938 240 243949
rect 291760 244227 293430 244238
rect 291760 244109 293221 244227
rect 293339 244109 293430 244227
rect 291760 244067 293430 244109
rect 291760 243949 293221 244067
rect 293339 243949 293430 244067
rect 291760 243938 293430 243949
rect -1468 243937 -1168 243938
rect 293130 243937 293430 243938
rect -3818 240638 -3518 240639
rect 295480 240638 295780 240639
rect -4288 240627 240 240638
rect -4288 240509 -3727 240627
rect -3609 240509 240 240627
rect -4288 240467 240 240509
rect -4288 240349 -3727 240467
rect -3609 240349 240 240467
rect -4288 240338 240 240349
rect 291760 240627 296250 240638
rect 291760 240509 295571 240627
rect 295689 240509 296250 240627
rect 291760 240467 296250 240509
rect 291760 240349 295571 240467
rect 295689 240349 296250 240467
rect 291760 240338 296250 240349
rect -3818 240337 -3518 240338
rect 295480 240337 295780 240338
rect -2878 238838 -2578 238839
rect 294540 238838 294840 238839
rect -3348 238827 240 238838
rect -3348 238709 -2787 238827
rect -2669 238709 240 238827
rect -3348 238667 240 238709
rect -3348 238549 -2787 238667
rect -2669 238549 240 238667
rect -3348 238538 240 238549
rect 291760 238827 295310 238838
rect 291760 238709 294631 238827
rect 294749 238709 295310 238827
rect 291760 238667 295310 238709
rect 291760 238549 294631 238667
rect 294749 238549 295310 238667
rect 291760 238538 295310 238549
rect -2878 238537 -2578 238538
rect 294540 238537 294840 238538
rect -1938 237038 -1638 237039
rect 293600 237038 293900 237039
rect -2408 237027 240 237038
rect -2408 236909 -1847 237027
rect -1729 236909 240 237027
rect -2408 236867 240 236909
rect -2408 236749 -1847 236867
rect -1729 236749 240 236867
rect -2408 236738 240 236749
rect 291760 237027 294370 237038
rect 291760 236909 293691 237027
rect 293809 236909 294370 237027
rect 291760 236867 294370 236909
rect 291760 236749 293691 236867
rect 293809 236749 294370 236867
rect 291760 236738 294370 236749
rect -1938 236737 -1638 236738
rect 293600 236737 293900 236738
rect -998 235238 -698 235239
rect 292660 235238 292960 235239
rect -1468 235227 240 235238
rect -1468 235109 -907 235227
rect -789 235109 240 235227
rect -1468 235067 240 235109
rect -1468 234949 -907 235067
rect -789 234949 240 235067
rect -1468 234938 240 234949
rect 291760 235227 293430 235238
rect 291760 235109 292751 235227
rect 292869 235109 293430 235227
rect 291760 235067 293430 235109
rect 291760 234949 292751 235067
rect 292869 234949 293430 235067
rect 291760 234938 293430 234949
rect -998 234937 -698 234938
rect 292660 234937 292960 234938
rect -4288 231638 -3988 231639
rect 295950 231638 296250 231639
rect -4288 231627 240 231638
rect -4288 231509 -4197 231627
rect -4079 231509 240 231627
rect -4288 231467 240 231509
rect -4288 231349 -4197 231467
rect -4079 231349 240 231467
rect -4288 231338 240 231349
rect 291760 231627 296250 231638
rect 291760 231509 296041 231627
rect 296159 231509 296250 231627
rect 291760 231467 296250 231509
rect 291760 231349 296041 231467
rect 296159 231349 296250 231467
rect 291760 231338 296250 231349
rect -4288 231337 -3988 231338
rect 295950 231337 296250 231338
rect -3348 229838 -3048 229839
rect 295010 229838 295310 229839
rect -3348 229827 240 229838
rect -3348 229709 -3257 229827
rect -3139 229709 240 229827
rect -3348 229667 240 229709
rect -3348 229549 -3257 229667
rect -3139 229549 240 229667
rect -3348 229538 240 229549
rect 291760 229827 295310 229838
rect 291760 229709 295101 229827
rect 295219 229709 295310 229827
rect 291760 229667 295310 229709
rect 291760 229549 295101 229667
rect 295219 229549 295310 229667
rect 291760 229538 295310 229549
rect -3348 229537 -3048 229538
rect 295010 229537 295310 229538
rect -2408 228038 -2108 228039
rect 294070 228038 294370 228039
rect -2408 228027 240 228038
rect -2408 227909 -2317 228027
rect -2199 227909 240 228027
rect -2408 227867 240 227909
rect -2408 227749 -2317 227867
rect -2199 227749 240 227867
rect -2408 227738 240 227749
rect 291760 228027 294370 228038
rect 291760 227909 294161 228027
rect 294279 227909 294370 228027
rect 291760 227867 294370 227909
rect 291760 227749 294161 227867
rect 294279 227749 294370 227867
rect 291760 227738 294370 227749
rect -2408 227737 -2108 227738
rect 294070 227737 294370 227738
rect -1468 226238 -1168 226239
rect 293130 226238 293430 226239
rect -1468 226227 240 226238
rect -1468 226109 -1377 226227
rect -1259 226109 240 226227
rect -1468 226067 240 226109
rect -1468 225949 -1377 226067
rect -1259 225949 240 226067
rect -1468 225938 240 225949
rect 291760 226227 293430 226238
rect 291760 226109 293221 226227
rect 293339 226109 293430 226227
rect 291760 226067 293430 226109
rect 291760 225949 293221 226067
rect 293339 225949 293430 226067
rect 291760 225938 293430 225949
rect -1468 225937 -1168 225938
rect 293130 225937 293430 225938
rect -3818 222638 -3518 222639
rect 295480 222638 295780 222639
rect -4288 222627 240 222638
rect -4288 222509 -3727 222627
rect -3609 222509 240 222627
rect -4288 222467 240 222509
rect -4288 222349 -3727 222467
rect -3609 222349 240 222467
rect -4288 222338 240 222349
rect 291760 222627 296250 222638
rect 291760 222509 295571 222627
rect 295689 222509 296250 222627
rect 291760 222467 296250 222509
rect 291760 222349 295571 222467
rect 295689 222349 296250 222467
rect 291760 222338 296250 222349
rect -3818 222337 -3518 222338
rect 295480 222337 295780 222338
rect -2878 220838 -2578 220839
rect 294540 220838 294840 220839
rect -3348 220827 240 220838
rect -3348 220709 -2787 220827
rect -2669 220709 240 220827
rect -3348 220667 240 220709
rect -3348 220549 -2787 220667
rect -2669 220549 240 220667
rect -3348 220538 240 220549
rect 291760 220827 295310 220838
rect 291760 220709 294631 220827
rect 294749 220709 295310 220827
rect 291760 220667 295310 220709
rect 291760 220549 294631 220667
rect 294749 220549 295310 220667
rect 291760 220538 295310 220549
rect -2878 220537 -2578 220538
rect 294540 220537 294840 220538
rect -1938 219038 -1638 219039
rect 293600 219038 293900 219039
rect -2408 219027 240 219038
rect -2408 218909 -1847 219027
rect -1729 218909 240 219027
rect -2408 218867 240 218909
rect -2408 218749 -1847 218867
rect -1729 218749 240 218867
rect -2408 218738 240 218749
rect 291760 219027 294370 219038
rect 291760 218909 293691 219027
rect 293809 218909 294370 219027
rect 291760 218867 294370 218909
rect 291760 218749 293691 218867
rect 293809 218749 294370 218867
rect 291760 218738 294370 218749
rect -1938 218737 -1638 218738
rect 293600 218737 293900 218738
rect -998 217238 -698 217239
rect 292660 217238 292960 217239
rect -1468 217227 240 217238
rect -1468 217109 -907 217227
rect -789 217109 240 217227
rect -1468 217067 240 217109
rect -1468 216949 -907 217067
rect -789 216949 240 217067
rect -1468 216938 240 216949
rect 291760 217227 293430 217238
rect 291760 217109 292751 217227
rect 292869 217109 293430 217227
rect 291760 217067 293430 217109
rect 291760 216949 292751 217067
rect 292869 216949 293430 217067
rect 291760 216938 293430 216949
rect -998 216937 -698 216938
rect 292660 216937 292960 216938
rect -4288 213638 -3988 213639
rect 295950 213638 296250 213639
rect -4288 213627 240 213638
rect -4288 213509 -4197 213627
rect -4079 213509 240 213627
rect -4288 213467 240 213509
rect -4288 213349 -4197 213467
rect -4079 213349 240 213467
rect -4288 213338 240 213349
rect 291760 213627 296250 213638
rect 291760 213509 296041 213627
rect 296159 213509 296250 213627
rect 291760 213467 296250 213509
rect 291760 213349 296041 213467
rect 296159 213349 296250 213467
rect 291760 213338 296250 213349
rect -4288 213337 -3988 213338
rect 295950 213337 296250 213338
rect -3348 211838 -3048 211839
rect 295010 211838 295310 211839
rect -3348 211827 240 211838
rect -3348 211709 -3257 211827
rect -3139 211709 240 211827
rect -3348 211667 240 211709
rect -3348 211549 -3257 211667
rect -3139 211549 240 211667
rect -3348 211538 240 211549
rect 291760 211827 295310 211838
rect 291760 211709 295101 211827
rect 295219 211709 295310 211827
rect 291760 211667 295310 211709
rect 291760 211549 295101 211667
rect 295219 211549 295310 211667
rect 291760 211538 295310 211549
rect -3348 211537 -3048 211538
rect 295010 211537 295310 211538
rect -2408 210038 -2108 210039
rect 294070 210038 294370 210039
rect -2408 210027 240 210038
rect -2408 209909 -2317 210027
rect -2199 209909 240 210027
rect -2408 209867 240 209909
rect -2408 209749 -2317 209867
rect -2199 209749 240 209867
rect -2408 209738 240 209749
rect 291760 210027 294370 210038
rect 291760 209909 294161 210027
rect 294279 209909 294370 210027
rect 291760 209867 294370 209909
rect 291760 209749 294161 209867
rect 294279 209749 294370 209867
rect 291760 209738 294370 209749
rect -2408 209737 -2108 209738
rect 294070 209737 294370 209738
rect -1468 208238 -1168 208239
rect 293130 208238 293430 208239
rect -1468 208227 240 208238
rect -1468 208109 -1377 208227
rect -1259 208109 240 208227
rect -1468 208067 240 208109
rect -1468 207949 -1377 208067
rect -1259 207949 240 208067
rect -1468 207938 240 207949
rect 291760 208227 293430 208238
rect 291760 208109 293221 208227
rect 293339 208109 293430 208227
rect 291760 208067 293430 208109
rect 291760 207949 293221 208067
rect 293339 207949 293430 208067
rect 291760 207938 293430 207949
rect -1468 207937 -1168 207938
rect 293130 207937 293430 207938
rect -3818 204638 -3518 204639
rect 295480 204638 295780 204639
rect -4288 204627 240 204638
rect -4288 204509 -3727 204627
rect -3609 204509 240 204627
rect -4288 204467 240 204509
rect -4288 204349 -3727 204467
rect -3609 204349 240 204467
rect -4288 204338 240 204349
rect 291760 204627 296250 204638
rect 291760 204509 295571 204627
rect 295689 204509 296250 204627
rect 291760 204467 296250 204509
rect 291760 204349 295571 204467
rect 295689 204349 296250 204467
rect 291760 204338 296250 204349
rect -3818 204337 -3518 204338
rect 295480 204337 295780 204338
rect -2878 202838 -2578 202839
rect 294540 202838 294840 202839
rect -3348 202827 240 202838
rect -3348 202709 -2787 202827
rect -2669 202709 240 202827
rect -3348 202667 240 202709
rect -3348 202549 -2787 202667
rect -2669 202549 240 202667
rect -3348 202538 240 202549
rect 291760 202827 295310 202838
rect 291760 202709 294631 202827
rect 294749 202709 295310 202827
rect 291760 202667 295310 202709
rect 291760 202549 294631 202667
rect 294749 202549 295310 202667
rect 291760 202538 295310 202549
rect -2878 202537 -2578 202538
rect 294540 202537 294840 202538
rect -1938 201038 -1638 201039
rect 293600 201038 293900 201039
rect -2408 201027 240 201038
rect -2408 200909 -1847 201027
rect -1729 200909 240 201027
rect -2408 200867 240 200909
rect -2408 200749 -1847 200867
rect -1729 200749 240 200867
rect -2408 200738 240 200749
rect 291760 201027 294370 201038
rect 291760 200909 293691 201027
rect 293809 200909 294370 201027
rect 291760 200867 294370 200909
rect 291760 200749 293691 200867
rect 293809 200749 294370 200867
rect 291760 200738 294370 200749
rect -1938 200737 -1638 200738
rect 293600 200737 293900 200738
rect -998 199238 -698 199239
rect 292660 199238 292960 199239
rect -1468 199227 240 199238
rect -1468 199109 -907 199227
rect -789 199109 240 199227
rect -1468 199067 240 199109
rect -1468 198949 -907 199067
rect -789 198949 240 199067
rect -1468 198938 240 198949
rect 291760 199227 293430 199238
rect 291760 199109 292751 199227
rect 292869 199109 293430 199227
rect 291760 199067 293430 199109
rect 291760 198949 292751 199067
rect 292869 198949 293430 199067
rect 291760 198938 293430 198949
rect -998 198937 -698 198938
rect 292660 198937 292960 198938
rect -4288 195638 -3988 195639
rect 295950 195638 296250 195639
rect -4288 195627 240 195638
rect -4288 195509 -4197 195627
rect -4079 195509 240 195627
rect -4288 195467 240 195509
rect -4288 195349 -4197 195467
rect -4079 195349 240 195467
rect -4288 195338 240 195349
rect 291760 195627 296250 195638
rect 291760 195509 296041 195627
rect 296159 195509 296250 195627
rect 291760 195467 296250 195509
rect 291760 195349 296041 195467
rect 296159 195349 296250 195467
rect 291760 195338 296250 195349
rect -4288 195337 -3988 195338
rect 295950 195337 296250 195338
rect -3348 193838 -3048 193839
rect 295010 193838 295310 193839
rect -3348 193827 240 193838
rect -3348 193709 -3257 193827
rect -3139 193709 240 193827
rect -3348 193667 240 193709
rect -3348 193549 -3257 193667
rect -3139 193549 240 193667
rect -3348 193538 240 193549
rect 291760 193827 295310 193838
rect 291760 193709 295101 193827
rect 295219 193709 295310 193827
rect 291760 193667 295310 193709
rect 291760 193549 295101 193667
rect 295219 193549 295310 193667
rect 291760 193538 295310 193549
rect -3348 193537 -3048 193538
rect 295010 193537 295310 193538
rect -2408 192038 -2108 192039
rect 294070 192038 294370 192039
rect -2408 192027 240 192038
rect -2408 191909 -2317 192027
rect -2199 191909 240 192027
rect -2408 191867 240 191909
rect -2408 191749 -2317 191867
rect -2199 191749 240 191867
rect -2408 191738 240 191749
rect 291760 192027 294370 192038
rect 291760 191909 294161 192027
rect 294279 191909 294370 192027
rect 291760 191867 294370 191909
rect 291760 191749 294161 191867
rect 294279 191749 294370 191867
rect 291760 191738 294370 191749
rect -2408 191737 -2108 191738
rect 294070 191737 294370 191738
rect -1468 190238 -1168 190239
rect 293130 190238 293430 190239
rect -1468 190227 240 190238
rect -1468 190109 -1377 190227
rect -1259 190109 240 190227
rect -1468 190067 240 190109
rect -1468 189949 -1377 190067
rect -1259 189949 240 190067
rect -1468 189938 240 189949
rect 291760 190227 293430 190238
rect 291760 190109 293221 190227
rect 293339 190109 293430 190227
rect 291760 190067 293430 190109
rect 291760 189949 293221 190067
rect 293339 189949 293430 190067
rect 291760 189938 293430 189949
rect -1468 189937 -1168 189938
rect 293130 189937 293430 189938
rect -3818 186638 -3518 186639
rect 295480 186638 295780 186639
rect -4288 186627 240 186638
rect -4288 186509 -3727 186627
rect -3609 186509 240 186627
rect -4288 186467 240 186509
rect -4288 186349 -3727 186467
rect -3609 186349 240 186467
rect -4288 186338 240 186349
rect 291760 186627 296250 186638
rect 291760 186509 295571 186627
rect 295689 186509 296250 186627
rect 291760 186467 296250 186509
rect 291760 186349 295571 186467
rect 295689 186349 296250 186467
rect 291760 186338 296250 186349
rect -3818 186337 -3518 186338
rect 295480 186337 295780 186338
rect -2878 184838 -2578 184839
rect 294540 184838 294840 184839
rect -3348 184827 240 184838
rect -3348 184709 -2787 184827
rect -2669 184709 240 184827
rect -3348 184667 240 184709
rect -3348 184549 -2787 184667
rect -2669 184549 240 184667
rect -3348 184538 240 184549
rect 291760 184827 295310 184838
rect 291760 184709 294631 184827
rect 294749 184709 295310 184827
rect 291760 184667 295310 184709
rect 291760 184549 294631 184667
rect 294749 184549 295310 184667
rect 291760 184538 295310 184549
rect -2878 184537 -2578 184538
rect 294540 184537 294840 184538
rect -1938 183038 -1638 183039
rect 293600 183038 293900 183039
rect -2408 183027 240 183038
rect -2408 182909 -1847 183027
rect -1729 182909 240 183027
rect -2408 182867 240 182909
rect -2408 182749 -1847 182867
rect -1729 182749 240 182867
rect -2408 182738 240 182749
rect 291760 183027 294370 183038
rect 291760 182909 293691 183027
rect 293809 182909 294370 183027
rect 291760 182867 294370 182909
rect 291760 182749 293691 182867
rect 293809 182749 294370 182867
rect 291760 182738 294370 182749
rect -1938 182737 -1638 182738
rect 293600 182737 293900 182738
rect -998 181238 -698 181239
rect 292660 181238 292960 181239
rect -1468 181227 240 181238
rect -1468 181109 -907 181227
rect -789 181109 240 181227
rect -1468 181067 240 181109
rect -1468 180949 -907 181067
rect -789 180949 240 181067
rect -1468 180938 240 180949
rect 291760 181227 293430 181238
rect 291760 181109 292751 181227
rect 292869 181109 293430 181227
rect 291760 181067 293430 181109
rect 291760 180949 292751 181067
rect 292869 180949 293430 181067
rect 291760 180938 293430 180949
rect -998 180937 -698 180938
rect 292660 180937 292960 180938
rect -4288 177638 -3988 177639
rect 295950 177638 296250 177639
rect -4288 177627 240 177638
rect -4288 177509 -4197 177627
rect -4079 177509 240 177627
rect -4288 177467 240 177509
rect -4288 177349 -4197 177467
rect -4079 177349 240 177467
rect -4288 177338 240 177349
rect 291760 177627 296250 177638
rect 291760 177509 296041 177627
rect 296159 177509 296250 177627
rect 291760 177467 296250 177509
rect 291760 177349 296041 177467
rect 296159 177349 296250 177467
rect 291760 177338 296250 177349
rect -4288 177337 -3988 177338
rect 295950 177337 296250 177338
rect -3348 175838 -3048 175839
rect 295010 175838 295310 175839
rect -3348 175827 240 175838
rect -3348 175709 -3257 175827
rect -3139 175709 240 175827
rect -3348 175667 240 175709
rect -3348 175549 -3257 175667
rect -3139 175549 240 175667
rect -3348 175538 240 175549
rect 291760 175827 295310 175838
rect 291760 175709 295101 175827
rect 295219 175709 295310 175827
rect 291760 175667 295310 175709
rect 291760 175549 295101 175667
rect 295219 175549 295310 175667
rect 291760 175538 295310 175549
rect -3348 175537 -3048 175538
rect 295010 175537 295310 175538
rect -2408 174038 -2108 174039
rect 294070 174038 294370 174039
rect -2408 174027 240 174038
rect -2408 173909 -2317 174027
rect -2199 173909 240 174027
rect -2408 173867 240 173909
rect -2408 173749 -2317 173867
rect -2199 173749 240 173867
rect -2408 173738 240 173749
rect 291760 174027 294370 174038
rect 291760 173909 294161 174027
rect 294279 173909 294370 174027
rect 291760 173867 294370 173909
rect 291760 173749 294161 173867
rect 294279 173749 294370 173867
rect 291760 173738 294370 173749
rect -2408 173737 -2108 173738
rect 294070 173737 294370 173738
rect -1468 172238 -1168 172239
rect 293130 172238 293430 172239
rect -1468 172227 240 172238
rect -1468 172109 -1377 172227
rect -1259 172109 240 172227
rect -1468 172067 240 172109
rect -1468 171949 -1377 172067
rect -1259 171949 240 172067
rect -1468 171938 240 171949
rect 291760 172227 293430 172238
rect 291760 172109 293221 172227
rect 293339 172109 293430 172227
rect 291760 172067 293430 172109
rect 291760 171949 293221 172067
rect 293339 171949 293430 172067
rect 291760 171938 293430 171949
rect -1468 171937 -1168 171938
rect 293130 171937 293430 171938
rect -3818 168638 -3518 168639
rect 295480 168638 295780 168639
rect -4288 168627 240 168638
rect -4288 168509 -3727 168627
rect -3609 168509 240 168627
rect -4288 168467 240 168509
rect -4288 168349 -3727 168467
rect -3609 168349 240 168467
rect -4288 168338 240 168349
rect 291760 168627 296250 168638
rect 291760 168509 295571 168627
rect 295689 168509 296250 168627
rect 291760 168467 296250 168509
rect 291760 168349 295571 168467
rect 295689 168349 296250 168467
rect 291760 168338 296250 168349
rect -3818 168337 -3518 168338
rect 295480 168337 295780 168338
rect -2878 166838 -2578 166839
rect 294540 166838 294840 166839
rect -3348 166827 240 166838
rect -3348 166709 -2787 166827
rect -2669 166709 240 166827
rect -3348 166667 240 166709
rect -3348 166549 -2787 166667
rect -2669 166549 240 166667
rect -3348 166538 240 166549
rect 291760 166827 295310 166838
rect 291760 166709 294631 166827
rect 294749 166709 295310 166827
rect 291760 166667 295310 166709
rect 291760 166549 294631 166667
rect 294749 166549 295310 166667
rect 291760 166538 295310 166549
rect -2878 166537 -2578 166538
rect 294540 166537 294840 166538
rect -1938 165038 -1638 165039
rect 293600 165038 293900 165039
rect -2408 165027 240 165038
rect -2408 164909 -1847 165027
rect -1729 164909 240 165027
rect -2408 164867 240 164909
rect -2408 164749 -1847 164867
rect -1729 164749 240 164867
rect -2408 164738 240 164749
rect 291760 165027 294370 165038
rect 291760 164909 293691 165027
rect 293809 164909 294370 165027
rect 291760 164867 294370 164909
rect 291760 164749 293691 164867
rect 293809 164749 294370 164867
rect 291760 164738 294370 164749
rect -1938 164737 -1638 164738
rect 293600 164737 293900 164738
rect -998 163238 -698 163239
rect 292660 163238 292960 163239
rect -1468 163227 240 163238
rect -1468 163109 -907 163227
rect -789 163109 240 163227
rect -1468 163067 240 163109
rect -1468 162949 -907 163067
rect -789 162949 240 163067
rect -1468 162938 240 162949
rect 291760 163227 293430 163238
rect 291760 163109 292751 163227
rect 292869 163109 293430 163227
rect 291760 163067 293430 163109
rect 291760 162949 292751 163067
rect 292869 162949 293430 163067
rect 291760 162938 293430 162949
rect -998 162937 -698 162938
rect 292660 162937 292960 162938
rect -4288 159638 -3988 159639
rect 295950 159638 296250 159639
rect -4288 159627 240 159638
rect -4288 159509 -4197 159627
rect -4079 159509 240 159627
rect -4288 159467 240 159509
rect -4288 159349 -4197 159467
rect -4079 159349 240 159467
rect -4288 159338 240 159349
rect 291760 159627 296250 159638
rect 291760 159509 296041 159627
rect 296159 159509 296250 159627
rect 291760 159467 296250 159509
rect 291760 159349 296041 159467
rect 296159 159349 296250 159467
rect 291760 159338 296250 159349
rect -4288 159337 -3988 159338
rect 295950 159337 296250 159338
rect -3348 157838 -3048 157839
rect 295010 157838 295310 157839
rect -3348 157827 240 157838
rect -3348 157709 -3257 157827
rect -3139 157709 240 157827
rect -3348 157667 240 157709
rect -3348 157549 -3257 157667
rect -3139 157549 240 157667
rect -3348 157538 240 157549
rect 291760 157827 295310 157838
rect 291760 157709 295101 157827
rect 295219 157709 295310 157827
rect 291760 157667 295310 157709
rect 291760 157549 295101 157667
rect 295219 157549 295310 157667
rect 291760 157538 295310 157549
rect -3348 157537 -3048 157538
rect 295010 157537 295310 157538
rect -2408 156038 -2108 156039
rect 294070 156038 294370 156039
rect -2408 156027 240 156038
rect -2408 155909 -2317 156027
rect -2199 155909 240 156027
rect -2408 155867 240 155909
rect -2408 155749 -2317 155867
rect -2199 155749 240 155867
rect -2408 155738 240 155749
rect 291760 156027 294370 156038
rect 291760 155909 294161 156027
rect 294279 155909 294370 156027
rect 291760 155867 294370 155909
rect 291760 155749 294161 155867
rect 294279 155749 294370 155867
rect 291760 155738 294370 155749
rect -2408 155737 -2108 155738
rect 294070 155737 294370 155738
rect -1468 154238 -1168 154239
rect 293130 154238 293430 154239
rect -1468 154227 240 154238
rect -1468 154109 -1377 154227
rect -1259 154109 240 154227
rect -1468 154067 240 154109
rect -1468 153949 -1377 154067
rect -1259 153949 240 154067
rect -1468 153938 240 153949
rect 291760 154227 293430 154238
rect 291760 154109 293221 154227
rect 293339 154109 293430 154227
rect 291760 154067 293430 154109
rect 291760 153949 293221 154067
rect 293339 153949 293430 154067
rect 291760 153938 293430 153949
rect -1468 153937 -1168 153938
rect 293130 153937 293430 153938
rect -3818 150638 -3518 150639
rect 295480 150638 295780 150639
rect -4288 150627 240 150638
rect -4288 150509 -3727 150627
rect -3609 150509 240 150627
rect -4288 150467 240 150509
rect -4288 150349 -3727 150467
rect -3609 150349 240 150467
rect -4288 150338 240 150349
rect 291760 150627 296250 150638
rect 291760 150509 295571 150627
rect 295689 150509 296250 150627
rect 291760 150467 296250 150509
rect 291760 150349 295571 150467
rect 295689 150349 296250 150467
rect 291760 150338 296250 150349
rect -3818 150337 -3518 150338
rect 295480 150337 295780 150338
rect -2878 148838 -2578 148839
rect 294540 148838 294840 148839
rect -3348 148827 240 148838
rect -3348 148709 -2787 148827
rect -2669 148709 240 148827
rect -3348 148667 240 148709
rect -3348 148549 -2787 148667
rect -2669 148549 240 148667
rect -3348 148538 240 148549
rect 291760 148827 295310 148838
rect 291760 148709 294631 148827
rect 294749 148709 295310 148827
rect 291760 148667 295310 148709
rect 291760 148549 294631 148667
rect 294749 148549 295310 148667
rect 291760 148538 295310 148549
rect -2878 148537 -2578 148538
rect 294540 148537 294840 148538
rect -1938 147038 -1638 147039
rect 293600 147038 293900 147039
rect -2408 147027 240 147038
rect -2408 146909 -1847 147027
rect -1729 146909 240 147027
rect -2408 146867 240 146909
rect -2408 146749 -1847 146867
rect -1729 146749 240 146867
rect -2408 146738 240 146749
rect 291760 147027 294370 147038
rect 291760 146909 293691 147027
rect 293809 146909 294370 147027
rect 291760 146867 294370 146909
rect 291760 146749 293691 146867
rect 293809 146749 294370 146867
rect 291760 146738 294370 146749
rect -1938 146737 -1638 146738
rect 293600 146737 293900 146738
rect -998 145238 -698 145239
rect 292660 145238 292960 145239
rect -1468 145227 240 145238
rect -1468 145109 -907 145227
rect -789 145109 240 145227
rect -1468 145067 240 145109
rect -1468 144949 -907 145067
rect -789 144949 240 145067
rect -1468 144938 240 144949
rect 291760 145227 293430 145238
rect 291760 145109 292751 145227
rect 292869 145109 293430 145227
rect 291760 145067 293430 145109
rect 291760 144949 292751 145067
rect 292869 144949 293430 145067
rect 291760 144938 293430 144949
rect -998 144937 -698 144938
rect 292660 144937 292960 144938
rect -4288 141638 -3988 141639
rect 295950 141638 296250 141639
rect -4288 141627 240 141638
rect -4288 141509 -4197 141627
rect -4079 141509 240 141627
rect -4288 141467 240 141509
rect -4288 141349 -4197 141467
rect -4079 141349 240 141467
rect -4288 141338 240 141349
rect 291760 141627 296250 141638
rect 291760 141509 296041 141627
rect 296159 141509 296250 141627
rect 291760 141467 296250 141509
rect 291760 141349 296041 141467
rect 296159 141349 296250 141467
rect 291760 141338 296250 141349
rect -4288 141337 -3988 141338
rect 295950 141337 296250 141338
rect -3348 139838 -3048 139839
rect 295010 139838 295310 139839
rect -3348 139827 240 139838
rect -3348 139709 -3257 139827
rect -3139 139709 240 139827
rect -3348 139667 240 139709
rect -3348 139549 -3257 139667
rect -3139 139549 240 139667
rect -3348 139538 240 139549
rect 291760 139827 295310 139838
rect 291760 139709 295101 139827
rect 295219 139709 295310 139827
rect 291760 139667 295310 139709
rect 291760 139549 295101 139667
rect 295219 139549 295310 139667
rect 291760 139538 295310 139549
rect -3348 139537 -3048 139538
rect 295010 139537 295310 139538
rect -2408 138038 -2108 138039
rect 294070 138038 294370 138039
rect -2408 138027 240 138038
rect -2408 137909 -2317 138027
rect -2199 137909 240 138027
rect -2408 137867 240 137909
rect -2408 137749 -2317 137867
rect -2199 137749 240 137867
rect -2408 137738 240 137749
rect 291760 138027 294370 138038
rect 291760 137909 294161 138027
rect 294279 137909 294370 138027
rect 291760 137867 294370 137909
rect 291760 137749 294161 137867
rect 294279 137749 294370 137867
rect 291760 137738 294370 137749
rect -2408 137737 -2108 137738
rect 294070 137737 294370 137738
rect -1468 136238 -1168 136239
rect 293130 136238 293430 136239
rect -1468 136227 240 136238
rect -1468 136109 -1377 136227
rect -1259 136109 240 136227
rect -1468 136067 240 136109
rect -1468 135949 -1377 136067
rect -1259 135949 240 136067
rect -1468 135938 240 135949
rect 291760 136227 293430 136238
rect 291760 136109 293221 136227
rect 293339 136109 293430 136227
rect 291760 136067 293430 136109
rect 291760 135949 293221 136067
rect 293339 135949 293430 136067
rect 291760 135938 293430 135949
rect -1468 135937 -1168 135938
rect 293130 135937 293430 135938
rect -3818 132638 -3518 132639
rect 295480 132638 295780 132639
rect -4288 132627 240 132638
rect -4288 132509 -3727 132627
rect -3609 132509 240 132627
rect -4288 132467 240 132509
rect -4288 132349 -3727 132467
rect -3609 132349 240 132467
rect -4288 132338 240 132349
rect 291760 132627 296250 132638
rect 291760 132509 295571 132627
rect 295689 132509 296250 132627
rect 291760 132467 296250 132509
rect 291760 132349 295571 132467
rect 295689 132349 296250 132467
rect 291760 132338 296250 132349
rect -3818 132337 -3518 132338
rect 295480 132337 295780 132338
rect -2878 130838 -2578 130839
rect 294540 130838 294840 130839
rect -3348 130827 240 130838
rect -3348 130709 -2787 130827
rect -2669 130709 240 130827
rect -3348 130667 240 130709
rect -3348 130549 -2787 130667
rect -2669 130549 240 130667
rect -3348 130538 240 130549
rect 291760 130827 295310 130838
rect 291760 130709 294631 130827
rect 294749 130709 295310 130827
rect 291760 130667 295310 130709
rect 291760 130549 294631 130667
rect 294749 130549 295310 130667
rect 291760 130538 295310 130549
rect -2878 130537 -2578 130538
rect 294540 130537 294840 130538
rect -1938 129038 -1638 129039
rect 293600 129038 293900 129039
rect -2408 129027 240 129038
rect -2408 128909 -1847 129027
rect -1729 128909 240 129027
rect -2408 128867 240 128909
rect -2408 128749 -1847 128867
rect -1729 128749 240 128867
rect -2408 128738 240 128749
rect 291760 129027 294370 129038
rect 291760 128909 293691 129027
rect 293809 128909 294370 129027
rect 291760 128867 294370 128909
rect 291760 128749 293691 128867
rect 293809 128749 294370 128867
rect 291760 128738 294370 128749
rect -1938 128737 -1638 128738
rect 293600 128737 293900 128738
rect -998 127238 -698 127239
rect 292660 127238 292960 127239
rect -1468 127227 240 127238
rect -1468 127109 -907 127227
rect -789 127109 240 127227
rect -1468 127067 240 127109
rect -1468 126949 -907 127067
rect -789 126949 240 127067
rect -1468 126938 240 126949
rect 291760 127227 293430 127238
rect 291760 127109 292751 127227
rect 292869 127109 293430 127227
rect 291760 127067 293430 127109
rect 291760 126949 292751 127067
rect 292869 126949 293430 127067
rect 291760 126938 293430 126949
rect -998 126937 -698 126938
rect 292660 126937 292960 126938
rect -4288 123638 -3988 123639
rect 295950 123638 296250 123639
rect -4288 123627 240 123638
rect -4288 123509 -4197 123627
rect -4079 123509 240 123627
rect -4288 123467 240 123509
rect -4288 123349 -4197 123467
rect -4079 123349 240 123467
rect -4288 123338 240 123349
rect 291760 123627 296250 123638
rect 291760 123509 296041 123627
rect 296159 123509 296250 123627
rect 291760 123467 296250 123509
rect 291760 123349 296041 123467
rect 296159 123349 296250 123467
rect 291760 123338 296250 123349
rect -4288 123337 -3988 123338
rect 295950 123337 296250 123338
rect -3348 121838 -3048 121839
rect 295010 121838 295310 121839
rect -3348 121827 240 121838
rect -3348 121709 -3257 121827
rect -3139 121709 240 121827
rect -3348 121667 240 121709
rect -3348 121549 -3257 121667
rect -3139 121549 240 121667
rect -3348 121538 240 121549
rect 291760 121827 295310 121838
rect 291760 121709 295101 121827
rect 295219 121709 295310 121827
rect 291760 121667 295310 121709
rect 291760 121549 295101 121667
rect 295219 121549 295310 121667
rect 291760 121538 295310 121549
rect -3348 121537 -3048 121538
rect 295010 121537 295310 121538
rect -2408 120038 -2108 120039
rect 294070 120038 294370 120039
rect -2408 120027 240 120038
rect -2408 119909 -2317 120027
rect -2199 119909 240 120027
rect -2408 119867 240 119909
rect -2408 119749 -2317 119867
rect -2199 119749 240 119867
rect -2408 119738 240 119749
rect 291760 120027 294370 120038
rect 291760 119909 294161 120027
rect 294279 119909 294370 120027
rect 291760 119867 294370 119909
rect 291760 119749 294161 119867
rect 294279 119749 294370 119867
rect 291760 119738 294370 119749
rect -2408 119737 -2108 119738
rect 294070 119737 294370 119738
rect -1468 118238 -1168 118239
rect 293130 118238 293430 118239
rect -1468 118227 240 118238
rect -1468 118109 -1377 118227
rect -1259 118109 240 118227
rect -1468 118067 240 118109
rect -1468 117949 -1377 118067
rect -1259 117949 240 118067
rect -1468 117938 240 117949
rect 291760 118227 293430 118238
rect 291760 118109 293221 118227
rect 293339 118109 293430 118227
rect 291760 118067 293430 118109
rect 291760 117949 293221 118067
rect 293339 117949 293430 118067
rect 291760 117938 293430 117949
rect -1468 117937 -1168 117938
rect 293130 117937 293430 117938
rect -3818 114638 -3518 114639
rect 295480 114638 295780 114639
rect -4288 114627 240 114638
rect -4288 114509 -3727 114627
rect -3609 114509 240 114627
rect -4288 114467 240 114509
rect -4288 114349 -3727 114467
rect -3609 114349 240 114467
rect -4288 114338 240 114349
rect 291760 114627 296250 114638
rect 291760 114509 295571 114627
rect 295689 114509 296250 114627
rect 291760 114467 296250 114509
rect 291760 114349 295571 114467
rect 295689 114349 296250 114467
rect 291760 114338 296250 114349
rect -3818 114337 -3518 114338
rect 295480 114337 295780 114338
rect -2878 112838 -2578 112839
rect 294540 112838 294840 112839
rect -3348 112827 240 112838
rect -3348 112709 -2787 112827
rect -2669 112709 240 112827
rect -3348 112667 240 112709
rect -3348 112549 -2787 112667
rect -2669 112549 240 112667
rect -3348 112538 240 112549
rect 291760 112827 295310 112838
rect 291760 112709 294631 112827
rect 294749 112709 295310 112827
rect 291760 112667 295310 112709
rect 291760 112549 294631 112667
rect 294749 112549 295310 112667
rect 291760 112538 295310 112549
rect -2878 112537 -2578 112538
rect 294540 112537 294840 112538
rect -1938 111038 -1638 111039
rect 293600 111038 293900 111039
rect -2408 111027 240 111038
rect -2408 110909 -1847 111027
rect -1729 110909 240 111027
rect -2408 110867 240 110909
rect -2408 110749 -1847 110867
rect -1729 110749 240 110867
rect -2408 110738 240 110749
rect 291760 111027 294370 111038
rect 291760 110909 293691 111027
rect 293809 110909 294370 111027
rect 291760 110867 294370 110909
rect 291760 110749 293691 110867
rect 293809 110749 294370 110867
rect 291760 110738 294370 110749
rect -1938 110737 -1638 110738
rect 293600 110737 293900 110738
rect -998 109238 -698 109239
rect 292660 109238 292960 109239
rect -1468 109227 240 109238
rect -1468 109109 -907 109227
rect -789 109109 240 109227
rect -1468 109067 240 109109
rect -1468 108949 -907 109067
rect -789 108949 240 109067
rect -1468 108938 240 108949
rect 291760 109227 293430 109238
rect 291760 109109 292751 109227
rect 292869 109109 293430 109227
rect 291760 109067 293430 109109
rect 291760 108949 292751 109067
rect 292869 108949 293430 109067
rect 291760 108938 293430 108949
rect -998 108937 -698 108938
rect 292660 108937 292960 108938
rect -4288 105638 -3988 105639
rect 295950 105638 296250 105639
rect -4288 105627 240 105638
rect -4288 105509 -4197 105627
rect -4079 105509 240 105627
rect -4288 105467 240 105509
rect -4288 105349 -4197 105467
rect -4079 105349 240 105467
rect -4288 105338 240 105349
rect 291760 105627 296250 105638
rect 291760 105509 296041 105627
rect 296159 105509 296250 105627
rect 291760 105467 296250 105509
rect 291760 105349 296041 105467
rect 296159 105349 296250 105467
rect 291760 105338 296250 105349
rect -4288 105337 -3988 105338
rect 295950 105337 296250 105338
rect -3348 103838 -3048 103839
rect 295010 103838 295310 103839
rect -3348 103827 240 103838
rect -3348 103709 -3257 103827
rect -3139 103709 240 103827
rect -3348 103667 240 103709
rect -3348 103549 -3257 103667
rect -3139 103549 240 103667
rect -3348 103538 240 103549
rect 291760 103827 295310 103838
rect 291760 103709 295101 103827
rect 295219 103709 295310 103827
rect 291760 103667 295310 103709
rect 291760 103549 295101 103667
rect 295219 103549 295310 103667
rect 291760 103538 295310 103549
rect -3348 103537 -3048 103538
rect 295010 103537 295310 103538
rect -2408 102038 -2108 102039
rect 294070 102038 294370 102039
rect -2408 102027 240 102038
rect -2408 101909 -2317 102027
rect -2199 101909 240 102027
rect -2408 101867 240 101909
rect -2408 101749 -2317 101867
rect -2199 101749 240 101867
rect -2408 101738 240 101749
rect 291760 102027 294370 102038
rect 291760 101909 294161 102027
rect 294279 101909 294370 102027
rect 291760 101867 294370 101909
rect 291760 101749 294161 101867
rect 294279 101749 294370 101867
rect 291760 101738 294370 101749
rect -2408 101737 -2108 101738
rect 294070 101737 294370 101738
rect -1468 100238 -1168 100239
rect 293130 100238 293430 100239
rect -1468 100227 240 100238
rect -1468 100109 -1377 100227
rect -1259 100109 240 100227
rect -1468 100067 240 100109
rect -1468 99949 -1377 100067
rect -1259 99949 240 100067
rect -1468 99938 240 99949
rect 291760 100227 293430 100238
rect 291760 100109 293221 100227
rect 293339 100109 293430 100227
rect 291760 100067 293430 100109
rect 291760 99949 293221 100067
rect 293339 99949 293430 100067
rect 291760 99938 293430 99949
rect -1468 99937 -1168 99938
rect 293130 99937 293430 99938
rect -3818 96638 -3518 96639
rect 295480 96638 295780 96639
rect -4288 96627 240 96638
rect -4288 96509 -3727 96627
rect -3609 96509 240 96627
rect -4288 96467 240 96509
rect -4288 96349 -3727 96467
rect -3609 96349 240 96467
rect -4288 96338 240 96349
rect 291760 96627 296250 96638
rect 291760 96509 295571 96627
rect 295689 96509 296250 96627
rect 291760 96467 296250 96509
rect 291760 96349 295571 96467
rect 295689 96349 296250 96467
rect 291760 96338 296250 96349
rect -3818 96337 -3518 96338
rect 295480 96337 295780 96338
rect -2878 94838 -2578 94839
rect 294540 94838 294840 94839
rect -3348 94827 240 94838
rect -3348 94709 -2787 94827
rect -2669 94709 240 94827
rect -3348 94667 240 94709
rect -3348 94549 -2787 94667
rect -2669 94549 240 94667
rect -3348 94538 240 94549
rect 291760 94827 295310 94838
rect 291760 94709 294631 94827
rect 294749 94709 295310 94827
rect 291760 94667 295310 94709
rect 291760 94549 294631 94667
rect 294749 94549 295310 94667
rect 291760 94538 295310 94549
rect -2878 94537 -2578 94538
rect 294540 94537 294840 94538
rect -1938 93038 -1638 93039
rect 293600 93038 293900 93039
rect -2408 93027 240 93038
rect -2408 92909 -1847 93027
rect -1729 92909 240 93027
rect -2408 92867 240 92909
rect -2408 92749 -1847 92867
rect -1729 92749 240 92867
rect -2408 92738 240 92749
rect 291760 93027 294370 93038
rect 291760 92909 293691 93027
rect 293809 92909 294370 93027
rect 291760 92867 294370 92909
rect 291760 92749 293691 92867
rect 293809 92749 294370 92867
rect 291760 92738 294370 92749
rect -1938 92737 -1638 92738
rect 293600 92737 293900 92738
rect -998 91238 -698 91239
rect 292660 91238 292960 91239
rect -1468 91227 240 91238
rect -1468 91109 -907 91227
rect -789 91109 240 91227
rect -1468 91067 240 91109
rect -1468 90949 -907 91067
rect -789 90949 240 91067
rect -1468 90938 240 90949
rect 291760 91227 293430 91238
rect 291760 91109 292751 91227
rect 292869 91109 293430 91227
rect 291760 91067 293430 91109
rect 291760 90949 292751 91067
rect 292869 90949 293430 91067
rect 291760 90938 293430 90949
rect -998 90937 -698 90938
rect 292660 90937 292960 90938
rect -4288 87638 -3988 87639
rect 295950 87638 296250 87639
rect -4288 87627 240 87638
rect -4288 87509 -4197 87627
rect -4079 87509 240 87627
rect -4288 87467 240 87509
rect -4288 87349 -4197 87467
rect -4079 87349 240 87467
rect -4288 87338 240 87349
rect 291760 87627 296250 87638
rect 291760 87509 296041 87627
rect 296159 87509 296250 87627
rect 291760 87467 296250 87509
rect 291760 87349 296041 87467
rect 296159 87349 296250 87467
rect 291760 87338 296250 87349
rect -4288 87337 -3988 87338
rect 295950 87337 296250 87338
rect -3348 85838 -3048 85839
rect 295010 85838 295310 85839
rect -3348 85827 240 85838
rect -3348 85709 -3257 85827
rect -3139 85709 240 85827
rect -3348 85667 240 85709
rect -3348 85549 -3257 85667
rect -3139 85549 240 85667
rect -3348 85538 240 85549
rect 291760 85827 295310 85838
rect 291760 85709 295101 85827
rect 295219 85709 295310 85827
rect 291760 85667 295310 85709
rect 291760 85549 295101 85667
rect 295219 85549 295310 85667
rect 291760 85538 295310 85549
rect -3348 85537 -3048 85538
rect 295010 85537 295310 85538
rect -2408 84038 -2108 84039
rect 294070 84038 294370 84039
rect -2408 84027 240 84038
rect -2408 83909 -2317 84027
rect -2199 83909 240 84027
rect -2408 83867 240 83909
rect -2408 83749 -2317 83867
rect -2199 83749 240 83867
rect -2408 83738 240 83749
rect 291760 84027 294370 84038
rect 291760 83909 294161 84027
rect 294279 83909 294370 84027
rect 291760 83867 294370 83909
rect 291760 83749 294161 83867
rect 294279 83749 294370 83867
rect 291760 83738 294370 83749
rect -2408 83737 -2108 83738
rect 294070 83737 294370 83738
rect -1468 82238 -1168 82239
rect 293130 82238 293430 82239
rect -1468 82227 240 82238
rect -1468 82109 -1377 82227
rect -1259 82109 240 82227
rect -1468 82067 240 82109
rect -1468 81949 -1377 82067
rect -1259 81949 240 82067
rect -1468 81938 240 81949
rect 291760 82227 293430 82238
rect 291760 82109 293221 82227
rect 293339 82109 293430 82227
rect 291760 82067 293430 82109
rect 291760 81949 293221 82067
rect 293339 81949 293430 82067
rect 291760 81938 293430 81949
rect -1468 81937 -1168 81938
rect 293130 81937 293430 81938
rect -3818 78638 -3518 78639
rect 295480 78638 295780 78639
rect -4288 78627 240 78638
rect -4288 78509 -3727 78627
rect -3609 78509 240 78627
rect -4288 78467 240 78509
rect -4288 78349 -3727 78467
rect -3609 78349 240 78467
rect -4288 78338 240 78349
rect 291760 78627 296250 78638
rect 291760 78509 295571 78627
rect 295689 78509 296250 78627
rect 291760 78467 296250 78509
rect 291760 78349 295571 78467
rect 295689 78349 296250 78467
rect 291760 78338 296250 78349
rect -3818 78337 -3518 78338
rect 295480 78337 295780 78338
rect -2878 76838 -2578 76839
rect 294540 76838 294840 76839
rect -3348 76827 240 76838
rect -3348 76709 -2787 76827
rect -2669 76709 240 76827
rect -3348 76667 240 76709
rect -3348 76549 -2787 76667
rect -2669 76549 240 76667
rect -3348 76538 240 76549
rect 291760 76827 295310 76838
rect 291760 76709 294631 76827
rect 294749 76709 295310 76827
rect 291760 76667 295310 76709
rect 291760 76549 294631 76667
rect 294749 76549 295310 76667
rect 291760 76538 295310 76549
rect -2878 76537 -2578 76538
rect 294540 76537 294840 76538
rect -1938 75038 -1638 75039
rect 293600 75038 293900 75039
rect -2408 75027 240 75038
rect -2408 74909 -1847 75027
rect -1729 74909 240 75027
rect -2408 74867 240 74909
rect -2408 74749 -1847 74867
rect -1729 74749 240 74867
rect -2408 74738 240 74749
rect 291760 75027 294370 75038
rect 291760 74909 293691 75027
rect 293809 74909 294370 75027
rect 291760 74867 294370 74909
rect 291760 74749 293691 74867
rect 293809 74749 294370 74867
rect 291760 74738 294370 74749
rect -1938 74737 -1638 74738
rect 293600 74737 293900 74738
rect -998 73238 -698 73239
rect 292660 73238 292960 73239
rect -1468 73227 240 73238
rect -1468 73109 -907 73227
rect -789 73109 240 73227
rect -1468 73067 240 73109
rect -1468 72949 -907 73067
rect -789 72949 240 73067
rect -1468 72938 240 72949
rect 291760 73227 293430 73238
rect 291760 73109 292751 73227
rect 292869 73109 293430 73227
rect 291760 73067 293430 73109
rect 291760 72949 292751 73067
rect 292869 72949 293430 73067
rect 291760 72938 293430 72949
rect -998 72937 -698 72938
rect 292660 72937 292960 72938
rect -4288 69638 -3988 69639
rect 295950 69638 296250 69639
rect -4288 69627 240 69638
rect -4288 69509 -4197 69627
rect -4079 69509 240 69627
rect -4288 69467 240 69509
rect -4288 69349 -4197 69467
rect -4079 69349 240 69467
rect -4288 69338 240 69349
rect 291760 69627 296250 69638
rect 291760 69509 296041 69627
rect 296159 69509 296250 69627
rect 291760 69467 296250 69509
rect 291760 69349 296041 69467
rect 296159 69349 296250 69467
rect 291760 69338 296250 69349
rect -4288 69337 -3988 69338
rect 295950 69337 296250 69338
rect -3348 67838 -3048 67839
rect 295010 67838 295310 67839
rect -3348 67827 240 67838
rect -3348 67709 -3257 67827
rect -3139 67709 240 67827
rect -3348 67667 240 67709
rect -3348 67549 -3257 67667
rect -3139 67549 240 67667
rect -3348 67538 240 67549
rect 291760 67827 295310 67838
rect 291760 67709 295101 67827
rect 295219 67709 295310 67827
rect 291760 67667 295310 67709
rect 291760 67549 295101 67667
rect 295219 67549 295310 67667
rect 291760 67538 295310 67549
rect -3348 67537 -3048 67538
rect 295010 67537 295310 67538
rect -2408 66038 -2108 66039
rect 294070 66038 294370 66039
rect -2408 66027 240 66038
rect -2408 65909 -2317 66027
rect -2199 65909 240 66027
rect -2408 65867 240 65909
rect -2408 65749 -2317 65867
rect -2199 65749 240 65867
rect -2408 65738 240 65749
rect 291760 66027 294370 66038
rect 291760 65909 294161 66027
rect 294279 65909 294370 66027
rect 291760 65867 294370 65909
rect 291760 65749 294161 65867
rect 294279 65749 294370 65867
rect 291760 65738 294370 65749
rect -2408 65737 -2108 65738
rect 294070 65737 294370 65738
rect -1468 64238 -1168 64239
rect 293130 64238 293430 64239
rect -1468 64227 240 64238
rect -1468 64109 -1377 64227
rect -1259 64109 240 64227
rect -1468 64067 240 64109
rect -1468 63949 -1377 64067
rect -1259 63949 240 64067
rect -1468 63938 240 63949
rect 291760 64227 293430 64238
rect 291760 64109 293221 64227
rect 293339 64109 293430 64227
rect 291760 64067 293430 64109
rect 291760 63949 293221 64067
rect 293339 63949 293430 64067
rect 291760 63938 293430 63949
rect -1468 63937 -1168 63938
rect 293130 63937 293430 63938
rect -3818 60638 -3518 60639
rect 295480 60638 295780 60639
rect -4288 60627 240 60638
rect -4288 60509 -3727 60627
rect -3609 60509 240 60627
rect -4288 60467 240 60509
rect -4288 60349 -3727 60467
rect -3609 60349 240 60467
rect -4288 60338 240 60349
rect 291760 60627 296250 60638
rect 291760 60509 295571 60627
rect 295689 60509 296250 60627
rect 291760 60467 296250 60509
rect 291760 60349 295571 60467
rect 295689 60349 296250 60467
rect 291760 60338 296250 60349
rect -3818 60337 -3518 60338
rect 295480 60337 295780 60338
rect -2878 58838 -2578 58839
rect 294540 58838 294840 58839
rect -3348 58827 240 58838
rect -3348 58709 -2787 58827
rect -2669 58709 240 58827
rect -3348 58667 240 58709
rect -3348 58549 -2787 58667
rect -2669 58549 240 58667
rect -3348 58538 240 58549
rect 291760 58827 295310 58838
rect 291760 58709 294631 58827
rect 294749 58709 295310 58827
rect 291760 58667 295310 58709
rect 291760 58549 294631 58667
rect 294749 58549 295310 58667
rect 291760 58538 295310 58549
rect -2878 58537 -2578 58538
rect 294540 58537 294840 58538
rect -1938 57038 -1638 57039
rect 293600 57038 293900 57039
rect -2408 57027 240 57038
rect -2408 56909 -1847 57027
rect -1729 56909 240 57027
rect -2408 56867 240 56909
rect -2408 56749 -1847 56867
rect -1729 56749 240 56867
rect -2408 56738 240 56749
rect 291760 57027 294370 57038
rect 291760 56909 293691 57027
rect 293809 56909 294370 57027
rect 291760 56867 294370 56909
rect 291760 56749 293691 56867
rect 293809 56749 294370 56867
rect 291760 56738 294370 56749
rect -1938 56737 -1638 56738
rect 293600 56737 293900 56738
rect -998 55238 -698 55239
rect 292660 55238 292960 55239
rect -1468 55227 240 55238
rect -1468 55109 -907 55227
rect -789 55109 240 55227
rect -1468 55067 240 55109
rect -1468 54949 -907 55067
rect -789 54949 240 55067
rect -1468 54938 240 54949
rect 291760 55227 293430 55238
rect 291760 55109 292751 55227
rect 292869 55109 293430 55227
rect 291760 55067 293430 55109
rect 291760 54949 292751 55067
rect 292869 54949 293430 55067
rect 291760 54938 293430 54949
rect -998 54937 -698 54938
rect 292660 54937 292960 54938
rect -4288 51638 -3988 51639
rect 295950 51638 296250 51639
rect -4288 51627 240 51638
rect -4288 51509 -4197 51627
rect -4079 51509 240 51627
rect -4288 51467 240 51509
rect -4288 51349 -4197 51467
rect -4079 51349 240 51467
rect -4288 51338 240 51349
rect 291760 51627 296250 51638
rect 291760 51509 296041 51627
rect 296159 51509 296250 51627
rect 291760 51467 296250 51509
rect 291760 51349 296041 51467
rect 296159 51349 296250 51467
rect 291760 51338 296250 51349
rect -4288 51337 -3988 51338
rect 295950 51337 296250 51338
rect -3348 49838 -3048 49839
rect 295010 49838 295310 49839
rect -3348 49827 240 49838
rect -3348 49709 -3257 49827
rect -3139 49709 240 49827
rect -3348 49667 240 49709
rect -3348 49549 -3257 49667
rect -3139 49549 240 49667
rect -3348 49538 240 49549
rect 291760 49827 295310 49838
rect 291760 49709 295101 49827
rect 295219 49709 295310 49827
rect 291760 49667 295310 49709
rect 291760 49549 295101 49667
rect 295219 49549 295310 49667
rect 291760 49538 295310 49549
rect -3348 49537 -3048 49538
rect 295010 49537 295310 49538
rect -2408 48038 -2108 48039
rect 294070 48038 294370 48039
rect -2408 48027 240 48038
rect -2408 47909 -2317 48027
rect -2199 47909 240 48027
rect -2408 47867 240 47909
rect -2408 47749 -2317 47867
rect -2199 47749 240 47867
rect -2408 47738 240 47749
rect 291760 48027 294370 48038
rect 291760 47909 294161 48027
rect 294279 47909 294370 48027
rect 291760 47867 294370 47909
rect 291760 47749 294161 47867
rect 294279 47749 294370 47867
rect 291760 47738 294370 47749
rect -2408 47737 -2108 47738
rect 294070 47737 294370 47738
rect -1468 46238 -1168 46239
rect 293130 46238 293430 46239
rect -1468 46227 240 46238
rect -1468 46109 -1377 46227
rect -1259 46109 240 46227
rect -1468 46067 240 46109
rect -1468 45949 -1377 46067
rect -1259 45949 240 46067
rect -1468 45938 240 45949
rect 291760 46227 293430 46238
rect 291760 46109 293221 46227
rect 293339 46109 293430 46227
rect 291760 46067 293430 46109
rect 291760 45949 293221 46067
rect 293339 45949 293430 46067
rect 291760 45938 293430 45949
rect -1468 45937 -1168 45938
rect 293130 45937 293430 45938
rect -3818 42638 -3518 42639
rect 295480 42638 295780 42639
rect -4288 42627 240 42638
rect -4288 42509 -3727 42627
rect -3609 42509 240 42627
rect -4288 42467 240 42509
rect -4288 42349 -3727 42467
rect -3609 42349 240 42467
rect -4288 42338 240 42349
rect 291760 42627 296250 42638
rect 291760 42509 295571 42627
rect 295689 42509 296250 42627
rect 291760 42467 296250 42509
rect 291760 42349 295571 42467
rect 295689 42349 296250 42467
rect 291760 42338 296250 42349
rect -3818 42337 -3518 42338
rect 295480 42337 295780 42338
rect -2878 40838 -2578 40839
rect 294540 40838 294840 40839
rect -3348 40827 240 40838
rect -3348 40709 -2787 40827
rect -2669 40709 240 40827
rect -3348 40667 240 40709
rect -3348 40549 -2787 40667
rect -2669 40549 240 40667
rect -3348 40538 240 40549
rect 291760 40827 295310 40838
rect 291760 40709 294631 40827
rect 294749 40709 295310 40827
rect 291760 40667 295310 40709
rect 291760 40549 294631 40667
rect 294749 40549 295310 40667
rect 291760 40538 295310 40549
rect -2878 40537 -2578 40538
rect 294540 40537 294840 40538
rect -1938 39038 -1638 39039
rect 293600 39038 293900 39039
rect -2408 39027 240 39038
rect -2408 38909 -1847 39027
rect -1729 38909 240 39027
rect -2408 38867 240 38909
rect -2408 38749 -1847 38867
rect -1729 38749 240 38867
rect -2408 38738 240 38749
rect 291760 39027 294370 39038
rect 291760 38909 293691 39027
rect 293809 38909 294370 39027
rect 291760 38867 294370 38909
rect 291760 38749 293691 38867
rect 293809 38749 294370 38867
rect 291760 38738 294370 38749
rect -1938 38737 -1638 38738
rect 293600 38737 293900 38738
rect -998 37238 -698 37239
rect 292660 37238 292960 37239
rect -1468 37227 240 37238
rect -1468 37109 -907 37227
rect -789 37109 240 37227
rect -1468 37067 240 37109
rect -1468 36949 -907 37067
rect -789 36949 240 37067
rect -1468 36938 240 36949
rect 291760 37227 293430 37238
rect 291760 37109 292751 37227
rect 292869 37109 293430 37227
rect 291760 37067 293430 37109
rect 291760 36949 292751 37067
rect 292869 36949 293430 37067
rect 291760 36938 293430 36949
rect -998 36937 -698 36938
rect 292660 36937 292960 36938
rect -4288 33638 -3988 33639
rect 295950 33638 296250 33639
rect -4288 33627 240 33638
rect -4288 33509 -4197 33627
rect -4079 33509 240 33627
rect -4288 33467 240 33509
rect -4288 33349 -4197 33467
rect -4079 33349 240 33467
rect -4288 33338 240 33349
rect 291760 33627 296250 33638
rect 291760 33509 296041 33627
rect 296159 33509 296250 33627
rect 291760 33467 296250 33509
rect 291760 33349 296041 33467
rect 296159 33349 296250 33467
rect 291760 33338 296250 33349
rect -4288 33337 -3988 33338
rect 295950 33337 296250 33338
rect -3348 31838 -3048 31839
rect 295010 31838 295310 31839
rect -3348 31827 240 31838
rect -3348 31709 -3257 31827
rect -3139 31709 240 31827
rect -3348 31667 240 31709
rect -3348 31549 -3257 31667
rect -3139 31549 240 31667
rect -3348 31538 240 31549
rect 291760 31827 295310 31838
rect 291760 31709 295101 31827
rect 295219 31709 295310 31827
rect 291760 31667 295310 31709
rect 291760 31549 295101 31667
rect 295219 31549 295310 31667
rect 291760 31538 295310 31549
rect -3348 31537 -3048 31538
rect 295010 31537 295310 31538
rect -2408 30038 -2108 30039
rect 294070 30038 294370 30039
rect -2408 30027 240 30038
rect -2408 29909 -2317 30027
rect -2199 29909 240 30027
rect -2408 29867 240 29909
rect -2408 29749 -2317 29867
rect -2199 29749 240 29867
rect -2408 29738 240 29749
rect 291760 30027 294370 30038
rect 291760 29909 294161 30027
rect 294279 29909 294370 30027
rect 291760 29867 294370 29909
rect 291760 29749 294161 29867
rect 294279 29749 294370 29867
rect 291760 29738 294370 29749
rect -2408 29737 -2108 29738
rect 294070 29737 294370 29738
rect -1468 28238 -1168 28239
rect 293130 28238 293430 28239
rect -1468 28227 240 28238
rect -1468 28109 -1377 28227
rect -1259 28109 240 28227
rect -1468 28067 240 28109
rect -1468 27949 -1377 28067
rect -1259 27949 240 28067
rect -1468 27938 240 27949
rect 291760 28227 293430 28238
rect 291760 28109 293221 28227
rect 293339 28109 293430 28227
rect 291760 28067 293430 28109
rect 291760 27949 293221 28067
rect 293339 27949 293430 28067
rect 291760 27938 293430 27949
rect -1468 27937 -1168 27938
rect 293130 27937 293430 27938
rect -3818 24638 -3518 24639
rect 295480 24638 295780 24639
rect -4288 24627 240 24638
rect -4288 24509 -3727 24627
rect -3609 24509 240 24627
rect -4288 24467 240 24509
rect -4288 24349 -3727 24467
rect -3609 24349 240 24467
rect -4288 24338 240 24349
rect 291760 24627 296250 24638
rect 291760 24509 295571 24627
rect 295689 24509 296250 24627
rect 291760 24467 296250 24509
rect 291760 24349 295571 24467
rect 295689 24349 296250 24467
rect 291760 24338 296250 24349
rect -3818 24337 -3518 24338
rect 295480 24337 295780 24338
rect -2878 22838 -2578 22839
rect 294540 22838 294840 22839
rect -3348 22827 240 22838
rect -3348 22709 -2787 22827
rect -2669 22709 240 22827
rect -3348 22667 240 22709
rect -3348 22549 -2787 22667
rect -2669 22549 240 22667
rect -3348 22538 240 22549
rect 291760 22827 295310 22838
rect 291760 22709 294631 22827
rect 294749 22709 295310 22827
rect 291760 22667 295310 22709
rect 291760 22549 294631 22667
rect 294749 22549 295310 22667
rect 291760 22538 295310 22549
rect -2878 22537 -2578 22538
rect 294540 22537 294840 22538
rect -1938 21038 -1638 21039
rect 293600 21038 293900 21039
rect -2408 21027 240 21038
rect -2408 20909 -1847 21027
rect -1729 20909 240 21027
rect -2408 20867 240 20909
rect -2408 20749 -1847 20867
rect -1729 20749 240 20867
rect -2408 20738 240 20749
rect 291760 21027 294370 21038
rect 291760 20909 293691 21027
rect 293809 20909 294370 21027
rect 291760 20867 294370 20909
rect 291760 20749 293691 20867
rect 293809 20749 294370 20867
rect 291760 20738 294370 20749
rect -1938 20737 -1638 20738
rect 293600 20737 293900 20738
rect -998 19238 -698 19239
rect 292660 19238 292960 19239
rect -1468 19227 240 19238
rect -1468 19109 -907 19227
rect -789 19109 240 19227
rect -1468 19067 240 19109
rect -1468 18949 -907 19067
rect -789 18949 240 19067
rect -1468 18938 240 18949
rect 291760 19227 293430 19238
rect 291760 19109 292751 19227
rect 292869 19109 293430 19227
rect 291760 19067 293430 19109
rect 291760 18949 292751 19067
rect 292869 18949 293430 19067
rect 291760 18938 293430 18949
rect -998 18937 -698 18938
rect 292660 18937 292960 18938
rect -4288 15638 -3988 15639
rect 295950 15638 296250 15639
rect -4288 15627 240 15638
rect -4288 15509 -4197 15627
rect -4079 15509 240 15627
rect -4288 15467 240 15509
rect -4288 15349 -4197 15467
rect -4079 15349 240 15467
rect -4288 15338 240 15349
rect 291760 15627 296250 15638
rect 291760 15509 296041 15627
rect 296159 15509 296250 15627
rect 291760 15467 296250 15509
rect 291760 15349 296041 15467
rect 296159 15349 296250 15467
rect 291760 15338 296250 15349
rect -4288 15337 -3988 15338
rect 295950 15337 296250 15338
rect -3348 13838 -3048 13839
rect 295010 13838 295310 13839
rect -3348 13827 240 13838
rect -3348 13709 -3257 13827
rect -3139 13709 240 13827
rect -3348 13667 240 13709
rect -3348 13549 -3257 13667
rect -3139 13549 240 13667
rect -3348 13538 240 13549
rect 291760 13827 295310 13838
rect 291760 13709 295101 13827
rect 295219 13709 295310 13827
rect 291760 13667 295310 13709
rect 291760 13549 295101 13667
rect 295219 13549 295310 13667
rect 291760 13538 295310 13549
rect -3348 13537 -3048 13538
rect 295010 13537 295310 13538
rect -2408 12038 -2108 12039
rect 294070 12038 294370 12039
rect -2408 12027 240 12038
rect -2408 11909 -2317 12027
rect -2199 11909 240 12027
rect -2408 11867 240 11909
rect -2408 11749 -2317 11867
rect -2199 11749 240 11867
rect -2408 11738 240 11749
rect 291760 12027 294370 12038
rect 291760 11909 294161 12027
rect 294279 11909 294370 12027
rect 291760 11867 294370 11909
rect 291760 11749 294161 11867
rect 294279 11749 294370 11867
rect 291760 11738 294370 11749
rect -2408 11737 -2108 11738
rect 294070 11737 294370 11738
rect -1468 10238 -1168 10239
rect 293130 10238 293430 10239
rect -1468 10227 240 10238
rect -1468 10109 -1377 10227
rect -1259 10109 240 10227
rect -1468 10067 240 10109
rect -1468 9949 -1377 10067
rect -1259 9949 240 10067
rect -1468 9938 240 9949
rect 291760 10227 293430 10238
rect 291760 10109 293221 10227
rect 293339 10109 293430 10227
rect 291760 10067 293430 10109
rect 291760 9949 293221 10067
rect 293339 9949 293430 10067
rect 291760 9938 293430 9949
rect -1468 9937 -1168 9938
rect 293130 9937 293430 9938
rect -3818 6638 -3518 6639
rect 295480 6638 295780 6639
rect -4288 6627 240 6638
rect -4288 6509 -3727 6627
rect -3609 6509 240 6627
rect -4288 6467 240 6509
rect -4288 6349 -3727 6467
rect -3609 6349 240 6467
rect -4288 6338 240 6349
rect 291760 6627 296250 6638
rect 291760 6509 295571 6627
rect 295689 6509 296250 6627
rect 291760 6467 296250 6509
rect 291760 6349 295571 6467
rect 295689 6349 296250 6467
rect 291760 6338 296250 6349
rect -3818 6337 -3518 6338
rect 295480 6337 295780 6338
rect -2878 4838 -2578 4839
rect 294540 4838 294840 4839
rect -3348 4827 240 4838
rect -3348 4709 -2787 4827
rect -2669 4709 240 4827
rect -3348 4667 240 4709
rect -3348 4549 -2787 4667
rect -2669 4549 240 4667
rect -3348 4538 240 4549
rect 291760 4827 295310 4838
rect 291760 4709 294631 4827
rect 294749 4709 295310 4827
rect 291760 4667 295310 4709
rect 291760 4549 294631 4667
rect 294749 4549 295310 4667
rect 291760 4538 295310 4549
rect -2878 4537 -2578 4538
rect 294540 4537 294840 4538
rect -1938 3038 -1638 3039
rect 293600 3038 293900 3039
rect -2408 3027 240 3038
rect -2408 2909 -1847 3027
rect -1729 2909 240 3027
rect -2408 2867 240 2909
rect -2408 2749 -1847 2867
rect -1729 2749 240 2867
rect -2408 2738 240 2749
rect 291760 3027 294370 3038
rect 291760 2909 293691 3027
rect 293809 2909 294370 3027
rect 291760 2867 294370 2909
rect 291760 2749 293691 2867
rect 293809 2749 294370 2867
rect 291760 2738 294370 2749
rect -1938 2737 -1638 2738
rect 293600 2737 293900 2738
rect -998 1238 -698 1239
rect 292660 1238 292960 1239
rect -1468 1227 240 1238
rect -1468 1109 -907 1227
rect -789 1109 240 1227
rect -1468 1067 240 1109
rect -1468 949 -907 1067
rect -789 949 240 1067
rect -1468 938 240 949
rect 291760 1227 293430 1238
rect 291760 1109 292751 1227
rect 292869 1109 293430 1227
rect 291760 1067 293430 1109
rect 291760 949 292751 1067
rect 292869 949 293430 1067
rect 291760 938 293430 949
rect -998 937 -698 938
rect 292660 937 292960 938
rect -998 -162 -698 -161
rect 402 -162 702 -161
rect 18402 -162 18702 -161
rect 36402 -162 36702 -161
rect 54402 -162 54702 -161
rect 72402 -162 72702 -161
rect 90402 -162 90702 -161
rect 108402 -162 108702 -161
rect 126402 -162 126702 -161
rect 144402 -162 144702 -161
rect 162402 -162 162702 -161
rect 180402 -162 180702 -161
rect 198402 -162 198702 -161
rect 216402 -162 216702 -161
rect 234402 -162 234702 -161
rect 252402 -162 252702 -161
rect 270402 -162 270702 -161
rect 288402 -162 288702 -161
rect 292660 -162 292960 -161
rect -998 -173 292960 -162
rect -998 -291 -907 -173
rect -789 -291 493 -173
rect 611 -291 18493 -173
rect 18611 -291 36493 -173
rect 36611 -291 54493 -173
rect 54611 -291 72493 -173
rect 72611 -291 90493 -173
rect 90611 -291 108493 -173
rect 108611 -291 126493 -173
rect 126611 -291 144493 -173
rect 144611 -291 162493 -173
rect 162611 -291 180493 -173
rect 180611 -291 198493 -173
rect 198611 -291 216493 -173
rect 216611 -291 234493 -173
rect 234611 -291 252493 -173
rect 252611 -291 270493 -173
rect 270611 -291 288493 -173
rect 288611 -291 292751 -173
rect 292869 -291 292960 -173
rect -998 -333 292960 -291
rect -998 -451 -907 -333
rect -789 -451 493 -333
rect 611 -451 18493 -333
rect 18611 -451 36493 -333
rect 36611 -451 54493 -333
rect 54611 -451 72493 -333
rect 72611 -451 90493 -333
rect 90611 -451 108493 -333
rect 108611 -451 126493 -333
rect 126611 -451 144493 -333
rect 144611 -451 162493 -333
rect 162611 -451 180493 -333
rect 180611 -451 198493 -333
rect 198611 -451 216493 -333
rect 216611 -451 234493 -333
rect 234611 -451 252493 -333
rect 252611 -451 270493 -333
rect 270611 -451 288493 -333
rect 288611 -451 292751 -333
rect 292869 -451 292960 -333
rect -998 -462 292960 -451
rect -998 -463 -698 -462
rect 402 -463 702 -462
rect 18402 -463 18702 -462
rect 36402 -463 36702 -462
rect 54402 -463 54702 -462
rect 72402 -463 72702 -462
rect 90402 -463 90702 -462
rect 108402 -463 108702 -462
rect 126402 -463 126702 -462
rect 144402 -463 144702 -462
rect 162402 -463 162702 -462
rect 180402 -463 180702 -462
rect 198402 -463 198702 -462
rect 216402 -463 216702 -462
rect 234402 -463 234702 -462
rect 252402 -463 252702 -462
rect 270402 -463 270702 -462
rect 288402 -463 288702 -462
rect 292660 -463 292960 -462
rect -1468 -632 -1168 -631
rect 9402 -632 9702 -631
rect 27402 -632 27702 -631
rect 45402 -632 45702 -631
rect 63402 -632 63702 -631
rect 81402 -632 81702 -631
rect 99402 -632 99702 -631
rect 117402 -632 117702 -631
rect 135402 -632 135702 -631
rect 153402 -632 153702 -631
rect 171402 -632 171702 -631
rect 189402 -632 189702 -631
rect 207402 -632 207702 -631
rect 225402 -632 225702 -631
rect 243402 -632 243702 -631
rect 261402 -632 261702 -631
rect 279402 -632 279702 -631
rect 293130 -632 293430 -631
rect -1468 -643 293430 -632
rect -1468 -761 -1377 -643
rect -1259 -761 9493 -643
rect 9611 -761 27493 -643
rect 27611 -761 45493 -643
rect 45611 -761 63493 -643
rect 63611 -761 81493 -643
rect 81611 -761 99493 -643
rect 99611 -761 117493 -643
rect 117611 -761 135493 -643
rect 135611 -761 153493 -643
rect 153611 -761 171493 -643
rect 171611 -761 189493 -643
rect 189611 -761 207493 -643
rect 207611 -761 225493 -643
rect 225611 -761 243493 -643
rect 243611 -761 261493 -643
rect 261611 -761 279493 -643
rect 279611 -761 293221 -643
rect 293339 -761 293430 -643
rect -1468 -803 293430 -761
rect -1468 -921 -1377 -803
rect -1259 -921 9493 -803
rect 9611 -921 27493 -803
rect 27611 -921 45493 -803
rect 45611 -921 63493 -803
rect 63611 -921 81493 -803
rect 81611 -921 99493 -803
rect 99611 -921 117493 -803
rect 117611 -921 135493 -803
rect 135611 -921 153493 -803
rect 153611 -921 171493 -803
rect 171611 -921 189493 -803
rect 189611 -921 207493 -803
rect 207611 -921 225493 -803
rect 225611 -921 243493 -803
rect 243611 -921 261493 -803
rect 261611 -921 279493 -803
rect 279611 -921 293221 -803
rect 293339 -921 293430 -803
rect -1468 -932 293430 -921
rect -1468 -933 -1168 -932
rect 9402 -933 9702 -932
rect 27402 -933 27702 -932
rect 45402 -933 45702 -932
rect 63402 -933 63702 -932
rect 81402 -933 81702 -932
rect 99402 -933 99702 -932
rect 117402 -933 117702 -932
rect 135402 -933 135702 -932
rect 153402 -933 153702 -932
rect 171402 -933 171702 -932
rect 189402 -933 189702 -932
rect 207402 -933 207702 -932
rect 225402 -933 225702 -932
rect 243402 -933 243702 -932
rect 261402 -933 261702 -932
rect 279402 -933 279702 -932
rect 293130 -933 293430 -932
rect -1938 -1102 -1638 -1101
rect 2202 -1102 2502 -1101
rect 20202 -1102 20502 -1101
rect 38202 -1102 38502 -1101
rect 56202 -1102 56502 -1101
rect 74202 -1102 74502 -1101
rect 92202 -1102 92502 -1101
rect 110202 -1102 110502 -1101
rect 128202 -1102 128502 -1101
rect 146202 -1102 146502 -1101
rect 164202 -1102 164502 -1101
rect 182202 -1102 182502 -1101
rect 200202 -1102 200502 -1101
rect 218202 -1102 218502 -1101
rect 236202 -1102 236502 -1101
rect 254202 -1102 254502 -1101
rect 272202 -1102 272502 -1101
rect 290202 -1102 290502 -1101
rect 293600 -1102 293900 -1101
rect -1938 -1113 293900 -1102
rect -1938 -1231 -1847 -1113
rect -1729 -1231 2293 -1113
rect 2411 -1231 20293 -1113
rect 20411 -1231 38293 -1113
rect 38411 -1231 56293 -1113
rect 56411 -1231 74293 -1113
rect 74411 -1231 92293 -1113
rect 92411 -1231 110293 -1113
rect 110411 -1231 128293 -1113
rect 128411 -1231 146293 -1113
rect 146411 -1231 164293 -1113
rect 164411 -1231 182293 -1113
rect 182411 -1231 200293 -1113
rect 200411 -1231 218293 -1113
rect 218411 -1231 236293 -1113
rect 236411 -1231 254293 -1113
rect 254411 -1231 272293 -1113
rect 272411 -1231 290293 -1113
rect 290411 -1231 293691 -1113
rect 293809 -1231 293900 -1113
rect -1938 -1273 293900 -1231
rect -1938 -1391 -1847 -1273
rect -1729 -1391 2293 -1273
rect 2411 -1391 20293 -1273
rect 20411 -1391 38293 -1273
rect 38411 -1391 56293 -1273
rect 56411 -1391 74293 -1273
rect 74411 -1391 92293 -1273
rect 92411 -1391 110293 -1273
rect 110411 -1391 128293 -1273
rect 128411 -1391 146293 -1273
rect 146411 -1391 164293 -1273
rect 164411 -1391 182293 -1273
rect 182411 -1391 200293 -1273
rect 200411 -1391 218293 -1273
rect 218411 -1391 236293 -1273
rect 236411 -1391 254293 -1273
rect 254411 -1391 272293 -1273
rect 272411 -1391 290293 -1273
rect 290411 -1391 293691 -1273
rect 293809 -1391 293900 -1273
rect -1938 -1402 293900 -1391
rect -1938 -1403 -1638 -1402
rect 2202 -1403 2502 -1402
rect 20202 -1403 20502 -1402
rect 38202 -1403 38502 -1402
rect 56202 -1403 56502 -1402
rect 74202 -1403 74502 -1402
rect 92202 -1403 92502 -1402
rect 110202 -1403 110502 -1402
rect 128202 -1403 128502 -1402
rect 146202 -1403 146502 -1402
rect 164202 -1403 164502 -1402
rect 182202 -1403 182502 -1402
rect 200202 -1403 200502 -1402
rect 218202 -1403 218502 -1402
rect 236202 -1403 236502 -1402
rect 254202 -1403 254502 -1402
rect 272202 -1403 272502 -1402
rect 290202 -1403 290502 -1402
rect 293600 -1403 293900 -1402
rect -2408 -1572 -2108 -1571
rect 11202 -1572 11502 -1571
rect 29202 -1572 29502 -1571
rect 47202 -1572 47502 -1571
rect 65202 -1572 65502 -1571
rect 83202 -1572 83502 -1571
rect 101202 -1572 101502 -1571
rect 119202 -1572 119502 -1571
rect 137202 -1572 137502 -1571
rect 155202 -1572 155502 -1571
rect 173202 -1572 173502 -1571
rect 191202 -1572 191502 -1571
rect 209202 -1572 209502 -1571
rect 227202 -1572 227502 -1571
rect 245202 -1572 245502 -1571
rect 263202 -1572 263502 -1571
rect 281202 -1572 281502 -1571
rect 294070 -1572 294370 -1571
rect -2408 -1583 294370 -1572
rect -2408 -1701 -2317 -1583
rect -2199 -1701 11293 -1583
rect 11411 -1701 29293 -1583
rect 29411 -1701 47293 -1583
rect 47411 -1701 65293 -1583
rect 65411 -1701 83293 -1583
rect 83411 -1701 101293 -1583
rect 101411 -1701 119293 -1583
rect 119411 -1701 137293 -1583
rect 137411 -1701 155293 -1583
rect 155411 -1701 173293 -1583
rect 173411 -1701 191293 -1583
rect 191411 -1701 209293 -1583
rect 209411 -1701 227293 -1583
rect 227411 -1701 245293 -1583
rect 245411 -1701 263293 -1583
rect 263411 -1701 281293 -1583
rect 281411 -1701 294161 -1583
rect 294279 -1701 294370 -1583
rect -2408 -1743 294370 -1701
rect -2408 -1861 -2317 -1743
rect -2199 -1861 11293 -1743
rect 11411 -1861 29293 -1743
rect 29411 -1861 47293 -1743
rect 47411 -1861 65293 -1743
rect 65411 -1861 83293 -1743
rect 83411 -1861 101293 -1743
rect 101411 -1861 119293 -1743
rect 119411 -1861 137293 -1743
rect 137411 -1861 155293 -1743
rect 155411 -1861 173293 -1743
rect 173411 -1861 191293 -1743
rect 191411 -1861 209293 -1743
rect 209411 -1861 227293 -1743
rect 227411 -1861 245293 -1743
rect 245411 -1861 263293 -1743
rect 263411 -1861 281293 -1743
rect 281411 -1861 294161 -1743
rect 294279 -1861 294370 -1743
rect -2408 -1872 294370 -1861
rect -2408 -1873 -2108 -1872
rect 11202 -1873 11502 -1872
rect 29202 -1873 29502 -1872
rect 47202 -1873 47502 -1872
rect 65202 -1873 65502 -1872
rect 83202 -1873 83502 -1872
rect 101202 -1873 101502 -1872
rect 119202 -1873 119502 -1872
rect 137202 -1873 137502 -1872
rect 155202 -1873 155502 -1872
rect 173202 -1873 173502 -1872
rect 191202 -1873 191502 -1872
rect 209202 -1873 209502 -1872
rect 227202 -1873 227502 -1872
rect 245202 -1873 245502 -1872
rect 263202 -1873 263502 -1872
rect 281202 -1873 281502 -1872
rect 294070 -1873 294370 -1872
rect -2878 -2042 -2578 -2041
rect 4002 -2042 4302 -2041
rect 22002 -2042 22302 -2041
rect 40002 -2042 40302 -2041
rect 58002 -2042 58302 -2041
rect 76002 -2042 76302 -2041
rect 94002 -2042 94302 -2041
rect 112002 -2042 112302 -2041
rect 130002 -2042 130302 -2041
rect 148002 -2042 148302 -2041
rect 166002 -2042 166302 -2041
rect 184002 -2042 184302 -2041
rect 202002 -2042 202302 -2041
rect 220002 -2042 220302 -2041
rect 238002 -2042 238302 -2041
rect 256002 -2042 256302 -2041
rect 274002 -2042 274302 -2041
rect 294540 -2042 294840 -2041
rect -2878 -2053 294840 -2042
rect -2878 -2171 -2787 -2053
rect -2669 -2171 4093 -2053
rect 4211 -2171 22093 -2053
rect 22211 -2171 40093 -2053
rect 40211 -2171 58093 -2053
rect 58211 -2171 76093 -2053
rect 76211 -2171 94093 -2053
rect 94211 -2171 112093 -2053
rect 112211 -2171 130093 -2053
rect 130211 -2171 148093 -2053
rect 148211 -2171 166093 -2053
rect 166211 -2171 184093 -2053
rect 184211 -2171 202093 -2053
rect 202211 -2171 220093 -2053
rect 220211 -2171 238093 -2053
rect 238211 -2171 256093 -2053
rect 256211 -2171 274093 -2053
rect 274211 -2171 294631 -2053
rect 294749 -2171 294840 -2053
rect -2878 -2213 294840 -2171
rect -2878 -2331 -2787 -2213
rect -2669 -2331 4093 -2213
rect 4211 -2331 22093 -2213
rect 22211 -2331 40093 -2213
rect 40211 -2331 58093 -2213
rect 58211 -2331 76093 -2213
rect 76211 -2331 94093 -2213
rect 94211 -2331 112093 -2213
rect 112211 -2331 130093 -2213
rect 130211 -2331 148093 -2213
rect 148211 -2331 166093 -2213
rect 166211 -2331 184093 -2213
rect 184211 -2331 202093 -2213
rect 202211 -2331 220093 -2213
rect 220211 -2331 238093 -2213
rect 238211 -2331 256093 -2213
rect 256211 -2331 274093 -2213
rect 274211 -2331 294631 -2213
rect 294749 -2331 294840 -2213
rect -2878 -2342 294840 -2331
rect -2878 -2343 -2578 -2342
rect 4002 -2343 4302 -2342
rect 22002 -2343 22302 -2342
rect 40002 -2343 40302 -2342
rect 58002 -2343 58302 -2342
rect 76002 -2343 76302 -2342
rect 94002 -2343 94302 -2342
rect 112002 -2343 112302 -2342
rect 130002 -2343 130302 -2342
rect 148002 -2343 148302 -2342
rect 166002 -2343 166302 -2342
rect 184002 -2343 184302 -2342
rect 202002 -2343 202302 -2342
rect 220002 -2343 220302 -2342
rect 238002 -2343 238302 -2342
rect 256002 -2343 256302 -2342
rect 274002 -2343 274302 -2342
rect 294540 -2343 294840 -2342
rect -3348 -2512 -3048 -2511
rect 13002 -2512 13302 -2511
rect 31002 -2512 31302 -2511
rect 49002 -2512 49302 -2511
rect 67002 -2512 67302 -2511
rect 85002 -2512 85302 -2511
rect 103002 -2512 103302 -2511
rect 121002 -2512 121302 -2511
rect 139002 -2512 139302 -2511
rect 157002 -2512 157302 -2511
rect 175002 -2512 175302 -2511
rect 193002 -2512 193302 -2511
rect 211002 -2512 211302 -2511
rect 229002 -2512 229302 -2511
rect 247002 -2512 247302 -2511
rect 265002 -2512 265302 -2511
rect 283002 -2512 283302 -2511
rect 295010 -2512 295310 -2511
rect -3348 -2523 295310 -2512
rect -3348 -2641 -3257 -2523
rect -3139 -2641 13093 -2523
rect 13211 -2641 31093 -2523
rect 31211 -2641 49093 -2523
rect 49211 -2641 67093 -2523
rect 67211 -2641 85093 -2523
rect 85211 -2641 103093 -2523
rect 103211 -2641 121093 -2523
rect 121211 -2641 139093 -2523
rect 139211 -2641 157093 -2523
rect 157211 -2641 175093 -2523
rect 175211 -2641 193093 -2523
rect 193211 -2641 211093 -2523
rect 211211 -2641 229093 -2523
rect 229211 -2641 247093 -2523
rect 247211 -2641 265093 -2523
rect 265211 -2641 283093 -2523
rect 283211 -2641 295101 -2523
rect 295219 -2641 295310 -2523
rect -3348 -2683 295310 -2641
rect -3348 -2801 -3257 -2683
rect -3139 -2801 13093 -2683
rect 13211 -2801 31093 -2683
rect 31211 -2801 49093 -2683
rect 49211 -2801 67093 -2683
rect 67211 -2801 85093 -2683
rect 85211 -2801 103093 -2683
rect 103211 -2801 121093 -2683
rect 121211 -2801 139093 -2683
rect 139211 -2801 157093 -2683
rect 157211 -2801 175093 -2683
rect 175211 -2801 193093 -2683
rect 193211 -2801 211093 -2683
rect 211211 -2801 229093 -2683
rect 229211 -2801 247093 -2683
rect 247211 -2801 265093 -2683
rect 265211 -2801 283093 -2683
rect 283211 -2801 295101 -2683
rect 295219 -2801 295310 -2683
rect -3348 -2812 295310 -2801
rect -3348 -2813 -3048 -2812
rect 13002 -2813 13302 -2812
rect 31002 -2813 31302 -2812
rect 49002 -2813 49302 -2812
rect 67002 -2813 67302 -2812
rect 85002 -2813 85302 -2812
rect 103002 -2813 103302 -2812
rect 121002 -2813 121302 -2812
rect 139002 -2813 139302 -2812
rect 157002 -2813 157302 -2812
rect 175002 -2813 175302 -2812
rect 193002 -2813 193302 -2812
rect 211002 -2813 211302 -2812
rect 229002 -2813 229302 -2812
rect 247002 -2813 247302 -2812
rect 265002 -2813 265302 -2812
rect 283002 -2813 283302 -2812
rect 295010 -2813 295310 -2812
rect -3818 -2982 -3518 -2981
rect 5802 -2982 6102 -2981
rect 23802 -2982 24102 -2981
rect 41802 -2982 42102 -2981
rect 59802 -2982 60102 -2981
rect 77802 -2982 78102 -2981
rect 95802 -2982 96102 -2981
rect 113802 -2982 114102 -2981
rect 131802 -2982 132102 -2981
rect 149802 -2982 150102 -2981
rect 167802 -2982 168102 -2981
rect 185802 -2982 186102 -2981
rect 203802 -2982 204102 -2981
rect 221802 -2982 222102 -2981
rect 239802 -2982 240102 -2981
rect 257802 -2982 258102 -2981
rect 275802 -2982 276102 -2981
rect 295480 -2982 295780 -2981
rect -3818 -2993 295780 -2982
rect -3818 -3111 -3727 -2993
rect -3609 -3111 5893 -2993
rect 6011 -3111 23893 -2993
rect 24011 -3111 41893 -2993
rect 42011 -3111 59893 -2993
rect 60011 -3111 77893 -2993
rect 78011 -3111 95893 -2993
rect 96011 -3111 113893 -2993
rect 114011 -3111 131893 -2993
rect 132011 -3111 149893 -2993
rect 150011 -3111 167893 -2993
rect 168011 -3111 185893 -2993
rect 186011 -3111 203893 -2993
rect 204011 -3111 221893 -2993
rect 222011 -3111 239893 -2993
rect 240011 -3111 257893 -2993
rect 258011 -3111 275893 -2993
rect 276011 -3111 295571 -2993
rect 295689 -3111 295780 -2993
rect -3818 -3153 295780 -3111
rect -3818 -3271 -3727 -3153
rect -3609 -3271 5893 -3153
rect 6011 -3271 23893 -3153
rect 24011 -3271 41893 -3153
rect 42011 -3271 59893 -3153
rect 60011 -3271 77893 -3153
rect 78011 -3271 95893 -3153
rect 96011 -3271 113893 -3153
rect 114011 -3271 131893 -3153
rect 132011 -3271 149893 -3153
rect 150011 -3271 167893 -3153
rect 168011 -3271 185893 -3153
rect 186011 -3271 203893 -3153
rect 204011 -3271 221893 -3153
rect 222011 -3271 239893 -3153
rect 240011 -3271 257893 -3153
rect 258011 -3271 275893 -3153
rect 276011 -3271 295571 -3153
rect 295689 -3271 295780 -3153
rect -3818 -3282 295780 -3271
rect -3818 -3283 -3518 -3282
rect 5802 -3283 6102 -3282
rect 23802 -3283 24102 -3282
rect 41802 -3283 42102 -3282
rect 59802 -3283 60102 -3282
rect 77802 -3283 78102 -3282
rect 95802 -3283 96102 -3282
rect 113802 -3283 114102 -3282
rect 131802 -3283 132102 -3282
rect 149802 -3283 150102 -3282
rect 167802 -3283 168102 -3282
rect 185802 -3283 186102 -3282
rect 203802 -3283 204102 -3282
rect 221802 -3283 222102 -3282
rect 239802 -3283 240102 -3282
rect 257802 -3283 258102 -3282
rect 275802 -3283 276102 -3282
rect 295480 -3283 295780 -3282
rect -4288 -3452 -3988 -3451
rect 14802 -3452 15102 -3451
rect 32802 -3452 33102 -3451
rect 50802 -3452 51102 -3451
rect 68802 -3452 69102 -3451
rect 86802 -3452 87102 -3451
rect 104802 -3452 105102 -3451
rect 122802 -3452 123102 -3451
rect 140802 -3452 141102 -3451
rect 158802 -3452 159102 -3451
rect 176802 -3452 177102 -3451
rect 194802 -3452 195102 -3451
rect 212802 -3452 213102 -3451
rect 230802 -3452 231102 -3451
rect 248802 -3452 249102 -3451
rect 266802 -3452 267102 -3451
rect 284802 -3452 285102 -3451
rect 295950 -3452 296250 -3451
rect -4288 -3463 296250 -3452
rect -4288 -3581 -4197 -3463
rect -4079 -3581 14893 -3463
rect 15011 -3581 32893 -3463
rect 33011 -3581 50893 -3463
rect 51011 -3581 68893 -3463
rect 69011 -3581 86893 -3463
rect 87011 -3581 104893 -3463
rect 105011 -3581 122893 -3463
rect 123011 -3581 140893 -3463
rect 141011 -3581 158893 -3463
rect 159011 -3581 176893 -3463
rect 177011 -3581 194893 -3463
rect 195011 -3581 212893 -3463
rect 213011 -3581 230893 -3463
rect 231011 -3581 248893 -3463
rect 249011 -3581 266893 -3463
rect 267011 -3581 284893 -3463
rect 285011 -3581 296041 -3463
rect 296159 -3581 296250 -3463
rect -4288 -3623 296250 -3581
rect -4288 -3741 -4197 -3623
rect -4079 -3741 14893 -3623
rect 15011 -3741 32893 -3623
rect 33011 -3741 50893 -3623
rect 51011 -3741 68893 -3623
rect 69011 -3741 86893 -3623
rect 87011 -3741 104893 -3623
rect 105011 -3741 122893 -3623
rect 123011 -3741 140893 -3623
rect 141011 -3741 158893 -3623
rect 159011 -3741 176893 -3623
rect 177011 -3741 194893 -3623
rect 195011 -3741 212893 -3623
rect 213011 -3741 230893 -3623
rect 231011 -3741 248893 -3623
rect 249011 -3741 266893 -3623
rect 267011 -3741 284893 -3623
rect 285011 -3741 296041 -3623
rect 296159 -3741 296250 -3623
rect -4288 -3752 296250 -3741
rect -4288 -3753 -3988 -3752
rect 14802 -3753 15102 -3752
rect 32802 -3753 33102 -3752
rect 50802 -3753 51102 -3752
rect 68802 -3753 69102 -3752
rect 86802 -3753 87102 -3752
rect 104802 -3753 105102 -3752
rect 122802 -3753 123102 -3752
rect 140802 -3753 141102 -3752
rect 158802 -3753 159102 -3752
rect 176802 -3753 177102 -3752
rect 194802 -3753 195102 -3752
rect 212802 -3753 213102 -3752
rect 230802 -3753 231102 -3752
rect 248802 -3753 249102 -3752
rect 266802 -3753 267102 -3752
rect 284802 -3753 285102 -3752
rect 295950 -3753 296250 -3752
<< labels >>
rlabel metal3 s 291760 2898 292480 3018 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 291760 237498 292480 237618 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 291760 260958 292480 261078 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 291760 284418 292480 284538 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 291760 307878 292480 307998 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 291760 331338 292480 331458 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 287909 351760 287965 352480 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 255479 351760 255535 352480 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 223049 351760 223105 352480 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 190573 351760 190629 352480 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 158143 351760 158199 352480 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 291760 26358 292480 26478 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 125713 351760 125769 352480 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 93237 351760 93293 352480 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 60807 351760 60863 352480 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 28377 351760 28433 352480 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -480 348270 240 348390 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -480 319506 240 319626 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -480 290810 240 290930 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -480 262046 240 262166 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -480 233350 240 233470 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -480 204586 240 204706 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 291760 49818 292480 49938 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -480 175890 240 176010 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 291760 73278 292480 73398 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 291760 96738 292480 96858 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 291760 120198 292480 120318 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 291760 143658 292480 143778 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 291760 167118 292480 167238 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 291760 190578 292480 190698 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 291760 214038 292480 214158 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 291760 8746 292480 8866 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 291760 243346 292480 243466 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 291760 266874 292480 266994 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 291760 290334 292480 290454 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 291760 313794 292480 313914 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 291760 337254 292480 337374 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 279813 351760 279869 352480 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 247383 351760 247439 352480 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 214907 351760 214963 352480 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 182477 351760 182533 352480 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 150047 351760 150103 352480 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 291760 32206 292480 32326 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 117571 351760 117627 352480 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 85141 351760 85197 352480 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 52711 351760 52767 352480 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 20235 351760 20291 352480 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -480 341062 240 341182 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -480 312366 240 312486 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -480 283602 240 283722 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -480 254906 240 255026 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -480 226142 240 226262 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -480 197446 240 197566 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 291760 55666 292480 55786 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -480 168682 240 168802 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -480 147126 240 147246 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -480 125570 240 125690 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -480 104014 240 104134 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -480 82458 240 82578 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -480 60970 240 61090 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -480 39414 240 39534 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -480 17858 240 17978 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 291760 79126 292480 79246 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 291760 102586 292480 102706 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 291760 126046 292480 126166 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 291760 149506 292480 149626 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 291760 172966 292480 173086 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 291760 196426 292480 196546 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 291760 219886 292480 220006 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 291760 20442 292480 20562 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 291760 255110 292480 255230 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 291760 278570 292480 278690 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 291760 302030 292480 302150 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 291760 325490 292480 325610 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 291760 348950 292480 349070 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 263575 351760 263631 352480 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 231145 351760 231201 352480 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 198715 351760 198771 352480 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 166239 351760 166295 352480 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 133809 351760 133865 352480 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 291760 43902 292480 44022 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 101379 351760 101435 352480 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 68903 351760 68959 352480 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 36473 351760 36529 352480 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 4043 351760 4099 352480 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -480 326714 240 326834 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -480 297950 240 298070 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -480 269254 240 269374 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -480 240490 240 240610 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -480 211794 240 211914 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -480 183030 240 183150 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 291760 67362 292480 67482 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -480 154334 240 154454 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -480 132778 240 132898 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -480 111222 240 111342 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -480 89666 240 89786 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -480 68110 240 68230 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -480 46554 240 46674 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -480 24998 240 25118 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -480 3510 240 3630 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 291760 90890 292480 91010 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 291760 114350 292480 114470 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 291760 137810 292480 137930 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 291760 161270 292480 161390 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 291760 184730 292480 184850 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 291760 208190 292480 208310 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 291760 231650 292480 231770 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 291760 14594 292480 14714 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 291760 249262 292480 249382 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 291760 272722 292480 272842 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 291760 296182 292480 296302 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 291760 319642 292480 319762 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 291760 343102 292480 343222 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 271717 351760 271773 352480 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 239241 351760 239297 352480 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 206811 351760 206867 352480 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 174381 351760 174437 352480 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 141905 351760 141961 352480 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 291760 38054 292480 38174 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 109475 351760 109531 352480 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 77045 351760 77101 352480 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 44569 351760 44625 352480 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 12139 351760 12195 352480 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -480 333922 240 334042 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -480 305158 240 305278 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -480 276462 240 276582 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -480 247698 240 247818 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -480 218934 240 219054 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -480 190238 240 190358 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 291760 61514 292480 61634 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -480 161474 240 161594 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -480 139986 240 140106 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -480 118430 240 118550 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -480 96874 240 96994 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -480 75318 240 75438 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -480 53762 240 53882 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -480 32206 240 32326 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -480 10650 240 10770 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 291760 84974 292480 85094 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 291760 108434 292480 108554 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 291760 131894 292480 132014 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 291760 155354 292480 155474 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 291760 178882 292480 179002 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 291760 202342 292480 202462 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 291760 225802 292480 225922 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 63291 -480 63347 240 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 241725 -480 241781 240 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 243473 -480 243529 240 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 245267 -480 245323 240 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 247061 -480 247117 240 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 248855 -480 248911 240 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 250603 -480 250659 240 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 252397 -480 252453 240 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 254191 -480 254247 240 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 255985 -480 256041 240 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 257779 -480 257835 240 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 81139 -480 81195 240 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 259527 -480 259583 240 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 261321 -480 261377 240 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 263115 -480 263171 240 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 264909 -480 264965 240 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 266703 -480 266759 240 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 268451 -480 268507 240 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 270245 -480 270301 240 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 272039 -480 272095 240 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 273833 -480 273889 240 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 275581 -480 275637 240 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 82933 -480 82989 240 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 277375 -480 277431 240 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 279169 -480 279225 240 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 280963 -480 281019 240 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 282757 -480 282813 240 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 284505 -480 284561 240 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 286299 -480 286355 240 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 288093 -480 288149 240 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 289887 -480 289943 240 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 84681 -480 84737 240 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 86475 -480 86531 240 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 88269 -480 88325 240 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 90063 -480 90119 240 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 91857 -480 91913 240 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 93605 -480 93661 240 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 95399 -480 95455 240 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 97193 -480 97249 240 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 65085 -480 65141 240 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 98987 -480 99043 240 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 100735 -480 100791 240 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 102529 -480 102585 240 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 104323 -480 104379 240 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 106117 -480 106173 240 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 107911 -480 107967 240 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 109659 -480 109715 240 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 111453 -480 111509 240 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 113247 -480 113303 240 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 115041 -480 115097 240 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 66879 -480 66935 240 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 116835 -480 116891 240 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 118583 -480 118639 240 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 120377 -480 120433 240 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 122171 -480 122227 240 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 123965 -480 124021 240 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 125713 -480 125769 240 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 127507 -480 127563 240 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 129301 -480 129357 240 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 131095 -480 131151 240 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 132889 -480 132945 240 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 68627 -480 68683 240 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 134637 -480 134693 240 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 136431 -480 136487 240 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 138225 -480 138281 240 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 140019 -480 140075 240 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 141813 -480 141869 240 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 143561 -480 143617 240 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 145355 -480 145411 240 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 147149 -480 147205 240 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 148943 -480 148999 240 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 150691 -480 150747 240 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 70421 -480 70477 240 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 152485 -480 152541 240 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 154279 -480 154335 240 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 156073 -480 156129 240 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 157867 -480 157923 240 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 159615 -480 159671 240 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 161409 -480 161465 240 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 163203 -480 163259 240 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 164997 -480 165053 240 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 166791 -480 166847 240 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 168539 -480 168595 240 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 72215 -480 72271 240 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 170333 -480 170389 240 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 172127 -480 172183 240 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 173921 -480 173977 240 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 175669 -480 175725 240 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 177463 -480 177519 240 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 179257 -480 179313 240 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 181051 -480 181107 240 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 182845 -480 182901 240 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 184593 -480 184649 240 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 186387 -480 186443 240 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 74009 -480 74065 240 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 188181 -480 188237 240 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 189975 -480 190031 240 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 191769 -480 191825 240 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 193517 -480 193573 240 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 195311 -480 195367 240 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 197105 -480 197161 240 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 198899 -480 198955 240 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 200647 -480 200703 240 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 202441 -480 202497 240 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 204235 -480 204291 240 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 75757 -480 75813 240 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 206029 -480 206085 240 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 207823 -480 207879 240 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 209571 -480 209627 240 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 211365 -480 211421 240 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 213159 -480 213215 240 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 214953 -480 215009 240 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 216747 -480 216803 240 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 218495 -480 218551 240 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 220289 -480 220345 240 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 222083 -480 222139 240 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 77551 -480 77607 240 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 223877 -480 223933 240 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 225625 -480 225681 240 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 227419 -480 227475 240 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 229213 -480 229269 240 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 231007 -480 231063 240 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 232801 -480 232857 240 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 234549 -480 234605 240 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 236343 -480 236399 240 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 238137 -480 238193 240 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 239931 -480 239987 240 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 79345 -480 79401 240 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 63889 -480 63945 240 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 242277 -480 242333 240 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 244071 -480 244127 240 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 245865 -480 245921 240 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 247659 -480 247715 240 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 249453 -480 249509 240 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 251201 -480 251257 240 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 252995 -480 253051 240 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 254789 -480 254845 240 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 256583 -480 256639 240 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 258377 -480 258433 240 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 81737 -480 81793 240 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 260125 -480 260181 240 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 261919 -480 261975 240 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 263713 -480 263769 240 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 265507 -480 265563 240 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 267255 -480 267311 240 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 269049 -480 269105 240 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 270843 -480 270899 240 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 272637 -480 272693 240 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 274431 -480 274487 240 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 276179 -480 276235 240 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 83531 -480 83587 240 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 277973 -480 278029 240 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 279767 -480 279823 240 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 281561 -480 281617 240 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 283355 -480 283411 240 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 285103 -480 285159 240 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 286897 -480 286953 240 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 288691 -480 288747 240 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 290485 -480 290541 240 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 85279 -480 85335 240 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 87073 -480 87129 240 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 88867 -480 88923 240 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 90661 -480 90717 240 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 92409 -480 92465 240 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 94203 -480 94259 240 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 95997 -480 96053 240 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 97791 -480 97847 240 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 65683 -480 65739 240 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 99585 -480 99641 240 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 101333 -480 101389 240 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 103127 -480 103183 240 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 104921 -480 104977 240 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 106715 -480 106771 240 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 108509 -480 108565 240 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 110257 -480 110313 240 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 112051 -480 112107 240 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 113845 -480 113901 240 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 115639 -480 115695 240 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 67431 -480 67487 240 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 117387 -480 117443 240 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 119181 -480 119237 240 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 120975 -480 121031 240 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 122769 -480 122825 240 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 124563 -480 124619 240 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 126311 -480 126367 240 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 128105 -480 128161 240 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 129899 -480 129955 240 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 131693 -480 131749 240 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 133487 -480 133543 240 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 69225 -480 69281 240 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 135235 -480 135291 240 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 137029 -480 137085 240 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 138823 -480 138879 240 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 140617 -480 140673 240 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 142365 -480 142421 240 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 144159 -480 144215 240 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 145953 -480 146009 240 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 147747 -480 147803 240 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 149541 -480 149597 240 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 151289 -480 151345 240 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 71019 -480 71075 240 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 153083 -480 153139 240 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 154877 -480 154933 240 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 156671 -480 156727 240 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 158465 -480 158521 240 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 160213 -480 160269 240 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 162007 -480 162063 240 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 163801 -480 163857 240 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 165595 -480 165651 240 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 167343 -480 167399 240 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 169137 -480 169193 240 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 72813 -480 72869 240 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 170931 -480 170987 240 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 172725 -480 172781 240 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 174519 -480 174575 240 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 176267 -480 176323 240 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 178061 -480 178117 240 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 179855 -480 179911 240 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 181649 -480 181705 240 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 183443 -480 183499 240 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 185191 -480 185247 240 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 186985 -480 187041 240 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 74607 -480 74663 240 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 188779 -480 188835 240 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 190573 -480 190629 240 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 192321 -480 192377 240 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 194115 -480 194171 240 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 195909 -480 195965 240 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 197703 -480 197759 240 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 199497 -480 199553 240 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 201245 -480 201301 240 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 203039 -480 203095 240 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 204833 -480 204889 240 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 76355 -480 76411 240 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 206627 -480 206683 240 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 208421 -480 208477 240 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 210169 -480 210225 240 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 211963 -480 212019 240 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 213757 -480 213813 240 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 215551 -480 215607 240 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 217299 -480 217355 240 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 219093 -480 219149 240 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 220887 -480 220943 240 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 222681 -480 222737 240 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 78149 -480 78205 240 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 224475 -480 224531 240 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 226223 -480 226279 240 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 228017 -480 228073 240 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 229811 -480 229867 240 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 231605 -480 231661 240 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 233399 -480 233455 240 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 235147 -480 235203 240 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 236941 -480 236997 240 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 238735 -480 238791 240 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 240529 -480 240585 240 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 79943 -480 79999 240 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 64487 -480 64543 240 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 242875 -480 242931 240 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 244669 -480 244725 240 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 246463 -480 246519 240 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 248257 -480 248313 240 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 250051 -480 250107 240 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 251799 -480 251855 240 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 253593 -480 253649 240 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 255387 -480 255443 240 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 257181 -480 257237 240 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 258929 -480 258985 240 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 82335 -480 82391 240 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 260723 -480 260779 240 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 262517 -480 262573 240 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 264311 -480 264367 240 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 266105 -480 266161 240 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 267853 -480 267909 240 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 269647 -480 269703 240 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 271441 -480 271497 240 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 273235 -480 273291 240 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 275029 -480 275085 240 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 276777 -480 276833 240 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 84083 -480 84139 240 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 278571 -480 278627 240 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 280365 -480 280421 240 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 282159 -480 282215 240 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 283907 -480 283963 240 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 285701 -480 285757 240 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 287495 -480 287551 240 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 289289 -480 289345 240 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 291083 -480 291139 240 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 85877 -480 85933 240 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 87671 -480 87727 240 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 89465 -480 89521 240 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 91259 -480 91315 240 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 93007 -480 93063 240 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 94801 -480 94857 240 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 96595 -480 96651 240 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 98389 -480 98445 240 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 66281 -480 66337 240 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 100183 -480 100239 240 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 101931 -480 101987 240 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 103725 -480 103781 240 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 105519 -480 105575 240 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 107313 -480 107369 240 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 109061 -480 109117 240 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 110855 -480 110911 240 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 112649 -480 112705 240 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 114443 -480 114499 240 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 116237 -480 116293 240 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 68029 -480 68085 240 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 117985 -480 118041 240 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 119779 -480 119835 240 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 121573 -480 121629 240 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 123367 -480 123423 240 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 125161 -480 125217 240 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 126909 -480 126965 240 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 128703 -480 128759 240 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 130497 -480 130553 240 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 132291 -480 132347 240 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 134039 -480 134095 240 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 69823 -480 69879 240 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 135833 -480 135889 240 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 137627 -480 137683 240 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 139421 -480 139477 240 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 141215 -480 141271 240 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 142963 -480 143019 240 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 144757 -480 144813 240 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 146551 -480 146607 240 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 148345 -480 148401 240 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 150139 -480 150195 240 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 151887 -480 151943 240 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 71617 -480 71673 240 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 153681 -480 153737 240 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 155475 -480 155531 240 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 157269 -480 157325 240 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 159017 -480 159073 240 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 160811 -480 160867 240 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 162605 -480 162661 240 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 164399 -480 164455 240 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 166193 -480 166249 240 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 167941 -480 167997 240 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 169735 -480 169791 240 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 73411 -480 73467 240 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 171529 -480 171585 240 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 173323 -480 173379 240 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 175117 -480 175173 240 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 176865 -480 176921 240 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 178659 -480 178715 240 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 180453 -480 180509 240 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 182247 -480 182303 240 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 183995 -480 184051 240 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 185789 -480 185845 240 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 187583 -480 187639 240 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 75205 -480 75261 240 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 189377 -480 189433 240 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 191171 -480 191227 240 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 192919 -480 192975 240 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 194713 -480 194769 240 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 196507 -480 196563 240 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 198301 -480 198357 240 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 200095 -480 200151 240 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 201843 -480 201899 240 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 203637 -480 203693 240 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 205431 -480 205487 240 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 76953 -480 77009 240 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 207225 -480 207281 240 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 208973 -480 209029 240 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 210767 -480 210823 240 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 212561 -480 212617 240 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 214355 -480 214411 240 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 216149 -480 216205 240 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 217897 -480 217953 240 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 219691 -480 219747 240 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 221485 -480 221541 240 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 223279 -480 223335 240 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 78747 -480 78803 240 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 225073 -480 225129 240 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 226821 -480 226877 240 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 228615 -480 228671 240 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 230409 -480 230465 240 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 232203 -480 232259 240 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 233951 -480 234007 240 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 235745 -480 235801 240 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 237539 -480 237595 240 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 239333 -480 239389 240 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 241127 -480 241183 240 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 80541 -480 80597 240 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 291681 -480 291737 240 8 user_clock2
port 529 nsew default input
rlabel metal2 s 271 -480 327 240 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 823 -480 879 240 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 1421 -480 1477 240 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 3813 -480 3869 240 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 24053 -480 24109 240 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 25801 -480 25857 240 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 27595 -480 27651 240 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 29389 -480 29445 240 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 31183 -480 31239 240 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 32977 -480 33033 240 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 34725 -480 34781 240 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 36519 -480 36575 240 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 38313 -480 38369 240 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 40107 -480 40163 240 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 6205 -480 6261 240 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 41901 -480 41957 240 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 43649 -480 43705 240 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 45443 -480 45499 240 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 47237 -480 47293 240 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 49031 -480 49087 240 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 50779 -480 50835 240 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 52573 -480 52629 240 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 54367 -480 54423 240 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 56161 -480 56217 240 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 57955 -480 58011 240 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 8597 -480 8653 240 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 59703 -480 59759 240 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 61497 -480 61553 240 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 10943 -480 10999 240 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 13335 -480 13391 240 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 15129 -480 15185 240 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 16923 -480 16979 240 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 18671 -480 18727 240 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 20465 -480 20521 240 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 22259 -480 22315 240 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 2019 -480 2075 240 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 4411 -480 4467 240 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 24651 -480 24707 240 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 26399 -480 26455 240 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 28193 -480 28249 240 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 29987 -480 30043 240 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 31781 -480 31837 240 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 33575 -480 33631 240 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 35323 -480 35379 240 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 37117 -480 37173 240 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 38911 -480 38967 240 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 40705 -480 40761 240 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 6803 -480 6859 240 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 42453 -480 42509 240 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 44247 -480 44303 240 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 46041 -480 46097 240 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 47835 -480 47891 240 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 49629 -480 49685 240 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 51377 -480 51433 240 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 53171 -480 53227 240 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 54965 -480 55021 240 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 56759 -480 56815 240 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 58553 -480 58609 240 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 9149 -480 9205 240 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 60301 -480 60357 240 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 62095 -480 62151 240 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 11541 -480 11597 240 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 13933 -480 13989 240 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 15727 -480 15783 240 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 17475 -480 17531 240 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 19269 -480 19325 240 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 21063 -480 21119 240 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 22857 -480 22913 240 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 5009 -480 5065 240 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 25249 -480 25305 240 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 26997 -480 27053 240 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 28791 -480 28847 240 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 30585 -480 30641 240 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 32379 -480 32435 240 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 34127 -480 34183 240 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 35921 -480 35977 240 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 37715 -480 37771 240 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 39509 -480 39565 240 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 41303 -480 41359 240 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 7401 -480 7457 240 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 43051 -480 43107 240 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 44845 -480 44901 240 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 46639 -480 46695 240 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 48433 -480 48489 240 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 50227 -480 50283 240 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 51975 -480 52031 240 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 53769 -480 53825 240 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 55563 -480 55619 240 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 57357 -480 57413 240 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 59105 -480 59161 240 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 9747 -480 9803 240 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 60899 -480 60955 240 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 62693 -480 62749 240 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 12139 -480 12195 240 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 14531 -480 14587 240 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 16325 -480 16381 240 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 18073 -480 18129 240 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 19867 -480 19923 240 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 21661 -480 21717 240 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 23455 -480 23511 240 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 5607 -480 5663 240 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 7999 -480 8055 240 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 10345 -480 10401 240 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 12737 -480 12793 240 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 2617 -480 2673 240 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 3215 -480 3271 240 8 wbs_we_i
port 635 nsew default input
rlabel metal4 s 288402 351760 288702 352900 6 vccd1
port 636 nsew default input
rlabel metal4 s 270402 351760 270702 352900 6 vccd1
port 637 nsew default input
rlabel metal4 s 252402 351760 252702 352900 6 vccd1
port 638 nsew default input
rlabel metal4 s 234402 351760 234702 352900 6 vccd1
port 639 nsew default input
rlabel metal4 s 216402 351760 216702 352900 6 vccd1
port 640 nsew default input
rlabel metal4 s 198402 351760 198702 352900 6 vccd1
port 641 nsew default input
rlabel metal4 s 180402 351760 180702 352900 6 vccd1
port 642 nsew default input
rlabel metal4 s 162402 351760 162702 352900 6 vccd1
port 643 nsew default input
rlabel metal4 s 144402 351760 144702 352900 6 vccd1
port 644 nsew default input
rlabel metal4 s 126402 351760 126702 352900 6 vccd1
port 645 nsew default input
rlabel metal4 s 108402 351760 108702 352900 6 vccd1
port 646 nsew default input
rlabel metal4 s 90402 351760 90702 352900 6 vccd1
port 647 nsew default input
rlabel metal4 s 72402 351760 72702 352900 6 vccd1
port 648 nsew default input
rlabel metal4 s 54402 351760 54702 352900 6 vccd1
port 649 nsew default input
rlabel metal4 s 36402 351760 36702 352900 6 vccd1
port 650 nsew default input
rlabel metal4 s 18402 351760 18702 352900 6 vccd1
port 651 nsew default input
rlabel metal4 s 402 351760 702 352900 6 vccd1
port 652 nsew default input
rlabel metal4 s 292660 -462 292960 352430 6 vccd1
port 653 nsew default input
rlabel metal4 s -998 -462 -698 352430 4 vccd1
port 654 nsew default input
rlabel metal4 s 288402 -932 288702 240 8 vccd1
port 655 nsew default input
rlabel metal4 s 270402 -932 270702 240 8 vccd1
port 656 nsew default input
rlabel metal4 s 252402 -932 252702 240 8 vccd1
port 657 nsew default input
rlabel metal4 s 234402 -932 234702 240 8 vccd1
port 658 nsew default input
rlabel metal4 s 216402 -932 216702 240 8 vccd1
port 659 nsew default input
rlabel metal4 s 198402 -932 198702 240 8 vccd1
port 660 nsew default input
rlabel metal4 s 180402 -932 180702 240 8 vccd1
port 661 nsew default input
rlabel metal4 s 162402 -932 162702 240 8 vccd1
port 662 nsew default input
rlabel metal4 s 144402 -932 144702 240 8 vccd1
port 663 nsew default input
rlabel metal4 s 126402 -932 126702 240 8 vccd1
port 664 nsew default input
rlabel metal4 s 108402 -932 108702 240 8 vccd1
port 665 nsew default input
rlabel metal4 s 90402 -932 90702 240 8 vccd1
port 666 nsew default input
rlabel metal4 s 72402 -932 72702 240 8 vccd1
port 667 nsew default input
rlabel metal4 s 54402 -932 54702 240 8 vccd1
port 668 nsew default input
rlabel metal4 s 36402 -932 36702 240 8 vccd1
port 669 nsew default input
rlabel metal4 s 18402 -932 18702 240 8 vccd1
port 670 nsew default input
rlabel metal4 s 402 -932 702 240 8 vccd1
port 671 nsew default input
rlabel metal5 s -998 352130 292960 352430 6 vccd1
port 672 nsew default input
rlabel metal5 s 291760 342938 293430 343238 6 vccd1
port 673 nsew default input
rlabel metal5 s -1468 342938 240 343238 4 vccd1
port 674 nsew default input
rlabel metal5 s 291760 324938 293430 325238 6 vccd1
port 675 nsew default input
rlabel metal5 s -1468 324938 240 325238 4 vccd1
port 676 nsew default input
rlabel metal5 s 291760 306938 293430 307238 6 vccd1
port 677 nsew default input
rlabel metal5 s -1468 306938 240 307238 4 vccd1
port 678 nsew default input
rlabel metal5 s 291760 288938 293430 289238 6 vccd1
port 679 nsew default input
rlabel metal5 s -1468 288938 240 289238 4 vccd1
port 680 nsew default input
rlabel metal5 s 291760 270938 293430 271238 6 vccd1
port 681 nsew default input
rlabel metal5 s -1468 270938 240 271238 4 vccd1
port 682 nsew default input
rlabel metal5 s 291760 252938 293430 253238 6 vccd1
port 683 nsew default input
rlabel metal5 s -1468 252938 240 253238 4 vccd1
port 684 nsew default input
rlabel metal5 s 291760 234938 293430 235238 6 vccd1
port 685 nsew default input
rlabel metal5 s -1468 234938 240 235238 4 vccd1
port 686 nsew default input
rlabel metal5 s 291760 216938 293430 217238 6 vccd1
port 687 nsew default input
rlabel metal5 s -1468 216938 240 217238 4 vccd1
port 688 nsew default input
rlabel metal5 s 291760 198938 293430 199238 6 vccd1
port 689 nsew default input
rlabel metal5 s -1468 198938 240 199238 4 vccd1
port 690 nsew default input
rlabel metal5 s 291760 180938 293430 181238 6 vccd1
port 691 nsew default input
rlabel metal5 s -1468 180938 240 181238 4 vccd1
port 692 nsew default input
rlabel metal5 s 291760 162938 293430 163238 6 vccd1
port 693 nsew default input
rlabel metal5 s -1468 162938 240 163238 4 vccd1
port 694 nsew default input
rlabel metal5 s 291760 144938 293430 145238 6 vccd1
port 695 nsew default input
rlabel metal5 s -1468 144938 240 145238 4 vccd1
port 696 nsew default input
rlabel metal5 s 291760 126938 293430 127238 6 vccd1
port 697 nsew default input
rlabel metal5 s -1468 126938 240 127238 4 vccd1
port 698 nsew default input
rlabel metal5 s 291760 108938 293430 109238 6 vccd1
port 699 nsew default input
rlabel metal5 s -1468 108938 240 109238 4 vccd1
port 700 nsew default input
rlabel metal5 s 291760 90938 293430 91238 6 vccd1
port 701 nsew default input
rlabel metal5 s -1468 90938 240 91238 4 vccd1
port 702 nsew default input
rlabel metal5 s 291760 72938 293430 73238 6 vccd1
port 703 nsew default input
rlabel metal5 s -1468 72938 240 73238 4 vccd1
port 704 nsew default input
rlabel metal5 s 291760 54938 293430 55238 6 vccd1
port 705 nsew default input
rlabel metal5 s -1468 54938 240 55238 4 vccd1
port 706 nsew default input
rlabel metal5 s 291760 36938 293430 37238 6 vccd1
port 707 nsew default input
rlabel metal5 s -1468 36938 240 37238 4 vccd1
port 708 nsew default input
rlabel metal5 s 291760 18938 293430 19238 6 vccd1
port 709 nsew default input
rlabel metal5 s -1468 18938 240 19238 4 vccd1
port 710 nsew default input
rlabel metal5 s 291760 938 293430 1238 6 vccd1
port 711 nsew default input
rlabel metal5 s -1468 938 240 1238 4 vccd1
port 712 nsew default input
rlabel metal5 s -998 -462 292960 -162 8 vccd1
port 713 nsew default input
rlabel metal4 s 293130 -932 293430 352900 6 vssd1
port 714 nsew default input
rlabel metal4 s 279402 351760 279702 352900 6 vssd1
port 715 nsew default input
rlabel metal4 s 261402 351760 261702 352900 6 vssd1
port 716 nsew default input
rlabel metal4 s 243402 351760 243702 352900 6 vssd1
port 717 nsew default input
rlabel metal4 s 225402 351760 225702 352900 6 vssd1
port 718 nsew default input
rlabel metal4 s 207402 351760 207702 352900 6 vssd1
port 719 nsew default input
rlabel metal4 s 189402 351760 189702 352900 6 vssd1
port 720 nsew default input
rlabel metal4 s 171402 351760 171702 352900 6 vssd1
port 721 nsew default input
rlabel metal4 s 153402 351760 153702 352900 6 vssd1
port 722 nsew default input
rlabel metal4 s 135402 351760 135702 352900 6 vssd1
port 723 nsew default input
rlabel metal4 s 117402 351760 117702 352900 6 vssd1
port 724 nsew default input
rlabel metal4 s 99402 351760 99702 352900 6 vssd1
port 725 nsew default input
rlabel metal4 s 81402 351760 81702 352900 6 vssd1
port 726 nsew default input
rlabel metal4 s 63402 351760 63702 352900 6 vssd1
port 727 nsew default input
rlabel metal4 s 45402 351760 45702 352900 6 vssd1
port 728 nsew default input
rlabel metal4 s 27402 351760 27702 352900 6 vssd1
port 729 nsew default input
rlabel metal4 s 9402 351760 9702 352900 6 vssd1
port 730 nsew default input
rlabel metal4 s -1468 -932 -1168 352900 4 vssd1
port 731 nsew default input
rlabel metal4 s 279402 -932 279702 240 8 vssd1
port 732 nsew default input
rlabel metal4 s 261402 -932 261702 240 8 vssd1
port 733 nsew default input
rlabel metal4 s 243402 -932 243702 240 8 vssd1
port 734 nsew default input
rlabel metal4 s 225402 -932 225702 240 8 vssd1
port 735 nsew default input
rlabel metal4 s 207402 -932 207702 240 8 vssd1
port 736 nsew default input
rlabel metal4 s 189402 -932 189702 240 8 vssd1
port 737 nsew default input
rlabel metal4 s 171402 -932 171702 240 8 vssd1
port 738 nsew default input
rlabel metal4 s 153402 -932 153702 240 8 vssd1
port 739 nsew default input
rlabel metal4 s 135402 -932 135702 240 8 vssd1
port 740 nsew default input
rlabel metal4 s 117402 -932 117702 240 8 vssd1
port 741 nsew default input
rlabel metal4 s 99402 -932 99702 240 8 vssd1
port 742 nsew default input
rlabel metal4 s 81402 -932 81702 240 8 vssd1
port 743 nsew default input
rlabel metal4 s 63402 -932 63702 240 8 vssd1
port 744 nsew default input
rlabel metal4 s 45402 -932 45702 240 8 vssd1
port 745 nsew default input
rlabel metal4 s 27402 -932 27702 240 8 vssd1
port 746 nsew default input
rlabel metal4 s 9402 -932 9702 240 8 vssd1
port 747 nsew default input
rlabel metal5 s -1468 352600 293430 352900 6 vssd1
port 748 nsew default input
rlabel metal5 s 291760 333938 293430 334238 6 vssd1
port 749 nsew default input
rlabel metal5 s -1468 333938 240 334238 4 vssd1
port 750 nsew default input
rlabel metal5 s 291760 315938 293430 316238 6 vssd1
port 751 nsew default input
rlabel metal5 s -1468 315938 240 316238 4 vssd1
port 752 nsew default input
rlabel metal5 s 291760 297938 293430 298238 6 vssd1
port 753 nsew default input
rlabel metal5 s -1468 297938 240 298238 4 vssd1
port 754 nsew default input
rlabel metal5 s 291760 279938 293430 280238 6 vssd1
port 755 nsew default input
rlabel metal5 s -1468 279938 240 280238 4 vssd1
port 756 nsew default input
rlabel metal5 s 291760 261938 293430 262238 6 vssd1
port 757 nsew default input
rlabel metal5 s -1468 261938 240 262238 4 vssd1
port 758 nsew default input
rlabel metal5 s 291760 243938 293430 244238 6 vssd1
port 759 nsew default input
rlabel metal5 s -1468 243938 240 244238 4 vssd1
port 760 nsew default input
rlabel metal5 s 291760 225938 293430 226238 6 vssd1
port 761 nsew default input
rlabel metal5 s -1468 225938 240 226238 4 vssd1
port 762 nsew default input
rlabel metal5 s 291760 207938 293430 208238 6 vssd1
port 763 nsew default input
rlabel metal5 s -1468 207938 240 208238 4 vssd1
port 764 nsew default input
rlabel metal5 s 291760 189938 293430 190238 6 vssd1
port 765 nsew default input
rlabel metal5 s -1468 189938 240 190238 4 vssd1
port 766 nsew default input
rlabel metal5 s 291760 171938 293430 172238 6 vssd1
port 767 nsew default input
rlabel metal5 s -1468 171938 240 172238 4 vssd1
port 768 nsew default input
rlabel metal5 s 291760 153938 293430 154238 6 vssd1
port 769 nsew default input
rlabel metal5 s -1468 153938 240 154238 4 vssd1
port 770 nsew default input
rlabel metal5 s 291760 135938 293430 136238 6 vssd1
port 771 nsew default input
rlabel metal5 s -1468 135938 240 136238 4 vssd1
port 772 nsew default input
rlabel metal5 s 291760 117938 293430 118238 6 vssd1
port 773 nsew default input
rlabel metal5 s -1468 117938 240 118238 4 vssd1
port 774 nsew default input
rlabel metal5 s 291760 99938 293430 100238 6 vssd1
port 775 nsew default input
rlabel metal5 s -1468 99938 240 100238 4 vssd1
port 776 nsew default input
rlabel metal5 s 291760 81938 293430 82238 6 vssd1
port 777 nsew default input
rlabel metal5 s -1468 81938 240 82238 4 vssd1
port 778 nsew default input
rlabel metal5 s 291760 63938 293430 64238 6 vssd1
port 779 nsew default input
rlabel metal5 s -1468 63938 240 64238 4 vssd1
port 780 nsew default input
rlabel metal5 s 291760 45938 293430 46238 6 vssd1
port 781 nsew default input
rlabel metal5 s -1468 45938 240 46238 4 vssd1
port 782 nsew default input
rlabel metal5 s 291760 27938 293430 28238 6 vssd1
port 783 nsew default input
rlabel metal5 s -1468 27938 240 28238 4 vssd1
port 784 nsew default input
rlabel metal5 s 291760 9938 293430 10238 6 vssd1
port 785 nsew default input
rlabel metal5 s -1468 9938 240 10238 4 vssd1
port 786 nsew default input
rlabel metal5 s -1468 -932 293430 -632 8 vssd1
port 787 nsew default input
rlabel metal4 s 290202 351760 290502 353840 6 vccd2
port 788 nsew default input
rlabel metal4 s 272202 351760 272502 353840 6 vccd2
port 789 nsew default input
rlabel metal4 s 254202 351760 254502 353840 6 vccd2
port 790 nsew default input
rlabel metal4 s 236202 351760 236502 353840 6 vccd2
port 791 nsew default input
rlabel metal4 s 218202 351760 218502 353840 6 vccd2
port 792 nsew default input
rlabel metal4 s 200202 351760 200502 353840 6 vccd2
port 793 nsew default input
rlabel metal4 s 182202 351760 182502 353840 6 vccd2
port 794 nsew default input
rlabel metal4 s 164202 351760 164502 353840 6 vccd2
port 795 nsew default input
rlabel metal4 s 146202 351760 146502 353840 6 vccd2
port 796 nsew default input
rlabel metal4 s 128202 351760 128502 353840 6 vccd2
port 797 nsew default input
rlabel metal4 s 110202 351760 110502 353840 6 vccd2
port 798 nsew default input
rlabel metal4 s 92202 351760 92502 353840 6 vccd2
port 799 nsew default input
rlabel metal4 s 74202 351760 74502 353840 6 vccd2
port 800 nsew default input
rlabel metal4 s 56202 351760 56502 353840 6 vccd2
port 801 nsew default input
rlabel metal4 s 38202 351760 38502 353840 6 vccd2
port 802 nsew default input
rlabel metal4 s 20202 351760 20502 353840 6 vccd2
port 803 nsew default input
rlabel metal4 s 2202 351760 2502 353840 6 vccd2
port 804 nsew default input
rlabel metal4 s 293600 -1402 293900 353370 6 vccd2
port 805 nsew default input
rlabel metal4 s -1938 -1402 -1638 353370 4 vccd2
port 806 nsew default input
rlabel metal4 s 290202 -1872 290502 240 8 vccd2
port 807 nsew default input
rlabel metal4 s 272202 -1872 272502 240 8 vccd2
port 808 nsew default input
rlabel metal4 s 254202 -1872 254502 240 8 vccd2
port 809 nsew default input
rlabel metal4 s 236202 -1872 236502 240 8 vccd2
port 810 nsew default input
rlabel metal4 s 218202 -1872 218502 240 8 vccd2
port 811 nsew default input
rlabel metal4 s 200202 -1872 200502 240 8 vccd2
port 812 nsew default input
rlabel metal4 s 182202 -1872 182502 240 8 vccd2
port 813 nsew default input
rlabel metal4 s 164202 -1872 164502 240 8 vccd2
port 814 nsew default input
rlabel metal4 s 146202 -1872 146502 240 8 vccd2
port 815 nsew default input
rlabel metal4 s 128202 -1872 128502 240 8 vccd2
port 816 nsew default input
rlabel metal4 s 110202 -1872 110502 240 8 vccd2
port 817 nsew default input
rlabel metal4 s 92202 -1872 92502 240 8 vccd2
port 818 nsew default input
rlabel metal4 s 74202 -1872 74502 240 8 vccd2
port 819 nsew default input
rlabel metal4 s 56202 -1872 56502 240 8 vccd2
port 820 nsew default input
rlabel metal4 s 38202 -1872 38502 240 8 vccd2
port 821 nsew default input
rlabel metal4 s 20202 -1872 20502 240 8 vccd2
port 822 nsew default input
rlabel metal4 s 2202 -1872 2502 240 8 vccd2
port 823 nsew default input
rlabel metal5 s -1938 353070 293900 353370 6 vccd2
port 824 nsew default input
rlabel metal5 s 291760 344738 294370 345038 6 vccd2
port 825 nsew default input
rlabel metal5 s -2408 344738 240 345038 4 vccd2
port 826 nsew default input
rlabel metal5 s 291760 326738 294370 327038 6 vccd2
port 827 nsew default input
rlabel metal5 s -2408 326738 240 327038 4 vccd2
port 828 nsew default input
rlabel metal5 s 291760 308738 294370 309038 6 vccd2
port 829 nsew default input
rlabel metal5 s -2408 308738 240 309038 4 vccd2
port 830 nsew default input
rlabel metal5 s 291760 290738 294370 291038 6 vccd2
port 831 nsew default input
rlabel metal5 s -2408 290738 240 291038 4 vccd2
port 832 nsew default input
rlabel metal5 s 291760 272738 294370 273038 6 vccd2
port 833 nsew default input
rlabel metal5 s -2408 272738 240 273038 4 vccd2
port 834 nsew default input
rlabel metal5 s 291760 254738 294370 255038 6 vccd2
port 835 nsew default input
rlabel metal5 s -2408 254738 240 255038 4 vccd2
port 836 nsew default input
rlabel metal5 s 291760 236738 294370 237038 6 vccd2
port 837 nsew default input
rlabel metal5 s -2408 236738 240 237038 4 vccd2
port 838 nsew default input
rlabel metal5 s 291760 218738 294370 219038 6 vccd2
port 839 nsew default input
rlabel metal5 s -2408 218738 240 219038 4 vccd2
port 840 nsew default input
rlabel metal5 s 291760 200738 294370 201038 6 vccd2
port 841 nsew default input
rlabel metal5 s -2408 200738 240 201038 4 vccd2
port 842 nsew default input
rlabel metal5 s 291760 182738 294370 183038 6 vccd2
port 843 nsew default input
rlabel metal5 s -2408 182738 240 183038 4 vccd2
port 844 nsew default input
rlabel metal5 s 291760 164738 294370 165038 6 vccd2
port 845 nsew default input
rlabel metal5 s -2408 164738 240 165038 4 vccd2
port 846 nsew default input
rlabel metal5 s 291760 146738 294370 147038 6 vccd2
port 847 nsew default input
rlabel metal5 s -2408 146738 240 147038 4 vccd2
port 848 nsew default input
rlabel metal5 s 291760 128738 294370 129038 6 vccd2
port 849 nsew default input
rlabel metal5 s -2408 128738 240 129038 4 vccd2
port 850 nsew default input
rlabel metal5 s 291760 110738 294370 111038 6 vccd2
port 851 nsew default input
rlabel metal5 s -2408 110738 240 111038 4 vccd2
port 852 nsew default input
rlabel metal5 s 291760 92738 294370 93038 6 vccd2
port 853 nsew default input
rlabel metal5 s -2408 92738 240 93038 4 vccd2
port 854 nsew default input
rlabel metal5 s 291760 74738 294370 75038 6 vccd2
port 855 nsew default input
rlabel metal5 s -2408 74738 240 75038 4 vccd2
port 856 nsew default input
rlabel metal5 s 291760 56738 294370 57038 6 vccd2
port 857 nsew default input
rlabel metal5 s -2408 56738 240 57038 4 vccd2
port 858 nsew default input
rlabel metal5 s 291760 38738 294370 39038 6 vccd2
port 859 nsew default input
rlabel metal5 s -2408 38738 240 39038 4 vccd2
port 860 nsew default input
rlabel metal5 s 291760 20738 294370 21038 6 vccd2
port 861 nsew default input
rlabel metal5 s -2408 20738 240 21038 4 vccd2
port 862 nsew default input
rlabel metal5 s 291760 2738 294370 3038 6 vccd2
port 863 nsew default input
rlabel metal5 s -2408 2738 240 3038 4 vccd2
port 864 nsew default input
rlabel metal5 s -1938 -1402 293900 -1102 8 vccd2
port 865 nsew default input
rlabel metal4 s 294070 -1872 294370 353840 6 vssd2
port 866 nsew default input
rlabel metal4 s 281202 351760 281502 353840 6 vssd2
port 867 nsew default input
rlabel metal4 s 263202 351760 263502 353840 6 vssd2
port 868 nsew default input
rlabel metal4 s 245202 351760 245502 353840 6 vssd2
port 869 nsew default input
rlabel metal4 s 227202 351760 227502 353840 6 vssd2
port 870 nsew default input
rlabel metal4 s 209202 351760 209502 353840 6 vssd2
port 871 nsew default input
rlabel metal4 s 191202 351760 191502 353840 6 vssd2
port 872 nsew default input
rlabel metal4 s 173202 351760 173502 353840 6 vssd2
port 873 nsew default input
rlabel metal4 s 155202 351760 155502 353840 6 vssd2
port 874 nsew default input
rlabel metal4 s 137202 351760 137502 353840 6 vssd2
port 875 nsew default input
rlabel metal4 s 119202 351760 119502 353840 6 vssd2
port 876 nsew default input
rlabel metal4 s 101202 351760 101502 353840 6 vssd2
port 877 nsew default input
rlabel metal4 s 83202 351760 83502 353840 6 vssd2
port 878 nsew default input
rlabel metal4 s 65202 351760 65502 353840 6 vssd2
port 879 nsew default input
rlabel metal4 s 47202 351760 47502 353840 6 vssd2
port 880 nsew default input
rlabel metal4 s 29202 351760 29502 353840 6 vssd2
port 881 nsew default input
rlabel metal4 s 11202 351760 11502 353840 6 vssd2
port 882 nsew default input
rlabel metal4 s -2408 -1872 -2108 353840 4 vssd2
port 883 nsew default input
rlabel metal4 s 281202 -1872 281502 240 8 vssd2
port 884 nsew default input
rlabel metal4 s 263202 -1872 263502 240 8 vssd2
port 885 nsew default input
rlabel metal4 s 245202 -1872 245502 240 8 vssd2
port 886 nsew default input
rlabel metal4 s 227202 -1872 227502 240 8 vssd2
port 887 nsew default input
rlabel metal4 s 209202 -1872 209502 240 8 vssd2
port 888 nsew default input
rlabel metal4 s 191202 -1872 191502 240 8 vssd2
port 889 nsew default input
rlabel metal4 s 173202 -1872 173502 240 8 vssd2
port 890 nsew default input
rlabel metal4 s 155202 -1872 155502 240 8 vssd2
port 891 nsew default input
rlabel metal4 s 137202 -1872 137502 240 8 vssd2
port 892 nsew default input
rlabel metal4 s 119202 -1872 119502 240 8 vssd2
port 893 nsew default input
rlabel metal4 s 101202 -1872 101502 240 8 vssd2
port 894 nsew default input
rlabel metal4 s 83202 -1872 83502 240 8 vssd2
port 895 nsew default input
rlabel metal4 s 65202 -1872 65502 240 8 vssd2
port 896 nsew default input
rlabel metal4 s 47202 -1872 47502 240 8 vssd2
port 897 nsew default input
rlabel metal4 s 29202 -1872 29502 240 8 vssd2
port 898 nsew default input
rlabel metal4 s 11202 -1872 11502 240 8 vssd2
port 899 nsew default input
rlabel metal5 s -2408 353540 294370 353840 6 vssd2
port 900 nsew default input
rlabel metal5 s 291760 335738 294370 336038 6 vssd2
port 901 nsew default input
rlabel metal5 s -2408 335738 240 336038 4 vssd2
port 902 nsew default input
rlabel metal5 s 291760 317738 294370 318038 6 vssd2
port 903 nsew default input
rlabel metal5 s -2408 317738 240 318038 4 vssd2
port 904 nsew default input
rlabel metal5 s 291760 299738 294370 300038 6 vssd2
port 905 nsew default input
rlabel metal5 s -2408 299738 240 300038 4 vssd2
port 906 nsew default input
rlabel metal5 s 291760 281738 294370 282038 6 vssd2
port 907 nsew default input
rlabel metal5 s -2408 281738 240 282038 4 vssd2
port 908 nsew default input
rlabel metal5 s 291760 263738 294370 264038 6 vssd2
port 909 nsew default input
rlabel metal5 s -2408 263738 240 264038 4 vssd2
port 910 nsew default input
rlabel metal5 s 291760 245738 294370 246038 6 vssd2
port 911 nsew default input
rlabel metal5 s -2408 245738 240 246038 4 vssd2
port 912 nsew default input
rlabel metal5 s 291760 227738 294370 228038 6 vssd2
port 913 nsew default input
rlabel metal5 s -2408 227738 240 228038 4 vssd2
port 914 nsew default input
rlabel metal5 s 291760 209738 294370 210038 6 vssd2
port 915 nsew default input
rlabel metal5 s -2408 209738 240 210038 4 vssd2
port 916 nsew default input
rlabel metal5 s 291760 191738 294370 192038 6 vssd2
port 917 nsew default input
rlabel metal5 s -2408 191738 240 192038 4 vssd2
port 918 nsew default input
rlabel metal5 s 291760 173738 294370 174038 6 vssd2
port 919 nsew default input
rlabel metal5 s -2408 173738 240 174038 4 vssd2
port 920 nsew default input
rlabel metal5 s 291760 155738 294370 156038 6 vssd2
port 921 nsew default input
rlabel metal5 s -2408 155738 240 156038 4 vssd2
port 922 nsew default input
rlabel metal5 s 291760 137738 294370 138038 6 vssd2
port 923 nsew default input
rlabel metal5 s -2408 137738 240 138038 4 vssd2
port 924 nsew default input
rlabel metal5 s 291760 119738 294370 120038 6 vssd2
port 925 nsew default input
rlabel metal5 s -2408 119738 240 120038 4 vssd2
port 926 nsew default input
rlabel metal5 s 291760 101738 294370 102038 6 vssd2
port 927 nsew default input
rlabel metal5 s -2408 101738 240 102038 4 vssd2
port 928 nsew default input
rlabel metal5 s 291760 83738 294370 84038 6 vssd2
port 929 nsew default input
rlabel metal5 s -2408 83738 240 84038 4 vssd2
port 930 nsew default input
rlabel metal5 s 291760 65738 294370 66038 6 vssd2
port 931 nsew default input
rlabel metal5 s -2408 65738 240 66038 4 vssd2
port 932 nsew default input
rlabel metal5 s 291760 47738 294370 48038 6 vssd2
port 933 nsew default input
rlabel metal5 s -2408 47738 240 48038 4 vssd2
port 934 nsew default input
rlabel metal5 s 291760 29738 294370 30038 6 vssd2
port 935 nsew default input
rlabel metal5 s -2408 29738 240 30038 4 vssd2
port 936 nsew default input
rlabel metal5 s 291760 11738 294370 12038 6 vssd2
port 937 nsew default input
rlabel metal5 s -2408 11738 240 12038 4 vssd2
port 938 nsew default input
rlabel metal5 s -2408 -1872 294370 -1572 8 vssd2
port 939 nsew default input
rlabel metal4 s 274002 351760 274302 354780 6 vdda1
port 940 nsew default input
rlabel metal4 s 256002 351760 256302 354780 6 vdda1
port 941 nsew default input
rlabel metal4 s 238002 351760 238302 354780 6 vdda1
port 942 nsew default input
rlabel metal4 s 220002 351760 220302 354780 6 vdda1
port 943 nsew default input
rlabel metal4 s 202002 351760 202302 354780 6 vdda1
port 944 nsew default input
rlabel metal4 s 184002 351760 184302 354780 6 vdda1
port 945 nsew default input
rlabel metal4 s 166002 351760 166302 354780 6 vdda1
port 946 nsew default input
rlabel metal4 s 148002 351760 148302 354780 6 vdda1
port 947 nsew default input
rlabel metal4 s 130002 351760 130302 354780 6 vdda1
port 948 nsew default input
rlabel metal4 s 112002 351760 112302 354780 6 vdda1
port 949 nsew default input
rlabel metal4 s 94002 351760 94302 354780 6 vdda1
port 950 nsew default input
rlabel metal4 s 76002 351760 76302 354780 6 vdda1
port 951 nsew default input
rlabel metal4 s 58002 351760 58302 354780 6 vdda1
port 952 nsew default input
rlabel metal4 s 40002 351760 40302 354780 6 vdda1
port 953 nsew default input
rlabel metal4 s 22002 351760 22302 354780 6 vdda1
port 954 nsew default input
rlabel metal4 s 4002 351760 4302 354780 6 vdda1
port 955 nsew default input
rlabel metal4 s 294540 -2342 294840 354310 6 vdda1
port 956 nsew default input
rlabel metal4 s -2878 -2342 -2578 354310 4 vdda1
port 957 nsew default input
rlabel metal4 s 274002 -2812 274302 240 8 vdda1
port 958 nsew default input
rlabel metal4 s 256002 -2812 256302 240 8 vdda1
port 959 nsew default input
rlabel metal4 s 238002 -2812 238302 240 8 vdda1
port 960 nsew default input
rlabel metal4 s 220002 -2812 220302 240 8 vdda1
port 961 nsew default input
rlabel metal4 s 202002 -2812 202302 240 8 vdda1
port 962 nsew default input
rlabel metal4 s 184002 -2812 184302 240 8 vdda1
port 963 nsew default input
rlabel metal4 s 166002 -2812 166302 240 8 vdda1
port 964 nsew default input
rlabel metal4 s 148002 -2812 148302 240 8 vdda1
port 965 nsew default input
rlabel metal4 s 130002 -2812 130302 240 8 vdda1
port 966 nsew default input
rlabel metal4 s 112002 -2812 112302 240 8 vdda1
port 967 nsew default input
rlabel metal4 s 94002 -2812 94302 240 8 vdda1
port 968 nsew default input
rlabel metal4 s 76002 -2812 76302 240 8 vdda1
port 969 nsew default input
rlabel metal4 s 58002 -2812 58302 240 8 vdda1
port 970 nsew default input
rlabel metal4 s 40002 -2812 40302 240 8 vdda1
port 971 nsew default input
rlabel metal4 s 22002 -2812 22302 240 8 vdda1
port 972 nsew default input
rlabel metal4 s 4002 -2812 4302 240 8 vdda1
port 973 nsew default input
rlabel metal5 s -2878 354010 294840 354310 6 vdda1
port 974 nsew default input
rlabel metal5 s 291760 346538 295310 346838 6 vdda1
port 975 nsew default input
rlabel metal5 s -3348 346538 240 346838 4 vdda1
port 976 nsew default input
rlabel metal5 s 291760 328538 295310 328838 6 vdda1
port 977 nsew default input
rlabel metal5 s -3348 328538 240 328838 4 vdda1
port 978 nsew default input
rlabel metal5 s 291760 310538 295310 310838 6 vdda1
port 979 nsew default input
rlabel metal5 s -3348 310538 240 310838 4 vdda1
port 980 nsew default input
rlabel metal5 s 291760 292538 295310 292838 6 vdda1
port 981 nsew default input
rlabel metal5 s -3348 292538 240 292838 4 vdda1
port 982 nsew default input
rlabel metal5 s 291760 274538 295310 274838 6 vdda1
port 983 nsew default input
rlabel metal5 s -3348 274538 240 274838 4 vdda1
port 984 nsew default input
rlabel metal5 s 291760 256538 295310 256838 6 vdda1
port 985 nsew default input
rlabel metal5 s -3348 256538 240 256838 4 vdda1
port 986 nsew default input
rlabel metal5 s 291760 238538 295310 238838 6 vdda1
port 987 nsew default input
rlabel metal5 s -3348 238538 240 238838 4 vdda1
port 988 nsew default input
rlabel metal5 s 291760 220538 295310 220838 6 vdda1
port 989 nsew default input
rlabel metal5 s -3348 220538 240 220838 4 vdda1
port 990 nsew default input
rlabel metal5 s 291760 202538 295310 202838 6 vdda1
port 991 nsew default input
rlabel metal5 s -3348 202538 240 202838 4 vdda1
port 992 nsew default input
rlabel metal5 s 291760 184538 295310 184838 6 vdda1
port 993 nsew default input
rlabel metal5 s -3348 184538 240 184838 4 vdda1
port 994 nsew default input
rlabel metal5 s 291760 166538 295310 166838 6 vdda1
port 995 nsew default input
rlabel metal5 s -3348 166538 240 166838 4 vdda1
port 996 nsew default input
rlabel metal5 s 291760 148538 295310 148838 6 vdda1
port 997 nsew default input
rlabel metal5 s -3348 148538 240 148838 4 vdda1
port 998 nsew default input
rlabel metal5 s 291760 130538 295310 130838 6 vdda1
port 999 nsew default input
rlabel metal5 s -3348 130538 240 130838 4 vdda1
port 1000 nsew default input
rlabel metal5 s 291760 112538 295310 112838 6 vdda1
port 1001 nsew default input
rlabel metal5 s -3348 112538 240 112838 4 vdda1
port 1002 nsew default input
rlabel metal5 s 291760 94538 295310 94838 6 vdda1
port 1003 nsew default input
rlabel metal5 s -3348 94538 240 94838 4 vdda1
port 1004 nsew default input
rlabel metal5 s 291760 76538 295310 76838 6 vdda1
port 1005 nsew default input
rlabel metal5 s -3348 76538 240 76838 4 vdda1
port 1006 nsew default input
rlabel metal5 s 291760 58538 295310 58838 6 vdda1
port 1007 nsew default input
rlabel metal5 s -3348 58538 240 58838 4 vdda1
port 1008 nsew default input
rlabel metal5 s 291760 40538 295310 40838 6 vdda1
port 1009 nsew default input
rlabel metal5 s -3348 40538 240 40838 4 vdda1
port 1010 nsew default input
rlabel metal5 s 291760 22538 295310 22838 6 vdda1
port 1011 nsew default input
rlabel metal5 s -3348 22538 240 22838 4 vdda1
port 1012 nsew default input
rlabel metal5 s 291760 4538 295310 4838 6 vdda1
port 1013 nsew default input
rlabel metal5 s -3348 4538 240 4838 4 vdda1
port 1014 nsew default input
rlabel metal5 s -2878 -2342 294840 -2042 8 vdda1
port 1015 nsew default input
rlabel metal4 s 295010 -2812 295310 354780 6 vssa1
port 1016 nsew default input
rlabel metal4 s 283002 351760 283302 354780 6 vssa1
port 1017 nsew default input
rlabel metal4 s 265002 351760 265302 354780 6 vssa1
port 1018 nsew default input
rlabel metal4 s 247002 351760 247302 354780 6 vssa1
port 1019 nsew default input
rlabel metal4 s 229002 351760 229302 354780 6 vssa1
port 1020 nsew default input
rlabel metal4 s 211002 351760 211302 354780 6 vssa1
port 1021 nsew default input
rlabel metal4 s 193002 351760 193302 354780 6 vssa1
port 1022 nsew default input
rlabel metal4 s 175002 351760 175302 354780 6 vssa1
port 1023 nsew default input
rlabel metal4 s 157002 351760 157302 354780 6 vssa1
port 1024 nsew default input
rlabel metal4 s 139002 351760 139302 354780 6 vssa1
port 1025 nsew default input
rlabel metal4 s 121002 351760 121302 354780 6 vssa1
port 1026 nsew default input
rlabel metal4 s 103002 351760 103302 354780 6 vssa1
port 1027 nsew default input
rlabel metal4 s 85002 351760 85302 354780 6 vssa1
port 1028 nsew default input
rlabel metal4 s 67002 351760 67302 354780 6 vssa1
port 1029 nsew default input
rlabel metal4 s 49002 351760 49302 354780 6 vssa1
port 1030 nsew default input
rlabel metal4 s 31002 351760 31302 354780 6 vssa1
port 1031 nsew default input
rlabel metal4 s 13002 351760 13302 354780 6 vssa1
port 1032 nsew default input
rlabel metal4 s -3348 -2812 -3048 354780 4 vssa1
port 1033 nsew default input
rlabel metal4 s 283002 -2812 283302 240 8 vssa1
port 1034 nsew default input
rlabel metal4 s 265002 -2812 265302 240 8 vssa1
port 1035 nsew default input
rlabel metal4 s 247002 -2812 247302 240 8 vssa1
port 1036 nsew default input
rlabel metal4 s 229002 -2812 229302 240 8 vssa1
port 1037 nsew default input
rlabel metal4 s 211002 -2812 211302 240 8 vssa1
port 1038 nsew default input
rlabel metal4 s 193002 -2812 193302 240 8 vssa1
port 1039 nsew default input
rlabel metal4 s 175002 -2812 175302 240 8 vssa1
port 1040 nsew default input
rlabel metal4 s 157002 -2812 157302 240 8 vssa1
port 1041 nsew default input
rlabel metal4 s 139002 -2812 139302 240 8 vssa1
port 1042 nsew default input
rlabel metal4 s 121002 -2812 121302 240 8 vssa1
port 1043 nsew default input
rlabel metal4 s 103002 -2812 103302 240 8 vssa1
port 1044 nsew default input
rlabel metal4 s 85002 -2812 85302 240 8 vssa1
port 1045 nsew default input
rlabel metal4 s 67002 -2812 67302 240 8 vssa1
port 1046 nsew default input
rlabel metal4 s 49002 -2812 49302 240 8 vssa1
port 1047 nsew default input
rlabel metal4 s 31002 -2812 31302 240 8 vssa1
port 1048 nsew default input
rlabel metal4 s 13002 -2812 13302 240 8 vssa1
port 1049 nsew default input
rlabel metal5 s -3348 354480 295310 354780 6 vssa1
port 1050 nsew default input
rlabel metal5 s 291760 337538 295310 337838 6 vssa1
port 1051 nsew default input
rlabel metal5 s -3348 337538 240 337838 4 vssa1
port 1052 nsew default input
rlabel metal5 s 291760 319538 295310 319838 6 vssa1
port 1053 nsew default input
rlabel metal5 s -3348 319538 240 319838 4 vssa1
port 1054 nsew default input
rlabel metal5 s 291760 301538 295310 301838 6 vssa1
port 1055 nsew default input
rlabel metal5 s -3348 301538 240 301838 4 vssa1
port 1056 nsew default input
rlabel metal5 s 291760 283538 295310 283838 6 vssa1
port 1057 nsew default input
rlabel metal5 s -3348 283538 240 283838 4 vssa1
port 1058 nsew default input
rlabel metal5 s 291760 265538 295310 265838 6 vssa1
port 1059 nsew default input
rlabel metal5 s -3348 265538 240 265838 4 vssa1
port 1060 nsew default input
rlabel metal5 s 291760 247538 295310 247838 6 vssa1
port 1061 nsew default input
rlabel metal5 s -3348 247538 240 247838 4 vssa1
port 1062 nsew default input
rlabel metal5 s 291760 229538 295310 229838 6 vssa1
port 1063 nsew default input
rlabel metal5 s -3348 229538 240 229838 4 vssa1
port 1064 nsew default input
rlabel metal5 s 291760 211538 295310 211838 6 vssa1
port 1065 nsew default input
rlabel metal5 s -3348 211538 240 211838 4 vssa1
port 1066 nsew default input
rlabel metal5 s 291760 193538 295310 193838 6 vssa1
port 1067 nsew default input
rlabel metal5 s -3348 193538 240 193838 4 vssa1
port 1068 nsew default input
rlabel metal5 s 291760 175538 295310 175838 6 vssa1
port 1069 nsew default input
rlabel metal5 s -3348 175538 240 175838 4 vssa1
port 1070 nsew default input
rlabel metal5 s 291760 157538 295310 157838 6 vssa1
port 1071 nsew default input
rlabel metal5 s -3348 157538 240 157838 4 vssa1
port 1072 nsew default input
rlabel metal5 s 291760 139538 295310 139838 6 vssa1
port 1073 nsew default input
rlabel metal5 s -3348 139538 240 139838 4 vssa1
port 1074 nsew default input
rlabel metal5 s 291760 121538 295310 121838 6 vssa1
port 1075 nsew default input
rlabel metal5 s -3348 121538 240 121838 4 vssa1
port 1076 nsew default input
rlabel metal5 s 291760 103538 295310 103838 6 vssa1
port 1077 nsew default input
rlabel metal5 s -3348 103538 240 103838 4 vssa1
port 1078 nsew default input
rlabel metal5 s 291760 85538 295310 85838 6 vssa1
port 1079 nsew default input
rlabel metal5 s -3348 85538 240 85838 4 vssa1
port 1080 nsew default input
rlabel metal5 s 291760 67538 295310 67838 6 vssa1
port 1081 nsew default input
rlabel metal5 s -3348 67538 240 67838 4 vssa1
port 1082 nsew default input
rlabel metal5 s 291760 49538 295310 49838 6 vssa1
port 1083 nsew default input
rlabel metal5 s -3348 49538 240 49838 4 vssa1
port 1084 nsew default input
rlabel metal5 s 291760 31538 295310 31838 6 vssa1
port 1085 nsew default input
rlabel metal5 s -3348 31538 240 31838 4 vssa1
port 1086 nsew default input
rlabel metal5 s 291760 13538 295310 13838 6 vssa1
port 1087 nsew default input
rlabel metal5 s -3348 13538 240 13838 4 vssa1
port 1088 nsew default input
rlabel metal5 s -3348 -2812 295310 -2512 8 vssa1
port 1089 nsew default input
rlabel metal4 s 275802 351760 276102 355720 6 vdda2
port 1090 nsew default input
rlabel metal4 s 257802 351760 258102 355720 6 vdda2
port 1091 nsew default input
rlabel metal4 s 239802 351760 240102 355720 6 vdda2
port 1092 nsew default input
rlabel metal4 s 221802 351760 222102 355720 6 vdda2
port 1093 nsew default input
rlabel metal4 s 203802 351760 204102 355720 6 vdda2
port 1094 nsew default input
rlabel metal4 s 185802 351760 186102 355720 6 vdda2
port 1095 nsew default input
rlabel metal4 s 167802 351760 168102 355720 6 vdda2
port 1096 nsew default input
rlabel metal4 s 149802 351760 150102 355720 6 vdda2
port 1097 nsew default input
rlabel metal4 s 131802 351760 132102 355720 6 vdda2
port 1098 nsew default input
rlabel metal4 s 113802 351760 114102 355720 6 vdda2
port 1099 nsew default input
rlabel metal4 s 95802 351760 96102 355720 6 vdda2
port 1100 nsew default input
rlabel metal4 s 77802 351760 78102 355720 6 vdda2
port 1101 nsew default input
rlabel metal4 s 59802 351760 60102 355720 6 vdda2
port 1102 nsew default input
rlabel metal4 s 41802 351760 42102 355720 6 vdda2
port 1103 nsew default input
rlabel metal4 s 23802 351760 24102 355720 6 vdda2
port 1104 nsew default input
rlabel metal4 s 5802 351760 6102 355720 6 vdda2
port 1105 nsew default input
rlabel metal4 s 295480 -3282 295780 355250 6 vdda2
port 1106 nsew default input
rlabel metal4 s -3818 -3282 -3518 355250 4 vdda2
port 1107 nsew default input
rlabel metal4 s 275802 -3752 276102 240 8 vdda2
port 1108 nsew default input
rlabel metal4 s 257802 -3752 258102 240 8 vdda2
port 1109 nsew default input
rlabel metal4 s 239802 -3752 240102 240 8 vdda2
port 1110 nsew default input
rlabel metal4 s 221802 -3752 222102 240 8 vdda2
port 1111 nsew default input
rlabel metal4 s 203802 -3752 204102 240 8 vdda2
port 1112 nsew default input
rlabel metal4 s 185802 -3752 186102 240 8 vdda2
port 1113 nsew default input
rlabel metal4 s 167802 -3752 168102 240 8 vdda2
port 1114 nsew default input
rlabel metal4 s 149802 -3752 150102 240 8 vdda2
port 1115 nsew default input
rlabel metal4 s 131802 -3752 132102 240 8 vdda2
port 1116 nsew default input
rlabel metal4 s 113802 -3752 114102 240 8 vdda2
port 1117 nsew default input
rlabel metal4 s 95802 -3752 96102 240 8 vdda2
port 1118 nsew default input
rlabel metal4 s 77802 -3752 78102 240 8 vdda2
port 1119 nsew default input
rlabel metal4 s 59802 -3752 60102 240 8 vdda2
port 1120 nsew default input
rlabel metal4 s 41802 -3752 42102 240 8 vdda2
port 1121 nsew default input
rlabel metal4 s 23802 -3752 24102 240 8 vdda2
port 1122 nsew default input
rlabel metal4 s 5802 -3752 6102 240 8 vdda2
port 1123 nsew default input
rlabel metal5 s -3818 354950 295780 355250 6 vdda2
port 1124 nsew default input
rlabel metal5 s 291760 348338 296250 348638 6 vdda2
port 1125 nsew default input
rlabel metal5 s -4288 348338 240 348638 4 vdda2
port 1126 nsew default input
rlabel metal5 s 291760 330338 296250 330638 6 vdda2
port 1127 nsew default input
rlabel metal5 s -4288 330338 240 330638 4 vdda2
port 1128 nsew default input
rlabel metal5 s 291760 312338 296250 312638 6 vdda2
port 1129 nsew default input
rlabel metal5 s -4288 312338 240 312638 4 vdda2
port 1130 nsew default input
rlabel metal5 s 291760 294338 296250 294638 6 vdda2
port 1131 nsew default input
rlabel metal5 s -4288 294338 240 294638 4 vdda2
port 1132 nsew default input
rlabel metal5 s 291760 276338 296250 276638 6 vdda2
port 1133 nsew default input
rlabel metal5 s -4288 276338 240 276638 4 vdda2
port 1134 nsew default input
rlabel metal5 s 291760 258338 296250 258638 6 vdda2
port 1135 nsew default input
rlabel metal5 s -4288 258338 240 258638 4 vdda2
port 1136 nsew default input
rlabel metal5 s 291760 240338 296250 240638 6 vdda2
port 1137 nsew default input
rlabel metal5 s -4288 240338 240 240638 4 vdda2
port 1138 nsew default input
rlabel metal5 s 291760 222338 296250 222638 6 vdda2
port 1139 nsew default input
rlabel metal5 s -4288 222338 240 222638 4 vdda2
port 1140 nsew default input
rlabel metal5 s 291760 204338 296250 204638 6 vdda2
port 1141 nsew default input
rlabel metal5 s -4288 204338 240 204638 4 vdda2
port 1142 nsew default input
rlabel metal5 s 291760 186338 296250 186638 6 vdda2
port 1143 nsew default input
rlabel metal5 s -4288 186338 240 186638 4 vdda2
port 1144 nsew default input
rlabel metal5 s 291760 168338 296250 168638 6 vdda2
port 1145 nsew default input
rlabel metal5 s -4288 168338 240 168638 4 vdda2
port 1146 nsew default input
rlabel metal5 s 291760 150338 296250 150638 6 vdda2
port 1147 nsew default input
rlabel metal5 s -4288 150338 240 150638 4 vdda2
port 1148 nsew default input
rlabel metal5 s 291760 132338 296250 132638 6 vdda2
port 1149 nsew default input
rlabel metal5 s -4288 132338 240 132638 4 vdda2
port 1150 nsew default input
rlabel metal5 s 291760 114338 296250 114638 6 vdda2
port 1151 nsew default input
rlabel metal5 s -4288 114338 240 114638 4 vdda2
port 1152 nsew default input
rlabel metal5 s 291760 96338 296250 96638 6 vdda2
port 1153 nsew default input
rlabel metal5 s -4288 96338 240 96638 4 vdda2
port 1154 nsew default input
rlabel metal5 s 291760 78338 296250 78638 6 vdda2
port 1155 nsew default input
rlabel metal5 s -4288 78338 240 78638 4 vdda2
port 1156 nsew default input
rlabel metal5 s 291760 60338 296250 60638 6 vdda2
port 1157 nsew default input
rlabel metal5 s -4288 60338 240 60638 4 vdda2
port 1158 nsew default input
rlabel metal5 s 291760 42338 296250 42638 6 vdda2
port 1159 nsew default input
rlabel metal5 s -4288 42338 240 42638 4 vdda2
port 1160 nsew default input
rlabel metal5 s 291760 24338 296250 24638 6 vdda2
port 1161 nsew default input
rlabel metal5 s -4288 24338 240 24638 4 vdda2
port 1162 nsew default input
rlabel metal5 s 291760 6338 296250 6638 6 vdda2
port 1163 nsew default input
rlabel metal5 s -4288 6338 240 6638 4 vdda2
port 1164 nsew default input
rlabel metal5 s -3818 -3282 295780 -2982 8 vdda2
port 1165 nsew default input
rlabel metal4 s 295950 -3752 296250 355720 6 vssa2
port 1166 nsew default input
rlabel metal4 s 284802 351760 285102 355720 6 vssa2
port 1167 nsew default input
rlabel metal4 s 266802 351760 267102 355720 6 vssa2
port 1168 nsew default input
rlabel metal4 s 248802 351760 249102 355720 6 vssa2
port 1169 nsew default input
rlabel metal4 s 230802 351760 231102 355720 6 vssa2
port 1170 nsew default input
rlabel metal4 s 212802 351760 213102 355720 6 vssa2
port 1171 nsew default input
rlabel metal4 s 194802 351760 195102 355720 6 vssa2
port 1172 nsew default input
rlabel metal4 s 176802 351760 177102 355720 6 vssa2
port 1173 nsew default input
rlabel metal4 s 158802 351760 159102 355720 6 vssa2
port 1174 nsew default input
rlabel metal4 s 140802 351760 141102 355720 6 vssa2
port 1175 nsew default input
rlabel metal4 s 122802 351760 123102 355720 6 vssa2
port 1176 nsew default input
rlabel metal4 s 104802 351760 105102 355720 6 vssa2
port 1177 nsew default input
rlabel metal4 s 86802 351760 87102 355720 6 vssa2
port 1178 nsew default input
rlabel metal4 s 68802 351760 69102 355720 6 vssa2
port 1179 nsew default input
rlabel metal4 s 50802 351760 51102 355720 6 vssa2
port 1180 nsew default input
rlabel metal4 s 32802 351760 33102 355720 6 vssa2
port 1181 nsew default input
rlabel metal4 s 14802 351760 15102 355720 6 vssa2
port 1182 nsew default input
rlabel metal4 s -4288 -3752 -3988 355720 4 vssa2
port 1183 nsew default input
rlabel metal4 s 284802 -3752 285102 240 8 vssa2
port 1184 nsew default input
rlabel metal4 s 266802 -3752 267102 240 8 vssa2
port 1185 nsew default input
rlabel metal4 s 248802 -3752 249102 240 8 vssa2
port 1186 nsew default input
rlabel metal4 s 230802 -3752 231102 240 8 vssa2
port 1187 nsew default input
rlabel metal4 s 212802 -3752 213102 240 8 vssa2
port 1188 nsew default input
rlabel metal4 s 194802 -3752 195102 240 8 vssa2
port 1189 nsew default input
rlabel metal4 s 176802 -3752 177102 240 8 vssa2
port 1190 nsew default input
rlabel metal4 s 158802 -3752 159102 240 8 vssa2
port 1191 nsew default input
rlabel metal4 s 140802 -3752 141102 240 8 vssa2
port 1192 nsew default input
rlabel metal4 s 122802 -3752 123102 240 8 vssa2
port 1193 nsew default input
rlabel metal4 s 104802 -3752 105102 240 8 vssa2
port 1194 nsew default input
rlabel metal4 s 86802 -3752 87102 240 8 vssa2
port 1195 nsew default input
rlabel metal4 s 68802 -3752 69102 240 8 vssa2
port 1196 nsew default input
rlabel metal4 s 50802 -3752 51102 240 8 vssa2
port 1197 nsew default input
rlabel metal4 s 32802 -3752 33102 240 8 vssa2
port 1198 nsew default input
rlabel metal4 s 14802 -3752 15102 240 8 vssa2
port 1199 nsew default input
rlabel metal5 s -4288 355420 296250 355720 6 vssa2
port 1200 nsew default input
rlabel metal5 s 291760 339338 296250 339638 6 vssa2
port 1201 nsew default input
rlabel metal5 s -4288 339338 240 339638 4 vssa2
port 1202 nsew default input
rlabel metal5 s 291760 321338 296250 321638 6 vssa2
port 1203 nsew default input
rlabel metal5 s -4288 321338 240 321638 4 vssa2
port 1204 nsew default input
rlabel metal5 s 291760 303338 296250 303638 6 vssa2
port 1205 nsew default input
rlabel metal5 s -4288 303338 240 303638 4 vssa2
port 1206 nsew default input
rlabel metal5 s 291760 285338 296250 285638 6 vssa2
port 1207 nsew default input
rlabel metal5 s -4288 285338 240 285638 4 vssa2
port 1208 nsew default input
rlabel metal5 s 291760 267338 296250 267638 6 vssa2
port 1209 nsew default input
rlabel metal5 s -4288 267338 240 267638 4 vssa2
port 1210 nsew default input
rlabel metal5 s 291760 249338 296250 249638 6 vssa2
port 1211 nsew default input
rlabel metal5 s -4288 249338 240 249638 4 vssa2
port 1212 nsew default input
rlabel metal5 s 291760 231338 296250 231638 6 vssa2
port 1213 nsew default input
rlabel metal5 s -4288 231338 240 231638 4 vssa2
port 1214 nsew default input
rlabel metal5 s 291760 213338 296250 213638 6 vssa2
port 1215 nsew default input
rlabel metal5 s -4288 213338 240 213638 4 vssa2
port 1216 nsew default input
rlabel metal5 s 291760 195338 296250 195638 6 vssa2
port 1217 nsew default input
rlabel metal5 s -4288 195338 240 195638 4 vssa2
port 1218 nsew default input
rlabel metal5 s 291760 177338 296250 177638 6 vssa2
port 1219 nsew default input
rlabel metal5 s -4288 177338 240 177638 4 vssa2
port 1220 nsew default input
rlabel metal5 s 291760 159338 296250 159638 6 vssa2
port 1221 nsew default input
rlabel metal5 s -4288 159338 240 159638 4 vssa2
port 1222 nsew default input
rlabel metal5 s 291760 141338 296250 141638 6 vssa2
port 1223 nsew default input
rlabel metal5 s -4288 141338 240 141638 4 vssa2
port 1224 nsew default input
rlabel metal5 s 291760 123338 296250 123638 6 vssa2
port 1225 nsew default input
rlabel metal5 s -4288 123338 240 123638 4 vssa2
port 1226 nsew default input
rlabel metal5 s 291760 105338 296250 105638 6 vssa2
port 1227 nsew default input
rlabel metal5 s -4288 105338 240 105638 4 vssa2
port 1228 nsew default input
rlabel metal5 s 291760 87338 296250 87638 6 vssa2
port 1229 nsew default input
rlabel metal5 s -4288 87338 240 87638 4 vssa2
port 1230 nsew default input
rlabel metal5 s 291760 69338 296250 69638 6 vssa2
port 1231 nsew default input
rlabel metal5 s -4288 69338 240 69638 4 vssa2
port 1232 nsew default input
rlabel metal5 s 291760 51338 296250 51638 6 vssa2
port 1233 nsew default input
rlabel metal5 s -4288 51338 240 51638 4 vssa2
port 1234 nsew default input
rlabel metal5 s 291760 33338 296250 33638 6 vssa2
port 1235 nsew default input
rlabel metal5 s -4288 33338 240 33638 4 vssa2
port 1236 nsew default input
rlabel metal5 s 291760 15338 296250 15638 6 vssa2
port 1237 nsew default input
rlabel metal5 s -4288 15338 240 15638 4 vssa2
port 1238 nsew default input
rlabel metal5 s -4288 -3752 296250 -3452 8 vssa2
port 1239 nsew default input
<< properties >>
string FIXED_BBOX 0 0 292000 352000
string GDS_FILE ../gds/user_project_wrapper_empty.gds
string GDS_END 370014
string GDS_START 130
<< end >>
