VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2924.580 BY 3520.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2845.350 35.940 2845.670 36.000 ;
        RECT 2893.190 35.940 2893.510 36.000 ;
        RECT 2845.350 35.800 2893.510 35.940 ;
        RECT 2845.350 35.740 2845.670 35.800 ;
        RECT 2893.190 35.740 2893.510 35.800 ;
        RECT 2404.210 34.920 2404.530 34.980 ;
        RECT 2417.550 34.920 2417.870 34.980 ;
        RECT 2404.210 34.780 2417.870 34.920 ;
        RECT 2404.210 34.720 2404.530 34.780 ;
        RECT 2417.550 34.720 2417.870 34.780 ;
        RECT 2790.150 34.920 2790.470 34.980 ;
        RECT 2837.990 34.920 2838.310 34.980 ;
        RECT 2790.150 34.780 2838.310 34.920 ;
        RECT 2790.150 34.720 2790.470 34.780 ;
        RECT 2837.990 34.720 2838.310 34.780 ;
        RECT 2120.390 33.900 2120.710 33.960 ;
        RECT 2144.770 33.900 2145.090 33.960 ;
        RECT 2120.390 33.760 2145.090 33.900 ;
        RECT 2120.390 33.700 2120.710 33.760 ;
        RECT 2144.770 33.700 2145.090 33.760 ;
        RECT 2266.210 33.560 2266.530 33.620 ;
        RECT 2313.590 33.560 2313.910 33.620 ;
        RECT 2266.210 33.420 2313.910 33.560 ;
        RECT 2266.210 33.360 2266.530 33.420 ;
        RECT 2313.590 33.360 2313.910 33.420 ;
      LAYER via ;
        RECT 2845.380 35.740 2845.640 36.000 ;
        RECT 2893.220 35.740 2893.480 36.000 ;
        RECT 2404.240 34.720 2404.500 34.980 ;
        RECT 2417.580 34.720 2417.840 34.980 ;
        RECT 2790.180 34.720 2790.440 34.980 ;
        RECT 2838.020 34.720 2838.280 34.980 ;
        RECT 2120.420 33.700 2120.680 33.960 ;
        RECT 2144.800 33.700 2145.060 33.960 ;
        RECT 2266.240 33.360 2266.500 33.620 ;
        RECT 2313.620 33.360 2313.880 33.620 ;
      LAYER met2 ;
        RECT 1148.040 35.885 1148.180 54.000 ;
        RECT 2919.430 38.915 2919.710 39.285 ;
        RECT 1275.390 37.555 1275.670 37.925 ;
        RECT 2555.110 37.555 2555.390 37.925 ;
        RECT 1162.230 36.875 1162.510 37.245 ;
        RECT 1147.970 35.515 1148.250 35.885 ;
        RECT 1161.770 35.515 1162.050 35.885 ;
        RECT 1161.840 35.090 1161.980 35.515 ;
        RECT 1162.300 35.090 1162.440 36.875 ;
        RECT 1275.460 35.885 1275.600 37.555 ;
        RECT 2058.310 36.875 2058.590 37.245 ;
        RECT 2065.210 36.875 2065.490 37.245 ;
        RECT 2058.380 35.885 2058.520 36.875 ;
        RECT 1275.390 35.515 1275.670 35.885 ;
        RECT 1299.770 35.515 1300.050 35.885 ;
        RECT 2058.310 35.515 2058.590 35.885 ;
        RECT 1161.840 34.950 1162.440 35.090 ;
        RECT 1299.840 33.845 1299.980 35.515 ;
        RECT 2065.280 35.205 2065.420 36.875 ;
        RECT 2555.180 35.885 2555.320 37.555 ;
        RECT 2734.510 36.875 2734.790 37.245 ;
        RECT 2144.790 35.515 2145.070 35.885 ;
        RECT 2403.840 35.630 2404.440 35.770 ;
        RECT 1347.610 34.835 1347.890 35.205 ;
        RECT 1830.610 34.835 1830.890 35.205 ;
        RECT 1949.290 34.835 1949.570 35.205 ;
        RECT 2065.210 34.835 2065.490 35.205 ;
        RECT 2120.410 34.835 2120.690 35.205 ;
        RECT 1347.680 33.845 1347.820 34.835 ;
        RECT 1299.770 33.475 1300.050 33.845 ;
        RECT 1347.610 33.475 1347.890 33.845 ;
        RECT 1830.680 33.165 1830.820 34.835 ;
        RECT 1949.360 33.165 1949.500 34.835 ;
        RECT 2120.480 33.990 2120.620 34.835 ;
        RECT 2144.860 33.990 2145.000 35.515 ;
        RECT 2403.840 35.205 2403.980 35.630 ;
        RECT 2266.230 34.835 2266.510 35.205 ;
        RECT 2313.610 34.835 2313.890 35.205 ;
        RECT 2403.770 34.835 2404.050 35.205 ;
        RECT 2404.300 35.010 2404.440 35.630 ;
        RECT 2555.110 35.515 2555.390 35.885 ;
        RECT 2673.330 35.770 2673.610 35.885 ;
        RECT 2672.480 35.630 2673.610 35.770 ;
        RECT 2672.480 35.205 2672.620 35.630 ;
        RECT 2673.330 35.515 2673.610 35.630 ;
        RECT 2734.580 35.205 2734.720 36.875 ;
        RECT 2790.170 35.515 2790.450 35.885 ;
        RECT 2845.380 35.710 2845.640 36.030 ;
        RECT 2893.220 35.885 2893.480 36.030 ;
        RECT 2919.500 35.885 2919.640 38.915 ;
        RECT 2120.420 33.670 2120.680 33.990 ;
        RECT 2144.800 33.670 2145.060 33.990 ;
        RECT 2266.300 33.650 2266.440 34.835 ;
        RECT 2313.680 33.650 2313.820 34.835 ;
        RECT 2404.240 34.690 2404.500 35.010 ;
        RECT 2417.570 34.835 2417.850 35.205 ;
        RECT 2603.410 34.835 2603.690 35.205 ;
        RECT 2672.410 34.835 2672.690 35.205 ;
        RECT 2734.510 34.835 2734.790 35.205 ;
        RECT 2790.240 35.010 2790.380 35.515 ;
        RECT 2845.440 35.205 2845.580 35.710 ;
        RECT 2893.210 35.515 2893.490 35.885 ;
        RECT 2919.430 35.515 2919.710 35.885 ;
        RECT 2417.580 34.690 2417.840 34.835 ;
        RECT 2603.480 34.525 2603.620 34.835 ;
        RECT 2790.180 34.690 2790.440 35.010 ;
        RECT 2838.010 34.835 2838.290 35.205 ;
        RECT 2845.370 34.835 2845.650 35.205 ;
        RECT 2838.020 34.690 2838.280 34.835 ;
        RECT 2603.410 34.155 2603.690 34.525 ;
        RECT 2266.240 33.330 2266.500 33.650 ;
        RECT 2313.620 33.330 2313.880 33.650 ;
        RECT 1830.610 32.795 1830.890 33.165 ;
        RECT 1949.290 32.795 1949.570 33.165 ;
      LAYER via2 ;
        RECT 2919.430 38.960 2919.710 39.240 ;
        RECT 1275.390 37.600 1275.670 37.880 ;
        RECT 2555.110 37.600 2555.390 37.880 ;
        RECT 1162.230 36.920 1162.510 37.200 ;
        RECT 1147.970 35.560 1148.250 35.840 ;
        RECT 1161.770 35.560 1162.050 35.840 ;
        RECT 2058.310 36.920 2058.590 37.200 ;
        RECT 2065.210 36.920 2065.490 37.200 ;
        RECT 1275.390 35.560 1275.670 35.840 ;
        RECT 1299.770 35.560 1300.050 35.840 ;
        RECT 2058.310 35.560 2058.590 35.840 ;
        RECT 2734.510 36.920 2734.790 37.200 ;
        RECT 2144.790 35.560 2145.070 35.840 ;
        RECT 1347.610 34.880 1347.890 35.160 ;
        RECT 1830.610 34.880 1830.890 35.160 ;
        RECT 1949.290 34.880 1949.570 35.160 ;
        RECT 2065.210 34.880 2065.490 35.160 ;
        RECT 2120.410 34.880 2120.690 35.160 ;
        RECT 1299.770 33.520 1300.050 33.800 ;
        RECT 1347.610 33.520 1347.890 33.800 ;
        RECT 2266.230 34.880 2266.510 35.160 ;
        RECT 2313.610 34.880 2313.890 35.160 ;
        RECT 2403.770 34.880 2404.050 35.160 ;
        RECT 2555.110 35.560 2555.390 35.840 ;
        RECT 2673.330 35.560 2673.610 35.840 ;
        RECT 2790.170 35.560 2790.450 35.840 ;
        RECT 2417.570 34.880 2417.850 35.160 ;
        RECT 2603.410 34.880 2603.690 35.160 ;
        RECT 2672.410 34.880 2672.690 35.160 ;
        RECT 2734.510 34.880 2734.790 35.160 ;
        RECT 2893.210 35.560 2893.490 35.840 ;
        RECT 2919.430 35.560 2919.710 35.840 ;
        RECT 2838.010 34.880 2838.290 35.160 ;
        RECT 2845.370 34.880 2845.650 35.160 ;
        RECT 2603.410 34.200 2603.690 34.480 ;
        RECT 1830.610 32.840 1830.890 33.120 ;
        RECT 1949.290 32.840 1949.570 33.120 ;
      LAYER met3 ;
        RECT 2919.405 39.250 2919.735 39.265 ;
        RECT 2920.080 39.250 2922.480 39.400 ;
        RECT 2919.405 38.950 2922.480 39.250 ;
        RECT 2919.405 38.935 2919.735 38.950 ;
        RECT 2920.080 38.800 2922.480 38.950 ;
        RECT 1251.190 37.890 1251.570 37.900 ;
        RECT 1275.365 37.890 1275.695 37.905 ;
        RECT 1251.190 37.590 1275.695 37.890 ;
        RECT 1251.190 37.580 1251.570 37.590 ;
        RECT 1275.365 37.575 1275.695 37.590 ;
        RECT 2506.990 37.890 2507.370 37.900 ;
        RECT 2555.085 37.890 2555.415 37.905 ;
        RECT 2506.990 37.590 2555.415 37.890 ;
        RECT 2506.990 37.580 2507.370 37.590 ;
        RECT 2555.085 37.575 2555.415 37.590 ;
        RECT 1162.205 37.210 1162.535 37.225 ;
        RECT 1968.790 37.210 1969.170 37.220 ;
        RECT 2058.285 37.210 2058.615 37.225 ;
        RECT 2065.185 37.210 2065.515 37.225 ;
        RECT 1162.205 36.910 1210.130 37.210 ;
        RECT 1162.205 36.895 1162.535 36.910 ;
        RECT 1209.830 36.530 1210.130 36.910 ;
        RECT 1968.790 36.910 2016.050 37.210 ;
        RECT 1968.790 36.900 1969.170 36.910 ;
        RECT 1251.190 36.530 1251.570 36.540 ;
        RECT 1209.830 36.230 1251.570 36.530 ;
        RECT 1251.190 36.220 1251.570 36.230 ;
        RECT 1540.990 36.530 1541.370 36.540 ;
        RECT 1540.990 36.230 1589.170 36.530 ;
        RECT 1540.990 36.220 1541.370 36.230 ;
        RECT 1147.945 35.850 1148.275 35.865 ;
        RECT 1161.745 35.850 1162.075 35.865 ;
        RECT 1147.945 35.550 1162.075 35.850 ;
        RECT 1147.945 35.535 1148.275 35.550 ;
        RECT 1161.745 35.535 1162.075 35.550 ;
        RECT 1275.365 35.850 1275.695 35.865 ;
        RECT 1299.745 35.850 1300.075 35.865 ;
        RECT 1464.630 35.850 1465.010 35.860 ;
        RECT 1275.365 35.550 1300.075 35.850 ;
        RECT 1275.365 35.535 1275.695 35.550 ;
        RECT 1299.745 35.535 1300.075 35.550 ;
        RECT 1444.430 35.550 1465.010 35.850 ;
        RECT 1347.585 35.170 1347.915 35.185 ;
        RECT 1444.430 35.170 1444.730 35.550 ;
        RECT 1464.630 35.540 1465.010 35.550 ;
        RECT 1465.550 35.850 1465.930 35.860 ;
        RECT 1499.590 35.850 1499.970 35.860 ;
        RECT 1465.550 35.550 1499.970 35.850 ;
        RECT 1465.550 35.540 1465.930 35.550 ;
        RECT 1499.590 35.540 1499.970 35.550 ;
        RECT 1347.585 34.870 1444.730 35.170 ;
        RECT 1588.870 35.170 1589.170 36.230 ;
        RECT 1596.230 36.230 1644.600 36.530 ;
        RECT 1596.230 35.170 1596.530 36.230 ;
        RECT 1588.870 34.870 1596.530 35.170 ;
        RECT 1644.300 35.170 1644.600 36.230 ;
        RECT 1830.830 36.230 1878.970 36.530 ;
        RECT 1830.830 35.185 1831.130 36.230 ;
        RECT 1878.670 35.860 1878.970 36.230 ;
        RECT 1878.630 35.540 1879.010 35.860 ;
        RECT 2015.750 35.850 2016.050 36.910 ;
        RECT 2058.285 36.910 2065.515 37.210 ;
        RECT 2058.285 36.895 2058.615 36.910 ;
        RECT 2065.185 36.895 2065.515 36.910 ;
        RECT 2686.390 37.210 2686.770 37.220 ;
        RECT 2734.485 37.210 2734.815 37.225 ;
        RECT 2686.390 36.910 2734.815 37.210 ;
        RECT 2686.390 36.900 2686.770 36.910 ;
        RECT 2734.485 36.895 2734.815 36.910 ;
        RECT 2506.990 36.530 2507.370 36.540 ;
        RECT 2479.430 36.230 2507.370 36.530 ;
        RECT 2058.285 35.850 2058.615 35.865 ;
        RECT 2015.750 35.550 2058.615 35.850 ;
        RECT 2058.285 35.535 2058.615 35.550 ;
        RECT 2144.765 35.850 2145.095 35.865 ;
        RECT 2217.190 35.850 2217.570 35.860 ;
        RECT 2144.765 35.550 2217.570 35.850 ;
        RECT 2144.765 35.535 2145.095 35.550 ;
        RECT 2217.190 35.540 2217.570 35.550 ;
        RECT 1733.270 35.170 1733.650 35.180 ;
        RECT 1644.300 34.870 1733.650 35.170 ;
        RECT 1347.585 34.855 1347.915 34.870 ;
        RECT 1733.270 34.860 1733.650 34.870 ;
        RECT 1734.190 35.170 1734.570 35.180 ;
        RECT 1830.585 35.170 1831.130 35.185 ;
        RECT 1734.190 34.870 1782.370 35.170 ;
        RECT 1830.180 34.870 1831.130 35.170 ;
        RECT 1949.265 35.170 1949.595 35.185 ;
        RECT 1968.790 35.170 1969.170 35.180 ;
        RECT 1949.265 34.870 1969.170 35.170 ;
        RECT 1734.190 34.860 1734.570 34.870 ;
        RECT 1500.510 34.490 1500.890 34.500 ;
        RECT 1540.990 34.490 1541.370 34.500 ;
        RECT 1500.510 34.190 1541.370 34.490 ;
        RECT 1782.070 34.490 1782.370 34.870 ;
        RECT 1830.585 34.855 1830.915 34.870 ;
        RECT 1949.265 34.855 1949.595 34.870 ;
        RECT 1968.790 34.860 1969.170 34.870 ;
        RECT 2065.185 35.170 2065.515 35.185 ;
        RECT 2120.385 35.170 2120.715 35.185 ;
        RECT 2266.205 35.170 2266.535 35.185 ;
        RECT 2065.185 34.870 2120.715 35.170 ;
        RECT 2065.185 34.855 2065.515 34.870 ;
        RECT 2120.385 34.855 2120.715 34.870 ;
        RECT 2265.070 34.870 2266.535 35.170 ;
        RECT 1879.550 34.490 1879.930 34.500 ;
        RECT 1913.590 34.490 1913.970 34.500 ;
        RECT 1782.070 34.190 1783.290 34.490 ;
        RECT 1500.510 34.180 1500.890 34.190 ;
        RECT 1540.990 34.180 1541.370 34.190 ;
        RECT 1299.745 33.810 1300.075 33.825 ;
        RECT 1347.585 33.810 1347.915 33.825 ;
        RECT 1299.745 33.510 1347.915 33.810 ;
        RECT 1299.745 33.495 1300.075 33.510 ;
        RECT 1347.585 33.495 1347.915 33.510 ;
        RECT 1733.270 33.810 1733.650 33.820 ;
        RECT 1734.190 33.810 1734.570 33.820 ;
        RECT 1733.270 33.510 1734.570 33.810 ;
        RECT 1733.270 33.500 1733.650 33.510 ;
        RECT 1734.190 33.500 1734.570 33.510 ;
        RECT 1782.990 33.130 1783.290 34.190 ;
        RECT 1879.550 34.190 1913.970 34.490 ;
        RECT 1879.550 34.180 1879.930 34.190 ;
        RECT 1913.590 34.180 1913.970 34.190 ;
        RECT 2217.190 34.490 2217.570 34.500 ;
        RECT 2265.070 34.490 2265.370 34.870 ;
        RECT 2266.205 34.855 2266.535 34.870 ;
        RECT 2313.585 35.170 2313.915 35.185 ;
        RECT 2403.745 35.170 2404.075 35.185 ;
        RECT 2313.585 34.870 2404.075 35.170 ;
        RECT 2313.585 34.855 2313.915 34.870 ;
        RECT 2403.745 34.855 2404.075 34.870 ;
        RECT 2417.545 35.170 2417.875 35.185 ;
        RECT 2479.430 35.170 2479.730 36.230 ;
        RECT 2506.990 36.220 2507.370 36.230 ;
        RECT 2555.085 35.850 2555.415 35.865 ;
        RECT 2673.305 35.850 2673.635 35.865 ;
        RECT 2686.390 35.850 2686.770 35.860 ;
        RECT 2790.145 35.850 2790.475 35.865 ;
        RECT 2555.085 35.550 2556.090 35.850 ;
        RECT 2555.085 35.535 2555.415 35.550 ;
        RECT 2417.545 34.870 2479.730 35.170 ;
        RECT 2417.545 34.855 2417.875 34.870 ;
        RECT 2217.190 34.190 2265.370 34.490 ;
        RECT 2555.790 34.490 2556.090 35.550 ;
        RECT 2673.305 35.550 2686.770 35.850 ;
        RECT 2673.305 35.535 2673.635 35.550 ;
        RECT 2686.390 35.540 2686.770 35.550 ;
        RECT 2768.310 35.550 2790.475 35.850 ;
        RECT 2603.385 35.170 2603.715 35.185 ;
        RECT 2672.385 35.170 2672.715 35.185 ;
        RECT 2603.385 34.870 2672.715 35.170 ;
        RECT 2603.385 34.855 2603.715 34.870 ;
        RECT 2672.385 34.855 2672.715 34.870 ;
        RECT 2734.485 35.170 2734.815 35.185 ;
        RECT 2768.310 35.170 2768.610 35.550 ;
        RECT 2790.145 35.535 2790.475 35.550 ;
        RECT 2893.185 35.850 2893.515 35.865 ;
        RECT 2919.405 35.850 2919.735 35.865 ;
        RECT 2893.185 35.550 2919.735 35.850 ;
        RECT 2893.185 35.535 2893.515 35.550 ;
        RECT 2919.405 35.535 2919.735 35.550 ;
        RECT 2734.485 34.870 2768.610 35.170 ;
        RECT 2837.985 35.170 2838.315 35.185 ;
        RECT 2845.345 35.170 2845.675 35.185 ;
        RECT 2837.985 34.870 2845.675 35.170 ;
        RECT 2734.485 34.855 2734.815 34.870 ;
        RECT 2837.985 34.855 2838.315 34.870 ;
        RECT 2845.345 34.855 2845.675 34.870 ;
        RECT 2603.385 34.490 2603.715 34.505 ;
        RECT 2555.790 34.190 2603.715 34.490 ;
        RECT 2217.190 34.180 2217.570 34.190 ;
        RECT 2603.385 34.175 2603.715 34.190 ;
        RECT 1830.585 33.130 1830.915 33.145 ;
        RECT 1782.990 32.830 1830.915 33.130 ;
        RECT 1830.585 32.815 1830.915 32.830 ;
        RECT 1913.590 33.130 1913.970 33.140 ;
        RECT 1949.265 33.130 1949.595 33.145 ;
        RECT 1913.590 32.830 1949.595 33.130 ;
        RECT 1913.590 32.820 1913.970 32.830 ;
        RECT 1949.265 32.815 1949.595 32.830 ;
      LAYER via3 ;
        RECT 1251.220 37.580 1251.540 37.900 ;
        RECT 2507.020 37.580 2507.340 37.900 ;
        RECT 1968.820 36.900 1969.140 37.220 ;
        RECT 1251.220 36.220 1251.540 36.540 ;
        RECT 1541.020 36.220 1541.340 36.540 ;
        RECT 1464.660 35.540 1464.980 35.860 ;
        RECT 1465.580 35.540 1465.900 35.860 ;
        RECT 1499.620 35.540 1499.940 35.860 ;
        RECT 1878.660 35.540 1878.980 35.860 ;
        RECT 2686.420 36.900 2686.740 37.220 ;
        RECT 2217.220 35.540 2217.540 35.860 ;
        RECT 1733.300 34.860 1733.620 35.180 ;
        RECT 1734.220 34.860 1734.540 35.180 ;
        RECT 1500.540 34.180 1500.860 34.500 ;
        RECT 1541.020 34.180 1541.340 34.500 ;
        RECT 1968.820 34.860 1969.140 35.180 ;
        RECT 1733.300 33.500 1733.620 33.820 ;
        RECT 1734.220 33.500 1734.540 33.820 ;
        RECT 1879.580 34.180 1879.900 34.500 ;
        RECT 1913.620 34.180 1913.940 34.500 ;
        RECT 2217.220 34.180 2217.540 34.500 ;
        RECT 2507.020 36.220 2507.340 36.540 ;
        RECT 2686.420 35.540 2686.740 35.860 ;
        RECT 1913.620 32.820 1913.940 33.140 ;
      LAYER met4 ;
        RECT 1251.215 37.575 1251.545 37.905 ;
        RECT 2507.015 37.575 2507.345 37.905 ;
        RECT 1251.230 36.545 1251.530 37.575 ;
        RECT 1968.815 36.895 1969.145 37.225 ;
        RECT 1251.215 36.215 1251.545 36.545 ;
        RECT 1541.015 36.215 1541.345 36.545 ;
        RECT 1464.655 35.850 1464.985 35.865 ;
        RECT 1465.575 35.850 1465.905 35.865 ;
        RECT 1464.655 35.550 1465.905 35.850 ;
        RECT 1464.655 35.535 1464.985 35.550 ;
        RECT 1465.575 35.535 1465.905 35.550 ;
        RECT 1499.615 35.850 1499.945 35.865 ;
        RECT 1499.615 35.550 1500.850 35.850 ;
        RECT 1499.615 35.535 1499.945 35.550 ;
        RECT 1500.550 34.505 1500.850 35.550 ;
        RECT 1541.030 34.505 1541.330 36.215 ;
        RECT 1878.655 35.850 1878.985 35.865 ;
        RECT 1878.655 35.550 1879.890 35.850 ;
        RECT 1878.655 35.535 1878.985 35.550 ;
        RECT 1733.295 34.855 1733.625 35.185 ;
        RECT 1734.215 34.855 1734.545 35.185 ;
        RECT 1500.535 34.175 1500.865 34.505 ;
        RECT 1541.015 34.175 1541.345 34.505 ;
        RECT 1733.310 33.825 1733.610 34.855 ;
        RECT 1734.230 33.825 1734.530 34.855 ;
        RECT 1879.590 34.505 1879.890 35.550 ;
        RECT 1968.830 35.185 1969.130 36.895 ;
        RECT 2507.030 36.545 2507.330 37.575 ;
        RECT 2686.415 36.895 2686.745 37.225 ;
        RECT 2507.015 36.215 2507.345 36.545 ;
        RECT 2686.430 35.865 2686.730 36.895 ;
        RECT 2217.215 35.535 2217.545 35.865 ;
        RECT 2686.415 35.535 2686.745 35.865 ;
        RECT 1968.815 34.855 1969.145 35.185 ;
        RECT 2217.230 34.505 2217.530 35.535 ;
        RECT 1879.575 34.175 1879.905 34.505 ;
        RECT 1913.615 34.175 1913.945 34.505 ;
        RECT 2217.215 34.175 2217.545 34.505 ;
        RECT 1733.295 33.495 1733.625 33.825 ;
        RECT 1734.215 33.495 1734.545 33.825 ;
        RECT 1913.630 33.145 1913.930 34.175 ;
        RECT 1913.615 32.815 1913.945 33.145 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2900.550 2380.580 2900.870 2380.640 ;
        RECT 2870.580 2380.440 2900.870 2380.580 ;
        RECT 2900.550 2380.380 2900.870 2380.440 ;
      LAYER via ;
        RECT 2900.580 2380.380 2900.840 2380.640 ;
      LAYER met2 ;
        RECT 2900.570 2384.915 2900.850 2385.285 ;
        RECT 2900.640 2380.670 2900.780 2384.915 ;
        RECT 2900.580 2380.350 2900.840 2380.670 ;
      LAYER via2 ;
        RECT 2900.570 2384.960 2900.850 2385.240 ;
      LAYER met3 ;
        RECT 2900.545 2385.250 2900.875 2385.265 ;
        RECT 2920.080 2385.250 2922.480 2385.400 ;
        RECT 2900.545 2384.950 2922.480 2385.250 ;
        RECT 2900.545 2384.935 2900.875 2384.950 ;
        RECT 2920.080 2384.800 2922.480 2384.950 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2900.550 2615.180 2900.870 2615.240 ;
        RECT 2870.580 2615.040 2900.870 2615.180 ;
        RECT 2900.550 2614.980 2900.870 2615.040 ;
      LAYER via ;
        RECT 2900.580 2614.980 2900.840 2615.240 ;
      LAYER met2 ;
        RECT 2900.570 2619.515 2900.850 2619.885 ;
        RECT 2900.640 2615.270 2900.780 2619.515 ;
        RECT 2900.580 2614.950 2900.840 2615.270 ;
      LAYER via2 ;
        RECT 2900.570 2619.560 2900.850 2619.840 ;
      LAYER met3 ;
        RECT 2900.545 2619.850 2900.875 2619.865 ;
        RECT 2920.080 2619.850 2922.480 2620.000 ;
        RECT 2900.545 2619.550 2922.480 2619.850 ;
        RECT 2900.545 2619.535 2900.875 2619.550 ;
        RECT 2920.080 2619.400 2922.480 2619.550 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2900.550 2849.780 2900.870 2849.840 ;
        RECT 2870.580 2849.640 2900.870 2849.780 ;
        RECT 2900.550 2849.580 2900.870 2849.640 ;
      LAYER via ;
        RECT 2900.580 2849.580 2900.840 2849.840 ;
      LAYER met2 ;
        RECT 2900.570 2854.115 2900.850 2854.485 ;
        RECT 2900.640 2849.870 2900.780 2854.115 ;
        RECT 2900.580 2849.550 2900.840 2849.870 ;
      LAYER via2 ;
        RECT 2900.570 2854.160 2900.850 2854.440 ;
      LAYER met3 ;
        RECT 2900.545 2854.450 2900.875 2854.465 ;
        RECT 2920.080 2854.450 2922.480 2854.600 ;
        RECT 2900.545 2854.150 2922.480 2854.450 ;
        RECT 2900.545 2854.135 2900.875 2854.150 ;
        RECT 2920.080 2854.000 2922.480 2854.150 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2900.550 3085.060 2900.870 3085.120 ;
        RECT 2870.580 3084.920 2900.870 3085.060 ;
        RECT 2900.550 3084.860 2900.870 3084.920 ;
      LAYER via ;
        RECT 2900.580 3084.860 2900.840 3085.120 ;
      LAYER met2 ;
        RECT 2900.570 3088.715 2900.850 3089.085 ;
        RECT 2900.640 3085.150 2900.780 3088.715 ;
        RECT 2900.580 3084.830 2900.840 3085.150 ;
      LAYER via2 ;
        RECT 2900.570 3088.760 2900.850 3089.040 ;
      LAYER met3 ;
        RECT 2900.545 3089.050 2900.875 3089.065 ;
        RECT 2920.080 3089.050 2922.480 3089.200 ;
        RECT 2900.545 3088.750 2922.480 3089.050 ;
        RECT 2900.545 3088.735 2900.875 3088.750 ;
        RECT 2920.080 3088.600 2922.480 3088.750 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2900.550 3318.980 2900.870 3319.040 ;
        RECT 2870.580 3318.840 2900.870 3318.980 ;
        RECT 2900.550 3318.780 2900.870 3318.840 ;
      LAYER via ;
        RECT 2900.580 3318.780 2900.840 3319.040 ;
      LAYER met2 ;
        RECT 2900.570 3323.315 2900.850 3323.685 ;
        RECT 2900.640 3319.070 2900.780 3323.315 ;
        RECT 2900.580 3318.750 2900.840 3319.070 ;
      LAYER via2 ;
        RECT 2900.570 3323.360 2900.850 3323.640 ;
      LAYER met3 ;
        RECT 2900.545 3323.650 2900.875 3323.665 ;
        RECT 2920.080 3323.650 2922.480 3323.800 ;
        RECT 2900.545 3323.350 2922.480 3323.650 ;
        RECT 2900.545 3323.335 2900.875 3323.350 ;
        RECT 2920.080 3323.200 2922.480 3323.350 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2867.910 3517.600 2868.190 3520.000 ;
        RECT 2867.980 3517.370 2868.120 3517.600 ;
        RECT 2867.060 3517.230 2868.120 3517.370 ;
        RECT 2867.060 3466.000 2867.200 3517.230 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2542.285 3466.000 2542.455 3477.435 ;
      LAYER mcon ;
        RECT 2542.285 3477.265 2542.455 3477.435 ;
      LAYER met1 ;
        RECT 2542.210 3477.420 2542.530 3477.480 ;
        RECT 2542.015 3477.280 2542.530 3477.420 ;
        RECT 2542.210 3477.220 2542.530 3477.280 ;
      LAYER via ;
        RECT 2542.240 3477.220 2542.500 3477.480 ;
      LAYER met2 ;
        RECT 2543.610 3517.600 2543.890 3520.000 ;
        RECT 2543.680 3511.930 2543.820 3517.600 ;
        RECT 2542.300 3511.790 2543.820 3511.930 ;
        RECT 2542.300 3477.510 2542.440 3511.790 ;
        RECT 2542.240 3477.190 2542.500 3477.510 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2219.310 3517.600 2219.590 3520.000 ;
        RECT 2219.380 3517.370 2219.520 3517.600 ;
        RECT 2218.460 3517.230 2219.520 3517.370 ;
        RECT 2218.460 3466.000 2218.600 3517.230 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1893.685 3466.000 1893.855 3477.435 ;
      LAYER mcon ;
        RECT 1893.685 3477.265 1893.855 3477.435 ;
      LAYER met1 ;
        RECT 1893.610 3477.420 1893.930 3477.480 ;
        RECT 1893.415 3477.280 1893.930 3477.420 ;
        RECT 1893.610 3477.220 1893.930 3477.280 ;
      LAYER via ;
        RECT 1893.640 3477.220 1893.900 3477.480 ;
      LAYER met2 ;
        RECT 1894.550 3517.600 1894.830 3520.000 ;
        RECT 1894.620 3511.930 1894.760 3517.600 ;
        RECT 1893.700 3511.790 1894.760 3511.930 ;
        RECT 1893.700 3477.510 1893.840 3511.790 ;
        RECT 1893.640 3477.190 1893.900 3477.510 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1570.250 3517.600 1570.530 3520.000 ;
        RECT 1570.320 3517.370 1570.460 3517.600 ;
        RECT 1569.860 3517.230 1570.460 3517.370 ;
        RECT 1569.860 3466.000 1570.000 3517.230 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2903.770 2291.160 2904.090 2291.220 ;
        RECT 2870.580 2291.020 2904.090 2291.160 ;
        RECT 2903.770 2290.960 2904.090 2291.020 ;
      LAYER via ;
        RECT 2903.800 2290.960 2904.060 2291.220 ;
      LAYER met2 ;
        RECT 2903.800 2290.930 2904.060 2291.250 ;
        RECT 2903.860 273.885 2904.000 2290.930 ;
        RECT 2903.790 273.515 2904.070 273.885 ;
      LAYER via2 ;
        RECT 2903.790 273.560 2904.070 273.840 ;
      LAYER met3 ;
        RECT 2903.765 273.850 2904.095 273.865 ;
        RECT 2920.080 273.850 2922.480 274.000 ;
        RECT 2903.765 273.550 2922.480 273.850 ;
        RECT 2903.765 273.535 2904.095 273.550 ;
        RECT 2920.080 273.400 2922.480 273.550 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1245.930 3504.620 1246.250 3504.680 ;
        RECT 1250.990 3504.620 1251.310 3504.680 ;
        RECT 1245.930 3504.480 1251.310 3504.620 ;
        RECT 1245.930 3504.420 1246.250 3504.480 ;
        RECT 1250.990 3504.420 1251.310 3504.480 ;
      LAYER via ;
        RECT 1245.960 3504.420 1246.220 3504.680 ;
        RECT 1251.020 3504.420 1251.280 3504.680 ;
      LAYER met2 ;
        RECT 1245.950 3517.600 1246.230 3520.000 ;
        RECT 1246.020 3504.710 1246.160 3517.600 ;
        RECT 1245.960 3504.390 1246.220 3504.710 ;
        RECT 1251.020 3504.390 1251.280 3504.710 ;
        RECT 1251.080 3466.000 1251.220 3504.390 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 921.170 3504.280 921.490 3504.340 ;
        RECT 926.690 3504.280 927.010 3504.340 ;
        RECT 921.170 3504.140 927.010 3504.280 ;
        RECT 921.170 3504.080 921.490 3504.140 ;
        RECT 926.690 3504.080 927.010 3504.140 ;
      LAYER via ;
        RECT 921.200 3504.080 921.460 3504.340 ;
        RECT 926.720 3504.080 926.980 3504.340 ;
      LAYER met2 ;
        RECT 921.190 3517.600 921.470 3520.000 ;
        RECT 921.260 3504.370 921.400 3517.600 ;
        RECT 921.200 3504.050 921.460 3504.370 ;
        RECT 926.720 3504.050 926.980 3504.370 ;
        RECT 926.780 3466.000 926.920 3504.050 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1461.745 3504.805 1462.835 3504.975 ;
      LAYER mcon ;
        RECT 1462.665 3504.805 1462.835 3504.975 ;
      LAYER met1 ;
        RECT 596.870 3504.960 597.190 3505.020 ;
        RECT 1461.685 3504.960 1461.975 3505.005 ;
        RECT 596.870 3504.820 1461.975 3504.960 ;
        RECT 596.870 3504.760 597.190 3504.820 ;
        RECT 1461.685 3504.775 1461.975 3504.820 ;
        RECT 1462.605 3504.960 1462.895 3505.005 ;
        RECT 1499.850 3504.960 1500.170 3505.020 ;
        RECT 1462.605 3504.820 1500.170 3504.960 ;
        RECT 1462.605 3504.775 1462.895 3504.820 ;
        RECT 1499.850 3504.760 1500.170 3504.820 ;
      LAYER via ;
        RECT 596.900 3504.760 597.160 3505.020 ;
        RECT 1499.880 3504.760 1500.140 3505.020 ;
      LAYER met2 ;
        RECT 596.890 3517.600 597.170 3520.000 ;
        RECT 596.960 3505.050 597.100 3517.600 ;
        RECT 596.900 3504.730 597.160 3505.050 ;
        RECT 1499.880 3504.730 1500.140 3505.050 ;
        RECT 1499.940 3466.000 1500.080 3504.730 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 272.570 3502.580 272.890 3502.640 ;
        RECT 1513.650 3502.580 1513.970 3502.640 ;
        RECT 272.570 3502.440 1513.970 3502.580 ;
        RECT 272.570 3502.380 272.890 3502.440 ;
        RECT 1513.650 3502.380 1513.970 3502.440 ;
      LAYER via ;
        RECT 272.600 3502.380 272.860 3502.640 ;
        RECT 1513.680 3502.380 1513.940 3502.640 ;
      LAYER met2 ;
        RECT 272.590 3517.600 272.870 3520.000 ;
        RECT 272.660 3502.670 272.800 3517.600 ;
        RECT 272.600 3502.350 272.860 3502.670 ;
        RECT 1513.680 3502.350 1513.940 3502.670 ;
        RECT 1513.740 3466.000 1513.880 3502.350 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.650 3471.300 18.970 3471.360 ;
        RECT 1527.910 3471.300 1528.230 3471.360 ;
        RECT 18.650 3471.160 1528.230 3471.300 ;
        RECT 18.650 3471.100 18.970 3471.160 ;
        RECT 1527.910 3471.100 1528.230 3471.160 ;
      LAYER via ;
        RECT 18.680 3471.100 18.940 3471.360 ;
        RECT 1527.940 3471.100 1528.200 3471.360 ;
      LAYER met2 ;
        RECT 18.670 3476.995 18.950 3477.365 ;
        RECT 18.740 3471.390 18.880 3476.995 ;
        RECT 18.680 3471.070 18.940 3471.390 ;
        RECT 1527.940 3471.070 1528.200 3471.390 ;
        RECT 1528.000 3466.000 1528.140 3471.070 ;
      LAYER via2 ;
        RECT 18.670 3477.040 18.950 3477.320 ;
      LAYER met3 ;
        RECT 2.480 3477.330 4.880 3477.480 ;
        RECT 18.645 3477.330 18.975 3477.345 ;
        RECT 2.480 3477.030 18.975 3477.330 ;
        RECT 2.480 3476.880 4.880 3477.030 ;
        RECT 18.645 3477.015 18.975 3477.030 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.730 3222.420 18.050 3222.480 ;
        RECT 17.730 3222.280 54.000 3222.420 ;
        RECT 17.730 3222.220 18.050 3222.280 ;
      LAYER via ;
        RECT 17.760 3222.220 18.020 3222.480 ;
      LAYER met2 ;
        RECT 17.750 3226.075 18.030 3226.445 ;
        RECT 17.820 3222.510 17.960 3226.075 ;
        RECT 17.760 3222.190 18.020 3222.510 ;
      LAYER via2 ;
        RECT 17.750 3226.120 18.030 3226.400 ;
      LAYER met3 ;
        RECT 2.480 3226.410 4.880 3226.560 ;
        RECT 17.725 3226.410 18.055 3226.425 ;
        RECT 2.480 3226.110 18.055 3226.410 ;
        RECT 2.480 3225.960 4.880 3226.110 ;
        RECT 17.725 3226.095 18.055 3226.110 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.570 2974.220 19.890 2974.280 ;
        RECT 19.570 2974.080 54.000 2974.220 ;
        RECT 19.570 2974.020 19.890 2974.080 ;
      LAYER via ;
        RECT 19.600 2974.020 19.860 2974.280 ;
      LAYER met2 ;
        RECT 19.590 2974.475 19.870 2974.845 ;
        RECT 19.660 2974.310 19.800 2974.475 ;
        RECT 19.600 2973.990 19.860 2974.310 ;
      LAYER via2 ;
        RECT 19.590 2974.520 19.870 2974.800 ;
      LAYER met3 ;
        RECT 2.480 2974.810 4.880 2974.960 ;
        RECT 19.565 2974.810 19.895 2974.825 ;
        RECT 2.480 2974.510 19.895 2974.810 ;
        RECT 2.480 2974.360 4.880 2974.510 ;
        RECT 19.565 2974.495 19.895 2974.510 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.190 2718.880 18.510 2718.940 ;
        RECT 18.190 2718.740 54.000 2718.880 ;
        RECT 18.190 2718.680 18.510 2718.740 ;
      LAYER via ;
        RECT 18.220 2718.680 18.480 2718.940 ;
      LAYER met2 ;
        RECT 18.210 2722.875 18.490 2723.245 ;
        RECT 18.280 2718.970 18.420 2722.875 ;
        RECT 18.220 2718.650 18.480 2718.970 ;
      LAYER via2 ;
        RECT 18.210 2722.920 18.490 2723.200 ;
      LAYER met3 ;
        RECT 2.480 2723.210 4.880 2723.360 ;
        RECT 18.185 2723.210 18.515 2723.225 ;
        RECT 2.480 2722.910 18.515 2723.210 ;
        RECT 2.480 2722.760 4.880 2722.910 ;
        RECT 18.185 2722.895 18.515 2722.910 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.650 2470.340 18.970 2470.400 ;
        RECT 18.650 2470.200 54.000 2470.340 ;
        RECT 18.650 2470.140 18.970 2470.200 ;
      LAYER via ;
        RECT 18.680 2470.140 18.940 2470.400 ;
      LAYER met2 ;
        RECT 18.670 2471.275 18.950 2471.645 ;
        RECT 18.740 2470.430 18.880 2471.275 ;
        RECT 18.680 2470.110 18.940 2470.430 ;
      LAYER via2 ;
        RECT 18.670 2471.320 18.950 2471.600 ;
      LAYER met3 ;
        RECT 2.480 2471.610 4.880 2471.760 ;
        RECT 18.645 2471.610 18.975 2471.625 ;
        RECT 2.480 2471.310 18.975 2471.610 ;
        RECT 2.480 2471.160 4.880 2471.310 ;
        RECT 18.645 2471.295 18.975 2471.310 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 33.830 2305.100 34.150 2305.160 ;
        RECT 33.830 2304.960 54.000 2305.100 ;
        RECT 33.830 2304.900 34.150 2304.960 ;
        RECT 18.190 2220.780 18.510 2220.840 ;
        RECT 33.830 2220.780 34.150 2220.840 ;
        RECT 18.190 2220.640 34.150 2220.780 ;
        RECT 18.190 2220.580 18.510 2220.640 ;
        RECT 33.830 2220.580 34.150 2220.640 ;
      LAYER via ;
        RECT 33.860 2304.900 34.120 2305.160 ;
        RECT 18.220 2220.580 18.480 2220.840 ;
        RECT 33.860 2220.580 34.120 2220.840 ;
      LAYER met2 ;
        RECT 33.860 2304.870 34.120 2305.190 ;
        RECT 33.920 2220.870 34.060 2304.870 ;
        RECT 18.220 2220.725 18.480 2220.870 ;
        RECT 18.210 2220.355 18.490 2220.725 ;
        RECT 33.860 2220.550 34.120 2220.870 ;
      LAYER via2 ;
        RECT 18.210 2220.400 18.490 2220.680 ;
      LAYER met3 ;
        RECT 2.480 2220.690 4.880 2220.840 ;
        RECT 18.185 2220.690 18.515 2220.705 ;
        RECT 2.480 2220.390 18.515 2220.690 ;
        RECT 2.480 2220.240 4.880 2220.390 ;
        RECT 18.185 2220.375 18.515 2220.390 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2920.080 508.450 2922.480 508.600 ;
        RECT 2919.190 508.150 2922.480 508.450 ;
        RECT 2919.190 505.050 2919.490 508.150 ;
        RECT 2920.080 508.000 2922.480 508.150 ;
        RECT 2870.580 504.750 2886.370 505.050 ;
        RECT 2886.070 504.370 2886.370 504.750 ;
        RECT 2886.990 504.750 2919.490 505.050 ;
        RECT 2886.990 504.370 2887.290 504.750 ;
        RECT 2886.070 504.070 2887.290 504.370 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.110 1973.260 19.430 1973.320 ;
        RECT 19.110 1973.120 54.000 1973.260 ;
        RECT 19.110 1973.060 19.430 1973.120 ;
      LAYER via ;
        RECT 19.140 1973.060 19.400 1973.320 ;
      LAYER met2 ;
        RECT 19.140 1973.030 19.400 1973.350 ;
        RECT 19.200 1969.125 19.340 1973.030 ;
        RECT 19.130 1968.755 19.410 1969.125 ;
      LAYER via2 ;
        RECT 19.130 1968.800 19.410 1969.080 ;
      LAYER met3 ;
        RECT 2.480 1969.090 4.880 1969.240 ;
        RECT 19.105 1969.090 19.435 1969.105 ;
        RECT 2.480 1968.790 19.435 1969.090 ;
        RECT 2.480 1968.640 4.880 1968.790 ;
        RECT 19.105 1968.775 19.435 1968.790 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.110 1717.920 19.430 1717.980 ;
        RECT 19.110 1717.780 54.000 1717.920 ;
        RECT 19.110 1717.720 19.430 1717.780 ;
      LAYER via ;
        RECT 19.140 1717.720 19.400 1717.980 ;
      LAYER met2 ;
        RECT 19.140 1717.690 19.400 1718.010 ;
        RECT 19.200 1717.525 19.340 1717.690 ;
        RECT 19.130 1717.155 19.410 1717.525 ;
      LAYER via2 ;
        RECT 19.130 1717.200 19.410 1717.480 ;
      LAYER met3 ;
        RECT 2.480 1717.490 4.880 1717.640 ;
        RECT 19.105 1717.490 19.435 1717.505 ;
        RECT 2.480 1717.190 19.435 1717.490 ;
        RECT 2.480 1717.040 4.880 1717.190 ;
        RECT 19.105 1717.175 19.435 1717.190 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 33.370 2291.840 33.690 2291.900 ;
        RECT 33.370 2291.700 54.000 2291.840 ;
        RECT 33.370 2291.640 33.690 2291.700 ;
        RECT 17.730 1469.380 18.050 1469.440 ;
        RECT 33.370 1469.380 33.690 1469.440 ;
        RECT 17.730 1469.240 33.690 1469.380 ;
        RECT 17.730 1469.180 18.050 1469.240 ;
        RECT 33.370 1469.180 33.690 1469.240 ;
      LAYER via ;
        RECT 33.400 2291.640 33.660 2291.900 ;
        RECT 17.760 1469.180 18.020 1469.440 ;
        RECT 33.400 1469.180 33.660 1469.440 ;
      LAYER met2 ;
        RECT 33.400 2291.610 33.660 2291.930 ;
        RECT 33.460 1469.470 33.600 2291.610 ;
        RECT 17.760 1469.150 18.020 1469.470 ;
        RECT 33.400 1469.150 33.660 1469.470 ;
        RECT 17.820 1466.605 17.960 1469.150 ;
        RECT 17.750 1466.235 18.030 1466.605 ;
      LAYER via2 ;
        RECT 17.750 1466.280 18.030 1466.560 ;
      LAYER met3 ;
        RECT 2.480 1466.570 4.880 1466.720 ;
        RECT 17.725 1466.570 18.055 1466.585 ;
        RECT 2.480 1466.270 18.055 1466.570 ;
        RECT 2.480 1466.120 4.880 1466.270 ;
        RECT 17.725 1466.255 18.055 1466.270 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.110 1220.840 19.430 1220.900 ;
        RECT 19.110 1220.700 54.000 1220.840 ;
        RECT 19.110 1220.640 19.430 1220.700 ;
      LAYER via ;
        RECT 19.140 1220.640 19.400 1220.900 ;
      LAYER met2 ;
        RECT 19.140 1220.610 19.400 1220.930 ;
        RECT 19.200 1215.005 19.340 1220.610 ;
        RECT 19.130 1214.635 19.410 1215.005 ;
      LAYER via2 ;
        RECT 19.130 1214.680 19.410 1214.960 ;
      LAYER met3 ;
        RECT 2.480 1214.970 4.880 1215.120 ;
        RECT 19.105 1214.970 19.435 1214.985 ;
        RECT 2.480 1214.670 19.435 1214.970 ;
        RECT 2.480 1214.520 4.880 1214.670 ;
        RECT 19.105 1214.655 19.435 1214.670 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 47.170 2291.500 47.490 2291.560 ;
        RECT 47.170 2291.360 54.000 2291.500 ;
        RECT 47.170 2291.300 47.490 2291.360 ;
        RECT 19.110 963.460 19.430 963.520 ;
        RECT 47.170 963.460 47.490 963.520 ;
        RECT 19.110 963.320 47.490 963.460 ;
        RECT 19.110 963.260 19.430 963.320 ;
        RECT 47.170 963.260 47.490 963.320 ;
      LAYER via ;
        RECT 47.200 2291.300 47.460 2291.560 ;
        RECT 19.140 963.260 19.400 963.520 ;
        RECT 47.200 963.260 47.460 963.520 ;
      LAYER met2 ;
        RECT 47.200 2291.270 47.460 2291.590 ;
        RECT 47.260 963.550 47.400 2291.270 ;
        RECT 19.140 963.405 19.400 963.550 ;
        RECT 19.130 963.035 19.410 963.405 ;
        RECT 47.200 963.230 47.460 963.550 ;
      LAYER via2 ;
        RECT 19.130 963.080 19.410 963.360 ;
      LAYER met3 ;
        RECT 2.480 963.370 4.880 963.520 ;
        RECT 19.105 963.370 19.435 963.385 ;
        RECT 2.480 963.070 19.435 963.370 ;
        RECT 2.480 962.920 4.880 963.070 ;
        RECT 19.105 963.055 19.435 963.070 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.030 717.640 20.350 717.700 ;
        RECT 20.030 717.500 54.000 717.640 ;
        RECT 20.030 717.440 20.350 717.500 ;
      LAYER via ;
        RECT 20.060 717.440 20.320 717.700 ;
      LAYER met2 ;
        RECT 20.060 717.410 20.320 717.730 ;
        RECT 20.120 711.805 20.260 717.410 ;
        RECT 20.050 711.435 20.330 711.805 ;
      LAYER via2 ;
        RECT 20.050 711.480 20.330 711.760 ;
      LAYER met3 ;
        RECT 2.480 711.770 4.880 711.920 ;
        RECT 20.025 711.770 20.355 711.785 ;
        RECT 2.480 711.470 20.355 711.770 ;
        RECT 2.480 711.320 4.880 711.470 ;
        RECT 20.025 711.455 20.355 711.470 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5.550 461.910 54.000 462.210 ;
        RECT 2.480 460.850 4.880 461.000 ;
        RECT 5.550 460.850 5.850 461.910 ;
        RECT 2.480 460.550 5.850 460.850 ;
        RECT 2.480 460.400 4.880 460.550 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.590 213.675 19.870 214.045 ;
        RECT 19.660 209.285 19.800 213.675 ;
        RECT 19.590 208.915 19.870 209.285 ;
      LAYER via2 ;
        RECT 19.590 213.720 19.870 214.000 ;
        RECT 19.590 208.960 19.870 209.240 ;
      LAYER met3 ;
        RECT 19.565 214.010 19.895 214.025 ;
        RECT 19.565 213.710 54.000 214.010 ;
        RECT 19.565 213.695 19.895 213.710 ;
        RECT 2.480 209.250 4.880 209.400 ;
        RECT 19.565 209.250 19.895 209.265 ;
        RECT 2.480 208.950 19.895 209.250 ;
        RECT 2.480 208.800 4.880 208.950 ;
        RECT 19.565 208.935 19.895 208.950 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2901.930 744.840 2902.250 744.900 ;
        RECT 2870.580 744.700 2902.250 744.840 ;
        RECT 2901.930 744.640 2902.250 744.700 ;
      LAYER via ;
        RECT 2901.960 744.640 2902.220 744.900 ;
      LAYER met2 ;
        RECT 2901.960 744.610 2902.220 744.930 ;
        RECT 2902.020 743.085 2902.160 744.610 ;
        RECT 2901.950 742.715 2902.230 743.085 ;
      LAYER via2 ;
        RECT 2901.950 742.760 2902.230 743.040 ;
      LAYER met3 ;
        RECT 2901.925 743.050 2902.255 743.065 ;
        RECT 2920.080 743.050 2922.480 743.200 ;
        RECT 2901.925 742.750 2922.480 743.050 ;
        RECT 2901.925 742.735 2902.255 742.750 ;
        RECT 2920.080 742.600 2922.480 742.750 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2903.310 979.780 2903.630 979.840 ;
        RECT 2870.580 979.640 2903.630 979.780 ;
        RECT 2903.310 979.580 2903.630 979.640 ;
      LAYER via ;
        RECT 2903.340 979.580 2903.600 979.840 ;
      LAYER met2 ;
        RECT 2903.340 979.550 2903.600 979.870 ;
        RECT 2903.400 977.685 2903.540 979.550 ;
        RECT 2903.330 977.315 2903.610 977.685 ;
      LAYER via2 ;
        RECT 2903.330 977.360 2903.610 977.640 ;
      LAYER met3 ;
        RECT 2903.305 977.650 2903.635 977.665 ;
        RECT 2920.080 977.650 2922.480 977.800 ;
        RECT 2903.305 977.350 2922.480 977.650 ;
        RECT 2903.305 977.335 2903.635 977.350 ;
        RECT 2920.080 977.200 2922.480 977.350 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2920.080 1212.250 2922.480 1212.400 ;
        RECT 2919.190 1211.950 2922.480 1212.250 ;
        RECT 2919.190 1208.850 2919.490 1211.950 ;
        RECT 2920.080 1211.800 2922.480 1211.950 ;
        RECT 2870.580 1208.550 2886.370 1208.850 ;
        RECT 2886.070 1208.170 2886.370 1208.550 ;
        RECT 2886.990 1208.550 2919.490 1208.850 ;
        RECT 2886.990 1208.170 2887.290 1208.550 ;
        RECT 2886.070 1207.870 2887.290 1208.170 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2903.310 1448.980 2903.630 1449.040 ;
        RECT 2870.580 1448.840 2903.630 1448.980 ;
        RECT 2903.310 1448.780 2903.630 1448.840 ;
      LAYER via ;
        RECT 2903.340 1448.780 2903.600 1449.040 ;
      LAYER met2 ;
        RECT 2903.340 1448.750 2903.600 1449.070 ;
        RECT 2903.400 1446.885 2903.540 1448.750 ;
        RECT 2903.330 1446.515 2903.610 1446.885 ;
      LAYER via2 ;
        RECT 2903.330 1446.560 2903.610 1446.840 ;
      LAYER met3 ;
        RECT 2903.305 1446.850 2903.635 1446.865 ;
        RECT 2920.080 1446.850 2922.480 1447.000 ;
        RECT 2903.305 1446.550 2922.480 1446.850 ;
        RECT 2903.305 1446.535 2903.635 1446.550 ;
        RECT 2920.080 1446.400 2922.480 1446.550 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2901.930 1683.240 2902.250 1683.300 ;
        RECT 2870.580 1683.100 2902.250 1683.240 ;
        RECT 2901.930 1683.040 2902.250 1683.100 ;
      LAYER via ;
        RECT 2901.960 1683.040 2902.220 1683.300 ;
      LAYER met2 ;
        RECT 2901.960 1683.010 2902.220 1683.330 ;
        RECT 2902.020 1681.485 2902.160 1683.010 ;
        RECT 2901.950 1681.115 2902.230 1681.485 ;
      LAYER via2 ;
        RECT 2901.950 1681.160 2902.230 1681.440 ;
      LAYER met3 ;
        RECT 2901.925 1681.450 2902.255 1681.465 ;
        RECT 2920.080 1681.450 2922.480 1681.600 ;
        RECT 2901.925 1681.150 2922.480 1681.450 ;
        RECT 2901.925 1681.135 2902.255 1681.150 ;
        RECT 2920.080 1681.000 2922.480 1681.150 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2903.310 1918.180 2903.630 1918.240 ;
        RECT 2870.580 1918.040 2903.630 1918.180 ;
        RECT 2903.310 1917.980 2903.630 1918.040 ;
      LAYER via ;
        RECT 2903.340 1917.980 2903.600 1918.240 ;
      LAYER met2 ;
        RECT 2903.340 1917.950 2903.600 1918.270 ;
        RECT 2903.400 1916.085 2903.540 1917.950 ;
        RECT 2903.330 1915.715 2903.610 1916.085 ;
      LAYER via2 ;
        RECT 2903.330 1915.760 2903.610 1916.040 ;
      LAYER met3 ;
        RECT 2903.305 1916.050 2903.635 1916.065 ;
        RECT 2920.080 1916.050 2922.480 1916.200 ;
        RECT 2903.305 1915.750 2922.480 1916.050 ;
        RECT 2903.305 1915.735 2903.635 1915.750 ;
        RECT 2920.080 1915.600 2922.480 1915.750 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2903.310 2152.780 2903.630 2152.840 ;
        RECT 2870.580 2152.640 2903.630 2152.780 ;
        RECT 2903.310 2152.580 2903.630 2152.640 ;
      LAYER via ;
        RECT 2903.340 2152.580 2903.600 2152.840 ;
      LAYER met2 ;
        RECT 2903.340 2152.550 2903.600 2152.870 ;
        RECT 2903.400 2150.685 2903.540 2152.550 ;
        RECT 2903.330 2150.315 2903.610 2150.685 ;
      LAYER via2 ;
        RECT 2903.330 2150.360 2903.610 2150.640 ;
      LAYER met3 ;
        RECT 2903.305 2150.650 2903.635 2150.665 ;
        RECT 2920.080 2150.650 2922.480 2150.800 ;
        RECT 2903.305 2150.350 2922.480 2150.650 ;
        RECT 2903.305 2150.335 2903.635 2150.350 ;
        RECT 2920.080 2150.200 2922.480 2150.350 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.080 195.650 2922.480 195.800 ;
        RECT 2919.190 195.350 2922.480 195.650 ;
        RECT 2919.190 194.290 2919.490 195.350 ;
        RECT 2920.080 195.200 2922.480 195.350 ;
        RECT 2870.580 193.990 2886.370 194.290 ;
        RECT 2886.070 193.610 2886.370 193.990 ;
        RECT 2886.990 193.990 2919.490 194.290 ;
        RECT 2886.990 193.610 2887.290 193.990 ;
        RECT 2886.070 193.310 2887.290 193.610 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.550 2539.360 2900.870 2539.420 ;
        RECT 2870.580 2539.220 2900.870 2539.360 ;
        RECT 2900.550 2539.160 2900.870 2539.220 ;
      LAYER via ;
        RECT 2900.580 2539.160 2900.840 2539.420 ;
      LAYER met2 ;
        RECT 2900.570 2541.315 2900.850 2541.685 ;
        RECT 2900.640 2539.450 2900.780 2541.315 ;
        RECT 2900.580 2539.130 2900.840 2539.450 ;
      LAYER via2 ;
        RECT 2900.570 2541.360 2900.850 2541.640 ;
      LAYER met3 ;
        RECT 2900.545 2541.650 2900.875 2541.665 ;
        RECT 2920.080 2541.650 2922.480 2541.800 ;
        RECT 2900.545 2541.350 2922.480 2541.650 ;
        RECT 2900.545 2541.335 2900.875 2541.350 ;
        RECT 2920.080 2541.200 2922.480 2541.350 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.550 2773.960 2900.870 2774.020 ;
        RECT 2870.580 2773.820 2900.870 2773.960 ;
        RECT 2900.550 2773.760 2900.870 2773.820 ;
      LAYER via ;
        RECT 2900.580 2773.760 2900.840 2774.020 ;
      LAYER met2 ;
        RECT 2900.570 2775.915 2900.850 2776.285 ;
        RECT 2900.640 2774.050 2900.780 2775.915 ;
        RECT 2900.580 2773.730 2900.840 2774.050 ;
      LAYER via2 ;
        RECT 2900.570 2775.960 2900.850 2776.240 ;
      LAYER met3 ;
        RECT 2900.545 2776.250 2900.875 2776.265 ;
        RECT 2920.080 2776.250 2922.480 2776.400 ;
        RECT 2900.545 2775.950 2922.480 2776.250 ;
        RECT 2900.545 2775.935 2900.875 2775.950 ;
        RECT 2920.080 2775.800 2922.480 2775.950 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.550 3008.900 2900.870 3008.960 ;
        RECT 2870.580 3008.760 2900.870 3008.900 ;
        RECT 2900.550 3008.700 2900.870 3008.760 ;
      LAYER via ;
        RECT 2900.580 3008.700 2900.840 3008.960 ;
      LAYER met2 ;
        RECT 2900.570 3010.515 2900.850 3010.885 ;
        RECT 2900.640 3008.990 2900.780 3010.515 ;
        RECT 2900.580 3008.670 2900.840 3008.990 ;
      LAYER via2 ;
        RECT 2900.570 3010.560 2900.850 3010.840 ;
      LAYER met3 ;
        RECT 2900.545 3010.850 2900.875 3010.865 ;
        RECT 2920.080 3010.850 2922.480 3011.000 ;
        RECT 2900.545 3010.550 2922.480 3010.850 ;
        RECT 2900.545 3010.535 2900.875 3010.550 ;
        RECT 2920.080 3010.400 2922.480 3010.550 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.550 3243.160 2900.870 3243.220 ;
        RECT 2870.580 3243.020 2900.870 3243.160 ;
        RECT 2900.550 3242.960 2900.870 3243.020 ;
      LAYER via ;
        RECT 2900.580 3242.960 2900.840 3243.220 ;
      LAYER met2 ;
        RECT 2900.570 3245.115 2900.850 3245.485 ;
        RECT 2900.640 3243.250 2900.780 3245.115 ;
        RECT 2900.580 3242.930 2900.840 3243.250 ;
      LAYER via2 ;
        RECT 2900.570 3245.160 2900.850 3245.440 ;
      LAYER met3 ;
        RECT 2900.545 3245.450 2900.875 3245.465 ;
        RECT 2920.080 3245.450 2922.480 3245.600 ;
        RECT 2900.545 3245.150 2922.480 3245.450 ;
        RECT 2900.545 3245.135 2900.875 3245.150 ;
        RECT 2920.080 3245.000 2922.480 3245.150 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1382.090 3477.760 1382.410 3477.820 ;
        RECT 2900.550 3477.760 2900.870 3477.820 ;
        RECT 1382.090 3477.620 2900.870 3477.760 ;
        RECT 1382.090 3477.560 1382.410 3477.620 ;
        RECT 2900.550 3477.560 2900.870 3477.620 ;
      LAYER via ;
        RECT 1382.120 3477.560 1382.380 3477.820 ;
        RECT 2900.580 3477.560 2900.840 3477.820 ;
      LAYER met2 ;
        RECT 2900.570 3479.715 2900.850 3480.085 ;
        RECT 2900.640 3477.850 2900.780 3479.715 ;
        RECT 1382.120 3477.530 1382.380 3477.850 ;
        RECT 2900.580 3477.530 2900.840 3477.850 ;
        RECT 1382.180 3466.000 1382.320 3477.530 ;
      LAYER via2 ;
        RECT 2900.570 3479.760 2900.850 3480.040 ;
      LAYER met3 ;
        RECT 2900.545 3480.050 2900.875 3480.065 ;
        RECT 2920.080 3480.050 2922.480 3480.200 ;
        RECT 2900.545 3479.750 2922.480 3480.050 ;
        RECT 2900.545 3479.735 2900.875 3479.750 ;
        RECT 2920.080 3479.600 2922.480 3479.750 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1402.790 3502.240 1403.110 3502.300 ;
        RECT 2651.690 3502.240 2652.010 3502.300 ;
        RECT 1402.790 3502.100 2652.010 3502.240 ;
        RECT 1402.790 3502.040 1403.110 3502.100 ;
        RECT 2651.690 3502.040 2652.010 3502.100 ;
      LAYER via ;
        RECT 1402.820 3502.040 1403.080 3502.300 ;
        RECT 2651.720 3502.040 2651.980 3502.300 ;
      LAYER met2 ;
        RECT 2651.710 3517.600 2651.990 3520.000 ;
        RECT 2651.780 3502.330 2651.920 3517.600 ;
        RECT 1402.820 3502.010 1403.080 3502.330 ;
        RECT 2651.720 3502.010 2651.980 3502.330 ;
        RECT 1402.880 3466.000 1403.020 3502.010 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1450.245 3499.365 1450.415 3505.655 ;
        RECT 1481.525 3504.465 1481.695 3505.655 ;
      LAYER mcon ;
        RECT 1450.245 3505.485 1450.415 3505.655 ;
        RECT 1481.525 3505.485 1481.695 3505.655 ;
      LAYER met1 ;
        RECT 1450.185 3505.640 1450.475 3505.685 ;
        RECT 1481.465 3505.640 1481.755 3505.685 ;
        RECT 1450.185 3505.500 1481.755 3505.640 ;
        RECT 1450.185 3505.455 1450.475 3505.500 ;
        RECT 1481.465 3505.455 1481.755 3505.500 ;
        RECT 1481.465 3504.620 1481.755 3504.665 ;
        RECT 2327.390 3504.620 2327.710 3504.680 ;
        RECT 1481.465 3504.480 2327.710 3504.620 ;
        RECT 1481.465 3504.435 1481.755 3504.480 ;
        RECT 2327.390 3504.420 2327.710 3504.480 ;
        RECT 1416.590 3499.520 1416.910 3499.580 ;
        RECT 1450.185 3499.520 1450.475 3499.565 ;
        RECT 1416.590 3499.380 1450.475 3499.520 ;
        RECT 1416.590 3499.320 1416.910 3499.380 ;
        RECT 1450.185 3499.335 1450.475 3499.380 ;
      LAYER via ;
        RECT 2327.420 3504.420 2327.680 3504.680 ;
        RECT 1416.620 3499.320 1416.880 3499.580 ;
      LAYER met2 ;
        RECT 2327.410 3517.600 2327.690 3520.000 ;
        RECT 2327.480 3504.710 2327.620 3517.600 ;
        RECT 2327.420 3504.390 2327.680 3504.710 ;
        RECT 1416.620 3499.290 1416.880 3499.610 ;
        RECT 1416.680 3466.000 1416.820 3499.290 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1443.805 3504.125 1443.975 3505.315 ;
        RECT 1481.065 3499.365 1481.235 3504.635 ;
      LAYER mcon ;
        RECT 1443.805 3505.145 1443.975 3505.315 ;
        RECT 1481.065 3504.465 1481.235 3504.635 ;
      LAYER met1 ;
        RECT 1443.745 3505.300 1444.035 3505.345 ;
        RECT 1443.745 3505.160 1462.360 3505.300 ;
        RECT 1443.745 3505.115 1444.035 3505.160 ;
        RECT 1462.220 3504.620 1462.360 3505.160 ;
        RECT 1481.005 3504.620 1481.295 3504.665 ;
        RECT 1462.220 3504.480 1481.295 3504.620 ;
        RECT 1481.005 3504.435 1481.295 3504.480 ;
        RECT 1430.390 3504.280 1430.710 3504.340 ;
        RECT 1443.745 3504.280 1444.035 3504.325 ;
        RECT 1430.390 3504.140 1444.035 3504.280 ;
        RECT 1430.390 3504.080 1430.710 3504.140 ;
        RECT 1443.745 3504.095 1444.035 3504.140 ;
        RECT 1481.005 3499.520 1481.295 3499.565 ;
        RECT 2003.090 3499.520 2003.410 3499.580 ;
        RECT 1481.005 3499.380 2003.410 3499.520 ;
        RECT 1481.005 3499.335 1481.295 3499.380 ;
        RECT 2003.090 3499.320 2003.410 3499.380 ;
      LAYER via ;
        RECT 1430.420 3504.080 1430.680 3504.340 ;
        RECT 2003.120 3499.320 2003.380 3499.580 ;
      LAYER met2 ;
        RECT 2003.110 3517.600 2003.390 3520.000 ;
        RECT 1430.420 3504.050 1430.680 3504.370 ;
        RECT 1430.480 3466.000 1430.620 3504.050 ;
        RECT 2003.180 3499.610 2003.320 3517.600 ;
        RECT 2003.120 3499.290 2003.380 3499.610 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1461.285 3504.125 1462.375 3504.295 ;
        RECT 1462.205 3500.045 1462.375 3504.125 ;
        RECT 1480.605 3499.025 1480.775 3500.215 ;
      LAYER mcon ;
        RECT 1480.605 3500.045 1480.775 3500.215 ;
      LAYER met1 ;
        RECT 1444.190 3504.280 1444.510 3504.340 ;
        RECT 1461.225 3504.280 1461.515 3504.325 ;
        RECT 1444.190 3504.140 1461.515 3504.280 ;
        RECT 1444.190 3504.080 1444.510 3504.140 ;
        RECT 1461.225 3504.095 1461.515 3504.140 ;
        RECT 1462.145 3500.200 1462.435 3500.245 ;
        RECT 1480.545 3500.200 1480.835 3500.245 ;
        RECT 1462.145 3500.060 1480.835 3500.200 ;
        RECT 1462.145 3500.015 1462.435 3500.060 ;
        RECT 1480.545 3500.015 1480.835 3500.060 ;
        RECT 1480.545 3499.180 1480.835 3499.225 ;
        RECT 1678.330 3499.180 1678.650 3499.240 ;
        RECT 1480.545 3499.040 1678.650 3499.180 ;
        RECT 1480.545 3498.995 1480.835 3499.040 ;
        RECT 1678.330 3498.980 1678.650 3499.040 ;
      LAYER via ;
        RECT 1444.220 3504.080 1444.480 3504.340 ;
        RECT 1678.360 3498.980 1678.620 3499.240 ;
      LAYER met2 ;
        RECT 1678.350 3517.600 1678.630 3520.000 ;
        RECT 1444.220 3504.050 1444.480 3504.370 ;
        RECT 1444.280 3466.000 1444.420 3504.050 ;
        RECT 1678.420 3499.270 1678.560 3517.600 ;
        RECT 1678.360 3498.950 1678.620 3499.270 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1393.205 3498.345 1393.375 3499.535 ;
        RECT 1444.265 3498.685 1445.355 3498.855 ;
        RECT 1444.265 3498.345 1444.435 3498.685 ;
      LAYER mcon ;
        RECT 1393.205 3499.365 1393.375 3499.535 ;
        RECT 1445.185 3498.685 1445.355 3498.855 ;
      LAYER met1 ;
        RECT 1354.030 3499.860 1354.350 3499.920 ;
        RECT 1354.030 3499.720 1392.440 3499.860 ;
        RECT 1354.030 3499.660 1354.350 3499.720 ;
        RECT 1392.300 3499.520 1392.440 3499.720 ;
        RECT 1393.145 3499.520 1393.435 3499.565 ;
        RECT 1392.300 3499.380 1393.435 3499.520 ;
        RECT 1393.145 3499.335 1393.435 3499.380 ;
        RECT 1445.125 3498.840 1445.415 3498.885 ;
        RECT 1458.910 3498.840 1459.230 3498.900 ;
        RECT 1445.125 3498.700 1459.230 3498.840 ;
        RECT 1445.125 3498.655 1445.415 3498.700 ;
        RECT 1458.910 3498.640 1459.230 3498.700 ;
        RECT 1393.145 3498.500 1393.435 3498.545 ;
        RECT 1444.205 3498.500 1444.495 3498.545 ;
        RECT 1393.145 3498.360 1444.495 3498.500 ;
        RECT 1393.145 3498.315 1393.435 3498.360 ;
        RECT 1444.205 3498.315 1444.495 3498.360 ;
      LAYER via ;
        RECT 1354.060 3499.660 1354.320 3499.920 ;
        RECT 1458.940 3498.640 1459.200 3498.900 ;
      LAYER met2 ;
        RECT 1354.050 3517.600 1354.330 3520.000 ;
        RECT 1354.120 3499.950 1354.260 3517.600 ;
        RECT 1354.060 3499.630 1354.320 3499.950 ;
        RECT 1458.940 3498.610 1459.200 3498.930 ;
        RECT 1459.000 3466.000 1459.140 3498.610 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2903.310 434.760 2903.630 434.820 ;
        RECT 2870.580 434.620 2903.630 434.760 ;
        RECT 2903.310 434.560 2903.630 434.620 ;
      LAYER via ;
        RECT 2903.340 434.560 2903.600 434.820 ;
      LAYER met2 ;
        RECT 2903.340 434.530 2903.600 434.850 ;
        RECT 2903.400 430.285 2903.540 434.530 ;
        RECT 2903.330 429.915 2903.610 430.285 ;
      LAYER via2 ;
        RECT 2903.330 429.960 2903.610 430.240 ;
      LAYER met3 ;
        RECT 2903.305 430.250 2903.635 430.265 ;
        RECT 2920.080 430.250 2922.480 430.400 ;
        RECT 2903.305 429.950 2922.480 430.250 ;
        RECT 2903.305 429.935 2903.635 429.950 ;
        RECT 2920.080 429.800 2922.480 429.950 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1472.250 3499.520 1472.570 3499.580 ;
        RECT 1450.720 3499.380 1472.570 3499.520 ;
        RECT 1029.730 3499.180 1030.050 3499.240 ;
        RECT 1450.720 3499.180 1450.860 3499.380 ;
        RECT 1472.250 3499.320 1472.570 3499.380 ;
        RECT 1029.730 3499.040 1450.860 3499.180 ;
        RECT 1029.730 3498.980 1030.050 3499.040 ;
      LAYER via ;
        RECT 1029.760 3498.980 1030.020 3499.240 ;
        RECT 1472.280 3499.320 1472.540 3499.580 ;
      LAYER met2 ;
        RECT 1029.750 3517.600 1030.030 3520.000 ;
        RECT 1029.820 3499.270 1029.960 3517.600 ;
        RECT 1472.280 3499.290 1472.540 3499.610 ;
        RECT 1029.760 3498.950 1030.020 3499.270 ;
        RECT 1472.340 3466.000 1472.480 3499.290 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1461.285 3499.195 1461.455 3501.235 ;
        RECT 1461.285 3499.025 1463.295 3499.195 ;
      LAYER mcon ;
        RECT 1461.285 3501.065 1461.455 3501.235 ;
        RECT 1463.125 3499.025 1463.295 3499.195 ;
      LAYER met1 ;
        RECT 704.970 3501.220 705.290 3501.280 ;
        RECT 1461.225 3501.220 1461.515 3501.265 ;
        RECT 704.970 3501.080 1461.515 3501.220 ;
        RECT 704.970 3501.020 705.290 3501.080 ;
        RECT 1461.225 3501.035 1461.515 3501.080 ;
        RECT 1463.065 3499.180 1463.355 3499.225 ;
        RECT 1463.065 3499.040 1480.300 3499.180 ;
        RECT 1463.065 3498.995 1463.355 3499.040 ;
        RECT 1480.160 3498.840 1480.300 3499.040 ;
        RECT 1486.050 3498.840 1486.370 3498.900 ;
        RECT 1480.160 3498.700 1486.370 3498.840 ;
        RECT 1486.050 3498.640 1486.370 3498.700 ;
      LAYER via ;
        RECT 705.000 3501.020 705.260 3501.280 ;
        RECT 1486.080 3498.640 1486.340 3498.900 ;
      LAYER met2 ;
        RECT 704.990 3517.600 705.270 3520.000 ;
        RECT 705.060 3501.310 705.200 3517.600 ;
        RECT 705.000 3500.990 705.260 3501.310 ;
        RECT 1486.080 3498.610 1486.340 3498.930 ;
        RECT 1486.140 3466.000 1486.280 3498.610 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 380.670 3502.920 380.990 3502.980 ;
        RECT 1507.210 3502.920 1507.530 3502.980 ;
        RECT 380.670 3502.780 1507.530 3502.920 ;
        RECT 380.670 3502.720 380.990 3502.780 ;
        RECT 1507.210 3502.720 1507.530 3502.780 ;
      LAYER via ;
        RECT 380.700 3502.720 380.960 3502.980 ;
        RECT 1507.240 3502.720 1507.500 3502.980 ;
      LAYER met2 ;
        RECT 380.690 3517.600 380.970 3520.000 ;
        RECT 380.760 3503.010 380.900 3517.600 ;
        RECT 380.700 3502.690 380.960 3503.010 ;
        RECT 1507.240 3502.690 1507.500 3503.010 ;
        RECT 1507.300 3466.000 1507.440 3502.690 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.390 3517.600 56.670 3520.000 ;
        RECT 56.460 3501.845 56.600 3517.600 ;
        RECT 56.390 3501.475 56.670 3501.845 ;
        RECT 1520.570 3501.475 1520.850 3501.845 ;
        RECT 1520.640 3466.000 1520.780 3501.475 ;
      LAYER via2 ;
        RECT 56.390 3501.520 56.670 3501.800 ;
        RECT 1520.570 3501.520 1520.850 3501.800 ;
      LAYER met3 ;
        RECT 56.365 3501.810 56.695 3501.825 ;
        RECT 1520.545 3501.810 1520.875 3501.825 ;
        RECT 56.365 3501.510 1520.875 3501.810 ;
        RECT 56.365 3501.495 56.695 3501.510 ;
        RECT 1520.545 3501.495 1520.875 3501.510 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.570 3305.380 19.890 3305.440 ;
        RECT 19.570 3305.240 54.000 3305.380 ;
        RECT 19.570 3305.180 19.890 3305.240 ;
      LAYER via ;
        RECT 19.600 3305.180 19.860 3305.440 ;
      LAYER met2 ;
        RECT 19.590 3309.715 19.870 3310.085 ;
        RECT 19.660 3305.470 19.800 3309.715 ;
        RECT 19.600 3305.150 19.860 3305.470 ;
      LAYER via2 ;
        RECT 19.590 3309.760 19.870 3310.040 ;
      LAYER met3 ;
        RECT 2.480 3310.050 4.880 3310.200 ;
        RECT 19.565 3310.050 19.895 3310.065 ;
        RECT 2.480 3309.750 19.895 3310.050 ;
        RECT 2.480 3309.600 4.880 3309.750 ;
        RECT 19.565 3309.735 19.895 3309.750 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.110 3056.840 19.430 3056.900 ;
        RECT 19.110 3056.700 54.000 3056.840 ;
        RECT 19.110 3056.640 19.430 3056.700 ;
      LAYER via ;
        RECT 19.140 3056.640 19.400 3056.900 ;
      LAYER met2 ;
        RECT 19.130 3058.115 19.410 3058.485 ;
        RECT 19.200 3056.930 19.340 3058.115 ;
        RECT 19.140 3056.610 19.400 3056.930 ;
      LAYER via2 ;
        RECT 19.130 3058.160 19.410 3058.440 ;
      LAYER met3 ;
        RECT 2.480 3058.450 4.880 3058.600 ;
        RECT 19.105 3058.450 19.435 3058.465 ;
        RECT 2.480 3058.150 19.435 3058.450 ;
        RECT 2.480 3058.000 4.880 3058.150 ;
        RECT 19.105 3058.135 19.435 3058.150 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.570 2802.180 19.890 2802.240 ;
        RECT 19.570 2802.040 54.000 2802.180 ;
        RECT 19.570 2801.980 19.890 2802.040 ;
      LAYER via ;
        RECT 19.600 2801.980 19.860 2802.240 ;
      LAYER met2 ;
        RECT 19.590 2806.515 19.870 2806.885 ;
        RECT 19.660 2802.270 19.800 2806.515 ;
        RECT 19.600 2801.950 19.860 2802.270 ;
      LAYER via2 ;
        RECT 19.590 2806.560 19.870 2806.840 ;
      LAYER met3 ;
        RECT 2.480 2806.850 4.880 2807.000 ;
        RECT 19.565 2806.850 19.895 2806.865 ;
        RECT 2.480 2806.550 19.895 2806.850 ;
        RECT 2.480 2806.400 4.880 2806.550 ;
        RECT 19.565 2806.535 19.895 2806.550 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.030 2553.300 20.350 2553.360 ;
        RECT 20.030 2553.160 54.000 2553.300 ;
        RECT 20.030 2553.100 20.350 2553.160 ;
      LAYER via ;
        RECT 20.060 2553.100 20.320 2553.360 ;
      LAYER met2 ;
        RECT 20.050 2555.595 20.330 2555.965 ;
        RECT 20.120 2553.390 20.260 2555.595 ;
        RECT 20.060 2553.070 20.320 2553.390 ;
      LAYER via2 ;
        RECT 20.050 2555.640 20.330 2555.920 ;
      LAYER met3 ;
        RECT 2.480 2555.930 4.880 2556.080 ;
        RECT 20.025 2555.930 20.355 2555.945 ;
        RECT 2.480 2555.630 20.355 2555.930 ;
        RECT 2.480 2555.480 4.880 2555.630 ;
        RECT 20.025 2555.615 20.355 2555.630 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 36.665 2297.465 36.835 2298.995 ;
        RECT 37.125 2297.805 37.295 2298.995 ;
      LAYER mcon ;
        RECT 36.665 2298.825 36.835 2298.995 ;
        RECT 37.125 2298.825 37.295 2298.995 ;
      LAYER met1 ;
        RECT 18.190 2298.980 18.510 2299.040 ;
        RECT 36.605 2298.980 36.895 2299.025 ;
        RECT 18.190 2298.840 36.895 2298.980 ;
        RECT 18.190 2298.780 18.510 2298.840 ;
        RECT 36.605 2298.795 36.895 2298.840 ;
        RECT 37.065 2298.980 37.355 2299.025 ;
        RECT 37.065 2298.840 54.000 2298.980 ;
        RECT 37.065 2298.795 37.355 2298.840 ;
        RECT 37.065 2297.775 37.355 2298.005 ;
        RECT 36.605 2297.620 36.895 2297.665 ;
        RECT 37.140 2297.620 37.280 2297.775 ;
        RECT 36.605 2297.480 37.280 2297.620 ;
        RECT 36.605 2297.435 36.895 2297.480 ;
      LAYER via ;
        RECT 18.220 2298.780 18.480 2299.040 ;
      LAYER met2 ;
        RECT 18.210 2303.995 18.490 2304.365 ;
        RECT 18.280 2299.070 18.420 2303.995 ;
        RECT 18.220 2298.750 18.480 2299.070 ;
      LAYER via2 ;
        RECT 18.210 2304.040 18.490 2304.320 ;
      LAYER met3 ;
        RECT 2.480 2304.330 4.880 2304.480 ;
        RECT 18.185 2304.330 18.515 2304.345 ;
        RECT 2.480 2304.030 18.515 2304.330 ;
        RECT 2.480 2303.880 4.880 2304.030 ;
        RECT 18.185 2304.015 18.515 2304.030 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.110 2055.880 19.430 2055.940 ;
        RECT 19.110 2055.740 54.000 2055.880 ;
        RECT 19.110 2055.680 19.430 2055.740 ;
      LAYER via ;
        RECT 19.140 2055.680 19.400 2055.940 ;
      LAYER met2 ;
        RECT 19.140 2055.650 19.400 2055.970 ;
        RECT 19.200 2052.765 19.340 2055.650 ;
        RECT 19.130 2052.395 19.410 2052.765 ;
      LAYER via2 ;
        RECT 19.130 2052.440 19.410 2052.720 ;
      LAYER met3 ;
        RECT 2.480 2052.730 4.880 2052.880 ;
        RECT 19.105 2052.730 19.435 2052.745 ;
        RECT 2.480 2052.430 19.435 2052.730 ;
        RECT 2.480 2052.280 4.880 2052.430 ;
        RECT 19.105 2052.415 19.435 2052.430 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.080 664.850 2922.480 665.000 ;
        RECT 2919.190 664.550 2922.480 664.850 ;
        RECT 2919.190 663.490 2919.490 664.550 ;
        RECT 2920.080 664.400 2922.480 664.550 ;
        RECT 2870.580 663.190 2886.370 663.490 ;
        RECT 2886.070 662.810 2886.370 663.190 ;
        RECT 2886.990 663.190 2919.490 663.490 ;
        RECT 2886.990 662.810 2887.290 663.190 ;
        RECT 2886.070 662.510 2887.290 662.810 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.110 1807.680 19.430 1807.740 ;
        RECT 19.110 1807.540 54.000 1807.680 ;
        RECT 19.110 1807.480 19.430 1807.540 ;
      LAYER via ;
        RECT 19.140 1807.480 19.400 1807.740 ;
      LAYER met2 ;
        RECT 19.140 1807.450 19.400 1807.770 ;
        RECT 19.200 1801.845 19.340 1807.450 ;
        RECT 19.130 1801.475 19.410 1801.845 ;
      LAYER via2 ;
        RECT 19.130 1801.520 19.410 1801.800 ;
      LAYER met3 ;
        RECT 2.480 1801.810 4.880 1801.960 ;
        RECT 19.105 1801.810 19.435 1801.825 ;
        RECT 2.480 1801.510 19.435 1801.810 ;
        RECT 2.480 1801.360 4.880 1801.510 ;
        RECT 19.105 1801.495 19.435 1801.510 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.190 1552.340 18.510 1552.400 ;
        RECT 18.190 1552.200 54.000 1552.340 ;
        RECT 18.190 1552.140 18.510 1552.200 ;
      LAYER via ;
        RECT 18.220 1552.140 18.480 1552.400 ;
      LAYER met2 ;
        RECT 18.220 1552.110 18.480 1552.430 ;
        RECT 18.280 1550.245 18.420 1552.110 ;
        RECT 18.210 1549.875 18.490 1550.245 ;
      LAYER via2 ;
        RECT 18.210 1549.920 18.490 1550.200 ;
      LAYER met3 ;
        RECT 2.480 1550.210 4.880 1550.360 ;
        RECT 18.185 1550.210 18.515 1550.225 ;
        RECT 2.480 1549.910 18.515 1550.210 ;
        RECT 2.480 1549.760 4.880 1549.910 ;
        RECT 18.185 1549.895 18.515 1549.910 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.110 1304.140 19.430 1304.200 ;
        RECT 19.110 1304.000 54.000 1304.140 ;
        RECT 19.110 1303.940 19.430 1304.000 ;
      LAYER via ;
        RECT 19.140 1303.940 19.400 1304.200 ;
      LAYER met2 ;
        RECT 19.140 1303.910 19.400 1304.230 ;
        RECT 19.200 1298.645 19.340 1303.910 ;
        RECT 19.130 1298.275 19.410 1298.645 ;
      LAYER via2 ;
        RECT 19.130 1298.320 19.410 1298.600 ;
      LAYER met3 ;
        RECT 2.480 1298.610 4.880 1298.760 ;
        RECT 19.105 1298.610 19.435 1298.625 ;
        RECT 2.480 1298.310 19.435 1298.610 ;
        RECT 2.480 1298.160 4.880 1298.310 ;
        RECT 19.105 1298.295 19.435 1298.310 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.650 1048.800 18.970 1048.860 ;
        RECT 18.650 1048.660 54.000 1048.800 ;
        RECT 18.650 1048.600 18.970 1048.660 ;
      LAYER via ;
        RECT 18.680 1048.600 18.940 1048.860 ;
      LAYER met2 ;
        RECT 18.680 1048.570 18.940 1048.890 ;
        RECT 18.740 1047.045 18.880 1048.570 ;
        RECT 18.670 1046.675 18.950 1047.045 ;
      LAYER via2 ;
        RECT 18.670 1046.720 18.950 1047.000 ;
      LAYER met3 ;
        RECT 2.480 1047.010 4.880 1047.160 ;
        RECT 18.645 1047.010 18.975 1047.025 ;
        RECT 2.480 1046.710 18.975 1047.010 ;
        RECT 2.480 1046.560 4.880 1046.710 ;
        RECT 18.645 1046.695 18.975 1046.710 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.030 2312.920 20.350 2312.980 ;
        RECT 20.030 2312.780 54.000 2312.920 ;
        RECT 20.030 2312.720 20.350 2312.780 ;
      LAYER via ;
        RECT 20.060 2312.720 20.320 2312.980 ;
      LAYER met2 ;
        RECT 20.060 2312.690 20.320 2313.010 ;
        RECT 20.120 796.125 20.260 2312.690 ;
        RECT 20.050 795.755 20.330 796.125 ;
      LAYER via2 ;
        RECT 20.050 795.800 20.330 796.080 ;
      LAYER met3 ;
        RECT 2.480 796.090 4.880 796.240 ;
        RECT 20.025 796.090 20.355 796.105 ;
        RECT 2.480 795.790 20.355 796.090 ;
        RECT 2.480 795.640 4.880 795.790 ;
        RECT 20.025 795.775 20.355 795.790 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.590 2312.155 19.870 2312.525 ;
        RECT 19.660 544.525 19.800 2312.155 ;
        RECT 19.590 544.155 19.870 544.525 ;
      LAYER via2 ;
        RECT 19.590 2312.200 19.870 2312.480 ;
        RECT 19.590 544.200 19.870 544.480 ;
      LAYER met3 ;
        RECT 19.565 2312.490 19.895 2312.505 ;
        RECT 19.565 2312.190 54.000 2312.490 ;
        RECT 19.565 2312.175 19.895 2312.190 ;
        RECT 2.480 544.490 4.880 544.640 ;
        RECT 19.565 544.490 19.895 544.505 ;
        RECT 2.480 544.190 19.895 544.490 ;
        RECT 2.480 544.040 4.880 544.190 ;
        RECT 19.565 544.175 19.895 544.190 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.190 296.040 18.510 296.100 ;
        RECT 18.190 295.900 54.000 296.040 ;
        RECT 18.190 295.840 18.510 295.900 ;
      LAYER via ;
        RECT 18.220 295.840 18.480 296.100 ;
      LAYER met2 ;
        RECT 18.220 295.810 18.480 296.130 ;
        RECT 18.280 292.925 18.420 295.810 ;
        RECT 18.210 292.555 18.490 292.925 ;
      LAYER via2 ;
        RECT 18.210 292.600 18.490 292.880 ;
      LAYER met3 ;
        RECT 2.480 292.890 4.880 293.040 ;
        RECT 18.185 292.890 18.515 292.905 ;
        RECT 2.480 292.590 18.515 292.890 ;
        RECT 2.480 292.440 4.880 292.590 ;
        RECT 18.185 292.575 18.515 292.590 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.590 47.755 19.870 48.125 ;
        RECT 19.660 42.005 19.800 47.755 ;
        RECT 19.590 41.635 19.870 42.005 ;
      LAYER via2 ;
        RECT 19.590 47.800 19.870 48.080 ;
        RECT 19.590 41.680 19.870 41.960 ;
      LAYER met3 ;
        RECT 19.565 48.090 19.895 48.105 ;
        RECT 1741.550 48.090 1741.930 48.100 ;
        RECT 19.565 47.790 1741.930 48.090 ;
        RECT 19.565 47.775 19.895 47.790 ;
        RECT 1741.550 47.780 1741.930 47.790 ;
        RECT 2.480 41.970 4.880 42.120 ;
        RECT 19.565 41.970 19.895 41.985 ;
        RECT 2.480 41.670 19.895 41.970 ;
        RECT 2.480 41.520 4.880 41.670 ;
        RECT 19.565 41.655 19.895 41.670 ;
      LAYER via3 ;
        RECT 1741.580 47.780 1741.900 48.100 ;
      LAYER met4 ;
        RECT 1741.590 48.105 1741.890 54.000 ;
        RECT 1741.575 47.775 1741.905 48.105 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.080 899.450 2922.480 899.600 ;
        RECT 2919.190 899.150 2922.480 899.450 ;
        RECT 2919.190 898.090 2919.490 899.150 ;
        RECT 2920.080 899.000 2922.480 899.150 ;
        RECT 2870.580 897.790 2886.370 898.090 ;
        RECT 2886.070 897.410 2886.370 897.790 ;
        RECT 2886.990 897.790 2919.490 898.090 ;
        RECT 2886.990 897.410 2887.290 897.790 ;
        RECT 2886.070 897.110 2887.290 897.410 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.080 1134.050 2922.480 1134.200 ;
        RECT 2919.190 1133.750 2922.480 1134.050 ;
        RECT 2919.190 1132.690 2919.490 1133.750 ;
        RECT 2920.080 1133.600 2922.480 1133.750 ;
        RECT 2870.580 1132.390 2886.370 1132.690 ;
        RECT 2886.070 1132.010 2886.370 1132.390 ;
        RECT 2886.990 1132.390 2919.490 1132.690 ;
        RECT 2886.990 1132.010 2887.290 1132.390 ;
        RECT 2886.070 1131.710 2887.290 1132.010 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2903.310 1373.160 2903.630 1373.220 ;
        RECT 2870.580 1373.020 2903.630 1373.160 ;
        RECT 2903.310 1372.960 2903.630 1373.020 ;
      LAYER via ;
        RECT 2903.340 1372.960 2903.600 1373.220 ;
      LAYER met2 ;
        RECT 2903.340 1372.930 2903.600 1373.250 ;
        RECT 2903.400 1368.685 2903.540 1372.930 ;
        RECT 2903.330 1368.315 2903.610 1368.685 ;
      LAYER via2 ;
        RECT 2903.330 1368.360 2903.610 1368.640 ;
      LAYER met3 ;
        RECT 2903.305 1368.650 2903.635 1368.665 ;
        RECT 2920.080 1368.650 2922.480 1368.800 ;
        RECT 2903.305 1368.350 2922.480 1368.650 ;
        RECT 2903.305 1368.335 2903.635 1368.350 ;
        RECT 2920.080 1368.200 2922.480 1368.350 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.080 1603.250 2922.480 1603.400 ;
        RECT 2919.190 1602.950 2922.480 1603.250 ;
        RECT 2919.190 1601.890 2919.490 1602.950 ;
        RECT 2920.080 1602.800 2922.480 1602.950 ;
        RECT 2870.580 1601.590 2886.370 1601.890 ;
        RECT 2886.070 1601.210 2886.370 1601.590 ;
        RECT 2886.990 1601.590 2919.490 1601.890 ;
        RECT 2886.990 1601.210 2887.290 1601.590 ;
        RECT 2886.070 1600.910 2887.290 1601.210 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2903.310 1842.360 2903.630 1842.420 ;
        RECT 2870.580 1842.220 2903.630 1842.360 ;
        RECT 2903.310 1842.160 2903.630 1842.220 ;
      LAYER via ;
        RECT 2903.340 1842.160 2903.600 1842.420 ;
      LAYER met2 ;
        RECT 2903.340 1842.130 2903.600 1842.450 ;
        RECT 2903.400 1837.885 2903.540 1842.130 ;
        RECT 2903.330 1837.515 2903.610 1837.885 ;
      LAYER via2 ;
        RECT 2903.330 1837.560 2903.610 1837.840 ;
      LAYER met3 ;
        RECT 2903.305 1837.850 2903.635 1837.865 ;
        RECT 2920.080 1837.850 2922.480 1838.000 ;
        RECT 2903.305 1837.550 2922.480 1837.850 ;
        RECT 2903.305 1837.535 2903.635 1837.550 ;
        RECT 2920.080 1837.400 2922.480 1837.550 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2903.310 2076.960 2903.630 2077.020 ;
        RECT 2870.580 2076.820 2903.630 2076.960 ;
        RECT 2903.310 2076.760 2903.630 2076.820 ;
      LAYER via ;
        RECT 2903.340 2076.760 2903.600 2077.020 ;
      LAYER met2 ;
        RECT 2903.340 2076.730 2903.600 2077.050 ;
        RECT 2903.400 2072.485 2903.540 2076.730 ;
        RECT 2903.330 2072.115 2903.610 2072.485 ;
      LAYER via2 ;
        RECT 2903.330 2072.160 2903.610 2072.440 ;
      LAYER met3 ;
        RECT 2903.305 2072.450 2903.635 2072.465 ;
        RECT 2920.080 2072.450 2922.480 2072.600 ;
        RECT 2903.305 2072.150 2922.480 2072.450 ;
        RECT 2903.305 2072.135 2903.635 2072.150 ;
        RECT 2920.080 2072.000 2922.480 2072.150 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2903.310 2304.760 2903.630 2304.820 ;
        RECT 2870.580 2304.620 2903.630 2304.760 ;
        RECT 2903.310 2304.560 2903.630 2304.620 ;
      LAYER via ;
        RECT 2903.340 2304.560 2903.600 2304.820 ;
      LAYER met2 ;
        RECT 2903.330 2306.715 2903.610 2307.085 ;
        RECT 2903.400 2304.850 2903.540 2306.715 ;
        RECT 2903.340 2304.530 2903.600 2304.850 ;
      LAYER via2 ;
        RECT 2903.330 2306.760 2903.610 2307.040 ;
      LAYER met3 ;
        RECT 2903.305 2307.050 2903.635 2307.065 ;
        RECT 2920.080 2307.050 2922.480 2307.200 ;
        RECT 2903.305 2306.750 2922.480 2307.050 ;
        RECT 2903.305 2306.735 2903.635 2306.750 ;
        RECT 2920.080 2306.600 2922.480 2306.750 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.080 117.450 2922.480 117.600 ;
        RECT 2870.580 117.150 2922.480 117.450 ;
        RECT 2920.080 117.000 2922.480 117.150 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.550 2463.540 2900.870 2463.600 ;
        RECT 2870.580 2463.400 2900.870 2463.540 ;
        RECT 2900.550 2463.340 2900.870 2463.400 ;
      LAYER via ;
        RECT 2900.580 2463.340 2900.840 2463.600 ;
      LAYER met2 ;
        RECT 2900.580 2463.485 2900.840 2463.630 ;
        RECT 2900.570 2463.115 2900.850 2463.485 ;
      LAYER via2 ;
        RECT 2900.570 2463.160 2900.850 2463.440 ;
      LAYER met3 ;
        RECT 2900.545 2463.450 2900.875 2463.465 ;
        RECT 2920.080 2463.450 2922.480 2463.600 ;
        RECT 2900.545 2463.150 2922.480 2463.450 ;
        RECT 2900.545 2463.135 2900.875 2463.150 ;
        RECT 2920.080 2463.000 2922.480 2463.150 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.550 2698.820 2900.870 2698.880 ;
        RECT 2870.580 2698.680 2900.870 2698.820 ;
        RECT 2900.550 2698.620 2900.870 2698.680 ;
      LAYER via ;
        RECT 2900.580 2698.620 2900.840 2698.880 ;
      LAYER met2 ;
        RECT 2900.580 2698.590 2900.840 2698.910 ;
        RECT 2900.640 2698.085 2900.780 2698.590 ;
        RECT 2900.570 2697.715 2900.850 2698.085 ;
      LAYER via2 ;
        RECT 2900.570 2697.760 2900.850 2698.040 ;
      LAYER met3 ;
        RECT 2900.545 2698.050 2900.875 2698.065 ;
        RECT 2920.080 2698.050 2922.480 2698.200 ;
        RECT 2900.545 2697.750 2922.480 2698.050 ;
        RECT 2900.545 2697.735 2900.875 2697.750 ;
        RECT 2920.080 2697.600 2922.480 2697.750 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.550 2932.740 2900.870 2932.800 ;
        RECT 2870.580 2932.600 2900.870 2932.740 ;
        RECT 2900.550 2932.540 2900.870 2932.600 ;
      LAYER via ;
        RECT 2900.580 2932.540 2900.840 2932.800 ;
      LAYER met2 ;
        RECT 2900.580 2932.685 2900.840 2932.830 ;
        RECT 2900.570 2932.315 2900.850 2932.685 ;
      LAYER via2 ;
        RECT 2900.570 2932.360 2900.850 2932.640 ;
      LAYER met3 ;
        RECT 2900.545 2932.650 2900.875 2932.665 ;
        RECT 2920.080 2932.650 2922.480 2932.800 ;
        RECT 2900.545 2932.350 2922.480 2932.650 ;
        RECT 2900.545 2932.335 2900.875 2932.350 ;
        RECT 2920.080 2932.200 2922.480 2932.350 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.550 3167.340 2900.870 3167.400 ;
        RECT 2870.580 3167.200 2900.870 3167.340 ;
        RECT 2900.550 3167.140 2900.870 3167.200 ;
      LAYER via ;
        RECT 2900.580 3167.140 2900.840 3167.400 ;
      LAYER met2 ;
        RECT 2900.580 3167.285 2900.840 3167.430 ;
        RECT 2900.570 3166.915 2900.850 3167.285 ;
      LAYER via2 ;
        RECT 2900.570 3166.960 2900.850 3167.240 ;
      LAYER met3 ;
        RECT 2900.545 3167.250 2900.875 3167.265 ;
        RECT 2920.080 3167.250 2922.480 3167.400 ;
        RECT 2900.545 3166.950 2922.480 3167.250 ;
        RECT 2900.545 3166.935 2900.875 3166.950 ;
        RECT 2920.080 3166.800 2922.480 3166.950 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.550 3401.940 2900.870 3402.000 ;
        RECT 2870.580 3401.800 2900.870 3401.940 ;
        RECT 2900.550 3401.740 2900.870 3401.800 ;
      LAYER via ;
        RECT 2900.580 3401.740 2900.840 3402.000 ;
      LAYER met2 ;
        RECT 2900.580 3401.885 2900.840 3402.030 ;
        RECT 2900.570 3401.515 2900.850 3401.885 ;
      LAYER via2 ;
        RECT 2900.570 3401.560 2900.850 3401.840 ;
      LAYER met3 ;
        RECT 2900.545 3401.850 2900.875 3401.865 ;
        RECT 2920.080 3401.850 2922.480 3402.000 ;
        RECT 2900.545 3401.550 2922.480 3401.850 ;
        RECT 2900.545 3401.535 2900.875 3401.550 ;
        RECT 2920.080 3401.400 2922.480 3401.550 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1402.330 3501.900 1402.650 3501.960 ;
        RECT 2759.790 3501.900 2760.110 3501.960 ;
        RECT 1402.330 3501.760 2760.110 3501.900 ;
        RECT 1402.330 3501.700 1402.650 3501.760 ;
        RECT 2759.790 3501.700 2760.110 3501.760 ;
      LAYER via ;
        RECT 1402.360 3501.700 1402.620 3501.960 ;
        RECT 2759.820 3501.700 2760.080 3501.960 ;
      LAYER met2 ;
        RECT 2759.810 3517.600 2760.090 3520.000 ;
        RECT 2759.880 3501.990 2760.020 3517.600 ;
        RECT 1402.360 3501.670 1402.620 3501.990 ;
        RECT 2759.820 3501.670 2760.080 3501.990 ;
        RECT 1402.420 3466.000 1402.560 3501.670 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1423.490 3504.620 1423.810 3504.680 ;
        RECT 1423.490 3504.480 1461.900 3504.620 ;
        RECT 1423.490 3504.420 1423.810 3504.480 ;
        RECT 1461.760 3504.280 1461.900 3504.480 ;
        RECT 2435.490 3504.280 2435.810 3504.340 ;
        RECT 1461.760 3504.140 2435.810 3504.280 ;
        RECT 2435.490 3504.080 2435.810 3504.140 ;
      LAYER via ;
        RECT 1423.520 3504.420 1423.780 3504.680 ;
        RECT 2435.520 3504.080 2435.780 3504.340 ;
      LAYER met2 ;
        RECT 2435.510 3517.600 2435.790 3520.000 ;
        RECT 1423.520 3504.390 1423.780 3504.710 ;
        RECT 1423.580 3466.000 1423.720 3504.390 ;
        RECT 2435.580 3504.370 2435.720 3517.600 ;
        RECT 2435.520 3504.050 2435.780 3504.370 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1472.785 3499.705 1473.875 3499.875 ;
      LAYER mcon ;
        RECT 1473.705 3499.705 1473.875 3499.875 ;
      LAYER met1 ;
        RECT 1437.290 3499.860 1437.610 3499.920 ;
        RECT 1472.725 3499.860 1473.015 3499.905 ;
        RECT 1437.290 3499.720 1473.015 3499.860 ;
        RECT 1437.290 3499.660 1437.610 3499.720 ;
        RECT 1472.725 3499.675 1473.015 3499.720 ;
        RECT 1473.645 3499.860 1473.935 3499.905 ;
        RECT 2111.190 3499.860 2111.510 3499.920 ;
        RECT 1473.645 3499.720 2111.510 3499.860 ;
        RECT 1473.645 3499.675 1473.935 3499.720 ;
        RECT 2111.190 3499.660 2111.510 3499.720 ;
      LAYER via ;
        RECT 1437.320 3499.660 1437.580 3499.920 ;
        RECT 2111.220 3499.660 2111.480 3499.920 ;
      LAYER met2 ;
        RECT 2111.210 3517.600 2111.490 3520.000 ;
        RECT 2111.280 3499.950 2111.420 3517.600 ;
        RECT 1437.320 3499.630 1437.580 3499.950 ;
        RECT 2111.220 3499.630 2111.480 3499.950 ;
        RECT 1437.380 3466.000 1437.520 3499.630 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1451.090 3499.180 1451.410 3499.240 ;
        RECT 1462.590 3499.180 1462.910 3499.240 ;
        RECT 1451.090 3499.040 1462.910 3499.180 ;
        RECT 1451.090 3498.980 1451.410 3499.040 ;
        RECT 1462.590 3498.980 1462.910 3499.040 ;
        RECT 1462.590 3498.500 1462.910 3498.560 ;
        RECT 1786.430 3498.500 1786.750 3498.560 ;
        RECT 1462.590 3498.360 1786.750 3498.500 ;
        RECT 1462.590 3498.300 1462.910 3498.360 ;
        RECT 1786.430 3498.300 1786.750 3498.360 ;
      LAYER via ;
        RECT 1451.120 3498.980 1451.380 3499.240 ;
        RECT 1462.620 3498.980 1462.880 3499.240 ;
        RECT 1462.620 3498.300 1462.880 3498.560 ;
        RECT 1786.460 3498.300 1786.720 3498.560 ;
      LAYER met2 ;
        RECT 1786.450 3517.600 1786.730 3520.000 ;
        RECT 1451.120 3498.950 1451.380 3499.270 ;
        RECT 1462.620 3498.950 1462.880 3499.270 ;
        RECT 1451.180 3466.000 1451.320 3498.950 ;
        RECT 1462.680 3498.590 1462.820 3498.950 ;
        RECT 1786.520 3498.590 1786.660 3517.600 ;
        RECT 1462.620 3498.270 1462.880 3498.590 ;
        RECT 1786.460 3498.270 1786.720 3498.590 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1458.450 3498.500 1458.770 3498.560 ;
        RECT 1462.130 3498.500 1462.450 3498.560 ;
        RECT 1458.450 3498.360 1462.450 3498.500 ;
        RECT 1458.450 3498.300 1458.770 3498.360 ;
        RECT 1462.130 3498.300 1462.450 3498.360 ;
      LAYER via ;
        RECT 1458.480 3498.300 1458.740 3498.560 ;
        RECT 1462.160 3498.300 1462.420 3498.560 ;
      LAYER met2 ;
        RECT 1462.150 3517.600 1462.430 3520.000 ;
        RECT 1462.220 3498.590 1462.360 3517.600 ;
        RECT 1458.480 3498.270 1458.740 3498.590 ;
        RECT 1462.160 3498.270 1462.420 3498.590 ;
        RECT 1458.540 3466.000 1458.680 3498.270 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.080 352.050 2922.480 352.200 ;
        RECT 2870.580 351.750 2922.480 352.050 ;
        RECT 2920.080 351.600 2922.480 351.750 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1148.025 3498.685 1148.195 3499.535 ;
        RECT 1196.325 3498.345 1196.495 3499.535 ;
        RECT 1296.145 3498.345 1296.315 3499.535 ;
        RECT 1320.525 3498.345 1320.695 3499.535 ;
        RECT 1392.745 3498.345 1392.915 3499.875 ;
        RECT 1436.905 3498.855 1437.075 3499.875 ;
        RECT 1436.905 3498.685 1437.535 3498.855 ;
        RECT 1458.065 3498.685 1459.615 3498.855 ;
        RECT 1458.065 3498.345 1458.235 3498.685 ;
      LAYER mcon ;
        RECT 1392.745 3499.705 1392.915 3499.875 ;
        RECT 1148.025 3499.365 1148.195 3499.535 ;
        RECT 1196.325 3499.365 1196.495 3499.535 ;
        RECT 1296.145 3499.365 1296.315 3499.535 ;
        RECT 1320.525 3499.365 1320.695 3499.535 ;
        RECT 1436.905 3499.705 1437.075 3499.875 ;
        RECT 1437.365 3498.685 1437.535 3498.855 ;
        RECT 1459.445 3498.685 1459.615 3498.855 ;
      LAYER met1 ;
        RECT 1392.685 3499.860 1392.975 3499.905 ;
        RECT 1436.845 3499.860 1437.135 3499.905 ;
        RECT 1392.685 3499.720 1437.135 3499.860 ;
        RECT 1392.685 3499.675 1392.975 3499.720 ;
        RECT 1436.845 3499.675 1437.135 3499.720 ;
        RECT 1147.965 3499.520 1148.255 3499.565 ;
        RECT 1196.265 3499.520 1196.555 3499.565 ;
        RECT 1147.965 3499.380 1196.555 3499.520 ;
        RECT 1147.965 3499.335 1148.255 3499.380 ;
        RECT 1196.265 3499.335 1196.555 3499.380 ;
        RECT 1296.085 3499.520 1296.375 3499.565 ;
        RECT 1320.465 3499.520 1320.755 3499.565 ;
        RECT 1296.085 3499.380 1320.755 3499.520 ;
        RECT 1296.085 3499.335 1296.375 3499.380 ;
        RECT 1320.465 3499.335 1320.755 3499.380 ;
        RECT 1137.830 3498.840 1138.150 3498.900 ;
        RECT 1147.965 3498.840 1148.255 3498.885 ;
        RECT 1137.830 3498.700 1148.255 3498.840 ;
        RECT 1137.830 3498.640 1138.150 3498.700 ;
        RECT 1147.965 3498.655 1148.255 3498.700 ;
        RECT 1437.305 3498.840 1437.595 3498.885 ;
        RECT 1459.385 3498.840 1459.675 3498.885 ;
        RECT 1479.610 3498.840 1479.930 3498.900 ;
        RECT 1437.305 3498.700 1444.880 3498.840 ;
        RECT 1437.305 3498.655 1437.595 3498.700 ;
        RECT 1196.265 3498.500 1196.555 3498.545 ;
        RECT 1296.085 3498.500 1296.375 3498.545 ;
        RECT 1196.265 3498.360 1296.375 3498.500 ;
        RECT 1196.265 3498.315 1196.555 3498.360 ;
        RECT 1296.085 3498.315 1296.375 3498.360 ;
        RECT 1320.465 3498.500 1320.755 3498.545 ;
        RECT 1392.685 3498.500 1392.975 3498.545 ;
        RECT 1320.465 3498.360 1392.975 3498.500 ;
        RECT 1444.740 3498.500 1444.880 3498.700 ;
        RECT 1459.385 3498.700 1479.930 3498.840 ;
        RECT 1459.385 3498.655 1459.675 3498.700 ;
        RECT 1479.610 3498.640 1479.930 3498.700 ;
        RECT 1458.005 3498.500 1458.295 3498.545 ;
        RECT 1444.740 3498.360 1458.295 3498.500 ;
        RECT 1320.465 3498.315 1320.755 3498.360 ;
        RECT 1392.685 3498.315 1392.975 3498.360 ;
        RECT 1458.005 3498.315 1458.295 3498.360 ;
      LAYER via ;
        RECT 1137.860 3498.640 1138.120 3498.900 ;
        RECT 1479.640 3498.640 1479.900 3498.900 ;
      LAYER met2 ;
        RECT 1137.850 3517.600 1138.130 3520.000 ;
        RECT 1137.920 3498.930 1138.060 3517.600 ;
        RECT 1137.860 3498.610 1138.120 3498.930 ;
        RECT 1479.640 3498.610 1479.900 3498.930 ;
        RECT 1479.700 3466.000 1479.840 3498.610 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1461.745 3500.045 1461.915 3501.235 ;
      LAYER mcon ;
        RECT 1461.745 3501.065 1461.915 3501.235 ;
      LAYER met1 ;
        RECT 1461.685 3501.220 1461.975 3501.265 ;
        RECT 1492.950 3501.220 1493.270 3501.280 ;
        RECT 1461.685 3501.080 1493.270 3501.220 ;
        RECT 1461.685 3501.035 1461.975 3501.080 ;
        RECT 1492.950 3501.020 1493.270 3501.080 ;
        RECT 813.070 3500.200 813.390 3500.260 ;
        RECT 1461.685 3500.200 1461.975 3500.245 ;
        RECT 813.070 3500.060 1461.975 3500.200 ;
        RECT 813.070 3500.000 813.390 3500.060 ;
        RECT 1461.685 3500.015 1461.975 3500.060 ;
      LAYER via ;
        RECT 1492.980 3501.020 1493.240 3501.280 ;
        RECT 813.100 3500.000 813.360 3500.260 ;
      LAYER met2 ;
        RECT 813.090 3517.600 813.370 3520.000 ;
        RECT 813.160 3500.290 813.300 3517.600 ;
        RECT 1492.980 3500.990 1493.240 3501.310 ;
        RECT 813.100 3499.970 813.360 3500.290 ;
        RECT 1493.040 3466.000 1493.180 3500.990 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 488.770 3503.940 489.090 3504.000 ;
        RECT 1506.750 3503.940 1507.070 3504.000 ;
        RECT 488.770 3503.800 1507.070 3503.940 ;
        RECT 488.770 3503.740 489.090 3503.800 ;
        RECT 1506.750 3503.740 1507.070 3503.800 ;
      LAYER via ;
        RECT 488.800 3503.740 489.060 3504.000 ;
        RECT 1506.780 3503.740 1507.040 3504.000 ;
      LAYER met2 ;
        RECT 488.790 3517.600 489.070 3520.000 ;
        RECT 488.860 3504.030 489.000 3517.600 ;
        RECT 488.800 3503.710 489.060 3504.030 ;
        RECT 1506.780 3503.710 1507.040 3504.030 ;
        RECT 1506.840 3466.000 1506.980 3503.710 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 164.470 3501.560 164.790 3501.620 ;
        RECT 1527.450 3501.560 1527.770 3501.620 ;
        RECT 164.470 3501.420 1527.770 3501.560 ;
        RECT 164.470 3501.360 164.790 3501.420 ;
        RECT 1527.450 3501.360 1527.770 3501.420 ;
      LAYER via ;
        RECT 164.500 3501.360 164.760 3501.620 ;
        RECT 1527.480 3501.360 1527.740 3501.620 ;
      LAYER met2 ;
        RECT 164.490 3517.600 164.770 3520.000 ;
        RECT 164.560 3501.650 164.700 3517.600 ;
        RECT 164.500 3501.330 164.760 3501.650 ;
        RECT 1527.480 3501.330 1527.740 3501.650 ;
        RECT 1527.540 3466.000 1527.680 3501.330 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.570 3388.000 19.890 3388.060 ;
        RECT 19.570 3387.860 54.000 3388.000 ;
        RECT 19.570 3387.800 19.890 3387.860 ;
      LAYER via ;
        RECT 19.600 3387.800 19.860 3388.060 ;
      LAYER met2 ;
        RECT 19.590 3393.355 19.870 3393.725 ;
        RECT 19.660 3388.090 19.800 3393.355 ;
        RECT 19.600 3387.770 19.860 3388.090 ;
      LAYER via2 ;
        RECT 19.590 3393.400 19.870 3393.680 ;
      LAYER met3 ;
        RECT 2.480 3393.690 4.880 3393.840 ;
        RECT 19.565 3393.690 19.895 3393.705 ;
        RECT 2.480 3393.390 19.895 3393.690 ;
        RECT 2.480 3393.240 4.880 3393.390 ;
        RECT 19.565 3393.375 19.895 3393.390 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.570 3139.800 19.890 3139.860 ;
        RECT 19.570 3139.660 54.000 3139.800 ;
        RECT 19.570 3139.600 19.890 3139.660 ;
      LAYER via ;
        RECT 19.600 3139.600 19.860 3139.860 ;
      LAYER met2 ;
        RECT 19.590 3141.755 19.870 3142.125 ;
        RECT 19.660 3139.890 19.800 3141.755 ;
        RECT 19.600 3139.570 19.860 3139.890 ;
      LAYER via2 ;
        RECT 19.590 3141.800 19.870 3142.080 ;
      LAYER met3 ;
        RECT 2.480 3142.090 4.880 3142.240 ;
        RECT 19.565 3142.090 19.895 3142.105 ;
        RECT 2.480 3141.790 19.895 3142.090 ;
        RECT 2.480 3141.640 4.880 3141.790 ;
        RECT 19.565 3141.775 19.895 3141.790 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.650 2884.460 18.970 2884.520 ;
        RECT 18.650 2884.320 54.000 2884.460 ;
        RECT 18.650 2884.260 18.970 2884.320 ;
      LAYER via ;
        RECT 18.680 2884.260 18.940 2884.520 ;
      LAYER met2 ;
        RECT 18.670 2890.835 18.950 2891.205 ;
        RECT 18.740 2884.550 18.880 2890.835 ;
        RECT 18.680 2884.230 18.940 2884.550 ;
      LAYER via2 ;
        RECT 18.670 2890.880 18.950 2891.160 ;
      LAYER met3 ;
        RECT 2.480 2891.170 4.880 2891.320 ;
        RECT 18.645 2891.170 18.975 2891.185 ;
        RECT 2.480 2890.870 18.975 2891.170 ;
        RECT 2.480 2890.720 4.880 2890.870 ;
        RECT 18.645 2890.855 18.975 2890.870 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.190 2636.260 18.510 2636.320 ;
        RECT 18.190 2636.120 54.000 2636.260 ;
        RECT 18.190 2636.060 18.510 2636.120 ;
      LAYER via ;
        RECT 18.220 2636.060 18.480 2636.320 ;
      LAYER met2 ;
        RECT 18.210 2639.235 18.490 2639.605 ;
        RECT 18.280 2636.350 18.420 2639.235 ;
        RECT 18.220 2636.030 18.480 2636.350 ;
      LAYER via2 ;
        RECT 18.210 2639.280 18.490 2639.560 ;
      LAYER met3 ;
        RECT 2.480 2639.570 4.880 2639.720 ;
        RECT 18.185 2639.570 18.515 2639.585 ;
        RECT 2.480 2639.270 18.515 2639.570 ;
        RECT 2.480 2639.120 4.880 2639.270 ;
        RECT 18.185 2639.255 18.515 2639.270 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.570 2387.720 19.890 2387.780 ;
        RECT 19.570 2387.580 54.000 2387.720 ;
        RECT 19.570 2387.520 19.890 2387.580 ;
      LAYER via ;
        RECT 19.600 2387.520 19.860 2387.780 ;
      LAYER met2 ;
        RECT 19.590 2387.635 19.870 2388.005 ;
        RECT 19.600 2387.490 19.860 2387.635 ;
      LAYER via2 ;
        RECT 19.590 2387.680 19.870 2387.960 ;
      LAYER met3 ;
        RECT 2.480 2387.970 4.880 2388.120 ;
        RECT 19.565 2387.970 19.895 2387.985 ;
        RECT 2.480 2387.670 19.895 2387.970 ;
        RECT 2.480 2387.520 4.880 2387.670 ;
        RECT 19.565 2387.655 19.895 2387.670 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.190 2138.840 18.510 2138.900 ;
        RECT 18.190 2138.700 54.000 2138.840 ;
        RECT 18.190 2138.640 18.510 2138.700 ;
      LAYER via ;
        RECT 18.220 2138.640 18.480 2138.900 ;
      LAYER met2 ;
        RECT 18.220 2138.610 18.480 2138.930 ;
        RECT 18.280 2136.405 18.420 2138.610 ;
        RECT 18.210 2136.035 18.490 2136.405 ;
      LAYER via2 ;
        RECT 18.210 2136.080 18.490 2136.360 ;
      LAYER met3 ;
        RECT 2.480 2136.370 4.880 2136.520 ;
        RECT 18.185 2136.370 18.515 2136.385 ;
        RECT 2.480 2136.070 18.515 2136.370 ;
        RECT 2.480 2135.920 4.880 2136.070 ;
        RECT 18.185 2136.055 18.515 2136.070 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.080 586.650 2922.480 586.800 ;
        RECT 2870.580 586.350 2922.480 586.650 ;
        RECT 2920.080 586.200 2922.480 586.350 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.730 1889.960 18.050 1890.020 ;
        RECT 17.730 1889.820 54.000 1889.960 ;
        RECT 17.730 1889.760 18.050 1889.820 ;
      LAYER via ;
        RECT 17.760 1889.760 18.020 1890.020 ;
      LAYER met2 ;
        RECT 17.760 1889.730 18.020 1890.050 ;
        RECT 17.820 1885.485 17.960 1889.730 ;
        RECT 17.750 1885.115 18.030 1885.485 ;
      LAYER via2 ;
        RECT 17.750 1885.160 18.030 1885.440 ;
      LAYER met3 ;
        RECT 2.480 1885.450 4.880 1885.600 ;
        RECT 17.725 1885.450 18.055 1885.465 ;
        RECT 2.480 1885.150 18.055 1885.450 ;
        RECT 2.480 1885.000 4.880 1885.150 ;
        RECT 17.725 1885.135 18.055 1885.150 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 21.870 2313.940 22.190 2314.000 ;
        RECT 21.870 2313.800 54.000 2313.940 ;
        RECT 21.870 2313.740 22.190 2313.800 ;
      LAYER via ;
        RECT 21.900 2313.740 22.160 2314.000 ;
      LAYER met2 ;
        RECT 21.900 2313.710 22.160 2314.030 ;
        RECT 21.960 1633.885 22.100 2313.710 ;
        RECT 21.890 1633.515 22.170 1633.885 ;
      LAYER via2 ;
        RECT 21.890 1633.560 22.170 1633.840 ;
      LAYER met3 ;
        RECT 2.480 1633.850 4.880 1634.000 ;
        RECT 21.865 1633.850 22.195 1633.865 ;
        RECT 2.480 1633.550 22.195 1633.850 ;
        RECT 2.480 1633.400 4.880 1633.550 ;
        RECT 21.865 1633.535 22.195 1633.550 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 21.410 2313.600 21.730 2313.660 ;
        RECT 21.410 2313.460 54.000 2313.600 ;
        RECT 21.410 2313.400 21.730 2313.460 ;
      LAYER via ;
        RECT 21.440 2313.400 21.700 2313.660 ;
      LAYER met2 ;
        RECT 21.440 2313.370 21.700 2313.690 ;
        RECT 21.500 1382.285 21.640 2313.370 ;
        RECT 21.430 1381.915 21.710 1382.285 ;
      LAYER via2 ;
        RECT 21.430 1381.960 21.710 1382.240 ;
      LAYER met3 ;
        RECT 2.480 1382.250 4.880 1382.400 ;
        RECT 21.405 1382.250 21.735 1382.265 ;
        RECT 2.480 1381.950 21.735 1382.250 ;
        RECT 2.480 1381.800 4.880 1381.950 ;
        RECT 21.405 1381.935 21.735 1381.950 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.950 2313.260 21.270 2313.320 ;
        RECT 20.950 2313.120 54.000 2313.260 ;
        RECT 20.950 2313.060 21.270 2313.120 ;
      LAYER via ;
        RECT 20.980 2313.060 21.240 2313.320 ;
      LAYER met2 ;
        RECT 20.980 2313.030 21.240 2313.350 ;
        RECT 21.040 1131.365 21.180 2313.030 ;
        RECT 20.970 1130.995 21.250 1131.365 ;
      LAYER via2 ;
        RECT 20.970 1131.040 21.250 1131.320 ;
      LAYER met3 ;
        RECT 2.480 1131.330 4.880 1131.480 ;
        RECT 20.945 1131.330 21.275 1131.345 ;
        RECT 2.480 1131.030 21.275 1131.330 ;
        RECT 2.480 1130.880 4.880 1131.030 ;
        RECT 20.945 1131.015 21.275 1131.030 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.490 2312.580 20.810 2312.640 ;
        RECT 20.490 2312.440 54.000 2312.580 ;
        RECT 20.490 2312.380 20.810 2312.440 ;
      LAYER via ;
        RECT 20.520 2312.380 20.780 2312.640 ;
      LAYER met2 ;
        RECT 20.520 2312.350 20.780 2312.670 ;
        RECT 20.580 879.765 20.720 2312.350 ;
        RECT 20.510 879.395 20.790 879.765 ;
      LAYER via2 ;
        RECT 20.510 879.440 20.790 879.720 ;
      LAYER met3 ;
        RECT 2.480 879.730 4.880 879.880 ;
        RECT 20.485 879.730 20.815 879.745 ;
        RECT 2.480 879.430 20.815 879.730 ;
        RECT 2.480 879.280 4.880 879.430 ;
        RECT 20.485 879.415 20.815 879.430 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 20.050 634.595 20.330 634.965 ;
        RECT 20.120 628.165 20.260 634.595 ;
        RECT 20.050 627.795 20.330 628.165 ;
      LAYER via2 ;
        RECT 20.050 634.640 20.330 634.920 ;
        RECT 20.050 627.840 20.330 628.120 ;
      LAYER met3 ;
        RECT 20.025 634.930 20.355 634.945 ;
        RECT 20.025 634.630 54.000 634.930 ;
        RECT 20.025 634.615 20.355 634.630 ;
        RECT 2.480 628.130 4.880 628.280 ;
        RECT 20.025 628.130 20.355 628.145 ;
        RECT 2.480 627.830 20.355 628.130 ;
        RECT 2.480 627.680 4.880 627.830 ;
        RECT 20.025 627.815 20.355 627.830 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5.550 378.950 54.000 379.250 ;
        RECT 2.480 376.530 4.880 376.680 ;
        RECT 5.550 376.530 5.850 378.950 ;
        RECT 2.480 376.230 5.850 376.530 ;
        RECT 2.480 376.080 4.880 376.230 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.570 131.140 19.890 131.200 ;
        RECT 19.570 131.000 54.000 131.140 ;
        RECT 19.570 130.940 19.890 131.000 ;
      LAYER via ;
        RECT 19.600 130.940 19.860 131.200 ;
      LAYER met2 ;
        RECT 19.600 130.910 19.860 131.230 ;
        RECT 19.660 125.645 19.800 130.910 ;
        RECT 19.590 125.275 19.870 125.645 ;
      LAYER via2 ;
        RECT 19.590 125.320 19.870 125.600 ;
      LAYER met3 ;
        RECT 2.480 125.610 4.880 125.760 ;
        RECT 19.565 125.610 19.895 125.625 ;
        RECT 2.480 125.310 19.895 125.610 ;
        RECT 2.480 125.160 4.880 125.310 ;
        RECT 19.565 125.295 19.895 125.310 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.080 821.250 2922.480 821.400 ;
        RECT 2870.580 820.950 2922.480 821.250 ;
        RECT 2920.080 820.800 2922.480 820.950 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.080 1055.850 2922.480 1056.000 ;
        RECT 2870.580 1055.550 2922.480 1055.850 ;
        RECT 2920.080 1055.400 2922.480 1055.550 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.080 1290.450 2922.480 1290.600 ;
        RECT 2870.580 1290.150 2922.480 1290.450 ;
        RECT 2920.080 1290.000 2922.480 1290.150 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.080 1525.050 2922.480 1525.200 ;
        RECT 2870.580 1524.750 2922.480 1525.050 ;
        RECT 2920.080 1524.600 2922.480 1524.750 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2903.310 1766.200 2903.630 1766.260 ;
        RECT 2870.580 1766.060 2903.630 1766.200 ;
        RECT 2903.310 1766.000 2903.630 1766.060 ;
      LAYER via ;
        RECT 2903.340 1766.000 2903.600 1766.260 ;
      LAYER met2 ;
        RECT 2903.340 1765.970 2903.600 1766.290 ;
        RECT 2903.400 1759.685 2903.540 1765.970 ;
        RECT 2903.330 1759.315 2903.610 1759.685 ;
      LAYER via2 ;
        RECT 2903.330 1759.360 2903.610 1759.640 ;
      LAYER met3 ;
        RECT 2903.305 1759.650 2903.635 1759.665 ;
        RECT 2920.080 1759.650 2922.480 1759.800 ;
        RECT 2903.305 1759.350 2922.480 1759.650 ;
        RECT 2903.305 1759.335 2903.635 1759.350 ;
        RECT 2920.080 1759.200 2922.480 1759.350 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2903.310 2000.800 2903.630 2000.860 ;
        RECT 2870.580 2000.660 2903.630 2000.800 ;
        RECT 2903.310 2000.600 2903.630 2000.660 ;
      LAYER via ;
        RECT 2903.340 2000.600 2903.600 2000.860 ;
      LAYER met2 ;
        RECT 2903.340 2000.570 2903.600 2000.890 ;
        RECT 2903.400 1994.285 2903.540 2000.570 ;
        RECT 2903.330 1993.915 2903.610 1994.285 ;
      LAYER via2 ;
        RECT 2903.330 1993.960 2903.610 1994.240 ;
      LAYER met3 ;
        RECT 2903.305 1994.250 2903.635 1994.265 ;
        RECT 2920.080 1994.250 2922.480 1994.400 ;
        RECT 2903.305 1993.950 2922.480 1994.250 ;
        RECT 2903.305 1993.935 2903.635 1993.950 ;
        RECT 2920.080 1993.800 2922.480 1993.950 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2903.310 2235.400 2903.630 2235.460 ;
        RECT 2870.580 2235.260 2903.630 2235.400 ;
        RECT 2903.310 2235.200 2903.630 2235.260 ;
      LAYER via ;
        RECT 2903.340 2235.200 2903.600 2235.460 ;
      LAYER met2 ;
        RECT 2903.340 2235.170 2903.600 2235.490 ;
        RECT 2903.400 2228.885 2903.540 2235.170 ;
        RECT 2903.330 2228.515 2903.610 2228.885 ;
      LAYER via2 ;
        RECT 2903.330 2228.560 2903.610 2228.840 ;
      LAYER met3 ;
        RECT 2903.305 2228.850 2903.635 2228.865 ;
        RECT 2920.080 2228.850 2922.480 2229.000 ;
        RECT 2903.305 2228.550 2922.480 2228.850 ;
        RECT 2903.305 2228.535 2903.635 2228.550 ;
        RECT 2920.080 2228.400 2922.480 2228.550 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 636.980 16.730 637.120 54.000 ;
        RECT 635.600 16.590 637.120 16.730 ;
        RECT 635.600 2.400 635.740 16.590 ;
        RECT 635.530 0.000 635.810 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2419.940 2.400 2420.080 54.000 ;
        RECT 2419.870 0.000 2420.150 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2431.350 35.940 2431.670 36.000 ;
        RECT 2437.330 35.940 2437.650 36.000 ;
        RECT 2431.350 35.800 2437.650 35.940 ;
        RECT 2431.350 35.740 2431.670 35.800 ;
        RECT 2437.330 35.740 2437.650 35.800 ;
      LAYER via ;
        RECT 2431.380 35.740 2431.640 36.000 ;
        RECT 2437.360 35.740 2437.620 36.000 ;
      LAYER met2 ;
        RECT 2431.440 36.030 2431.580 54.000 ;
        RECT 2431.380 35.710 2431.640 36.030 ;
        RECT 2437.360 35.710 2437.620 36.030 ;
        RECT 2437.420 2.400 2437.560 35.710 ;
        RECT 2437.350 0.000 2437.630 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2452.050 2.960 2452.370 3.020 ;
        RECT 2455.270 2.960 2455.590 3.020 ;
        RECT 2452.050 2.820 2455.590 2.960 ;
        RECT 2452.050 2.760 2452.370 2.820 ;
        RECT 2455.270 2.760 2455.590 2.820 ;
      LAYER via ;
        RECT 2452.080 2.760 2452.340 3.020 ;
        RECT 2455.300 2.760 2455.560 3.020 ;
      LAYER met2 ;
        RECT 2452.140 3.050 2452.280 54.000 ;
        RECT 2452.080 2.730 2452.340 3.050 ;
        RECT 2455.300 2.730 2455.560 3.050 ;
        RECT 2455.360 2.400 2455.500 2.730 ;
        RECT 2455.290 0.000 2455.570 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2472.840 2.960 2472.980 54.000 ;
        RECT 2472.840 2.820 2473.440 2.960 ;
        RECT 2473.300 2.400 2473.440 2.820 ;
        RECT 2473.230 0.000 2473.510 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2486.550 2.960 2486.870 3.020 ;
        RECT 2491.150 2.960 2491.470 3.020 ;
        RECT 2486.550 2.820 2491.470 2.960 ;
        RECT 2486.550 2.760 2486.870 2.820 ;
        RECT 2491.150 2.760 2491.470 2.820 ;
      LAYER via ;
        RECT 2486.580 2.760 2486.840 3.020 ;
        RECT 2491.180 2.760 2491.440 3.020 ;
      LAYER met2 ;
        RECT 2486.640 3.050 2486.780 54.000 ;
        RECT 2486.580 2.730 2486.840 3.050 ;
        RECT 2491.180 2.730 2491.440 3.050 ;
        RECT 2491.240 2.400 2491.380 2.730 ;
        RECT 2491.170 0.000 2491.450 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2507.250 2.960 2507.570 3.020 ;
        RECT 2508.630 2.960 2508.950 3.020 ;
        RECT 2507.250 2.820 2508.950 2.960 ;
        RECT 2507.250 2.760 2507.570 2.820 ;
        RECT 2508.630 2.760 2508.950 2.820 ;
      LAYER via ;
        RECT 2507.280 2.760 2507.540 3.020 ;
        RECT 2508.660 2.760 2508.920 3.020 ;
      LAYER met2 ;
        RECT 2507.340 3.050 2507.480 54.000 ;
        RECT 2507.280 2.730 2507.540 3.050 ;
        RECT 2508.660 2.730 2508.920 3.050 ;
        RECT 2508.720 2.400 2508.860 2.730 ;
        RECT 2508.650 0.000 2508.930 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2521.050 2.960 2521.370 3.020 ;
        RECT 2526.570 2.960 2526.890 3.020 ;
        RECT 2521.050 2.820 2526.890 2.960 ;
        RECT 2521.050 2.760 2521.370 2.820 ;
        RECT 2526.570 2.760 2526.890 2.820 ;
      LAYER via ;
        RECT 2521.080 2.760 2521.340 3.020 ;
        RECT 2526.600 2.760 2526.860 3.020 ;
      LAYER met2 ;
        RECT 2521.140 3.050 2521.280 54.000 ;
        RECT 2521.080 2.730 2521.340 3.050 ;
        RECT 2526.600 2.730 2526.860 3.050 ;
        RECT 2526.660 2.400 2526.800 2.730 ;
        RECT 2526.590 0.000 2526.870 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2541.750 2.960 2542.070 3.020 ;
        RECT 2544.510 2.960 2544.830 3.020 ;
        RECT 2541.750 2.820 2544.830 2.960 ;
        RECT 2541.750 2.760 2542.070 2.820 ;
        RECT 2544.510 2.760 2544.830 2.820 ;
      LAYER via ;
        RECT 2541.780 2.760 2542.040 3.020 ;
        RECT 2544.540 2.760 2544.800 3.020 ;
      LAYER met2 ;
        RECT 2541.840 3.050 2541.980 54.000 ;
        RECT 2541.780 2.730 2542.040 3.050 ;
        RECT 2544.540 2.730 2544.800 3.050 ;
        RECT 2544.600 2.400 2544.740 2.730 ;
        RECT 2544.530 0.000 2544.810 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2528.025 20.145 2528.195 25.075 ;
      LAYER mcon ;
        RECT 2528.025 24.905 2528.195 25.075 ;
      LAYER met1 ;
        RECT 1678.790 25.060 1679.110 25.120 ;
        RECT 2527.965 25.060 2528.255 25.105 ;
        RECT 1678.790 24.920 2528.255 25.060 ;
        RECT 1678.790 24.860 1679.110 24.920 ;
        RECT 2527.965 24.875 2528.255 24.920 ;
        RECT 2527.965 20.300 2528.255 20.345 ;
        RECT 2562.450 20.300 2562.770 20.360 ;
        RECT 2527.965 20.160 2562.770 20.300 ;
        RECT 2527.965 20.115 2528.255 20.160 ;
        RECT 2562.450 20.100 2562.770 20.160 ;
      LAYER via ;
        RECT 1678.820 24.860 1679.080 25.120 ;
        RECT 2562.480 20.100 2562.740 20.360 ;
      LAYER met2 ;
        RECT 1678.880 25.150 1679.020 54.000 ;
        RECT 1678.820 24.830 1679.080 25.150 ;
        RECT 2562.480 20.070 2562.740 20.390 ;
        RECT 2562.540 2.400 2562.680 20.070 ;
        RECT 2562.470 0.000 2562.750 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1727.165 23.205 1727.335 25.415 ;
        RECT 2528.945 19.805 2529.115 25.415 ;
      LAYER mcon ;
        RECT 1727.165 25.245 1727.335 25.415 ;
        RECT 2528.945 25.245 2529.115 25.415 ;
      LAYER met1 ;
        RECT 1727.105 25.400 1727.395 25.445 ;
        RECT 2528.885 25.400 2529.175 25.445 ;
        RECT 1727.105 25.260 2529.175 25.400 ;
        RECT 1727.105 25.215 1727.395 25.260 ;
        RECT 2528.885 25.215 2529.175 25.260 ;
        RECT 1685.690 23.360 1686.010 23.420 ;
        RECT 1727.105 23.360 1727.395 23.405 ;
        RECT 1685.690 23.220 1727.395 23.360 ;
        RECT 1685.690 23.160 1686.010 23.220 ;
        RECT 1727.105 23.175 1727.395 23.220 ;
        RECT 2528.885 19.960 2529.175 20.005 ;
        RECT 2580.390 19.960 2580.710 20.020 ;
        RECT 2528.885 19.820 2580.710 19.960 ;
        RECT 2528.885 19.775 2529.175 19.820 ;
        RECT 2580.390 19.760 2580.710 19.820 ;
      LAYER via ;
        RECT 1685.720 23.160 1685.980 23.420 ;
        RECT 2580.420 19.760 2580.680 20.020 ;
      LAYER met2 ;
        RECT 1685.780 23.450 1685.920 54.000 ;
        RECT 1685.720 23.130 1685.980 23.450 ;
        RECT 2580.420 19.730 2580.680 20.050 ;
        RECT 2580.480 2.400 2580.620 19.730 ;
        RECT 2580.410 0.000 2580.690 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 813.990 18.260 814.310 18.320 ;
        RECT 816.290 18.260 816.610 18.320 ;
        RECT 813.990 18.120 816.610 18.260 ;
        RECT 813.990 18.060 814.310 18.120 ;
        RECT 816.290 18.060 816.610 18.120 ;
      LAYER via ;
        RECT 814.020 18.060 814.280 18.320 ;
        RECT 816.320 18.060 816.580 18.320 ;
      LAYER met2 ;
        RECT 816.380 18.350 816.520 54.000 ;
        RECT 814.020 18.030 814.280 18.350 ;
        RECT 816.320 18.030 816.580 18.350 ;
        RECT 814.080 2.400 814.220 18.030 ;
        RECT 814.010 0.000 814.290 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1706.925 26.435 1707.095 26.775 ;
        RECT 1706.465 26.265 1707.095 26.435 ;
        RECT 1731.765 23.885 1731.935 26.775 ;
      LAYER mcon ;
        RECT 1706.925 26.605 1707.095 26.775 ;
        RECT 1731.765 26.605 1731.935 26.775 ;
      LAYER met1 ;
        RECT 1706.865 26.760 1707.155 26.805 ;
        RECT 1731.705 26.760 1731.995 26.805 ;
        RECT 1706.865 26.620 1731.995 26.760 ;
        RECT 1706.865 26.575 1707.155 26.620 ;
        RECT 1731.705 26.575 1731.995 26.620 ;
        RECT 1690.290 26.420 1690.610 26.480 ;
        RECT 1706.405 26.420 1706.695 26.465 ;
        RECT 1690.290 26.280 1706.695 26.420 ;
        RECT 1690.290 26.220 1690.610 26.280 ;
        RECT 1706.405 26.235 1706.695 26.280 ;
        RECT 1731.705 24.040 1731.995 24.085 ;
        RECT 2576.250 24.040 2576.570 24.100 ;
        RECT 1731.705 23.900 2576.570 24.040 ;
        RECT 1731.705 23.855 1731.995 23.900 ;
        RECT 2576.250 23.840 2576.570 23.900 ;
      LAYER via ;
        RECT 1690.320 26.220 1690.580 26.480 ;
        RECT 2576.280 23.840 2576.540 24.100 ;
      LAYER met2 ;
        RECT 1690.380 26.510 1690.520 54.000 ;
        RECT 1690.320 26.190 1690.580 26.510 ;
        RECT 2576.280 23.810 2576.540 24.130 ;
        RECT 2576.340 23.645 2576.480 23.810 ;
        RECT 2576.270 23.275 2576.550 23.645 ;
        RECT 2597.890 23.275 2598.170 23.645 ;
        RECT 2597.960 2.400 2598.100 23.275 ;
        RECT 2597.890 0.000 2598.170 2.400 ;
      LAYER via2 ;
        RECT 2576.270 23.320 2576.550 23.600 ;
        RECT 2597.890 23.320 2598.170 23.600 ;
      LAYER met3 ;
        RECT 2576.245 23.610 2576.575 23.625 ;
        RECT 2597.865 23.610 2598.195 23.625 ;
        RECT 2576.245 23.310 2598.195 23.610 ;
        RECT 2576.245 23.295 2576.575 23.310 ;
        RECT 2597.865 23.295 2598.195 23.310 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2576.325 20.655 2576.495 20.995 ;
        RECT 2576.325 20.485 2577.415 20.655 ;
      LAYER mcon ;
        RECT 2576.325 20.825 2576.495 20.995 ;
        RECT 2577.245 20.485 2577.415 20.655 ;
      LAYER met1 ;
        RECT 1692.130 20.980 1692.450 21.040 ;
        RECT 2576.265 20.980 2576.555 21.025 ;
        RECT 2615.810 20.980 2616.130 21.040 ;
        RECT 1692.130 20.840 2576.555 20.980 ;
        RECT 1692.130 20.780 1692.450 20.840 ;
        RECT 2576.265 20.795 2576.555 20.840 ;
        RECT 2580.940 20.840 2616.130 20.980 ;
        RECT 2577.185 20.640 2577.475 20.685 ;
        RECT 2580.940 20.640 2581.080 20.840 ;
        RECT 2615.810 20.780 2616.130 20.840 ;
        RECT 2577.185 20.500 2581.080 20.640 ;
        RECT 2577.185 20.455 2577.475 20.500 ;
      LAYER via ;
        RECT 1692.160 20.780 1692.420 21.040 ;
        RECT 2615.840 20.780 2616.100 21.040 ;
      LAYER met2 ;
        RECT 1692.220 21.070 1692.360 54.000 ;
        RECT 1692.160 20.750 1692.420 21.070 ;
        RECT 2615.840 20.750 2616.100 21.070 ;
        RECT 2615.900 2.400 2616.040 20.750 ;
        RECT 2615.830 0.000 2616.110 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1731.305 21.165 1731.475 24.055 ;
      LAYER mcon ;
        RECT 1731.305 23.885 1731.475 24.055 ;
      LAYER met1 ;
        RECT 1699.030 24.040 1699.350 24.100 ;
        RECT 1731.245 24.040 1731.535 24.085 ;
        RECT 1699.030 23.900 1731.535 24.040 ;
        RECT 1699.030 23.840 1699.350 23.900 ;
        RECT 1731.245 23.855 1731.535 23.900 ;
        RECT 2576.710 24.040 2577.030 24.100 ;
        RECT 2633.750 24.040 2634.070 24.100 ;
        RECT 2576.710 23.900 2634.070 24.040 ;
        RECT 2576.710 23.840 2577.030 23.900 ;
        RECT 2633.750 23.840 2634.070 23.900 ;
        RECT 1731.245 21.320 1731.535 21.365 ;
        RECT 2576.710 21.320 2577.030 21.380 ;
        RECT 1731.245 21.180 2577.030 21.320 ;
        RECT 1731.245 21.135 1731.535 21.180 ;
        RECT 2576.710 21.120 2577.030 21.180 ;
      LAYER via ;
        RECT 1699.060 23.840 1699.320 24.100 ;
        RECT 2576.740 23.840 2577.000 24.100 ;
        RECT 2633.780 23.840 2634.040 24.100 ;
        RECT 2576.740 21.120 2577.000 21.380 ;
      LAYER met2 ;
        RECT 1699.120 24.130 1699.260 54.000 ;
        RECT 1699.060 23.810 1699.320 24.130 ;
        RECT 2576.740 23.810 2577.000 24.130 ;
        RECT 2633.780 23.810 2634.040 24.130 ;
        RECT 2576.800 21.410 2576.940 23.810 ;
        RECT 2576.740 21.090 2577.000 21.410 ;
        RECT 2633.840 2.400 2633.980 23.810 ;
        RECT 2633.770 0.000 2634.050 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1730.845 21.165 1731.015 22.355 ;
      LAYER mcon ;
        RECT 1730.845 22.185 1731.015 22.355 ;
      LAYER met1 ;
        RECT 1730.785 22.340 1731.075 22.385 ;
        RECT 2651.690 22.340 2652.010 22.400 ;
        RECT 1730.785 22.200 2652.010 22.340 ;
        RECT 1730.785 22.155 1731.075 22.200 ;
        RECT 2651.690 22.140 2652.010 22.200 ;
        RECT 1697.190 21.320 1697.510 21.380 ;
        RECT 1730.785 21.320 1731.075 21.365 ;
        RECT 1697.190 21.180 1731.075 21.320 ;
        RECT 1697.190 21.120 1697.510 21.180 ;
        RECT 1730.785 21.135 1731.075 21.180 ;
      LAYER via ;
        RECT 2651.720 22.140 2651.980 22.400 ;
        RECT 1697.220 21.120 1697.480 21.380 ;
      LAYER met2 ;
        RECT 1697.280 21.410 1697.420 54.000 ;
        RECT 2651.720 22.110 2651.980 22.430 ;
        RECT 1697.220 21.090 1697.480 21.410 ;
        RECT 2651.780 2.400 2651.920 22.110 ;
        RECT 2651.710 0.000 2651.990 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1732.685 22.525 1732.855 46.835 ;
      LAYER mcon ;
        RECT 1732.685 46.665 1732.855 46.835 ;
      LAYER met1 ;
        RECT 1706.390 46.820 1706.710 46.880 ;
        RECT 1732.625 46.820 1732.915 46.865 ;
        RECT 1706.390 46.680 1732.915 46.820 ;
        RECT 1706.390 46.620 1706.710 46.680 ;
        RECT 1732.625 46.635 1732.915 46.680 ;
        RECT 1732.625 22.680 1732.915 22.725 ;
        RECT 2669.630 22.680 2669.950 22.740 ;
        RECT 1732.625 22.540 2669.950 22.680 ;
        RECT 1732.625 22.495 1732.915 22.540 ;
        RECT 2669.630 22.480 2669.950 22.540 ;
      LAYER via ;
        RECT 1706.420 46.620 1706.680 46.880 ;
        RECT 2669.660 22.480 2669.920 22.740 ;
      LAYER met2 ;
        RECT 1706.480 46.910 1706.620 54.000 ;
        RECT 1706.420 46.590 1706.680 46.910 ;
        RECT 2669.660 22.450 2669.920 22.770 ;
        RECT 2669.720 2.400 2669.860 22.450 ;
        RECT 2669.650 0.000 2669.930 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2648.085 21.165 2648.255 23.035 ;
      LAYER mcon ;
        RECT 2648.085 22.865 2648.255 23.035 ;
      LAYER met1 ;
        RECT 1704.550 23.700 1704.870 23.760 ;
        RECT 1704.550 23.560 1727.780 23.700 ;
        RECT 1704.550 23.500 1704.870 23.560 ;
        RECT 1727.640 23.020 1727.780 23.560 ;
        RECT 2648.025 23.020 2648.315 23.065 ;
        RECT 1727.640 22.880 2648.315 23.020 ;
        RECT 2648.025 22.835 2648.315 22.880 ;
        RECT 2648.025 21.320 2648.315 21.365 ;
        RECT 2687.110 21.320 2687.430 21.380 ;
        RECT 2648.025 21.180 2687.430 21.320 ;
        RECT 2648.025 21.135 2648.315 21.180 ;
        RECT 2687.110 21.120 2687.430 21.180 ;
      LAYER via ;
        RECT 1704.580 23.500 1704.840 23.760 ;
        RECT 2687.140 21.120 2687.400 21.380 ;
      LAYER met2 ;
        RECT 1703.720 48.805 1703.860 54.000 ;
        RECT 1703.650 48.435 1703.930 48.805 ;
        RECT 1704.570 48.435 1704.850 48.805 ;
        RECT 1704.640 23.790 1704.780 48.435 ;
        RECT 1704.580 23.470 1704.840 23.790 ;
        RECT 2687.140 21.090 2687.400 21.410 ;
        RECT 2687.200 2.400 2687.340 21.090 ;
        RECT 2687.130 0.000 2687.410 2.400 ;
      LAYER via2 ;
        RECT 1703.650 48.480 1703.930 48.760 ;
        RECT 1704.570 48.480 1704.850 48.760 ;
      LAYER met3 ;
        RECT 1703.625 48.770 1703.955 48.785 ;
        RECT 1704.545 48.770 1704.875 48.785 ;
        RECT 1703.625 48.470 1704.875 48.770 ;
        RECT 1703.625 48.455 1703.955 48.470 ;
        RECT 1704.545 48.455 1704.875 48.470 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1754.230 23.360 1754.550 23.420 ;
        RECT 1754.230 23.220 2648.700 23.360 ;
        RECT 1754.230 23.160 1754.550 23.220 ;
        RECT 2648.560 23.020 2648.700 23.220 ;
        RECT 2705.050 23.020 2705.370 23.080 ;
        RECT 2648.560 22.880 2705.370 23.020 ;
        RECT 2705.050 22.820 2705.370 22.880 ;
      LAYER via ;
        RECT 1754.260 23.160 1754.520 23.420 ;
        RECT 2705.080 22.820 2705.340 23.080 ;
      LAYER met2 ;
        RECT 1713.380 22.285 1713.520 54.000 ;
        RECT 1754.260 23.130 1754.520 23.450 ;
        RECT 1754.320 22.285 1754.460 23.130 ;
        RECT 2705.080 22.790 2705.340 23.110 ;
        RECT 1713.310 21.915 1713.590 22.285 ;
        RECT 1754.250 21.915 1754.530 22.285 ;
        RECT 2705.140 2.400 2705.280 22.790 ;
        RECT 2705.070 0.000 2705.350 2.400 ;
      LAYER via2 ;
        RECT 1713.310 21.960 1713.590 22.240 ;
        RECT 1754.250 21.960 1754.530 22.240 ;
      LAYER met3 ;
        RECT 1713.285 22.250 1713.615 22.265 ;
        RECT 1754.225 22.250 1754.555 22.265 ;
        RECT 1713.285 21.950 1754.555 22.250 ;
        RECT 1713.285 21.935 1713.615 21.950 ;
        RECT 1754.225 21.935 1754.555 21.950 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1712.830 25.400 1713.150 25.460 ;
        RECT 1726.630 25.400 1726.950 25.460 ;
        RECT 1712.830 25.260 1726.950 25.400 ;
        RECT 1712.830 25.200 1713.150 25.260 ;
        RECT 1726.630 25.200 1726.950 25.260 ;
        RECT 1754.690 23.700 1755.010 23.760 ;
        RECT 2722.990 23.700 2723.310 23.760 ;
        RECT 1754.690 23.560 2723.310 23.700 ;
        RECT 1754.690 23.500 1755.010 23.560 ;
        RECT 2722.990 23.500 2723.310 23.560 ;
      LAYER via ;
        RECT 1712.860 25.200 1713.120 25.460 ;
        RECT 1726.660 25.200 1726.920 25.460 ;
        RECT 1754.720 23.500 1754.980 23.760 ;
        RECT 2723.020 23.500 2723.280 23.760 ;
      LAYER met2 ;
        RECT 1712.920 25.490 1713.060 54.000 ;
        RECT 1712.860 25.170 1713.120 25.490 ;
        RECT 1726.660 25.170 1726.920 25.490 ;
        RECT 1726.720 22.965 1726.860 25.170 ;
        RECT 1754.720 23.470 1754.980 23.790 ;
        RECT 2723.020 23.470 2723.280 23.790 ;
        RECT 1754.780 22.965 1754.920 23.470 ;
        RECT 1726.650 22.595 1726.930 22.965 ;
        RECT 1754.710 22.595 1754.990 22.965 ;
        RECT 2723.080 2.400 2723.220 23.470 ;
        RECT 2723.010 0.000 2723.290 2.400 ;
      LAYER via2 ;
        RECT 1726.650 22.640 1726.930 22.920 ;
        RECT 1754.710 22.640 1754.990 22.920 ;
      LAYER met3 ;
        RECT 1726.625 22.930 1726.955 22.945 ;
        RECT 1754.685 22.930 1755.015 22.945 ;
        RECT 1726.625 22.630 1755.015 22.930 ;
        RECT 1726.625 22.615 1726.955 22.630 ;
        RECT 1754.685 22.615 1755.015 22.630 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1726.705 26.945 1732.395 27.115 ;
        RECT 1726.705 26.265 1726.875 26.945 ;
        RECT 1732.225 26.605 1732.395 26.945 ;
      LAYER met1 ;
        RECT 1732.165 26.760 1732.455 26.805 ;
        RECT 2740.930 26.760 2741.250 26.820 ;
        RECT 1732.165 26.620 2741.250 26.760 ;
        RECT 1732.165 26.575 1732.455 26.620 ;
        RECT 2740.930 26.560 2741.250 26.620 ;
        RECT 1717.890 26.420 1718.210 26.480 ;
        RECT 1726.645 26.420 1726.935 26.465 ;
        RECT 1717.890 26.280 1726.935 26.420 ;
        RECT 1717.890 26.220 1718.210 26.280 ;
        RECT 1726.645 26.235 1726.935 26.280 ;
      LAYER via ;
        RECT 2740.960 26.560 2741.220 26.820 ;
        RECT 1717.920 26.220 1718.180 26.480 ;
      LAYER met2 ;
        RECT 1717.980 26.510 1718.120 54.000 ;
        RECT 2740.960 26.530 2741.220 26.850 ;
        RECT 1717.920 26.190 1718.180 26.510 ;
        RECT 2741.020 2.400 2741.160 26.530 ;
        RECT 2740.950 0.000 2741.230 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2758.410 26.420 2758.730 26.480 ;
        RECT 1730.860 26.280 2758.730 26.420 ;
        RECT 1719.730 25.740 1720.050 25.800 ;
        RECT 1730.860 25.740 1731.000 26.280 ;
        RECT 2758.410 26.220 2758.730 26.280 ;
        RECT 1719.730 25.600 1731.000 25.740 ;
        RECT 1719.730 25.540 1720.050 25.600 ;
      LAYER via ;
        RECT 1719.760 25.540 1720.020 25.800 ;
        RECT 2758.440 26.220 2758.700 26.480 ;
      LAYER met2 ;
        RECT 1719.820 25.830 1719.960 54.000 ;
        RECT 2758.440 26.190 2758.700 26.510 ;
        RECT 1719.760 25.510 1720.020 25.830 ;
        RECT 2758.500 2.400 2758.640 26.190 ;
        RECT 2758.430 0.000 2758.710 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 831.930 18.260 832.250 18.320 ;
        RECT 836.070 18.260 836.390 18.320 ;
        RECT 831.930 18.120 836.390 18.260 ;
        RECT 831.930 18.060 832.250 18.120 ;
        RECT 836.070 18.060 836.390 18.120 ;
      LAYER via ;
        RECT 831.960 18.060 832.220 18.320 ;
        RECT 836.100 18.060 836.360 18.320 ;
      LAYER met2 ;
        RECT 831.960 18.030 832.220 18.350 ;
        RECT 836.100 18.090 836.360 18.350 ;
        RECT 837.080 18.090 837.220 54.000 ;
        RECT 836.100 18.030 837.220 18.090 ;
        RECT 832.020 2.400 832.160 18.030 ;
        RECT 836.160 17.950 837.220 18.030 ;
        RECT 831.950 0.000 832.230 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1730.385 25.755 1730.555 26.435 ;
        RECT 1730.385 25.585 1731.475 25.755 ;
      LAYER mcon ;
        RECT 1730.385 26.265 1730.555 26.435 ;
        RECT 1731.305 25.585 1731.475 25.755 ;
      LAYER met1 ;
        RECT 1727.090 26.420 1727.410 26.480 ;
        RECT 1730.325 26.420 1730.615 26.465 ;
        RECT 1727.090 26.280 1730.615 26.420 ;
        RECT 1727.090 26.220 1727.410 26.280 ;
        RECT 1730.325 26.235 1730.615 26.280 ;
        RECT 2776.350 26.080 2776.670 26.140 ;
        RECT 1731.780 25.940 2776.670 26.080 ;
        RECT 1731.245 25.740 1731.535 25.785 ;
        RECT 1731.780 25.740 1731.920 25.940 ;
        RECT 2776.350 25.880 2776.670 25.940 ;
        RECT 1731.245 25.600 1731.920 25.740 ;
        RECT 1731.245 25.555 1731.535 25.600 ;
      LAYER via ;
        RECT 1727.120 26.220 1727.380 26.480 ;
        RECT 2776.380 25.880 2776.640 26.140 ;
      LAYER met2 ;
        RECT 1727.180 26.510 1727.320 54.000 ;
        RECT 1727.120 26.190 1727.380 26.510 ;
        RECT 2776.380 25.850 2776.640 26.170 ;
        RECT 2776.440 2.400 2776.580 25.850 ;
        RECT 2776.370 0.000 2776.650 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1754.690 25.740 1755.010 25.800 ;
        RECT 2794.290 25.740 2794.610 25.800 ;
        RECT 1754.690 25.600 2794.610 25.740 ;
        RECT 1754.690 25.540 1755.010 25.600 ;
        RECT 2794.290 25.540 2794.610 25.600 ;
      LAYER via ;
        RECT 1754.720 25.540 1754.980 25.800 ;
        RECT 2794.320 25.540 2794.580 25.800 ;
      LAYER met2 ;
        RECT 1726.720 26.365 1726.860 54.000 ;
        RECT 1726.650 25.995 1726.930 26.365 ;
        RECT 1754.710 25.995 1754.990 26.365 ;
        RECT 1754.780 25.830 1754.920 25.995 ;
        RECT 1754.720 25.510 1754.980 25.830 ;
        RECT 2794.320 25.510 2794.580 25.830 ;
        RECT 2794.380 2.400 2794.520 25.510 ;
        RECT 2794.310 0.000 2794.590 2.400 ;
      LAYER via2 ;
        RECT 1726.650 26.040 1726.930 26.320 ;
        RECT 1754.710 26.040 1754.990 26.320 ;
      LAYER met3 ;
        RECT 1726.625 26.330 1726.955 26.345 ;
        RECT 1754.685 26.330 1755.015 26.345 ;
        RECT 1726.625 26.030 1755.015 26.330 ;
        RECT 1726.625 26.015 1726.955 26.030 ;
        RECT 1754.685 26.015 1755.015 26.030 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2529.405 25.245 2529.575 27.795 ;
      LAYER mcon ;
        RECT 2529.405 27.625 2529.575 27.795 ;
      LAYER met1 ;
        RECT 1854.510 27.780 1854.830 27.840 ;
        RECT 2529.345 27.780 2529.635 27.825 ;
        RECT 1854.510 27.640 2529.635 27.780 ;
        RECT 1854.510 27.580 1854.830 27.640 ;
        RECT 2529.345 27.595 2529.635 27.640 ;
        RECT 1733.990 25.740 1734.310 25.800 ;
        RECT 1754.230 25.740 1754.550 25.800 ;
        RECT 1733.990 25.600 1754.550 25.740 ;
        RECT 1733.990 25.540 1734.310 25.600 ;
        RECT 1754.230 25.540 1754.550 25.600 ;
        RECT 2529.345 25.400 2529.635 25.445 ;
        RECT 2812.230 25.400 2812.550 25.460 ;
        RECT 2529.345 25.260 2812.550 25.400 ;
        RECT 2529.345 25.215 2529.635 25.260 ;
        RECT 2812.230 25.200 2812.550 25.260 ;
      LAYER via ;
        RECT 1854.540 27.580 1854.800 27.840 ;
        RECT 1734.020 25.540 1734.280 25.800 ;
        RECT 1754.260 25.540 1754.520 25.800 ;
        RECT 2812.260 25.200 2812.520 25.460 ;
      LAYER met2 ;
        RECT 1734.080 25.830 1734.220 54.000 ;
        RECT 1854.540 27.550 1854.800 27.870 ;
        RECT 1734.020 25.510 1734.280 25.830 ;
        RECT 1754.260 25.685 1754.520 25.830 ;
        RECT 1854.600 25.685 1854.740 27.550 ;
        RECT 1754.250 25.315 1754.530 25.685 ;
        RECT 1854.530 25.315 1854.810 25.685 ;
        RECT 2812.260 25.170 2812.520 25.490 ;
        RECT 2812.320 2.400 2812.460 25.170 ;
        RECT 2812.250 0.000 2812.530 2.400 ;
      LAYER via2 ;
        RECT 1754.250 25.360 1754.530 25.640 ;
        RECT 1854.530 25.360 1854.810 25.640 ;
      LAYER met3 ;
        RECT 1754.225 25.650 1754.555 25.665 ;
        RECT 1854.505 25.650 1854.835 25.665 ;
        RECT 1754.225 25.350 1854.835 25.650 ;
        RECT 1754.225 25.335 1754.555 25.350 ;
        RECT 1854.505 25.335 1854.835 25.350 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2575.865 24.905 2576.035 28.135 ;
      LAYER mcon ;
        RECT 2575.865 27.965 2576.035 28.135 ;
      LAYER met1 ;
        RECT 1854.970 28.120 1855.290 28.180 ;
        RECT 2575.805 28.120 2576.095 28.165 ;
        RECT 1854.970 27.980 2576.095 28.120 ;
        RECT 1854.970 27.920 1855.290 27.980 ;
        RECT 2575.805 27.935 2576.095 27.980 ;
        RECT 2575.805 25.060 2576.095 25.105 ;
        RECT 2830.170 25.060 2830.490 25.120 ;
        RECT 2575.805 24.920 2830.490 25.060 ;
        RECT 2575.805 24.875 2576.095 24.920 ;
        RECT 2830.170 24.860 2830.490 24.920 ;
        RECT 1733.530 23.360 1733.850 23.420 ;
        RECT 1753.310 23.360 1753.630 23.420 ;
        RECT 1733.530 23.220 1753.630 23.360 ;
        RECT 1733.530 23.160 1733.850 23.220 ;
        RECT 1753.310 23.160 1753.630 23.220 ;
      LAYER via ;
        RECT 1855.000 27.920 1855.260 28.180 ;
        RECT 2830.200 24.860 2830.460 25.120 ;
        RECT 1733.560 23.160 1733.820 23.420 ;
        RECT 1753.340 23.160 1753.600 23.420 ;
      LAYER met2 ;
        RECT 1733.620 23.450 1733.760 54.000 ;
        RECT 1855.000 27.890 1855.260 28.210 ;
        RECT 1855.060 25.005 1855.200 27.890 ;
        RECT 1753.330 24.635 1753.610 25.005 ;
        RECT 1854.990 24.635 1855.270 25.005 ;
        RECT 2830.200 24.830 2830.460 25.150 ;
        RECT 1753.400 23.450 1753.540 24.635 ;
        RECT 1733.560 23.130 1733.820 23.450 ;
        RECT 1753.340 23.130 1753.600 23.450 ;
        RECT 2830.260 2.400 2830.400 24.830 ;
        RECT 2830.190 0.000 2830.470 2.400 ;
      LAYER via2 ;
        RECT 1753.330 24.680 1753.610 24.960 ;
        RECT 1854.990 24.680 1855.270 24.960 ;
      LAYER met3 ;
        RECT 1753.305 24.970 1753.635 24.985 ;
        RECT 1854.965 24.970 1855.295 24.985 ;
        RECT 1753.305 24.670 1855.295 24.970 ;
        RECT 1753.305 24.655 1753.635 24.670 ;
        RECT 1854.965 24.655 1855.295 24.670 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2528.485 20.485 2528.655 25.075 ;
        RECT 2575.405 20.485 2575.575 25.075 ;
        RECT 2647.625 21.165 2647.795 24.055 ;
        RECT 2672.925 23.205 2673.095 24.055 ;
        RECT 2797.125 23.545 2797.755 23.715 ;
        RECT 2693.625 22.185 2693.795 23.375 ;
        RECT 2749.285 23.035 2749.455 23.375 ;
        RECT 2741.465 22.185 2741.635 23.035 ;
        RECT 2748.825 22.865 2749.455 23.035 ;
      LAYER mcon ;
        RECT 2528.485 24.905 2528.655 25.075 ;
        RECT 2575.405 24.905 2575.575 25.075 ;
        RECT 2647.625 23.885 2647.795 24.055 ;
        RECT 2672.925 23.885 2673.095 24.055 ;
        RECT 2797.585 23.545 2797.755 23.715 ;
        RECT 2693.625 23.205 2693.795 23.375 ;
        RECT 2749.285 23.205 2749.455 23.375 ;
        RECT 2741.465 22.865 2741.635 23.035 ;
      LAYER met1 ;
        RECT 2528.425 25.060 2528.715 25.105 ;
        RECT 2575.345 25.060 2575.635 25.105 ;
        RECT 2528.425 24.920 2575.635 25.060 ;
        RECT 2528.425 24.875 2528.715 24.920 ;
        RECT 2575.345 24.875 2575.635 24.920 ;
        RECT 2647.565 24.040 2647.855 24.085 ;
        RECT 2672.865 24.040 2673.155 24.085 ;
        RECT 2647.565 23.900 2673.155 24.040 ;
        RECT 2647.565 23.855 2647.855 23.900 ;
        RECT 2672.865 23.855 2673.155 23.900 ;
        RECT 1739.510 23.700 1739.830 23.760 ;
        RECT 1752.850 23.700 1753.170 23.760 ;
        RECT 1739.510 23.560 1753.170 23.700 ;
        RECT 1739.510 23.500 1739.830 23.560 ;
        RECT 1752.850 23.500 1753.170 23.560 ;
        RECT 2797.065 23.515 2797.355 23.745 ;
        RECT 2797.525 23.700 2797.815 23.745 ;
        RECT 2847.650 23.700 2847.970 23.760 ;
        RECT 2797.525 23.560 2847.970 23.700 ;
        RECT 2797.525 23.515 2797.815 23.560 ;
        RECT 2672.865 23.360 2673.155 23.405 ;
        RECT 2693.565 23.360 2693.855 23.405 ;
        RECT 2672.865 23.220 2693.855 23.360 ;
        RECT 2672.865 23.175 2673.155 23.220 ;
        RECT 2693.565 23.175 2693.855 23.220 ;
        RECT 2749.225 23.360 2749.515 23.405 ;
        RECT 2797.140 23.360 2797.280 23.515 ;
        RECT 2847.650 23.500 2847.970 23.560 ;
        RECT 2749.225 23.220 2797.280 23.360 ;
        RECT 2749.225 23.175 2749.515 23.220 ;
        RECT 2741.405 23.020 2741.695 23.065 ;
        RECT 2748.765 23.020 2749.055 23.065 ;
        RECT 2741.405 22.880 2749.055 23.020 ;
        RECT 2741.405 22.835 2741.695 22.880 ;
        RECT 2748.765 22.835 2749.055 22.880 ;
        RECT 2693.565 22.340 2693.855 22.385 ;
        RECT 2741.405 22.340 2741.695 22.385 ;
        RECT 2693.565 22.200 2741.695 22.340 ;
        RECT 2693.565 22.155 2693.855 22.200 ;
        RECT 2741.405 22.155 2741.695 22.200 ;
        RECT 2647.565 21.320 2647.855 21.365 ;
        RECT 2577.260 21.180 2647.855 21.320 ;
        RECT 2577.260 20.980 2577.400 21.180 ;
        RECT 2647.565 21.135 2647.855 21.180 ;
        RECT 2576.800 20.840 2577.400 20.980 ;
        RECT 2094.170 20.640 2094.490 20.700 ;
        RECT 2528.425 20.640 2528.715 20.685 ;
        RECT 2094.170 20.500 2528.715 20.640 ;
        RECT 2094.170 20.440 2094.490 20.500 ;
        RECT 2528.425 20.455 2528.715 20.500 ;
        RECT 2575.345 20.640 2575.635 20.685 ;
        RECT 2576.800 20.640 2576.940 20.840 ;
        RECT 2575.345 20.500 2576.940 20.640 ;
        RECT 2575.345 20.455 2575.635 20.500 ;
      LAYER via ;
        RECT 1739.540 23.500 1739.800 23.760 ;
        RECT 1752.880 23.500 1753.140 23.760 ;
        RECT 2847.680 23.500 2847.940 23.760 ;
        RECT 2094.200 20.440 2094.460 20.700 ;
      LAYER met2 ;
        RECT 1739.600 23.790 1739.740 54.000 ;
        RECT 1752.870 23.955 1753.150 24.325 ;
        RECT 1752.940 23.790 1753.080 23.955 ;
        RECT 1739.540 23.470 1739.800 23.790 ;
        RECT 1752.880 23.470 1753.140 23.790 ;
        RECT 2094.190 23.275 2094.470 23.645 ;
        RECT 2847.680 23.470 2847.940 23.790 ;
        RECT 2094.260 20.730 2094.400 23.275 ;
        RECT 2094.200 20.410 2094.460 20.730 ;
        RECT 2847.740 2.400 2847.880 23.470 ;
        RECT 2847.670 0.000 2847.950 2.400 ;
      LAYER via2 ;
        RECT 1752.870 24.000 1753.150 24.280 ;
        RECT 2094.190 23.320 2094.470 23.600 ;
      LAYER met3 ;
        RECT 1752.845 24.290 1753.175 24.305 ;
        RECT 1752.845 23.990 1759.370 24.290 ;
        RECT 1752.845 23.975 1753.175 23.990 ;
        RECT 1759.070 23.610 1759.370 23.990 ;
        RECT 2094.165 23.610 2094.495 23.625 ;
        RECT 1759.070 23.310 2094.495 23.610 ;
        RECT 2094.165 23.295 2094.495 23.310 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1746.040 23.645 1746.180 54.000 ;
        RECT 1779.090 23.955 1779.370 24.325 ;
        RECT 2865.610 23.955 2865.890 24.325 ;
        RECT 1745.970 23.275 1746.250 23.645 ;
        RECT 1779.160 22.965 1779.300 23.955 ;
        RECT 1779.090 22.595 1779.370 22.965 ;
        RECT 2865.680 2.400 2865.820 23.955 ;
        RECT 2865.610 0.000 2865.890 2.400 ;
      LAYER via2 ;
        RECT 1779.090 24.000 1779.370 24.280 ;
        RECT 2865.610 24.000 2865.890 24.280 ;
        RECT 1745.970 23.320 1746.250 23.600 ;
        RECT 1779.090 22.640 1779.370 22.920 ;
      LAYER met3 ;
        RECT 1779.065 24.290 1779.395 24.305 ;
        RECT 2865.585 24.290 2865.915 24.305 ;
        RECT 1779.065 23.990 2865.915 24.290 ;
        RECT 1779.065 23.975 1779.395 23.990 ;
        RECT 2865.585 23.975 2865.915 23.990 ;
        RECT 1745.945 23.610 1746.275 23.625 ;
        RECT 1745.945 23.310 1758.450 23.610 ;
        RECT 1745.945 23.295 1746.275 23.310 ;
        RECT 1758.150 22.930 1758.450 23.310 ;
        RECT 1779.065 22.930 1779.395 22.945 ;
        RECT 1758.150 22.630 1779.395 22.930 ;
        RECT 1779.065 22.615 1779.395 22.630 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2879.850 1666.240 2880.170 1666.300 ;
        RECT 2870.580 1666.100 2880.170 1666.240 ;
        RECT 2879.850 1666.040 2880.170 1666.100 ;
        RECT 2879.850 62.120 2880.170 62.180 ;
        RECT 2883.530 62.120 2883.850 62.180 ;
        RECT 2879.850 61.980 2883.850 62.120 ;
        RECT 2879.850 61.920 2880.170 61.980 ;
        RECT 2883.530 61.920 2883.850 61.980 ;
      LAYER via ;
        RECT 2879.880 1666.040 2880.140 1666.300 ;
        RECT 2879.880 61.920 2880.140 62.180 ;
        RECT 2883.560 61.920 2883.820 62.180 ;
      LAYER met2 ;
        RECT 2879.880 1666.010 2880.140 1666.330 ;
        RECT 2879.940 62.210 2880.080 1666.010 ;
        RECT 2879.880 61.890 2880.140 62.210 ;
        RECT 2883.560 61.890 2883.820 62.210 ;
        RECT 2883.620 2.400 2883.760 61.890 ;
        RECT 2883.550 0.000 2883.830 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2896.870 1562.880 2897.190 1562.940 ;
        RECT 2870.580 1562.740 2897.190 1562.880 ;
        RECT 2896.870 1562.680 2897.190 1562.740 ;
        RECT 2896.870 20.640 2897.190 20.700 ;
        RECT 2901.470 20.640 2901.790 20.700 ;
        RECT 2896.870 20.500 2901.790 20.640 ;
        RECT 2896.870 20.440 2897.190 20.500 ;
        RECT 2901.470 20.440 2901.790 20.500 ;
      LAYER via ;
        RECT 2896.900 1562.680 2897.160 1562.940 ;
        RECT 2896.900 20.440 2897.160 20.700 ;
        RECT 2901.500 20.440 2901.760 20.700 ;
      LAYER met2 ;
        RECT 2896.900 1562.650 2897.160 1562.970 ;
        RECT 2896.960 20.730 2897.100 1562.650 ;
        RECT 2896.900 20.410 2897.160 20.730 ;
        RECT 2901.500 20.410 2901.760 20.730 ;
        RECT 2901.560 2.400 2901.700 20.410 ;
        RECT 2901.490 0.000 2901.770 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 849.410 2.960 849.730 3.020 ;
        RECT 849.870 2.960 850.190 3.020 ;
        RECT 849.410 2.820 850.190 2.960 ;
        RECT 849.410 2.760 849.730 2.820 ;
        RECT 849.870 2.760 850.190 2.820 ;
      LAYER via ;
        RECT 849.440 2.760 849.700 3.020 ;
        RECT 849.900 2.760 850.160 3.020 ;
      LAYER met2 ;
        RECT 848.580 48.805 848.720 54.000 ;
        RECT 848.510 48.435 848.790 48.805 ;
        RECT 849.430 48.435 849.710 48.805 ;
        RECT 849.500 48.010 849.640 48.435 ;
        RECT 849.500 47.870 850.100 48.010 ;
        RECT 849.960 3.050 850.100 47.870 ;
        RECT 849.440 2.730 849.700 3.050 ;
        RECT 849.900 2.730 850.160 3.050 ;
        RECT 849.500 2.400 849.640 2.730 ;
        RECT 849.430 0.000 849.710 2.400 ;
      LAYER via2 ;
        RECT 848.510 48.480 848.790 48.760 ;
        RECT 849.430 48.480 849.710 48.760 ;
      LAYER met3 ;
        RECT 848.485 48.770 848.815 48.785 ;
        RECT 849.405 48.770 849.735 48.785 ;
        RECT 848.485 48.470 849.735 48.770 ;
        RECT 848.485 48.455 848.815 48.470 ;
        RECT 849.405 48.455 849.735 48.470 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 867.350 2.960 867.670 3.020 ;
        RECT 871.490 2.960 871.810 3.020 ;
        RECT 867.350 2.820 871.810 2.960 ;
        RECT 867.350 2.760 867.670 2.820 ;
        RECT 871.490 2.760 871.810 2.820 ;
      LAYER via ;
        RECT 867.380 2.760 867.640 3.020 ;
        RECT 871.520 2.760 871.780 3.020 ;
      LAYER met2 ;
        RECT 871.580 3.050 871.720 54.000 ;
        RECT 867.380 2.730 867.640 3.050 ;
        RECT 871.520 2.730 871.780 3.050 ;
        RECT 867.440 2.400 867.580 2.730 ;
        RECT 867.370 0.000 867.650 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 885.380 2.400 885.520 54.000 ;
        RECT 885.310 0.000 885.590 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 903.230 2.960 903.550 3.020 ;
        RECT 905.990 2.960 906.310 3.020 ;
        RECT 903.230 2.820 906.310 2.960 ;
        RECT 903.230 2.760 903.550 2.820 ;
        RECT 905.990 2.760 906.310 2.820 ;
      LAYER via ;
        RECT 903.260 2.760 903.520 3.020 ;
        RECT 906.020 2.760 906.280 3.020 ;
      LAYER met2 ;
        RECT 906.080 3.050 906.220 54.000 ;
        RECT 903.260 2.730 903.520 3.050 ;
        RECT 906.020 2.730 906.280 3.050 ;
        RECT 903.320 2.400 903.460 2.730 ;
        RECT 903.250 0.000 903.530 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 921.170 42.060 921.490 42.120 ;
        RECT 926.690 42.060 927.010 42.120 ;
        RECT 921.170 41.920 927.010 42.060 ;
        RECT 921.170 41.860 921.490 41.920 ;
        RECT 926.690 41.860 927.010 41.920 ;
      LAYER via ;
        RECT 921.200 41.860 921.460 42.120 ;
        RECT 926.720 41.860 926.980 42.120 ;
      LAYER met2 ;
        RECT 926.780 42.150 926.920 54.000 ;
        RECT 921.200 41.830 921.460 42.150 ;
        RECT 926.720 41.830 926.980 42.150 ;
        RECT 921.260 2.400 921.400 41.830 ;
        RECT 921.190 0.000 921.470 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1343.540 24.325 1343.680 54.000 ;
        RECT 938.670 23.955 938.950 24.325 ;
        RECT 1343.470 23.955 1343.750 24.325 ;
        RECT 938.740 2.400 938.880 23.955 ;
        RECT 938.670 0.000 938.950 2.400 ;
      LAYER via2 ;
        RECT 938.670 24.000 938.950 24.280 ;
        RECT 1343.470 24.000 1343.750 24.280 ;
      LAYER met3 ;
        RECT 938.645 24.290 938.975 24.305 ;
        RECT 1343.445 24.290 1343.775 24.305 ;
        RECT 938.645 23.990 1343.775 24.290 ;
        RECT 938.645 23.975 938.975 23.990 ;
        RECT 1343.445 23.975 1343.775 23.990 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1320.985 26.945 1322.075 27.115 ;
        RECT 1320.985 26.605 1321.155 26.945 ;
        RECT 1321.905 26.775 1322.075 26.945 ;
        RECT 1321.905 26.605 1322.535 26.775 ;
        RECT 1322.365 22.525 1322.535 26.605 ;
      LAYER met1 ;
        RECT 956.590 26.760 956.910 26.820 ;
        RECT 1320.925 26.760 1321.215 26.805 ;
        RECT 956.590 26.620 1321.215 26.760 ;
        RECT 956.590 26.560 956.910 26.620 ;
        RECT 1320.925 26.575 1321.215 26.620 ;
        RECT 1322.305 22.680 1322.595 22.725 ;
        RECT 1348.510 22.680 1348.830 22.740 ;
        RECT 1322.305 22.540 1348.830 22.680 ;
        RECT 1322.305 22.495 1322.595 22.540 ;
        RECT 1348.510 22.480 1348.830 22.540 ;
      LAYER via ;
        RECT 956.620 26.560 956.880 26.820 ;
        RECT 1348.540 22.480 1348.800 22.740 ;
      LAYER met2 ;
        RECT 956.620 26.530 956.880 26.850 ;
        RECT 956.680 2.400 956.820 26.530 ;
        RECT 1348.600 22.770 1348.740 54.000 ;
        RECT 1348.540 22.450 1348.800 22.770 ;
        RECT 956.610 0.000 956.890 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1295.225 23.545 1295.395 31.875 ;
      LAYER mcon ;
        RECT 1295.225 31.705 1295.395 31.875 ;
      LAYER met1 ;
        RECT 1295.165 31.860 1295.455 31.905 ;
        RECT 1350.350 31.860 1350.670 31.920 ;
        RECT 1295.165 31.720 1350.670 31.860 ;
        RECT 1295.165 31.675 1295.455 31.720 ;
        RECT 1350.350 31.660 1350.670 31.720 ;
        RECT 974.990 23.700 975.310 23.760 ;
        RECT 1295.165 23.700 1295.455 23.745 ;
        RECT 974.990 23.560 1295.455 23.700 ;
        RECT 974.990 23.500 975.310 23.560 ;
        RECT 1295.165 23.515 1295.455 23.560 ;
      LAYER via ;
        RECT 1350.380 31.660 1350.640 31.920 ;
        RECT 975.020 23.500 975.280 23.760 ;
      LAYER met2 ;
        RECT 1350.440 31.950 1350.580 54.000 ;
        RECT 1350.380 31.630 1350.640 31.950 ;
        RECT 975.020 23.470 975.280 23.790 ;
        RECT 975.080 11.970 975.220 23.470 ;
        RECT 974.620 11.830 975.220 11.970 ;
        RECT 974.620 2.400 974.760 11.830 ;
        RECT 974.550 0.000 974.830 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 653.450 26.080 653.770 26.140 ;
        RECT 1224.310 26.080 1224.630 26.140 ;
        RECT 653.450 25.940 1224.630 26.080 ;
        RECT 653.450 25.880 653.770 25.940 ;
        RECT 1224.310 25.880 1224.630 25.940 ;
      LAYER via ;
        RECT 653.480 25.880 653.740 26.140 ;
        RECT 1224.340 25.880 1224.600 26.140 ;
      LAYER met2 ;
        RECT 1286.500 27.045 1286.640 54.000 ;
        RECT 1224.330 26.675 1224.610 27.045 ;
        RECT 1286.430 26.675 1286.710 27.045 ;
        RECT 1224.400 26.170 1224.540 26.675 ;
        RECT 653.480 25.850 653.740 26.170 ;
        RECT 1224.340 25.850 1224.600 26.170 ;
        RECT 653.540 2.400 653.680 25.850 ;
        RECT 653.470 0.000 653.750 2.400 ;
      LAYER via2 ;
        RECT 1224.330 26.720 1224.610 27.000 ;
        RECT 1286.430 26.720 1286.710 27.000 ;
      LAYER met3 ;
        RECT 1224.305 27.010 1224.635 27.025 ;
        RECT 1286.405 27.010 1286.735 27.025 ;
        RECT 1224.305 26.710 1286.735 27.010 ;
        RECT 1224.305 26.695 1224.635 26.710 ;
        RECT 1286.405 26.695 1286.735 26.710 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1337.545 22.185 1337.715 23.035 ;
      LAYER mcon ;
        RECT 1337.545 22.865 1337.715 23.035 ;
      LAYER met1 ;
        RECT 992.470 23.360 992.790 23.420 ;
        RECT 992.470 23.220 1322.060 23.360 ;
        RECT 992.470 23.160 992.790 23.220 ;
        RECT 1321.920 23.020 1322.060 23.220 ;
        RECT 1337.485 23.020 1337.775 23.065 ;
        RECT 1321.920 22.880 1337.775 23.020 ;
        RECT 1337.485 22.835 1337.775 22.880 ;
        RECT 1337.485 22.340 1337.775 22.385 ;
        RECT 1354.950 22.340 1355.270 22.400 ;
        RECT 1337.485 22.200 1355.270 22.340 ;
        RECT 1337.485 22.155 1337.775 22.200 ;
        RECT 1354.950 22.140 1355.270 22.200 ;
      LAYER via ;
        RECT 992.500 23.160 992.760 23.420 ;
        RECT 1354.980 22.140 1355.240 22.400 ;
      LAYER met2 ;
        RECT 992.500 23.130 992.760 23.450 ;
        RECT 992.560 2.400 992.700 23.130 ;
        RECT 1355.040 22.430 1355.180 54.000 ;
        RECT 1354.980 22.110 1355.240 22.430 ;
        RECT 992.490 0.000 992.770 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1337.085 20.485 1337.255 22.355 ;
      LAYER mcon ;
        RECT 1337.085 22.185 1337.255 22.355 ;
      LAYER met1 ;
        RECT 1009.950 23.020 1010.270 23.080 ;
        RECT 1321.370 23.020 1321.690 23.080 ;
        RECT 1009.950 22.880 1321.690 23.020 ;
        RECT 1009.950 22.820 1010.270 22.880 ;
        RECT 1321.370 22.820 1321.690 22.880 ;
        RECT 1321.370 22.340 1321.690 22.400 ;
        RECT 1337.025 22.340 1337.315 22.385 ;
        RECT 1321.370 22.200 1337.315 22.340 ;
        RECT 1321.370 22.140 1321.690 22.200 ;
        RECT 1337.025 22.155 1337.315 22.200 ;
        RECT 1356.790 20.980 1357.110 21.040 ;
        RECT 1344.920 20.840 1357.110 20.980 ;
        RECT 1337.025 20.640 1337.315 20.685 ;
        RECT 1344.920 20.640 1345.060 20.840 ;
        RECT 1356.790 20.780 1357.110 20.840 ;
        RECT 1337.025 20.500 1345.060 20.640 ;
        RECT 1337.025 20.455 1337.315 20.500 ;
      LAYER via ;
        RECT 1009.980 22.820 1010.240 23.080 ;
        RECT 1321.400 22.820 1321.660 23.080 ;
        RECT 1321.400 22.140 1321.660 22.400 ;
        RECT 1356.820 20.780 1357.080 21.040 ;
      LAYER met2 ;
        RECT 1356.880 48.690 1357.020 54.000 ;
        RECT 1356.880 48.550 1357.940 48.690 ;
        RECT 1357.800 48.010 1357.940 48.550 ;
        RECT 1356.880 47.870 1357.940 48.010 ;
        RECT 1009.980 22.790 1010.240 23.110 ;
        RECT 1321.400 22.790 1321.660 23.110 ;
        RECT 1010.040 2.400 1010.180 22.790 ;
        RECT 1321.460 22.430 1321.600 22.790 ;
        RECT 1321.400 22.110 1321.660 22.430 ;
        RECT 1356.880 21.070 1357.020 47.870 ;
        RECT 1356.820 20.750 1357.080 21.070 ;
        RECT 1009.970 0.000 1010.250 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1027.890 22.680 1028.210 22.740 ;
        RECT 1321.830 22.680 1322.150 22.740 ;
        RECT 1027.890 22.540 1322.150 22.680 ;
        RECT 1027.890 22.480 1028.210 22.540 ;
        RECT 1321.830 22.480 1322.150 22.540 ;
        RECT 1348.970 22.680 1349.290 22.740 ;
        RECT 1362.310 22.680 1362.630 22.740 ;
        RECT 1348.970 22.540 1362.630 22.680 ;
        RECT 1348.970 22.480 1349.290 22.540 ;
        RECT 1362.310 22.480 1362.630 22.540 ;
      LAYER via ;
        RECT 1027.920 22.480 1028.180 22.740 ;
        RECT 1321.860 22.480 1322.120 22.740 ;
        RECT 1349.000 22.480 1349.260 22.740 ;
        RECT 1362.340 22.480 1362.600 22.740 ;
      LAYER met2 ;
        RECT 1027.920 22.450 1028.180 22.770 ;
        RECT 1321.850 22.595 1322.130 22.965 ;
        RECT 1348.990 22.595 1349.270 22.965 ;
        RECT 1362.400 22.770 1362.540 54.000 ;
        RECT 1321.860 22.450 1322.120 22.595 ;
        RECT 1349.000 22.450 1349.260 22.595 ;
        RECT 1362.340 22.450 1362.600 22.770 ;
        RECT 1027.980 2.400 1028.120 22.450 ;
        RECT 1027.910 0.000 1028.190 2.400 ;
      LAYER via2 ;
        RECT 1321.850 22.640 1322.130 22.920 ;
        RECT 1348.990 22.640 1349.270 22.920 ;
      LAYER met3 ;
        RECT 1321.825 22.930 1322.155 22.945 ;
        RECT 1348.965 22.930 1349.295 22.945 ;
        RECT 1321.825 22.630 1349.295 22.930 ;
        RECT 1321.825 22.615 1322.155 22.630 ;
        RECT 1348.965 22.615 1349.295 22.630 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1045.830 22.340 1046.150 22.400 ;
        RECT 1320.910 22.340 1321.230 22.400 ;
        RECT 1045.830 22.200 1321.230 22.340 ;
        RECT 1045.830 22.140 1046.150 22.200 ;
        RECT 1320.910 22.140 1321.230 22.200 ;
      LAYER via ;
        RECT 1045.860 22.140 1046.120 22.400 ;
        RECT 1320.940 22.140 1321.200 22.400 ;
      LAYER met2 ;
        RECT 1045.860 22.110 1046.120 22.430 ;
        RECT 1320.940 22.285 1321.200 22.430 ;
        RECT 1364.700 22.285 1364.840 54.000 ;
        RECT 1045.920 2.400 1046.060 22.110 ;
        RECT 1320.930 21.915 1321.210 22.285 ;
        RECT 1364.630 21.915 1364.910 22.285 ;
        RECT 1045.850 0.000 1046.130 2.400 ;
      LAYER via2 ;
        RECT 1320.930 21.960 1321.210 22.240 ;
        RECT 1364.630 21.960 1364.910 22.240 ;
      LAYER met3 ;
        RECT 1320.905 22.250 1321.235 22.265 ;
        RECT 1364.605 22.250 1364.935 22.265 ;
        RECT 1320.905 21.950 1364.935 22.250 ;
        RECT 1320.905 21.935 1321.235 21.950 ;
        RECT 1364.605 21.935 1364.935 21.950 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1102.485 21.165 1103.575 21.335 ;
        RECT 1102.485 20.825 1102.655 21.165 ;
      LAYER mcon ;
        RECT 1103.405 21.165 1103.575 21.335 ;
      LAYER met1 ;
        RECT 1103.345 21.320 1103.635 21.365 ;
        RECT 1371.050 21.320 1371.370 21.380 ;
        RECT 1103.345 21.180 1371.370 21.320 ;
        RECT 1103.345 21.135 1103.635 21.180 ;
        RECT 1371.050 21.120 1371.370 21.180 ;
        RECT 1063.770 20.980 1064.090 21.040 ;
        RECT 1102.425 20.980 1102.715 21.025 ;
        RECT 1063.770 20.840 1102.715 20.980 ;
        RECT 1063.770 20.780 1064.090 20.840 ;
        RECT 1102.425 20.795 1102.715 20.840 ;
      LAYER via ;
        RECT 1371.080 21.120 1371.340 21.380 ;
        RECT 1063.800 20.780 1064.060 21.040 ;
      LAYER met2 ;
        RECT 1371.140 21.410 1371.280 54.000 ;
        RECT 1371.080 21.090 1371.340 21.410 ;
        RECT 1063.800 20.750 1064.060 21.070 ;
        RECT 1063.860 2.400 1064.000 20.750 ;
        RECT 1063.790 0.000 1064.070 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1344.445 20.825 1344.615 23.035 ;
      LAYER mcon ;
        RECT 1344.445 22.865 1344.615 23.035 ;
      LAYER met1 ;
        RECT 1344.385 23.020 1344.675 23.065 ;
        RECT 1370.590 23.020 1370.910 23.080 ;
        RECT 1344.385 22.880 1370.910 23.020 ;
        RECT 1344.385 22.835 1344.675 22.880 ;
        RECT 1370.590 22.820 1370.910 22.880 ;
        RECT 1093.210 21.320 1093.530 21.380 ;
        RECT 1093.210 21.180 1103.100 21.320 ;
        RECT 1093.210 21.120 1093.530 21.180 ;
        RECT 1102.960 20.980 1103.100 21.180 ;
        RECT 1344.385 20.980 1344.675 21.025 ;
        RECT 1102.960 20.840 1344.675 20.980 ;
        RECT 1344.385 20.795 1344.675 20.840 ;
      LAYER via ;
        RECT 1370.620 22.820 1370.880 23.080 ;
        RECT 1093.240 21.120 1093.500 21.380 ;
      LAYER met2 ;
        RECT 1370.680 23.110 1370.820 54.000 ;
        RECT 1370.620 22.790 1370.880 23.110 ;
        RECT 1081.730 21.235 1082.010 21.605 ;
        RECT 1093.230 21.235 1093.510 21.605 ;
        RECT 1081.800 2.400 1081.940 21.235 ;
        RECT 1093.240 21.090 1093.500 21.235 ;
        RECT 1081.730 0.000 1082.010 2.400 ;
      LAYER via2 ;
        RECT 1081.730 21.280 1082.010 21.560 ;
        RECT 1093.230 21.280 1093.510 21.560 ;
      LAYER met3 ;
        RECT 1081.705 21.570 1082.035 21.585 ;
        RECT 1093.205 21.570 1093.535 21.585 ;
        RECT 1081.705 21.270 1093.535 21.570 ;
        RECT 1081.705 21.255 1082.035 21.270 ;
        RECT 1093.205 21.255 1093.535 21.270 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1126.790 24.040 1127.110 24.100 ;
        RECT 1376.110 24.040 1376.430 24.100 ;
        RECT 1126.790 23.900 1376.430 24.040 ;
        RECT 1126.790 23.840 1127.110 23.900 ;
        RECT 1376.110 23.840 1376.430 23.900 ;
      LAYER via ;
        RECT 1126.820 23.840 1127.080 24.100 ;
        RECT 1376.140 23.840 1376.400 24.100 ;
      LAYER met2 ;
        RECT 1376.200 24.130 1376.340 54.000 ;
        RECT 1126.820 23.810 1127.080 24.130 ;
        RECT 1376.140 23.810 1376.400 24.130 ;
        RECT 1098.290 23.275 1098.570 23.645 ;
        RECT 1126.350 23.530 1126.630 23.645 ;
        RECT 1126.880 23.530 1127.020 23.810 ;
        RECT 1126.350 23.390 1127.020 23.530 ;
        RECT 1126.350 23.275 1126.630 23.390 ;
        RECT 1098.360 6.530 1098.500 23.275 ;
        RECT 1098.360 6.390 1099.420 6.530 ;
        RECT 1099.280 2.400 1099.420 6.390 ;
        RECT 1099.210 0.000 1099.490 2.400 ;
      LAYER via2 ;
        RECT 1098.290 23.320 1098.570 23.600 ;
        RECT 1126.350 23.320 1126.630 23.600 ;
      LAYER met3 ;
        RECT 1098.265 23.610 1098.595 23.625 ;
        RECT 1126.325 23.610 1126.655 23.625 ;
        RECT 1098.265 23.310 1126.655 23.610 ;
        RECT 1098.265 23.295 1098.595 23.310 ;
        RECT 1126.325 23.295 1126.655 23.310 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1147.105 13.005 1147.275 25.415 ;
      LAYER mcon ;
        RECT 1147.105 25.245 1147.275 25.415 ;
      LAYER met1 ;
        RECT 1147.045 25.400 1147.335 25.445 ;
        RECT 1378.410 25.400 1378.730 25.460 ;
        RECT 1147.045 25.260 1378.730 25.400 ;
        RECT 1147.045 25.215 1147.335 25.260 ;
        RECT 1378.410 25.200 1378.730 25.260 ;
        RECT 1117.130 13.160 1117.450 13.220 ;
        RECT 1147.045 13.160 1147.335 13.205 ;
        RECT 1117.130 13.020 1147.335 13.160 ;
        RECT 1117.130 12.960 1117.450 13.020 ;
        RECT 1147.045 12.975 1147.335 13.020 ;
      LAYER via ;
        RECT 1378.440 25.200 1378.700 25.460 ;
        RECT 1117.160 12.960 1117.420 13.220 ;
      LAYER met2 ;
        RECT 1378.500 25.490 1378.640 54.000 ;
        RECT 1378.440 25.170 1378.700 25.490 ;
        RECT 1117.160 12.930 1117.420 13.250 ;
        RECT 1117.220 2.400 1117.360 12.930 ;
        RECT 1117.150 0.000 1117.430 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1135.070 25.740 1135.390 25.800 ;
        RECT 1382.550 25.740 1382.870 25.800 ;
        RECT 1135.070 25.600 1382.870 25.740 ;
        RECT 1135.070 25.540 1135.390 25.600 ;
        RECT 1382.550 25.540 1382.870 25.600 ;
      LAYER via ;
        RECT 1135.100 25.540 1135.360 25.800 ;
        RECT 1382.580 25.540 1382.840 25.800 ;
      LAYER met2 ;
        RECT 1382.640 25.830 1382.780 54.000 ;
        RECT 1135.100 25.510 1135.360 25.830 ;
        RECT 1382.580 25.510 1382.840 25.830 ;
        RECT 1135.160 2.400 1135.300 25.510 ;
        RECT 1135.090 0.000 1135.370 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1153.010 25.060 1153.330 25.120 ;
        RECT 1384.850 25.060 1385.170 25.120 ;
        RECT 1153.010 24.920 1385.170 25.060 ;
        RECT 1153.010 24.860 1153.330 24.920 ;
        RECT 1384.850 24.860 1385.170 24.920 ;
      LAYER via ;
        RECT 1153.040 24.860 1153.300 25.120 ;
        RECT 1384.880 24.860 1385.140 25.120 ;
      LAYER met2 ;
        RECT 1384.940 25.150 1385.080 54.000 ;
        RECT 1153.040 24.830 1153.300 25.150 ;
        RECT 1384.880 24.830 1385.140 25.150 ;
        RECT 1153.100 2.400 1153.240 24.830 ;
        RECT 1153.030 0.000 1153.310 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 671.390 26.420 671.710 26.480 ;
        RECT 1223.850 26.420 1224.170 26.480 ;
        RECT 671.390 26.280 1224.170 26.420 ;
        RECT 671.390 26.220 671.710 26.280 ;
        RECT 1223.850 26.220 1224.170 26.280 ;
      LAYER via ;
        RECT 671.420 26.220 671.680 26.480 ;
        RECT 1223.880 26.220 1224.140 26.480 ;
      LAYER met2 ;
        RECT 1288.800 27.725 1288.940 54.000 ;
        RECT 1223.870 27.355 1224.150 27.725 ;
        RECT 1288.730 27.355 1289.010 27.725 ;
        RECT 1223.940 26.510 1224.080 27.355 ;
        RECT 671.420 26.190 671.680 26.510 ;
        RECT 1223.880 26.190 1224.140 26.510 ;
        RECT 671.480 2.400 671.620 26.190 ;
        RECT 671.410 0.000 671.690 2.400 ;
      LAYER via2 ;
        RECT 1223.870 27.400 1224.150 27.680 ;
        RECT 1288.730 27.400 1289.010 27.680 ;
      LAYER met3 ;
        RECT 1223.845 27.690 1224.175 27.705 ;
        RECT 1288.705 27.690 1289.035 27.705 ;
        RECT 1223.845 27.390 1289.035 27.690 ;
        RECT 1223.845 27.375 1224.175 27.390 ;
        RECT 1288.705 27.375 1289.035 27.390 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1176.085 2.805 1176.255 31.535 ;
        RECT 1225.305 26.265 1225.475 31.535 ;
        RECT 1270.845 26.265 1271.015 31.535 ;
      LAYER mcon ;
        RECT 1176.085 31.365 1176.255 31.535 ;
        RECT 1225.305 31.365 1225.475 31.535 ;
        RECT 1270.845 31.365 1271.015 31.535 ;
      LAYER met1 ;
        RECT 1176.025 31.520 1176.315 31.565 ;
        RECT 1225.245 31.520 1225.535 31.565 ;
        RECT 1176.025 31.380 1225.535 31.520 ;
        RECT 1176.025 31.335 1176.315 31.380 ;
        RECT 1225.245 31.335 1225.535 31.380 ;
        RECT 1270.785 31.520 1271.075 31.565 ;
        RECT 1319.990 31.520 1320.310 31.580 ;
        RECT 1270.785 31.380 1320.310 31.520 ;
        RECT 1270.785 31.335 1271.075 31.380 ;
        RECT 1319.990 31.320 1320.310 31.380 ;
        RECT 1225.245 26.420 1225.535 26.465 ;
        RECT 1270.785 26.420 1271.075 26.465 ;
        RECT 1225.245 26.280 1271.075 26.420 ;
        RECT 1225.245 26.235 1225.535 26.280 ;
        RECT 1270.785 26.235 1271.075 26.280 ;
        RECT 1319.990 26.420 1320.310 26.480 ;
        RECT 1391.290 26.420 1391.610 26.480 ;
        RECT 1319.990 26.280 1391.610 26.420 ;
        RECT 1319.990 26.220 1320.310 26.280 ;
        RECT 1391.290 26.220 1391.610 26.280 ;
        RECT 1170.950 2.960 1171.270 3.020 ;
        RECT 1176.025 2.960 1176.315 3.005 ;
        RECT 1170.950 2.820 1176.315 2.960 ;
        RECT 1170.950 2.760 1171.270 2.820 ;
        RECT 1176.025 2.775 1176.315 2.820 ;
      LAYER via ;
        RECT 1320.020 31.320 1320.280 31.580 ;
        RECT 1320.020 26.220 1320.280 26.480 ;
        RECT 1391.320 26.220 1391.580 26.480 ;
        RECT 1170.980 2.760 1171.240 3.020 ;
      LAYER met2 ;
        RECT 1320.020 31.290 1320.280 31.610 ;
        RECT 1320.080 26.510 1320.220 31.290 ;
        RECT 1391.380 26.510 1391.520 54.000 ;
        RECT 1320.020 26.190 1320.280 26.510 ;
        RECT 1391.320 26.190 1391.580 26.510 ;
        RECT 1170.980 2.730 1171.240 3.050 ;
        RECT 1171.040 2.400 1171.180 2.730 ;
        RECT 1170.970 0.000 1171.250 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1296.145 26.265 1297.235 26.435 ;
        RECT 1297.065 25.925 1297.235 26.265 ;
      LAYER met1 ;
        RECT 1392.210 34.580 1392.530 34.640 ;
        RECT 1393.590 34.580 1393.910 34.640 ;
        RECT 1392.210 34.440 1393.910 34.580 ;
        RECT 1392.210 34.380 1392.530 34.440 ;
        RECT 1393.590 34.380 1393.910 34.440 ;
        RECT 1296.085 26.420 1296.375 26.465 ;
        RECT 1271.320 26.280 1296.375 26.420 ;
        RECT 1224.770 26.080 1225.090 26.140 ;
        RECT 1271.320 26.080 1271.460 26.280 ;
        RECT 1296.085 26.235 1296.375 26.280 ;
        RECT 1224.770 25.940 1271.460 26.080 ;
        RECT 1297.005 26.080 1297.295 26.125 ;
        RECT 1393.590 26.080 1393.910 26.140 ;
        RECT 1297.005 25.940 1393.910 26.080 ;
        RECT 1224.770 25.880 1225.090 25.940 ;
        RECT 1297.005 25.895 1297.295 25.940 ;
        RECT 1393.590 25.880 1393.910 25.940 ;
      LAYER via ;
        RECT 1392.240 34.380 1392.500 34.640 ;
        RECT 1393.620 34.380 1393.880 34.640 ;
        RECT 1224.800 25.880 1225.060 26.140 ;
        RECT 1393.620 25.880 1393.880 26.140 ;
      LAYER met2 ;
        RECT 1392.300 34.670 1392.440 54.000 ;
        RECT 1392.240 34.350 1392.500 34.670 ;
        RECT 1393.620 34.350 1393.880 34.670 ;
        RECT 1188.450 25.995 1188.730 26.365 ;
        RECT 1224.790 25.995 1225.070 26.365 ;
        RECT 1393.680 26.170 1393.820 34.350 ;
        RECT 1188.520 2.400 1188.660 25.995 ;
        RECT 1224.800 25.850 1225.060 25.995 ;
        RECT 1393.620 25.850 1393.880 26.170 ;
        RECT 1188.450 0.000 1188.730 2.400 ;
      LAYER via2 ;
        RECT 1188.450 26.040 1188.730 26.320 ;
        RECT 1224.790 26.040 1225.070 26.320 ;
      LAYER met3 ;
        RECT 1188.425 26.330 1188.755 26.345 ;
        RECT 1224.765 26.330 1225.095 26.345 ;
        RECT 1188.425 26.030 1225.095 26.330 ;
        RECT 1188.425 26.015 1188.755 26.030 ;
        RECT 1224.765 26.015 1225.095 26.030 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1319.605 26.265 1320.235 26.435 ;
        RECT 1271.765 20.145 1271.935 26.095 ;
        RECT 1320.065 23.545 1320.235 26.265 ;
      LAYER mcon ;
        RECT 1271.765 25.925 1271.935 26.095 ;
      LAYER met1 ;
        RECT 1319.545 26.420 1319.835 26.465 ;
        RECT 1296.620 26.280 1319.835 26.420 ;
        RECT 1271.705 26.080 1271.995 26.125 ;
        RECT 1296.620 26.080 1296.760 26.280 ;
        RECT 1319.545 26.235 1319.835 26.280 ;
        RECT 1271.705 25.940 1296.760 26.080 ;
        RECT 1271.705 25.895 1271.995 25.940 ;
        RECT 1320.005 23.700 1320.295 23.745 ;
        RECT 1396.810 23.700 1397.130 23.760 ;
        RECT 1320.005 23.560 1397.130 23.700 ;
        RECT 1320.005 23.515 1320.295 23.560 ;
        RECT 1396.810 23.500 1397.130 23.560 ;
        RECT 1206.370 20.300 1206.690 20.360 ;
        RECT 1271.705 20.300 1271.995 20.345 ;
        RECT 1206.370 20.160 1271.995 20.300 ;
        RECT 1206.370 20.100 1206.690 20.160 ;
        RECT 1271.705 20.115 1271.995 20.160 ;
      LAYER via ;
        RECT 1396.840 23.500 1397.100 23.760 ;
        RECT 1206.400 20.100 1206.660 20.360 ;
      LAYER met2 ;
        RECT 1396.900 23.790 1397.040 54.000 ;
        RECT 1396.840 23.470 1397.100 23.790 ;
        RECT 1206.400 20.070 1206.660 20.390 ;
        RECT 1206.460 2.400 1206.600 20.070 ;
        RECT 1206.390 0.000 1206.670 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1224.310 20.640 1224.630 20.700 ;
        RECT 1230.290 20.640 1230.610 20.700 ;
        RECT 1224.310 20.500 1230.610 20.640 ;
        RECT 1224.310 20.440 1224.630 20.500 ;
        RECT 1230.290 20.440 1230.610 20.500 ;
      LAYER via ;
        RECT 1224.340 20.440 1224.600 20.700 ;
        RECT 1230.320 20.440 1230.580 20.700 ;
      LAYER met2 ;
        RECT 1230.380 20.730 1230.520 54.000 ;
        RECT 1224.340 20.410 1224.600 20.730 ;
        RECT 1230.320 20.410 1230.580 20.730 ;
        RECT 1224.400 2.400 1224.540 20.410 ;
        RECT 1224.330 0.000 1224.610 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1242.250 2.960 1242.570 3.020 ;
        RECT 1244.090 2.960 1244.410 3.020 ;
        RECT 1242.250 2.820 1244.410 2.960 ;
        RECT 1242.250 2.760 1242.570 2.820 ;
        RECT 1244.090 2.760 1244.410 2.820 ;
      LAYER via ;
        RECT 1242.280 2.760 1242.540 3.020 ;
        RECT 1244.120 2.760 1244.380 3.020 ;
      LAYER met2 ;
        RECT 1244.180 3.050 1244.320 54.000 ;
        RECT 1242.280 2.730 1242.540 3.050 ;
        RECT 1244.120 2.730 1244.380 3.050 ;
        RECT 1242.340 2.400 1242.480 2.730 ;
        RECT 1242.270 0.000 1242.550 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1259.730 20.640 1260.050 20.700 ;
        RECT 1264.790 20.640 1265.110 20.700 ;
        RECT 1259.730 20.500 1265.110 20.640 ;
        RECT 1259.730 20.440 1260.050 20.500 ;
        RECT 1264.790 20.440 1265.110 20.500 ;
      LAYER via ;
        RECT 1259.760 20.440 1260.020 20.700 ;
        RECT 1264.820 20.440 1265.080 20.700 ;
      LAYER met2 ;
        RECT 1264.880 20.730 1265.020 54.000 ;
        RECT 1259.760 20.410 1260.020 20.730 ;
        RECT 1264.820 20.410 1265.080 20.730 ;
        RECT 1259.820 2.400 1259.960 20.410 ;
        RECT 1259.750 0.000 1260.030 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1278.590 52.260 1278.910 52.320 ;
        RECT 1412.450 52.260 1412.770 52.320 ;
        RECT 1278.590 52.120 1412.770 52.260 ;
        RECT 1278.590 52.060 1278.910 52.120 ;
        RECT 1412.450 52.060 1412.770 52.120 ;
      LAYER via ;
        RECT 1278.620 52.060 1278.880 52.320 ;
        RECT 1412.480 52.060 1412.740 52.320 ;
      LAYER met2 ;
        RECT 1412.540 52.350 1412.680 54.000 ;
        RECT 1278.620 52.030 1278.880 52.350 ;
        RECT 1412.480 52.030 1412.740 52.350 ;
        RECT 1278.680 3.130 1278.820 52.030 ;
        RECT 1277.760 2.990 1278.820 3.130 ;
        RECT 1277.760 2.400 1277.900 2.990 ;
        RECT 1277.690 0.000 1277.970 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1319.605 20.485 1319.775 23.715 ;
        RECT 1321.445 20.485 1321.615 26.775 ;
      LAYER mcon ;
        RECT 1321.445 26.605 1321.615 26.775 ;
        RECT 1319.605 23.545 1319.775 23.715 ;
      LAYER met1 ;
        RECT 1321.385 26.760 1321.675 26.805 ;
        RECT 1417.970 26.760 1418.290 26.820 ;
        RECT 1321.385 26.620 1418.290 26.760 ;
        RECT 1321.385 26.575 1321.675 26.620 ;
        RECT 1417.970 26.560 1418.290 26.620 ;
        RECT 1295.610 23.700 1295.930 23.760 ;
        RECT 1319.545 23.700 1319.835 23.745 ;
        RECT 1295.610 23.560 1319.835 23.700 ;
        RECT 1295.610 23.500 1295.930 23.560 ;
        RECT 1319.545 23.515 1319.835 23.560 ;
        RECT 1319.545 20.640 1319.835 20.685 ;
        RECT 1321.385 20.640 1321.675 20.685 ;
        RECT 1319.545 20.500 1321.675 20.640 ;
        RECT 1319.545 20.455 1319.835 20.500 ;
        RECT 1321.385 20.455 1321.675 20.500 ;
      LAYER via ;
        RECT 1418.000 26.560 1418.260 26.820 ;
        RECT 1295.640 23.500 1295.900 23.760 ;
      LAYER met2 ;
        RECT 1418.060 26.850 1418.200 54.000 ;
        RECT 1418.000 26.530 1418.260 26.850 ;
        RECT 1295.640 23.470 1295.900 23.790 ;
        RECT 1295.700 2.400 1295.840 23.470 ;
        RECT 1295.630 0.000 1295.910 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1322.825 16.745 1322.995 23.375 ;
      LAYER mcon ;
        RECT 1322.825 23.205 1322.995 23.375 ;
      LAYER met1 ;
        RECT 1322.765 23.360 1323.055 23.405 ;
        RECT 1417.510 23.360 1417.830 23.420 ;
        RECT 1322.765 23.220 1417.830 23.360 ;
        RECT 1322.765 23.175 1323.055 23.220 ;
        RECT 1417.510 23.160 1417.830 23.220 ;
        RECT 1314.470 16.900 1314.790 16.960 ;
        RECT 1322.765 16.900 1323.055 16.945 ;
        RECT 1314.470 16.760 1323.055 16.900 ;
        RECT 1314.470 16.700 1314.790 16.760 ;
        RECT 1322.765 16.715 1323.055 16.760 ;
      LAYER via ;
        RECT 1417.540 23.160 1417.800 23.420 ;
        RECT 1314.500 16.700 1314.760 16.960 ;
      LAYER met2 ;
        RECT 1417.600 23.450 1417.740 54.000 ;
        RECT 1417.540 23.130 1417.800 23.450 ;
        RECT 1313.640 17.270 1314.700 17.410 ;
        RECT 1313.640 2.400 1313.780 17.270 ;
        RECT 1314.560 16.990 1314.700 17.270 ;
        RECT 1314.500 16.670 1314.760 16.990 ;
        RECT 1313.570 0.000 1313.850 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1331.490 19.620 1331.810 19.680 ;
        RECT 1420.270 19.620 1420.590 19.680 ;
        RECT 1331.490 19.480 1420.590 19.620 ;
        RECT 1331.490 19.420 1331.810 19.480 ;
        RECT 1420.270 19.420 1420.590 19.480 ;
      LAYER via ;
        RECT 1331.520 19.420 1331.780 19.680 ;
        RECT 1420.300 19.420 1420.560 19.680 ;
      LAYER met2 ;
        RECT 1420.820 21.490 1420.960 54.000 ;
        RECT 1420.360 21.350 1420.960 21.490 ;
        RECT 1420.360 19.710 1420.500 21.350 ;
        RECT 1331.520 19.390 1331.780 19.710 ;
        RECT 1420.300 19.390 1420.560 19.710 ;
        RECT 1331.580 2.400 1331.720 19.390 ;
        RECT 1331.510 0.000 1331.790 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 688.870 19.960 689.190 20.020 ;
        RECT 690.250 19.960 690.570 20.020 ;
        RECT 688.870 19.820 690.570 19.960 ;
        RECT 688.870 19.760 689.190 19.820 ;
        RECT 690.250 19.760 690.570 19.820 ;
      LAYER via ;
        RECT 688.900 19.760 689.160 20.020 ;
        RECT 690.280 19.760 690.540 20.020 ;
      LAYER met2 ;
        RECT 692.180 53.450 692.320 54.000 ;
        RECT 690.340 53.310 692.320 53.450 ;
        RECT 690.340 20.050 690.480 53.310 ;
        RECT 688.900 19.730 689.160 20.050 ;
        RECT 690.280 19.730 690.540 20.050 ;
        RECT 688.960 2.400 689.100 19.730 ;
        RECT 688.890 0.000 689.170 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1348.970 20.640 1349.290 20.700 ;
        RECT 1348.970 20.500 1420.500 20.640 ;
        RECT 1348.970 20.440 1349.290 20.500 ;
        RECT 1420.360 20.300 1420.500 20.500 ;
        RECT 1424.870 20.300 1425.190 20.360 ;
        RECT 1420.360 20.160 1425.190 20.300 ;
        RECT 1424.870 20.100 1425.190 20.160 ;
      LAYER via ;
        RECT 1349.000 20.440 1349.260 20.700 ;
        RECT 1424.900 20.100 1425.160 20.360 ;
      LAYER met2 ;
        RECT 1349.000 20.410 1349.260 20.730 ;
        RECT 1349.060 2.400 1349.200 20.410 ;
        RECT 1424.960 20.390 1425.100 54.000 ;
        RECT 1424.900 20.070 1425.160 20.390 ;
        RECT 1348.990 0.000 1349.270 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1366.910 17.920 1367.230 17.980 ;
        RECT 1392.210 17.920 1392.530 17.980 ;
        RECT 1366.910 17.780 1392.530 17.920 ;
        RECT 1366.910 17.720 1367.230 17.780 ;
        RECT 1392.210 17.720 1392.530 17.780 ;
      LAYER via ;
        RECT 1366.940 17.720 1367.200 17.980 ;
        RECT 1392.240 17.720 1392.500 17.980 ;
      LAYER met2 ;
        RECT 1366.940 17.690 1367.200 18.010 ;
        RECT 1392.240 17.920 1392.500 18.010 ;
        RECT 1392.760 17.920 1392.900 54.000 ;
        RECT 1392.240 17.780 1392.900 17.920 ;
        RECT 1392.240 17.690 1392.500 17.780 ;
        RECT 1367.000 2.400 1367.140 17.690 ;
        RECT 1366.930 0.000 1367.210 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1384.850 14.520 1385.170 14.580 ;
        RECT 1399.570 14.520 1399.890 14.580 ;
        RECT 1384.850 14.380 1399.890 14.520 ;
        RECT 1384.850 14.320 1385.170 14.380 ;
        RECT 1399.570 14.320 1399.890 14.380 ;
      LAYER via ;
        RECT 1384.880 14.320 1385.140 14.580 ;
        RECT 1399.600 14.320 1399.860 14.580 ;
      LAYER met2 ;
        RECT 1399.660 14.610 1399.800 54.000 ;
        RECT 1384.880 14.290 1385.140 14.610 ;
        RECT 1399.600 14.290 1399.860 14.610 ;
        RECT 1384.940 2.400 1385.080 14.290 ;
        RECT 1384.870 0.000 1385.150 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1402.790 14.520 1403.110 14.580 ;
        RECT 1419.810 14.520 1420.130 14.580 ;
        RECT 1402.790 14.380 1420.130 14.520 ;
        RECT 1402.790 14.320 1403.110 14.380 ;
        RECT 1419.810 14.320 1420.130 14.380 ;
      LAYER via ;
        RECT 1402.820 14.320 1403.080 14.580 ;
        RECT 1419.840 14.320 1420.100 14.580 ;
      LAYER met2 ;
        RECT 1420.360 22.170 1420.500 54.000 ;
        RECT 1419.900 22.030 1420.500 22.170 ;
        RECT 1419.900 14.610 1420.040 22.030 ;
        RECT 1402.820 14.290 1403.080 14.610 ;
        RECT 1419.840 14.290 1420.100 14.610 ;
        RECT 1402.880 2.400 1403.020 14.290 ;
        RECT 1402.810 0.000 1403.090 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1420.730 20.640 1421.050 20.700 ;
        RECT 1427.170 20.640 1427.490 20.700 ;
        RECT 1420.730 20.500 1427.490 20.640 ;
        RECT 1420.730 20.440 1421.050 20.500 ;
        RECT 1427.170 20.440 1427.490 20.500 ;
      LAYER via ;
        RECT 1420.760 20.440 1421.020 20.700 ;
        RECT 1427.200 20.440 1427.460 20.700 ;
      LAYER met2 ;
        RECT 1427.260 20.730 1427.400 54.000 ;
        RECT 1420.760 20.410 1421.020 20.730 ;
        RECT 1427.200 20.410 1427.460 20.730 ;
        RECT 1420.820 2.400 1420.960 20.410 ;
        RECT 1420.750 0.000 1421.030 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1444.190 21.120 1444.510 21.380 ;
        RECT 1444.280 20.980 1444.420 21.120 ;
        RECT 1443.820 20.840 1444.420 20.980 ;
        RECT 1438.210 20.640 1438.530 20.700 ;
        RECT 1443.820 20.640 1443.960 20.840 ;
        RECT 1438.210 20.500 1443.960 20.640 ;
        RECT 1438.210 20.440 1438.530 20.500 ;
      LAYER via ;
        RECT 1444.220 21.120 1444.480 21.380 ;
        RECT 1438.240 20.440 1438.500 20.700 ;
      LAYER met2 ;
        RECT 1444.280 21.410 1444.420 54.000 ;
        RECT 1444.220 21.090 1444.480 21.410 ;
        RECT 1438.240 20.410 1438.500 20.730 ;
        RECT 1438.300 2.400 1438.440 20.410 ;
        RECT 1438.230 0.000 1438.510 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1452.930 2.960 1453.250 3.020 ;
        RECT 1456.150 2.960 1456.470 3.020 ;
        RECT 1452.930 2.820 1456.470 2.960 ;
        RECT 1452.930 2.760 1453.250 2.820 ;
        RECT 1456.150 2.760 1456.470 2.820 ;
      LAYER via ;
        RECT 1452.960 2.760 1453.220 3.020 ;
        RECT 1456.180 2.760 1456.440 3.020 ;
      LAYER met2 ;
        RECT 1453.020 3.050 1453.160 54.000 ;
        RECT 1452.960 2.730 1453.220 3.050 ;
        RECT 1456.180 2.730 1456.440 3.050 ;
        RECT 1456.240 2.400 1456.380 2.730 ;
        RECT 1456.170 0.000 1456.450 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1457.990 14.860 1458.310 14.920 ;
        RECT 1474.090 14.860 1474.410 14.920 ;
        RECT 1457.990 14.720 1474.410 14.860 ;
        RECT 1457.990 14.660 1458.310 14.720 ;
        RECT 1474.090 14.660 1474.410 14.720 ;
      LAYER via ;
        RECT 1458.020 14.660 1458.280 14.920 ;
        RECT 1474.120 14.660 1474.380 14.920 ;
      LAYER met2 ;
        RECT 1458.080 14.950 1458.220 54.000 ;
        RECT 1458.020 14.630 1458.280 14.950 ;
        RECT 1474.120 14.630 1474.380 14.950 ;
        RECT 1474.180 2.400 1474.320 14.630 ;
        RECT 1474.110 0.000 1474.390 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1463.970 19.620 1464.290 19.680 ;
        RECT 1492.030 19.620 1492.350 19.680 ;
        RECT 1463.970 19.480 1492.350 19.620 ;
        RECT 1463.970 19.420 1464.290 19.480 ;
        RECT 1492.030 19.420 1492.350 19.480 ;
      LAYER via ;
        RECT 1464.000 19.420 1464.260 19.680 ;
        RECT 1492.060 19.420 1492.320 19.680 ;
      LAYER met2 ;
        RECT 1464.060 19.710 1464.200 54.000 ;
        RECT 1464.000 19.390 1464.260 19.710 ;
        RECT 1492.060 19.390 1492.320 19.710 ;
        RECT 1492.120 2.400 1492.260 19.390 ;
        RECT 1492.050 0.000 1492.330 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1464.890 14.520 1465.210 14.580 ;
        RECT 1509.510 14.520 1509.830 14.580 ;
        RECT 1464.890 14.380 1509.830 14.520 ;
        RECT 1464.890 14.320 1465.210 14.380 ;
        RECT 1509.510 14.320 1509.830 14.380 ;
      LAYER via ;
        RECT 1464.920 14.320 1465.180 14.580 ;
        RECT 1509.540 14.320 1509.800 14.580 ;
      LAYER met2 ;
        RECT 1464.980 14.610 1465.120 54.000 ;
        RECT 1464.920 14.290 1465.180 14.610 ;
        RECT 1509.540 14.290 1509.800 14.610 ;
        RECT 1509.600 2.400 1509.740 14.290 ;
        RECT 1509.530 0.000 1509.810 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 706.810 18.260 707.130 18.320 ;
        RECT 712.790 18.260 713.110 18.320 ;
        RECT 706.810 18.120 713.110 18.260 ;
        RECT 706.810 18.060 707.130 18.120 ;
        RECT 712.790 18.060 713.110 18.120 ;
      LAYER via ;
        RECT 706.840 18.060 707.100 18.320 ;
        RECT 712.820 18.060 713.080 18.320 ;
      LAYER met2 ;
        RECT 712.880 18.350 713.020 54.000 ;
        RECT 706.840 18.030 707.100 18.350 ;
        RECT 712.820 18.030 713.080 18.350 ;
        RECT 706.900 2.400 707.040 18.030 ;
        RECT 706.830 0.000 707.110 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1512.345 20.485 1513.435 20.655 ;
        RECT 1512.345 19.805 1512.515 20.485 ;
      LAYER mcon ;
        RECT 1513.265 20.485 1513.435 20.655 ;
      LAYER met1 ;
        RECT 1513.205 20.640 1513.495 20.685 ;
        RECT 1527.450 20.640 1527.770 20.700 ;
        RECT 1513.205 20.500 1527.770 20.640 ;
        RECT 1513.205 20.455 1513.495 20.500 ;
        RECT 1527.450 20.440 1527.770 20.500 ;
        RECT 1475.470 19.960 1475.790 20.020 ;
        RECT 1512.285 19.960 1512.575 20.005 ;
        RECT 1475.470 19.820 1512.575 19.960 ;
        RECT 1475.470 19.760 1475.790 19.820 ;
        RECT 1512.285 19.775 1512.575 19.820 ;
      LAYER via ;
        RECT 1527.480 20.440 1527.740 20.700 ;
        RECT 1475.500 19.760 1475.760 20.020 ;
      LAYER met2 ;
        RECT 1475.560 20.050 1475.700 54.000 ;
        RECT 1527.480 20.410 1527.740 20.730 ;
        RECT 1475.500 19.730 1475.760 20.050 ;
        RECT 1527.540 2.400 1527.680 20.410 ;
        RECT 1527.470 0.000 1527.750 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1541.325 48.365 1541.495 54.000 ;
        RECT 1545.465 2.805 1545.635 14.195 ;
      LAYER mcon ;
        RECT 1545.465 14.025 1545.635 14.195 ;
      LAYER met1 ;
        RECT 1541.250 48.520 1541.570 48.580 ;
        RECT 1541.055 48.380 1541.570 48.520 ;
        RECT 1541.250 48.320 1541.570 48.380 ;
        RECT 1541.250 14.180 1541.570 14.240 ;
        RECT 1545.405 14.180 1545.695 14.225 ;
        RECT 1541.250 14.040 1545.695 14.180 ;
        RECT 1541.250 13.980 1541.570 14.040 ;
        RECT 1545.405 13.995 1545.695 14.040 ;
        RECT 1545.390 2.960 1545.710 3.020 ;
        RECT 1545.195 2.820 1545.710 2.960 ;
        RECT 1545.390 2.760 1545.710 2.820 ;
      LAYER via ;
        RECT 1541.280 48.320 1541.540 48.580 ;
        RECT 1541.280 13.980 1541.540 14.240 ;
        RECT 1545.420 2.760 1545.680 3.020 ;
      LAYER met2 ;
        RECT 1541.280 48.290 1541.540 48.610 ;
        RECT 1541.340 14.270 1541.480 48.290 ;
        RECT 1541.280 13.950 1541.540 14.270 ;
        RECT 1545.420 2.730 1545.680 3.050 ;
        RECT 1545.480 2.400 1545.620 2.730 ;
        RECT 1545.410 0.000 1545.690 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1551.370 41.380 1551.690 41.440 ;
        RECT 1563.330 41.380 1563.650 41.440 ;
        RECT 1551.370 41.240 1563.650 41.380 ;
        RECT 1551.370 41.180 1551.690 41.240 ;
        RECT 1563.330 41.180 1563.650 41.240 ;
      LAYER via ;
        RECT 1551.400 41.180 1551.660 41.440 ;
        RECT 1563.360 41.180 1563.620 41.440 ;
      LAYER met2 ;
        RECT 1551.460 41.470 1551.600 54.000 ;
        RECT 1551.400 41.150 1551.660 41.470 ;
        RECT 1563.360 41.150 1563.620 41.470 ;
        RECT 1563.420 2.400 1563.560 41.150 ;
        RECT 1563.350 0.000 1563.630 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1580.900 32.370 1581.040 54.000 ;
        RECT 1580.900 32.230 1581.500 32.370 ;
        RECT 1581.360 2.400 1581.500 32.230 ;
        RECT 1581.290 0.000 1581.570 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1562.025 20.485 1562.195 23.715 ;
      LAYER mcon ;
        RECT 1562.025 23.545 1562.195 23.715 ;
      LAYER met1 ;
        RECT 1485.130 23.700 1485.450 23.760 ;
        RECT 1561.965 23.700 1562.255 23.745 ;
        RECT 1485.130 23.560 1562.255 23.700 ;
        RECT 1485.130 23.500 1485.450 23.560 ;
        RECT 1561.965 23.515 1562.255 23.560 ;
        RECT 1561.965 20.640 1562.255 20.685 ;
        RECT 1598.750 20.640 1599.070 20.700 ;
        RECT 1561.965 20.500 1599.070 20.640 ;
        RECT 1561.965 20.455 1562.255 20.500 ;
        RECT 1598.750 20.440 1599.070 20.500 ;
      LAYER via ;
        RECT 1485.160 23.500 1485.420 23.760 ;
        RECT 1598.780 20.440 1599.040 20.700 ;
      LAYER met2 ;
        RECT 1485.220 23.790 1485.360 54.000 ;
        RECT 1485.160 23.470 1485.420 23.790 ;
        RECT 1598.780 20.410 1599.040 20.730 ;
        RECT 1598.840 2.400 1598.980 20.410 ;
        RECT 1598.770 0.000 1599.050 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1505.445 20.485 1505.615 24.055 ;
      LAYER mcon ;
        RECT 1505.445 23.885 1505.615 24.055 ;
      LAYER met1 ;
        RECT 1484.670 24.040 1484.990 24.100 ;
        RECT 1505.385 24.040 1505.675 24.085 ;
        RECT 1484.670 23.900 1505.675 24.040 ;
        RECT 1484.670 23.840 1484.990 23.900 ;
        RECT 1505.385 23.855 1505.675 23.900 ;
        RECT 1616.690 20.980 1617.010 21.040 ;
        RECT 1512.820 20.840 1617.010 20.980 ;
        RECT 1505.385 20.640 1505.675 20.685 ;
        RECT 1512.820 20.640 1512.960 20.840 ;
        RECT 1616.690 20.780 1617.010 20.840 ;
        RECT 1505.385 20.500 1512.960 20.640 ;
        RECT 1505.385 20.455 1505.675 20.500 ;
      LAYER via ;
        RECT 1484.700 23.840 1484.960 24.100 ;
        RECT 1616.720 20.780 1616.980 21.040 ;
      LAYER met2 ;
        RECT 1484.760 24.130 1484.900 54.000 ;
        RECT 1484.700 23.810 1484.960 24.130 ;
        RECT 1616.720 20.750 1616.980 21.070 ;
        RECT 1616.780 2.400 1616.920 20.750 ;
        RECT 1616.710 0.000 1616.990 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1515.030 22.340 1515.350 22.400 ;
        RECT 1634.630 22.340 1634.950 22.400 ;
        RECT 1515.030 22.200 1634.950 22.340 ;
        RECT 1515.030 22.140 1515.350 22.200 ;
        RECT 1634.630 22.140 1634.950 22.200 ;
        RECT 1491.570 20.980 1491.890 21.040 ;
        RECT 1512.270 20.980 1512.590 21.040 ;
        RECT 1491.570 20.840 1512.590 20.980 ;
        RECT 1491.570 20.780 1491.890 20.840 ;
        RECT 1512.270 20.780 1512.590 20.840 ;
      LAYER via ;
        RECT 1515.060 22.140 1515.320 22.400 ;
        RECT 1634.660 22.140 1634.920 22.400 ;
        RECT 1491.600 20.780 1491.860 21.040 ;
        RECT 1512.300 20.780 1512.560 21.040 ;
      LAYER met2 ;
        RECT 1491.660 21.070 1491.800 54.000 ;
        RECT 1515.060 22.285 1515.320 22.430 ;
        RECT 1512.290 21.915 1512.570 22.285 ;
        RECT 1515.050 21.915 1515.330 22.285 ;
        RECT 1634.660 22.110 1634.920 22.430 ;
        RECT 1512.360 21.070 1512.500 21.915 ;
        RECT 1491.600 20.750 1491.860 21.070 ;
        RECT 1512.300 20.750 1512.560 21.070 ;
        RECT 1634.720 2.400 1634.860 22.110 ;
        RECT 1634.650 0.000 1634.930 2.400 ;
      LAYER via2 ;
        RECT 1512.290 21.960 1512.570 22.240 ;
        RECT 1515.050 21.960 1515.330 22.240 ;
      LAYER met3 ;
        RECT 1512.265 22.250 1512.595 22.265 ;
        RECT 1515.025 22.250 1515.355 22.265 ;
        RECT 1512.265 21.950 1515.355 22.250 ;
        RECT 1512.265 21.935 1512.595 21.950 ;
        RECT 1515.025 21.935 1515.355 21.950 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1652.570 23.020 1652.890 23.080 ;
        RECT 1514.660 22.880 1652.890 23.020 ;
        RECT 1492.490 22.340 1492.810 22.400 ;
        RECT 1514.660 22.340 1514.800 22.880 ;
        RECT 1652.570 22.820 1652.890 22.880 ;
        RECT 1492.490 22.200 1514.800 22.340 ;
        RECT 1492.490 22.140 1492.810 22.200 ;
      LAYER via ;
        RECT 1492.520 22.140 1492.780 22.400 ;
        RECT 1652.600 22.820 1652.860 23.080 ;
      LAYER met2 ;
        RECT 1492.580 22.430 1492.720 54.000 ;
        RECT 1652.600 22.790 1652.860 23.110 ;
        RECT 1492.520 22.110 1492.780 22.430 ;
        RECT 1652.660 2.400 1652.800 22.790 ;
        RECT 1652.590 0.000 1652.870 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1512.805 26.265 1512.975 28.135 ;
      LAYER mcon ;
        RECT 1512.805 27.965 1512.975 28.135 ;
      LAYER met1 ;
        RECT 1512.745 28.120 1513.035 28.165 ;
        RECT 1560.110 28.120 1560.430 28.180 ;
        RECT 1512.745 27.980 1560.430 28.120 ;
        RECT 1512.745 27.935 1513.035 27.980 ;
        RECT 1560.110 27.920 1560.430 27.980 ;
        RECT 1498.930 26.420 1499.250 26.480 ;
        RECT 1512.745 26.420 1513.035 26.465 ;
        RECT 1498.930 26.280 1513.035 26.420 ;
        RECT 1498.930 26.220 1499.250 26.280 ;
        RECT 1512.745 26.235 1513.035 26.280 ;
        RECT 1561.490 23.360 1561.810 23.420 ;
        RECT 1670.510 23.360 1670.830 23.420 ;
        RECT 1561.490 23.220 1670.830 23.360 ;
        RECT 1561.490 23.160 1561.810 23.220 ;
        RECT 1670.510 23.160 1670.830 23.220 ;
      LAYER via ;
        RECT 1560.140 27.920 1560.400 28.180 ;
        RECT 1498.960 26.220 1499.220 26.480 ;
        RECT 1561.520 23.160 1561.780 23.420 ;
        RECT 1670.540 23.160 1670.800 23.420 ;
      LAYER met2 ;
        RECT 1499.020 26.510 1499.160 54.000 ;
        RECT 1560.140 27.890 1560.400 28.210 ;
        RECT 1560.200 26.930 1560.340 27.890 ;
        RECT 1560.200 26.790 1561.720 26.930 ;
        RECT 1498.960 26.190 1499.220 26.510 ;
        RECT 1561.580 23.450 1561.720 26.790 ;
        RECT 1561.520 23.130 1561.780 23.450 ;
        RECT 1670.540 23.130 1670.800 23.450 ;
        RECT 1670.600 2.400 1670.740 23.130 ;
        RECT 1670.530 0.000 1670.810 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1514.185 23.035 1514.355 24.055 ;
        RECT 1513.725 22.865 1514.355 23.035 ;
      LAYER mcon ;
        RECT 1514.185 23.885 1514.355 24.055 ;
      LAYER met1 ;
        RECT 1514.125 24.040 1514.415 24.085 ;
        RECT 1609.790 24.040 1610.110 24.100 ;
        RECT 1514.125 23.900 1610.110 24.040 ;
        RECT 1514.125 23.855 1514.415 23.900 ;
        RECT 1609.790 23.840 1610.110 23.900 ;
        RECT 1610.710 24.040 1611.030 24.100 ;
        RECT 1687.990 24.040 1688.310 24.100 ;
        RECT 1610.710 23.900 1688.310 24.040 ;
        RECT 1610.710 23.840 1611.030 23.900 ;
        RECT 1687.990 23.840 1688.310 23.900 ;
        RECT 1498.470 23.020 1498.790 23.080 ;
        RECT 1513.665 23.020 1513.955 23.065 ;
        RECT 1498.470 22.880 1513.955 23.020 ;
        RECT 1498.470 22.820 1498.790 22.880 ;
        RECT 1513.665 22.835 1513.955 22.880 ;
      LAYER via ;
        RECT 1609.820 23.840 1610.080 24.100 ;
        RECT 1610.740 23.840 1611.000 24.100 ;
        RECT 1688.020 23.840 1688.280 24.100 ;
        RECT 1498.500 22.820 1498.760 23.080 ;
      LAYER met2 ;
        RECT 1498.560 23.110 1498.700 54.000 ;
        RECT 1609.820 23.810 1610.080 24.130 ;
        RECT 1610.740 23.810 1611.000 24.130 ;
        RECT 1688.020 23.810 1688.280 24.130 ;
        RECT 1609.880 23.645 1610.020 23.810 ;
        RECT 1610.800 23.645 1610.940 23.810 ;
        RECT 1609.810 23.275 1610.090 23.645 ;
        RECT 1610.730 23.275 1611.010 23.645 ;
        RECT 1498.500 22.790 1498.760 23.110 ;
        RECT 1688.080 2.400 1688.220 23.810 ;
        RECT 1688.010 0.000 1688.290 2.400 ;
      LAYER via2 ;
        RECT 1609.810 23.320 1610.090 23.600 ;
        RECT 1610.730 23.320 1611.010 23.600 ;
      LAYER met3 ;
        RECT 1609.785 23.610 1610.115 23.625 ;
        RECT 1610.705 23.610 1611.035 23.625 ;
        RECT 1609.785 23.310 1611.035 23.610 ;
        RECT 1609.785 23.295 1610.115 23.310 ;
        RECT 1610.705 23.295 1611.035 23.310 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 725.300 3.130 725.440 54.000 ;
        RECT 724.840 2.990 725.440 3.130 ;
        RECT 724.840 2.400 724.980 2.990 ;
        RECT 724.770 0.000 725.050 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1586.405 25.585 1586.575 26.775 ;
      LAYER mcon ;
        RECT 1586.405 26.605 1586.575 26.775 ;
      LAYER met1 ;
        RECT 1586.345 26.760 1586.635 26.805 ;
        RECT 1705.930 26.760 1706.250 26.820 ;
        RECT 1586.345 26.620 1706.250 26.760 ;
        RECT 1586.345 26.575 1586.635 26.620 ;
        RECT 1705.930 26.560 1706.250 26.620 ;
        RECT 1537.570 25.740 1537.890 25.800 ;
        RECT 1586.345 25.740 1586.635 25.785 ;
        RECT 1537.570 25.600 1586.635 25.740 ;
        RECT 1537.570 25.540 1537.890 25.600 ;
        RECT 1586.345 25.555 1586.635 25.600 ;
        RECT 1504.910 25.060 1505.230 25.120 ;
        RECT 1537.570 25.060 1537.890 25.120 ;
        RECT 1504.910 24.920 1537.890 25.060 ;
        RECT 1504.910 24.860 1505.230 24.920 ;
        RECT 1537.570 24.860 1537.890 24.920 ;
      LAYER via ;
        RECT 1705.960 26.560 1706.220 26.820 ;
        RECT 1537.600 25.540 1537.860 25.800 ;
        RECT 1504.940 24.860 1505.200 25.120 ;
        RECT 1537.600 24.860 1537.860 25.120 ;
      LAYER met2 ;
        RECT 1505.000 25.150 1505.140 54.000 ;
        RECT 1705.960 26.530 1706.220 26.850 ;
        RECT 1537.600 25.510 1537.860 25.830 ;
        RECT 1537.660 25.150 1537.800 25.510 ;
        RECT 1504.940 24.830 1505.200 25.150 ;
        RECT 1537.600 24.830 1537.860 25.150 ;
        RECT 1706.020 2.400 1706.160 26.530 ;
        RECT 1705.950 0.000 1706.230 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1561.105 26.605 1561.275 28.815 ;
        RECT 1563.405 26.265 1563.575 28.815 ;
        RECT 1585.485 25.415 1585.655 26.435 ;
        RECT 1586.865 25.415 1587.035 25.755 ;
        RECT 1585.485 25.245 1587.035 25.415 ;
        RECT 1661.845 22.865 1662.015 25.755 ;
      LAYER mcon ;
        RECT 1561.105 28.645 1561.275 28.815 ;
        RECT 1563.405 28.645 1563.575 28.815 ;
        RECT 1585.485 26.265 1585.655 26.435 ;
        RECT 1586.865 25.585 1587.035 25.755 ;
        RECT 1661.845 25.585 1662.015 25.755 ;
      LAYER met1 ;
        RECT 1561.045 28.800 1561.335 28.845 ;
        RECT 1563.345 28.800 1563.635 28.845 ;
        RECT 1561.045 28.660 1563.635 28.800 ;
        RECT 1561.045 28.615 1561.335 28.660 ;
        RECT 1563.345 28.615 1563.635 28.660 ;
        RECT 1505.370 26.760 1505.690 26.820 ;
        RECT 1561.045 26.760 1561.335 26.805 ;
        RECT 1505.370 26.620 1561.335 26.760 ;
        RECT 1505.370 26.560 1505.690 26.620 ;
        RECT 1561.045 26.575 1561.335 26.620 ;
        RECT 1563.345 26.420 1563.635 26.465 ;
        RECT 1585.425 26.420 1585.715 26.465 ;
        RECT 1563.345 26.280 1585.715 26.420 ;
        RECT 1563.345 26.235 1563.635 26.280 ;
        RECT 1585.425 26.235 1585.715 26.280 ;
        RECT 1586.805 25.740 1587.095 25.785 ;
        RECT 1661.785 25.740 1662.075 25.785 ;
        RECT 1586.805 25.600 1662.075 25.740 ;
        RECT 1586.805 25.555 1587.095 25.600 ;
        RECT 1661.785 25.555 1662.075 25.600 ;
        RECT 1661.785 23.020 1662.075 23.065 ;
        RECT 1723.870 23.020 1724.190 23.080 ;
        RECT 1661.785 22.880 1724.190 23.020 ;
        RECT 1661.785 22.835 1662.075 22.880 ;
        RECT 1723.870 22.820 1724.190 22.880 ;
      LAYER via ;
        RECT 1505.400 26.560 1505.660 26.820 ;
        RECT 1723.900 22.820 1724.160 23.080 ;
      LAYER met2 ;
        RECT 1505.460 26.850 1505.600 54.000 ;
        RECT 1505.400 26.530 1505.660 26.850 ;
        RECT 1723.900 22.790 1724.160 23.110 ;
        RECT 1723.960 2.400 1724.100 22.790 ;
        RECT 1723.890 0.000 1724.170 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1512.820 24.325 1512.960 54.000 ;
        RECT 1512.750 23.955 1513.030 24.325 ;
        RECT 1741.830 23.955 1742.110 24.325 ;
        RECT 1741.900 2.400 1742.040 23.955 ;
        RECT 1741.830 0.000 1742.110 2.400 ;
      LAYER via2 ;
        RECT 1512.750 24.000 1513.030 24.280 ;
        RECT 1741.830 24.000 1742.110 24.280 ;
      LAYER met3 ;
        RECT 1512.725 24.290 1513.055 24.305 ;
        RECT 1741.805 24.290 1742.135 24.305 ;
        RECT 1512.725 23.990 1742.135 24.290 ;
        RECT 1512.725 23.975 1513.055 23.990 ;
        RECT 1741.805 23.975 1742.135 23.990 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.620 48.805 1756.760 54.000 ;
        RECT 1756.550 48.435 1756.830 48.805 ;
        RECT 1757.930 48.435 1758.210 48.805 ;
        RECT 1758.000 24.210 1758.140 48.435 ;
        RECT 1758.000 24.070 1759.520 24.210 ;
        RECT 1759.380 2.400 1759.520 24.070 ;
        RECT 1759.310 0.000 1759.590 2.400 ;
      LAYER via2 ;
        RECT 1756.550 48.480 1756.830 48.760 ;
        RECT 1757.930 48.480 1758.210 48.760 ;
      LAYER met3 ;
        RECT 1756.525 48.770 1756.855 48.785 ;
        RECT 1757.905 48.770 1758.235 48.785 ;
        RECT 1756.525 48.470 1758.235 48.770 ;
        RECT 1756.525 48.455 1756.855 48.470 ;
        RECT 1757.905 48.455 1758.235 48.470 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1775.940 14.010 1776.080 54.000 ;
        RECT 1775.940 13.870 1776.540 14.010 ;
        RECT 1776.400 13.330 1776.540 13.870 ;
        RECT 1776.400 13.190 1777.460 13.330 ;
        RECT 1777.320 2.400 1777.460 13.190 ;
        RECT 1777.250 0.000 1777.530 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1790.110 13.160 1790.430 13.220 ;
        RECT 1795.170 13.160 1795.490 13.220 ;
        RECT 1790.110 13.020 1795.490 13.160 ;
        RECT 1790.110 12.960 1790.430 13.020 ;
        RECT 1795.170 12.960 1795.490 13.020 ;
      LAYER via ;
        RECT 1790.140 12.960 1790.400 13.220 ;
        RECT 1795.200 12.960 1795.460 13.220 ;
      LAYER met2 ;
        RECT 1789.740 37.810 1789.880 54.000 ;
        RECT 1789.740 37.670 1790.340 37.810 ;
        RECT 1790.200 13.250 1790.340 37.670 ;
        RECT 1790.140 12.930 1790.400 13.250 ;
        RECT 1795.200 12.930 1795.460 13.250 ;
        RECT 1795.260 2.400 1795.400 12.930 ;
        RECT 1795.190 0.000 1795.470 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1810.350 13.160 1810.670 13.220 ;
        RECT 1813.110 13.160 1813.430 13.220 ;
        RECT 1810.350 13.020 1813.430 13.160 ;
        RECT 1810.350 12.960 1810.670 13.020 ;
        RECT 1813.110 12.960 1813.430 13.020 ;
      LAYER via ;
        RECT 1810.380 12.960 1810.640 13.220 ;
        RECT 1813.140 12.960 1813.400 13.220 ;
      LAYER met2 ;
        RECT 1810.440 13.250 1810.580 54.000 ;
        RECT 1810.380 12.930 1810.640 13.250 ;
        RECT 1813.140 12.930 1813.400 13.250 ;
        RECT 1813.200 2.400 1813.340 12.930 ;
        RECT 1813.130 0.000 1813.410 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1831.140 2.400 1831.280 54.000 ;
        RECT 1831.070 0.000 1831.350 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1848.160 12.650 1848.300 54.000 ;
        RECT 1848.160 12.510 1848.760 12.650 ;
        RECT 1848.620 2.400 1848.760 12.510 ;
        RECT 1848.550 0.000 1848.830 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1865.625 41.905 1865.795 54.000 ;
      LAYER met1 ;
        RECT 1865.550 42.060 1865.870 42.120 ;
        RECT 1865.355 41.920 1865.870 42.060 ;
        RECT 1865.550 41.860 1865.870 41.920 ;
      LAYER via ;
        RECT 1865.580 41.860 1865.840 42.120 ;
      LAYER met2 ;
        RECT 1865.580 41.830 1865.840 42.150 ;
        RECT 1865.640 14.010 1865.780 41.830 ;
        RECT 1865.180 13.870 1865.780 14.010 ;
        RECT 1865.180 12.650 1865.320 13.870 ;
        RECT 1865.180 12.510 1866.700 12.650 ;
        RECT 1866.560 2.400 1866.700 12.510 ;
        RECT 1866.490 0.000 1866.770 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 742.690 18.260 743.010 18.320 ;
        RECT 747.290 18.260 747.610 18.320 ;
        RECT 742.690 18.120 747.610 18.260 ;
        RECT 742.690 18.060 743.010 18.120 ;
        RECT 747.290 18.060 747.610 18.120 ;
      LAYER via ;
        RECT 742.720 18.060 742.980 18.320 ;
        RECT 747.320 18.060 747.580 18.320 ;
      LAYER met2 ;
        RECT 747.380 18.350 747.520 54.000 ;
        RECT 742.720 18.030 742.980 18.350 ;
        RECT 747.320 18.030 747.580 18.350 ;
        RECT 742.780 2.400 742.920 18.030 ;
        RECT 742.710 0.000 742.990 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1538.950 30.840 1539.270 30.900 ;
        RECT 1851.750 30.840 1852.070 30.900 ;
        RECT 1538.950 30.700 1852.070 30.840 ;
        RECT 1538.950 30.640 1539.270 30.700 ;
        RECT 1851.750 30.640 1852.070 30.700 ;
      LAYER via ;
        RECT 1538.980 30.640 1539.240 30.900 ;
        RECT 1851.780 30.640 1852.040 30.900 ;
      LAYER met2 ;
        RECT 1539.040 30.930 1539.180 54.000 ;
        RECT 1538.980 30.610 1539.240 30.930 ;
        RECT 1851.780 30.610 1852.040 30.930 ;
        RECT 1851.840 29.765 1851.980 30.610 ;
        RECT 1851.770 29.395 1852.050 29.765 ;
        RECT 1884.430 29.395 1884.710 29.765 ;
        RECT 1884.500 2.400 1884.640 29.395 ;
        RECT 1884.430 0.000 1884.710 2.400 ;
      LAYER via2 ;
        RECT 1851.770 29.440 1852.050 29.720 ;
        RECT 1884.430 29.440 1884.710 29.720 ;
      LAYER met3 ;
        RECT 1851.745 29.730 1852.075 29.745 ;
        RECT 1884.405 29.730 1884.735 29.745 ;
        RECT 1851.745 29.430 1884.735 29.730 ;
        RECT 1851.745 29.415 1852.075 29.430 ;
        RECT 1884.405 29.415 1884.735 29.430 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1561.565 27.625 1561.735 30.515 ;
        RECT 1854.125 15.895 1854.295 27.795 ;
        RECT 1854.125 15.725 1873.615 15.895 ;
        RECT 1873.445 12.325 1873.615 15.725 ;
      LAYER mcon ;
        RECT 1561.565 30.345 1561.735 30.515 ;
        RECT 1854.125 27.625 1854.295 27.795 ;
      LAYER met1 ;
        RECT 1546.770 30.500 1547.090 30.560 ;
        RECT 1561.505 30.500 1561.795 30.545 ;
        RECT 1546.770 30.360 1561.795 30.500 ;
        RECT 1546.770 30.300 1547.090 30.360 ;
        RECT 1561.505 30.315 1561.795 30.360 ;
        RECT 1561.505 27.780 1561.795 27.825 ;
        RECT 1854.065 27.780 1854.355 27.825 ;
        RECT 1561.505 27.640 1854.355 27.780 ;
        RECT 1561.505 27.595 1561.795 27.640 ;
        RECT 1854.065 27.595 1854.355 27.640 ;
        RECT 1873.385 12.480 1873.675 12.525 ;
        RECT 1902.350 12.480 1902.670 12.540 ;
        RECT 1873.385 12.340 1902.670 12.480 ;
        RECT 1873.385 12.295 1873.675 12.340 ;
        RECT 1902.350 12.280 1902.670 12.340 ;
      LAYER via ;
        RECT 1546.800 30.300 1547.060 30.560 ;
        RECT 1902.380 12.280 1902.640 12.540 ;
      LAYER met2 ;
        RECT 1546.860 30.590 1547.000 54.000 ;
        RECT 1546.800 30.270 1547.060 30.590 ;
        RECT 1902.380 12.250 1902.640 12.570 ;
        RECT 1902.440 2.400 1902.580 12.250 ;
        RECT 1902.370 0.000 1902.650 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1853.665 27.965 1854.755 28.135 ;
        RECT 1854.585 16.235 1854.755 27.965 ;
        RECT 1854.585 16.065 1874.075 16.235 ;
        RECT 1873.905 11.985 1874.075 16.065 ;
      LAYER met1 ;
        RECT 1853.605 28.120 1853.895 28.165 ;
        RECT 1561.120 27.980 1853.895 28.120 ;
        RECT 1547.230 27.780 1547.550 27.840 ;
        RECT 1561.120 27.780 1561.260 27.980 ;
        RECT 1853.605 27.935 1853.895 27.980 ;
        RECT 1547.230 27.640 1561.260 27.780 ;
        RECT 1547.230 27.580 1547.550 27.640 ;
        RECT 1873.845 12.140 1874.135 12.185 ;
        RECT 1920.290 12.140 1920.610 12.200 ;
        RECT 1873.845 12.000 1920.610 12.140 ;
        RECT 1873.845 11.955 1874.135 12.000 ;
        RECT 1920.290 11.940 1920.610 12.000 ;
      LAYER via ;
        RECT 1547.260 27.580 1547.520 27.840 ;
        RECT 1920.320 11.940 1920.580 12.200 ;
      LAYER met2 ;
        RECT 1547.320 27.870 1547.460 54.000 ;
        RECT 1547.260 27.550 1547.520 27.870 ;
        RECT 1920.320 11.910 1920.580 12.230 ;
        RECT 1920.380 2.400 1920.520 11.910 ;
        RECT 1920.310 0.000 1920.590 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1573.065 28.305 1573.235 31.535 ;
      LAYER mcon ;
        RECT 1573.065 31.365 1573.235 31.535 ;
      LAYER met1 ;
        RECT 1554.130 31.520 1554.450 31.580 ;
        RECT 1573.005 31.520 1573.295 31.565 ;
        RECT 1554.130 31.380 1573.295 31.520 ;
        RECT 1554.130 31.320 1554.450 31.380 ;
        RECT 1573.005 31.335 1573.295 31.380 ;
        RECT 1573.005 28.460 1573.295 28.505 ;
        RECT 1937.770 28.460 1938.090 28.520 ;
        RECT 1573.005 28.320 1938.090 28.460 ;
        RECT 1573.005 28.275 1573.295 28.320 ;
        RECT 1937.770 28.260 1938.090 28.320 ;
      LAYER via ;
        RECT 1554.160 31.320 1554.420 31.580 ;
        RECT 1937.800 28.260 1938.060 28.520 ;
      LAYER met2 ;
        RECT 1554.220 31.610 1554.360 54.000 ;
        RECT 1554.160 31.290 1554.420 31.610 ;
        RECT 1937.800 28.230 1938.060 28.550 ;
        RECT 1937.860 2.400 1938.000 28.230 ;
        RECT 1937.790 0.000 1938.070 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1585.945 28.645 1586.115 31.875 ;
      LAYER mcon ;
        RECT 1585.945 31.705 1586.115 31.875 ;
      LAYER met1 ;
        RECT 1553.670 31.860 1553.990 31.920 ;
        RECT 1585.885 31.860 1586.175 31.905 ;
        RECT 1553.670 31.720 1586.175 31.860 ;
        RECT 1553.670 31.660 1553.990 31.720 ;
        RECT 1585.885 31.675 1586.175 31.720 ;
        RECT 1585.885 28.800 1586.175 28.845 ;
        RECT 1955.710 28.800 1956.030 28.860 ;
        RECT 1585.885 28.660 1956.030 28.800 ;
        RECT 1585.885 28.615 1586.175 28.660 ;
        RECT 1955.710 28.600 1956.030 28.660 ;
      LAYER via ;
        RECT 1553.700 31.660 1553.960 31.920 ;
        RECT 1955.740 28.600 1956.000 28.860 ;
      LAYER met2 ;
        RECT 1553.760 31.950 1553.900 54.000 ;
        RECT 1553.700 31.630 1553.960 31.950 ;
        RECT 1955.740 28.570 1956.000 28.890 ;
        RECT 1955.800 2.400 1955.940 28.570 ;
        RECT 1955.730 0.000 1956.010 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1560.570 29.280 1560.890 29.540 ;
        RECT 1560.660 29.140 1560.800 29.280 ;
        RECT 1973.650 29.140 1973.970 29.200 ;
        RECT 1560.660 29.000 1973.970 29.140 ;
        RECT 1973.650 28.940 1973.970 29.000 ;
      LAYER via ;
        RECT 1560.600 29.280 1560.860 29.540 ;
        RECT 1973.680 28.940 1973.940 29.200 ;
      LAYER met2 ;
        RECT 1560.660 29.570 1560.800 54.000 ;
        RECT 1560.600 29.250 1560.860 29.570 ;
        RECT 1973.680 28.910 1973.940 29.230 ;
        RECT 1973.740 2.400 1973.880 28.910 ;
        RECT 1973.670 0.000 1973.950 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1561.030 29.480 1561.350 29.540 ;
        RECT 1991.590 29.480 1991.910 29.540 ;
        RECT 1561.030 29.340 1991.910 29.480 ;
        RECT 1561.030 29.280 1561.350 29.340 ;
        RECT 1991.590 29.280 1991.910 29.340 ;
      LAYER via ;
        RECT 1561.060 29.280 1561.320 29.540 ;
        RECT 1991.620 29.280 1991.880 29.540 ;
      LAYER met2 ;
        RECT 1561.120 29.570 1561.260 54.000 ;
        RECT 1561.060 29.250 1561.320 29.570 ;
        RECT 1991.620 29.250 1991.880 29.570 ;
        RECT 1991.680 2.400 1991.820 29.250 ;
        RECT 1991.610 0.000 1991.890 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1567.930 32.200 1568.250 32.260 ;
        RECT 1567.930 32.060 1586.560 32.200 ;
        RECT 1567.930 32.000 1568.250 32.060 ;
        RECT 1586.420 31.860 1586.560 32.060 ;
        RECT 1594.150 31.860 1594.470 31.920 ;
        RECT 1586.420 31.720 1594.470 31.860 ;
        RECT 1594.150 31.660 1594.470 31.720 ;
        RECT 1609.790 30.500 1610.110 30.560 ;
        RECT 2009.070 30.500 2009.390 30.560 ;
        RECT 1609.790 30.360 2009.390 30.500 ;
        RECT 1609.790 30.300 1610.110 30.360 ;
        RECT 2009.070 30.300 2009.390 30.360 ;
      LAYER via ;
        RECT 1567.960 32.000 1568.220 32.260 ;
        RECT 1594.180 31.660 1594.440 31.920 ;
        RECT 1609.820 30.300 1610.080 30.560 ;
        RECT 2009.100 30.300 2009.360 30.560 ;
      LAYER met2 ;
        RECT 1568.020 32.290 1568.160 54.000 ;
        RECT 1567.960 31.970 1568.220 32.290 ;
        RECT 1594.180 31.805 1594.440 31.950 ;
        RECT 1594.170 31.435 1594.450 31.805 ;
        RECT 1609.810 31.435 1610.090 31.805 ;
        RECT 1609.880 30.590 1610.020 31.435 ;
        RECT 1609.820 30.270 1610.080 30.590 ;
        RECT 2009.100 30.270 2009.360 30.590 ;
        RECT 2009.160 2.400 2009.300 30.270 ;
        RECT 2009.090 0.000 2009.370 2.400 ;
      LAYER via2 ;
        RECT 1594.170 31.480 1594.450 31.760 ;
        RECT 1609.810 31.480 1610.090 31.760 ;
      LAYER met3 ;
        RECT 1594.145 31.770 1594.475 31.785 ;
        RECT 1609.785 31.770 1610.115 31.785 ;
        RECT 1594.145 31.470 1610.115 31.770 ;
        RECT 1594.145 31.455 1594.475 31.470 ;
        RECT 1609.785 31.455 1610.115 31.470 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1567.470 34.240 1567.790 34.300 ;
        RECT 2027.010 34.240 2027.330 34.300 ;
        RECT 1567.470 34.100 2027.330 34.240 ;
        RECT 1567.470 34.040 1567.790 34.100 ;
        RECT 2027.010 34.040 2027.330 34.100 ;
      LAYER via ;
        RECT 1567.500 34.040 1567.760 34.300 ;
        RECT 2027.040 34.040 2027.300 34.300 ;
      LAYER met2 ;
        RECT 1567.560 34.330 1567.700 54.000 ;
        RECT 1567.500 34.010 1567.760 34.330 ;
        RECT 2027.040 34.010 2027.300 34.330 ;
        RECT 2027.100 2.400 2027.240 34.010 ;
        RECT 2027.030 0.000 2027.310 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1574.830 33.900 1575.150 33.960 ;
        RECT 2044.950 33.900 2045.270 33.960 ;
        RECT 1574.830 33.760 2045.270 33.900 ;
        RECT 1574.830 33.700 1575.150 33.760 ;
        RECT 2044.950 33.700 2045.270 33.760 ;
      LAYER via ;
        RECT 1574.860 33.700 1575.120 33.960 ;
        RECT 2044.980 33.700 2045.240 33.960 ;
      LAYER met2 ;
        RECT 1574.920 33.990 1575.060 54.000 ;
        RECT 1574.860 33.670 1575.120 33.990 ;
        RECT 2044.980 33.670 2045.240 33.990 ;
        RECT 2045.040 2.400 2045.180 33.670 ;
        RECT 2044.970 0.000 2045.250 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 760.170 2.960 760.490 3.020 ;
        RECT 760.630 2.960 760.950 3.020 ;
        RECT 760.170 2.820 760.950 2.960 ;
        RECT 760.170 2.760 760.490 2.820 ;
        RECT 760.630 2.760 760.950 2.820 ;
      LAYER via ;
        RECT 760.200 2.760 760.460 3.020 ;
        RECT 760.660 2.760 760.920 3.020 ;
      LAYER met2 ;
        RECT 759.340 48.805 759.480 54.000 ;
        RECT 759.270 48.435 759.550 48.805 ;
        RECT 760.190 48.435 760.470 48.805 ;
        RECT 760.260 47.840 760.400 48.435 ;
        RECT 760.260 47.700 760.860 47.840 ;
        RECT 760.720 3.050 760.860 47.700 ;
        RECT 760.200 2.730 760.460 3.050 ;
        RECT 760.660 2.730 760.920 3.050 ;
        RECT 760.260 2.400 760.400 2.730 ;
        RECT 760.190 0.000 760.470 2.400 ;
      LAYER via2 ;
        RECT 759.270 48.480 759.550 48.760 ;
        RECT 760.190 48.480 760.470 48.760 ;
      LAYER met3 ;
        RECT 759.245 48.770 759.575 48.785 ;
        RECT 760.165 48.770 760.495 48.785 ;
        RECT 759.245 48.470 760.495 48.770 ;
        RECT 759.245 48.455 759.575 48.470 ;
        RECT 760.165 48.455 760.495 48.470 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1581.730 33.560 1582.050 33.620 ;
        RECT 2062.890 33.560 2063.210 33.620 ;
        RECT 1581.730 33.420 2063.210 33.560 ;
        RECT 1581.730 33.360 1582.050 33.420 ;
        RECT 2062.890 33.360 2063.210 33.420 ;
      LAYER via ;
        RECT 1581.760 33.360 1582.020 33.620 ;
        RECT 2062.920 33.360 2063.180 33.620 ;
      LAYER met2 ;
        RECT 1581.820 33.650 1581.960 54.000 ;
        RECT 1581.760 33.330 1582.020 33.650 ;
        RECT 2062.920 33.330 2063.180 33.650 ;
        RECT 2062.980 2.400 2063.120 33.330 ;
        RECT 2062.910 0.000 2063.190 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1581.270 33.220 1581.590 33.280 ;
        RECT 2080.830 33.220 2081.150 33.280 ;
        RECT 1581.270 33.080 2081.150 33.220 ;
        RECT 1581.270 33.020 1581.590 33.080 ;
        RECT 2080.830 33.020 2081.150 33.080 ;
      LAYER via ;
        RECT 1581.300 33.020 1581.560 33.280 ;
        RECT 2080.860 33.020 2081.120 33.280 ;
      LAYER met2 ;
        RECT 1581.360 33.310 1581.500 54.000 ;
        RECT 1581.300 32.990 1581.560 33.310 ;
        RECT 2080.860 32.990 2081.120 33.310 ;
        RECT 2080.920 2.400 2081.060 32.990 ;
        RECT 2080.850 0.000 2081.130 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1619.065 32.045 1619.235 36.295 ;
      LAYER mcon ;
        RECT 1619.065 36.125 1619.235 36.295 ;
      LAYER met1 ;
        RECT 1588.170 36.280 1588.490 36.340 ;
        RECT 1619.005 36.280 1619.295 36.325 ;
        RECT 1588.170 36.140 1619.295 36.280 ;
        RECT 1588.170 36.080 1588.490 36.140 ;
        RECT 1619.005 36.095 1619.295 36.140 ;
        RECT 1619.005 32.200 1619.295 32.245 ;
        RECT 2098.310 32.200 2098.630 32.260 ;
        RECT 1619.005 32.060 2098.630 32.200 ;
        RECT 1619.005 32.015 1619.295 32.060 ;
        RECT 2098.310 32.000 2098.630 32.060 ;
      LAYER via ;
        RECT 1588.200 36.080 1588.460 36.340 ;
        RECT 2098.340 32.000 2098.600 32.260 ;
      LAYER met2 ;
        RECT 1588.260 36.370 1588.400 54.000 ;
        RECT 1588.200 36.050 1588.460 36.370 ;
        RECT 2098.340 31.970 2098.600 32.290 ;
        RECT 2098.400 2.400 2098.540 31.970 ;
        RECT 2098.330 0.000 2098.610 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1609.405 31.875 1609.575 32.215 ;
        RECT 1609.405 31.705 1610.495 31.875 ;
        RECT 1789.725 31.705 1790.815 31.875 ;
      LAYER mcon ;
        RECT 1609.405 32.045 1609.575 32.215 ;
        RECT 1610.325 31.705 1610.495 31.875 ;
        RECT 1790.645 31.705 1790.815 31.875 ;
      LAYER met1 ;
        RECT 1588.630 32.200 1588.950 32.260 ;
        RECT 1609.345 32.200 1609.635 32.245 ;
        RECT 1588.630 32.060 1609.635 32.200 ;
        RECT 1588.630 32.000 1588.950 32.060 ;
        RECT 1609.345 32.015 1609.635 32.060 ;
        RECT 1610.265 31.860 1610.555 31.905 ;
        RECT 1789.665 31.860 1789.955 31.905 ;
        RECT 1610.265 31.720 1789.955 31.860 ;
        RECT 1610.265 31.675 1610.555 31.720 ;
        RECT 1789.665 31.675 1789.955 31.720 ;
        RECT 1790.585 31.860 1790.875 31.905 ;
        RECT 2116.250 31.860 2116.570 31.920 ;
        RECT 1790.585 31.720 2116.570 31.860 ;
        RECT 1790.585 31.675 1790.875 31.720 ;
        RECT 2116.250 31.660 2116.570 31.720 ;
      LAYER via ;
        RECT 1588.660 32.000 1588.920 32.260 ;
        RECT 2116.280 31.660 2116.540 31.920 ;
      LAYER met2 ;
        RECT 1588.720 32.290 1588.860 54.000 ;
        RECT 1588.660 31.970 1588.920 32.290 ;
        RECT 2116.280 31.630 2116.540 31.950 ;
        RECT 2116.340 2.400 2116.480 31.630 ;
        RECT 2116.270 0.000 2116.550 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1643.445 31.365 1644.535 31.535 ;
        RECT 1734.525 31.365 1735.155 31.535 ;
        RECT 2120.925 30.345 2121.095 31.535 ;
      LAYER mcon ;
        RECT 1644.365 31.365 1644.535 31.535 ;
        RECT 1734.985 31.365 1735.155 31.535 ;
        RECT 2120.925 31.365 2121.095 31.535 ;
      LAYER met1 ;
        RECT 1643.370 31.520 1643.690 31.580 ;
        RECT 1644.305 31.520 1644.595 31.565 ;
        RECT 1686.150 31.520 1686.470 31.580 ;
        RECT 1643.370 31.380 1643.885 31.520 ;
        RECT 1644.305 31.380 1686.470 31.520 ;
        RECT 1643.370 31.320 1643.690 31.380 ;
        RECT 1644.305 31.335 1644.595 31.380 ;
        RECT 1686.150 31.320 1686.470 31.380 ;
        RECT 1693.970 31.520 1694.290 31.580 ;
        RECT 1734.465 31.520 1734.755 31.565 ;
        RECT 1734.910 31.520 1735.230 31.580 ;
        RECT 1693.970 31.380 1735.230 31.520 ;
        RECT 1693.970 31.320 1694.290 31.380 ;
        RECT 1734.465 31.335 1734.755 31.380 ;
        RECT 1734.910 31.320 1735.230 31.380 ;
        RECT 1782.290 31.520 1782.610 31.580 ;
        RECT 2120.865 31.520 2121.155 31.565 ;
        RECT 1782.290 31.380 2121.155 31.520 ;
        RECT 1782.290 31.320 1782.610 31.380 ;
        RECT 2120.865 31.335 2121.155 31.380 ;
        RECT 2120.865 30.500 2121.155 30.545 ;
        RECT 2134.190 30.500 2134.510 30.560 ;
        RECT 2120.865 30.360 2134.510 30.500 ;
        RECT 2120.865 30.315 2121.155 30.360 ;
        RECT 2134.190 30.300 2134.510 30.360 ;
      LAYER via ;
        RECT 1643.400 31.320 1643.660 31.580 ;
        RECT 1686.180 31.320 1686.440 31.580 ;
        RECT 1694.000 31.320 1694.260 31.580 ;
        RECT 1734.940 31.320 1735.200 31.580 ;
        RECT 1782.320 31.320 1782.580 31.580 ;
        RECT 2134.220 30.300 2134.480 30.560 ;
      LAYER met2 ;
        RECT 1594.700 32.485 1594.840 54.000 ;
        RECT 1594.630 32.115 1594.910 32.485 ;
        RECT 1643.390 32.115 1643.670 32.485 ;
        RECT 1686.170 32.115 1686.450 32.485 ;
        RECT 1693.990 32.115 1694.270 32.485 ;
        RECT 1734.930 32.115 1735.210 32.485 ;
        RECT 1782.310 32.115 1782.590 32.485 ;
        RECT 1643.460 31.610 1643.600 32.115 ;
        RECT 1686.240 31.610 1686.380 32.115 ;
        RECT 1694.060 31.610 1694.200 32.115 ;
        RECT 1735.000 31.610 1735.140 32.115 ;
        RECT 1782.380 31.610 1782.520 32.115 ;
        RECT 1643.400 31.290 1643.660 31.610 ;
        RECT 1686.180 31.290 1686.440 31.610 ;
        RECT 1694.000 31.290 1694.260 31.610 ;
        RECT 1734.940 31.290 1735.200 31.610 ;
        RECT 1782.320 31.290 1782.580 31.610 ;
        RECT 2134.220 30.270 2134.480 30.590 ;
        RECT 2134.280 2.400 2134.420 30.270 ;
        RECT 2134.210 0.000 2134.490 2.400 ;
      LAYER via2 ;
        RECT 1594.630 32.160 1594.910 32.440 ;
        RECT 1643.390 32.160 1643.670 32.440 ;
        RECT 1686.170 32.160 1686.450 32.440 ;
        RECT 1693.990 32.160 1694.270 32.440 ;
        RECT 1734.930 32.160 1735.210 32.440 ;
        RECT 1782.310 32.160 1782.590 32.440 ;
      LAYER met3 ;
        RECT 1594.605 32.450 1594.935 32.465 ;
        RECT 1643.365 32.450 1643.695 32.465 ;
        RECT 1594.605 32.150 1643.695 32.450 ;
        RECT 1594.605 32.135 1594.935 32.150 ;
        RECT 1643.365 32.135 1643.695 32.150 ;
        RECT 1686.145 32.450 1686.475 32.465 ;
        RECT 1693.965 32.450 1694.295 32.465 ;
        RECT 1686.145 32.150 1694.295 32.450 ;
        RECT 1686.145 32.135 1686.475 32.150 ;
        RECT 1693.965 32.135 1694.295 32.150 ;
        RECT 1734.905 32.450 1735.235 32.465 ;
        RECT 1782.285 32.450 1782.615 32.465 ;
        RECT 1734.905 32.150 1782.615 32.450 ;
        RECT 1734.905 32.135 1735.235 32.150 ;
        RECT 1782.285 32.135 1782.615 32.150 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1595.070 31.520 1595.390 31.580 ;
        RECT 1595.070 31.380 1609.560 31.520 ;
        RECT 1595.070 31.320 1595.390 31.380 ;
        RECT 1609.420 31.180 1609.560 31.380 ;
        RECT 2152.130 31.180 2152.450 31.240 ;
        RECT 1609.420 31.040 2152.450 31.180 ;
        RECT 2152.130 30.980 2152.450 31.040 ;
      LAYER via ;
        RECT 1595.100 31.320 1595.360 31.580 ;
        RECT 2152.160 30.980 2152.420 31.240 ;
      LAYER met2 ;
        RECT 1595.160 31.610 1595.300 54.000 ;
        RECT 1595.100 31.290 1595.360 31.610 ;
        RECT 2152.160 30.950 2152.420 31.270 ;
        RECT 2152.220 2.400 2152.360 30.950 ;
        RECT 2152.150 0.000 2152.430 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1610.785 34.765 1610.955 35.955 ;
      LAYER mcon ;
        RECT 1610.785 35.785 1610.955 35.955 ;
      LAYER met1 ;
        RECT 1601.510 35.940 1601.830 36.000 ;
        RECT 1610.725 35.940 1611.015 35.985 ;
        RECT 1601.510 35.800 1611.015 35.940 ;
        RECT 1601.510 35.740 1601.830 35.800 ;
        RECT 1610.725 35.755 1611.015 35.800 ;
        RECT 1610.725 34.920 1611.015 34.965 ;
        RECT 1658.550 34.920 1658.870 34.980 ;
        RECT 1610.725 34.780 1658.870 34.920 ;
        RECT 1610.725 34.735 1611.015 34.780 ;
        RECT 1658.550 34.720 1658.870 34.780 ;
        RECT 1852.210 30.840 1852.530 30.900 ;
        RECT 2170.070 30.840 2170.390 30.900 ;
        RECT 1852.210 30.700 2170.390 30.840 ;
        RECT 1852.210 30.640 1852.530 30.700 ;
        RECT 2170.070 30.640 2170.390 30.700 ;
      LAYER via ;
        RECT 1601.540 35.740 1601.800 36.000 ;
        RECT 1658.580 34.720 1658.840 34.980 ;
        RECT 1852.240 30.640 1852.500 30.900 ;
        RECT 2170.100 30.640 2170.360 30.900 ;
      LAYER met2 ;
        RECT 1601.600 36.030 1601.740 54.000 ;
        RECT 1601.540 35.710 1601.800 36.030 ;
        RECT 1658.580 34.690 1658.840 35.010 ;
        RECT 1658.640 30.445 1658.780 34.690 ;
        RECT 1852.240 30.610 1852.500 30.930 ;
        RECT 2170.100 30.610 2170.360 30.930 ;
        RECT 1852.300 30.445 1852.440 30.610 ;
        RECT 1658.570 30.075 1658.850 30.445 ;
        RECT 1852.230 30.075 1852.510 30.445 ;
        RECT 2170.160 2.400 2170.300 30.610 ;
        RECT 2170.090 0.000 2170.370 2.400 ;
      LAYER via2 ;
        RECT 1658.570 30.120 1658.850 30.400 ;
        RECT 1852.230 30.120 1852.510 30.400 ;
      LAYER met3 ;
        RECT 1658.545 30.410 1658.875 30.425 ;
        RECT 1852.205 30.410 1852.535 30.425 ;
        RECT 1658.545 30.110 1852.535 30.410 ;
        RECT 1658.545 30.095 1658.875 30.110 ;
        RECT 1852.205 30.095 1852.535 30.110 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1602.060 31.125 1602.200 54.000 ;
        RECT 1601.990 30.755 1602.270 31.125 ;
        RECT 2187.570 30.755 2187.850 31.125 ;
        RECT 2187.640 2.400 2187.780 30.755 ;
        RECT 2187.570 0.000 2187.850 2.400 ;
      LAYER via2 ;
        RECT 1601.990 30.800 1602.270 31.080 ;
        RECT 2187.570 30.800 2187.850 31.080 ;
      LAYER met3 ;
        RECT 1601.965 31.090 1602.295 31.105 ;
        RECT 2187.545 31.090 2187.875 31.105 ;
        RECT 1601.965 30.790 2187.875 31.090 ;
        RECT 1601.965 30.775 1602.295 30.790 ;
        RECT 2187.545 30.775 2187.875 30.790 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2203.740 3.130 2203.880 54.000 ;
        RECT 2203.740 2.990 2205.260 3.130 ;
        RECT 2205.120 2.960 2205.260 2.990 ;
        RECT 2205.120 2.820 2205.720 2.960 ;
        RECT 2205.580 2.400 2205.720 2.820 ;
        RECT 2205.510 0.000 2205.790 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2217.910 2.960 2218.230 3.020 ;
        RECT 2223.430 2.960 2223.750 3.020 ;
        RECT 2217.910 2.820 2223.750 2.960 ;
        RECT 2217.910 2.760 2218.230 2.820 ;
        RECT 2223.430 2.760 2223.750 2.820 ;
      LAYER via ;
        RECT 2217.940 2.760 2218.200 3.020 ;
        RECT 2223.460 2.760 2223.720 3.020 ;
      LAYER met2 ;
        RECT 2218.000 3.050 2218.140 54.000 ;
        RECT 2217.940 2.730 2218.200 3.050 ;
        RECT 2223.460 2.730 2223.720 3.050 ;
        RECT 2223.520 2.400 2223.660 2.730 ;
        RECT 2223.450 0.000 2223.730 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 778.110 2.960 778.430 3.020 ;
        RECT 781.790 2.960 782.110 3.020 ;
        RECT 778.110 2.820 782.110 2.960 ;
        RECT 778.110 2.760 778.430 2.820 ;
        RECT 781.790 2.760 782.110 2.820 ;
      LAYER via ;
        RECT 778.140 2.760 778.400 3.020 ;
        RECT 781.820 2.760 782.080 3.020 ;
      LAYER met2 ;
        RECT 781.880 3.050 782.020 54.000 ;
        RECT 778.140 2.730 778.400 3.050 ;
        RECT 781.820 2.730 782.080 3.050 ;
        RECT 778.200 2.400 778.340 2.730 ;
        RECT 778.130 0.000 778.410 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2238.150 2.960 2238.470 3.020 ;
        RECT 2241.370 2.960 2241.690 3.020 ;
        RECT 2238.150 2.820 2241.690 2.960 ;
        RECT 2238.150 2.760 2238.470 2.820 ;
        RECT 2241.370 2.760 2241.690 2.820 ;
      LAYER via ;
        RECT 2238.180 2.760 2238.440 3.020 ;
        RECT 2241.400 2.760 2241.660 3.020 ;
      LAYER met2 ;
        RECT 2238.240 3.050 2238.380 54.000 ;
        RECT 2238.180 2.730 2238.440 3.050 ;
        RECT 2241.400 2.730 2241.660 3.050 ;
        RECT 2241.460 2.400 2241.600 2.730 ;
        RECT 2241.390 0.000 2241.670 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2258.940 2.400 2259.080 54.000 ;
        RECT 2258.870 0.000 2259.150 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2272.650 2.960 2272.970 3.020 ;
        RECT 2276.790 2.960 2277.110 3.020 ;
        RECT 2272.650 2.820 2277.110 2.960 ;
        RECT 2272.650 2.760 2272.970 2.820 ;
        RECT 2276.790 2.760 2277.110 2.820 ;
      LAYER via ;
        RECT 2272.680 2.760 2272.940 3.020 ;
        RECT 2276.820 2.760 2277.080 3.020 ;
      LAYER met2 ;
        RECT 2272.740 3.050 2272.880 54.000 ;
        RECT 2272.680 2.730 2272.940 3.050 ;
        RECT 2276.820 2.730 2277.080 3.050 ;
        RECT 2276.880 2.400 2277.020 2.730 ;
        RECT 2276.810 0.000 2277.090 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2293.440 3.130 2293.580 54.000 ;
        RECT 2293.440 2.990 2294.500 3.130 ;
        RECT 2294.360 2.960 2294.500 2.990 ;
        RECT 2294.360 2.820 2294.960 2.960 ;
        RECT 2294.820 2.400 2294.960 2.820 ;
        RECT 2294.750 0.000 2295.030 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2307.150 2.960 2307.470 3.020 ;
        RECT 2312.670 2.960 2312.990 3.020 ;
        RECT 2307.150 2.820 2312.990 2.960 ;
        RECT 2307.150 2.760 2307.470 2.820 ;
        RECT 2312.670 2.760 2312.990 2.820 ;
      LAYER via ;
        RECT 2307.180 2.760 2307.440 3.020 ;
        RECT 2312.700 2.760 2312.960 3.020 ;
      LAYER met2 ;
        RECT 2307.240 3.050 2307.380 54.000 ;
        RECT 2307.180 2.730 2307.440 3.050 ;
        RECT 2312.700 2.730 2312.960 3.050 ;
        RECT 2312.760 2.400 2312.900 2.730 ;
        RECT 2312.690 0.000 2312.970 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2327.850 2.960 2328.170 3.020 ;
        RECT 2330.610 2.960 2330.930 3.020 ;
        RECT 2327.850 2.820 2330.930 2.960 ;
        RECT 2327.850 2.760 2328.170 2.820 ;
        RECT 2330.610 2.760 2330.930 2.820 ;
      LAYER via ;
        RECT 2327.880 2.760 2328.140 3.020 ;
        RECT 2330.640 2.760 2330.900 3.020 ;
      LAYER met2 ;
        RECT 2327.940 3.050 2328.080 54.000 ;
        RECT 2327.880 2.730 2328.140 3.050 ;
        RECT 2330.640 2.730 2330.900 3.050 ;
        RECT 2330.700 2.400 2330.840 2.730 ;
        RECT 2330.630 0.000 2330.910 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2286.985 34.085 2287.155 39.015 ;
      LAYER mcon ;
        RECT 2286.985 38.845 2287.155 39.015 ;
      LAYER met1 ;
        RECT 1636.470 39.000 1636.790 39.060 ;
        RECT 2286.925 39.000 2287.215 39.045 ;
        RECT 1636.470 38.860 2287.215 39.000 ;
        RECT 1636.470 38.800 1636.790 38.860 ;
        RECT 2286.925 38.815 2287.215 38.860 ;
        RECT 2286.925 34.240 2287.215 34.285 ;
        RECT 2348.090 34.240 2348.410 34.300 ;
        RECT 2286.925 34.100 2348.410 34.240 ;
        RECT 2286.925 34.055 2287.215 34.100 ;
        RECT 2348.090 34.040 2348.410 34.100 ;
      LAYER via ;
        RECT 1636.500 38.800 1636.760 39.060 ;
        RECT 2348.120 34.040 2348.380 34.300 ;
      LAYER met2 ;
        RECT 1636.560 39.090 1636.700 54.000 ;
        RECT 1636.500 38.770 1636.760 39.090 ;
        RECT 2348.120 34.010 2348.380 34.330 ;
        RECT 2348.180 2.400 2348.320 34.010 ;
        RECT 2348.110 0.000 2348.390 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2286.525 33.745 2286.695 38.675 ;
      LAYER mcon ;
        RECT 2286.525 38.505 2286.695 38.675 ;
      LAYER met1 ;
        RECT 1643.370 38.660 1643.690 38.720 ;
        RECT 2286.465 38.660 2286.755 38.705 ;
        RECT 1643.370 38.520 2286.755 38.660 ;
        RECT 1643.370 38.460 1643.690 38.520 ;
        RECT 2286.465 38.475 2286.755 38.520 ;
        RECT 2286.465 33.900 2286.755 33.945 ;
        RECT 2366.030 33.900 2366.350 33.960 ;
        RECT 2286.465 33.760 2366.350 33.900 ;
        RECT 2286.465 33.715 2286.755 33.760 ;
        RECT 2366.030 33.700 2366.350 33.760 ;
      LAYER via ;
        RECT 1643.400 38.460 1643.660 38.720 ;
        RECT 2366.060 33.700 2366.320 33.960 ;
      LAYER met2 ;
        RECT 1643.460 38.750 1643.600 54.000 ;
        RECT 1643.400 38.430 1643.660 38.750 ;
        RECT 2366.060 33.670 2366.320 33.990 ;
        RECT 2366.120 2.400 2366.260 33.670 ;
        RECT 2366.050 0.000 2366.330 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1642.910 34.580 1643.230 34.640 ;
        RECT 2383.970 34.580 2384.290 34.640 ;
        RECT 1642.910 34.440 2384.290 34.580 ;
        RECT 1642.910 34.380 1643.230 34.440 ;
        RECT 2383.970 34.380 2384.290 34.440 ;
      LAYER via ;
        RECT 1642.940 34.380 1643.200 34.640 ;
        RECT 2384.000 34.380 2384.260 34.640 ;
      LAYER met2 ;
        RECT 1643.000 34.670 1643.140 54.000 ;
        RECT 1642.940 34.350 1643.200 34.670 ;
        RECT 2384.000 34.350 2384.260 34.670 ;
        RECT 2384.060 2.400 2384.200 34.350 ;
        RECT 2383.990 0.000 2384.270 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1682.545 34.765 1682.715 39.355 ;
      LAYER mcon ;
        RECT 1682.545 39.185 1682.715 39.355 ;
      LAYER met1 ;
        RECT 1650.270 39.340 1650.590 39.400 ;
        RECT 1682.485 39.340 1682.775 39.385 ;
        RECT 1650.270 39.200 1682.775 39.340 ;
        RECT 1650.270 39.140 1650.590 39.200 ;
        RECT 1682.485 39.155 1682.775 39.200 ;
        RECT 1682.485 34.920 1682.775 34.965 ;
        RECT 2401.910 34.920 2402.230 34.980 ;
        RECT 1682.485 34.780 2402.230 34.920 ;
        RECT 1682.485 34.735 1682.775 34.780 ;
        RECT 2401.910 34.720 2402.230 34.780 ;
      LAYER via ;
        RECT 1650.300 39.140 1650.560 39.400 ;
        RECT 2401.940 34.720 2402.200 34.980 ;
      LAYER met2 ;
        RECT 1650.360 39.430 1650.500 54.000 ;
        RECT 1650.300 39.110 1650.560 39.430 ;
        RECT 2401.940 34.690 2402.200 35.010 ;
        RECT 2402.000 2.400 2402.140 34.690 ;
        RECT 2401.930 0.000 2402.210 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 796.050 18.260 796.370 18.320 ;
        RECT 802.490 18.260 802.810 18.320 ;
        RECT 796.050 18.120 802.810 18.260 ;
        RECT 796.050 18.060 796.370 18.120 ;
        RECT 802.490 18.060 802.810 18.120 ;
      LAYER via ;
        RECT 796.080 18.060 796.340 18.320 ;
        RECT 802.520 18.060 802.780 18.320 ;
      LAYER met2 ;
        RECT 802.580 18.350 802.720 54.000 ;
        RECT 796.080 18.030 796.340 18.350 ;
        RECT 802.520 18.030 802.780 18.350 ;
        RECT 796.140 2.400 796.280 18.030 ;
        RECT 796.070 0.000 796.350 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 641.490 17.580 641.810 17.640 ;
        RECT 643.790 17.580 644.110 17.640 ;
        RECT 641.490 17.440 644.110 17.580 ;
        RECT 641.490 17.380 641.810 17.440 ;
        RECT 643.790 17.380 644.110 17.440 ;
      LAYER via ;
        RECT 641.520 17.380 641.780 17.640 ;
        RECT 643.820 17.380 644.080 17.640 ;
      LAYER met2 ;
        RECT 643.880 17.670 644.020 54.000 ;
        RECT 641.520 17.350 641.780 17.670 ;
        RECT 643.820 17.350 644.080 17.670 ;
        RECT 641.580 2.400 641.720 17.350 ;
        RECT 641.510 0.000 641.790 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1650.730 35.940 1651.050 36.000 ;
        RECT 2369.250 35.940 2369.570 36.000 ;
        RECT 1650.730 35.800 2369.570 35.940 ;
        RECT 1650.730 35.740 1651.050 35.800 ;
        RECT 2369.250 35.740 2369.570 35.800 ;
        RECT 2371.090 35.940 2371.410 36.000 ;
        RECT 2425.370 35.940 2425.690 36.000 ;
        RECT 2371.090 35.800 2425.690 35.940 ;
        RECT 2371.090 35.740 2371.410 35.800 ;
        RECT 2425.370 35.740 2425.690 35.800 ;
      LAYER via ;
        RECT 1650.760 35.740 1651.020 36.000 ;
        RECT 2369.280 35.740 2369.540 36.000 ;
        RECT 2371.120 35.740 2371.380 36.000 ;
        RECT 2425.400 35.740 2425.660 36.000 ;
      LAYER met2 ;
        RECT 1650.820 36.030 1650.960 54.000 ;
        RECT 1650.760 35.710 1651.020 36.030 ;
        RECT 2369.280 35.885 2369.540 36.030 ;
        RECT 2371.120 35.885 2371.380 36.030 ;
        RECT 2369.270 35.515 2369.550 35.885 ;
        RECT 2371.110 35.515 2371.390 35.885 ;
        RECT 2425.400 35.710 2425.660 36.030 ;
        RECT 2425.460 2.400 2425.600 35.710 ;
        RECT 2425.390 0.000 2425.670 2.400 ;
      LAYER via2 ;
        RECT 2369.270 35.560 2369.550 35.840 ;
        RECT 2371.110 35.560 2371.390 35.840 ;
      LAYER met3 ;
        RECT 2369.245 35.850 2369.575 35.865 ;
        RECT 2371.085 35.850 2371.415 35.865 ;
        RECT 2369.245 35.550 2371.415 35.850 ;
        RECT 2369.245 35.535 2369.575 35.550 ;
        RECT 2371.085 35.535 2371.415 35.550 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2369.785 36.125 2370.875 36.295 ;
      LAYER mcon ;
        RECT 2370.705 36.125 2370.875 36.295 ;
      LAYER met1 ;
        RECT 1655.790 36.280 1656.110 36.340 ;
        RECT 2369.725 36.280 2370.015 36.325 ;
        RECT 1655.790 36.140 2370.015 36.280 ;
        RECT 1655.790 36.080 1656.110 36.140 ;
        RECT 2369.725 36.095 2370.015 36.140 ;
        RECT 2370.645 36.280 2370.935 36.325 ;
        RECT 2443.310 36.280 2443.630 36.340 ;
        RECT 2370.645 36.140 2443.630 36.280 ;
        RECT 2370.645 36.095 2370.935 36.140 ;
        RECT 2443.310 36.080 2443.630 36.140 ;
      LAYER via ;
        RECT 1655.820 36.080 1656.080 36.340 ;
        RECT 2443.340 36.080 2443.600 36.340 ;
      LAYER met2 ;
        RECT 1655.880 36.370 1656.020 54.000 ;
        RECT 1655.820 36.050 1656.080 36.370 ;
        RECT 2443.340 36.050 2443.600 36.370 ;
        RECT 2443.400 2.400 2443.540 36.050 ;
        RECT 2443.330 0.000 2443.610 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1657.170 36.620 1657.490 36.680 ;
        RECT 2461.250 36.620 2461.570 36.680 ;
        RECT 1657.170 36.480 2461.570 36.620 ;
        RECT 1657.170 36.420 1657.490 36.480 ;
        RECT 2461.250 36.420 2461.570 36.480 ;
      LAYER via ;
        RECT 1657.200 36.420 1657.460 36.680 ;
        RECT 2461.280 36.420 2461.540 36.680 ;
      LAYER met2 ;
        RECT 1657.260 53.990 1657.860 54.000 ;
        RECT 1657.260 36.710 1657.400 53.990 ;
        RECT 1657.200 36.390 1657.460 36.710 ;
        RECT 2461.280 36.390 2461.540 36.710 ;
        RECT 2461.340 2.400 2461.480 36.390 ;
        RECT 2461.270 0.000 2461.550 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1734.525 36.805 1735.155 36.975 ;
        RECT 2120.925 34.085 2121.095 36.975 ;
        RECT 2168.765 34.085 2168.935 36.975 ;
        RECT 2314.125 33.405 2314.295 36.975 ;
        RECT 2361.965 33.405 2362.135 36.975 ;
        RECT 2369.785 36.805 2370.875 36.975 ;
      LAYER mcon ;
        RECT 1734.985 36.805 1735.155 36.975 ;
        RECT 2120.925 36.805 2121.095 36.975 ;
        RECT 2168.765 36.805 2168.935 36.975 ;
        RECT 2314.125 36.805 2314.295 36.975 ;
        RECT 2361.965 36.805 2362.135 36.975 ;
        RECT 2370.705 36.805 2370.875 36.975 ;
      LAYER met1 ;
        RECT 1664.990 40.020 1665.310 40.080 ;
        RECT 1690.750 40.020 1691.070 40.080 ;
        RECT 1664.990 39.880 1691.070 40.020 ;
        RECT 1664.990 39.820 1665.310 39.880 ;
        RECT 1690.750 39.820 1691.070 39.880 ;
        RECT 1716.970 36.960 1717.290 37.020 ;
        RECT 1734.465 36.960 1734.755 37.005 ;
        RECT 1734.910 36.960 1735.230 37.020 ;
        RECT 1716.970 36.820 1735.230 36.960 ;
        RECT 1716.970 36.760 1717.290 36.820 ;
        RECT 1734.465 36.775 1734.755 36.820 ;
        RECT 1734.910 36.760 1735.230 36.820 ;
        RECT 1782.290 36.960 1782.610 37.020 ;
        RECT 2120.865 36.960 2121.155 37.005 ;
        RECT 1782.290 36.820 2121.155 36.960 ;
        RECT 1782.290 36.760 1782.610 36.820 ;
        RECT 2120.865 36.775 2121.155 36.820 ;
        RECT 2168.705 36.960 2168.995 37.005 ;
        RECT 2314.065 36.960 2314.355 37.005 ;
        RECT 2168.705 36.820 2314.355 36.960 ;
        RECT 2168.705 36.775 2168.995 36.820 ;
        RECT 2314.065 36.775 2314.355 36.820 ;
        RECT 2361.905 36.960 2362.195 37.005 ;
        RECT 2369.725 36.960 2370.015 37.005 ;
        RECT 2361.905 36.820 2370.015 36.960 ;
        RECT 2361.905 36.775 2362.195 36.820 ;
        RECT 2369.725 36.775 2370.015 36.820 ;
        RECT 2370.645 36.960 2370.935 37.005 ;
        RECT 2479.190 36.960 2479.510 37.020 ;
        RECT 2370.645 36.820 2479.510 36.960 ;
        RECT 2370.645 36.775 2370.935 36.820 ;
        RECT 2479.190 36.760 2479.510 36.820 ;
        RECT 2120.865 34.240 2121.155 34.285 ;
        RECT 2168.705 34.240 2168.995 34.285 ;
        RECT 2120.865 34.100 2168.995 34.240 ;
        RECT 2120.865 34.055 2121.155 34.100 ;
        RECT 2168.705 34.055 2168.995 34.100 ;
        RECT 2314.065 33.560 2314.355 33.605 ;
        RECT 2361.905 33.560 2362.195 33.605 ;
        RECT 2314.065 33.420 2362.195 33.560 ;
        RECT 2314.065 33.375 2314.355 33.420 ;
        RECT 2361.905 33.375 2362.195 33.420 ;
      LAYER via ;
        RECT 1665.020 39.820 1665.280 40.080 ;
        RECT 1690.780 39.820 1691.040 40.080 ;
        RECT 1717.000 36.760 1717.260 37.020 ;
        RECT 1734.940 36.760 1735.200 37.020 ;
        RECT 1782.320 36.760 1782.580 37.020 ;
        RECT 2479.220 36.760 2479.480 37.020 ;
      LAYER met2 ;
        RECT 1665.080 40.110 1665.220 54.000 ;
        RECT 1665.020 39.790 1665.280 40.110 ;
        RECT 1690.780 39.790 1691.040 40.110 ;
        RECT 1690.840 37.245 1690.980 39.790 ;
        RECT 1690.770 36.875 1691.050 37.245 ;
        RECT 1716.990 36.875 1717.270 37.245 ;
        RECT 1734.930 36.875 1735.210 37.245 ;
        RECT 1782.310 36.875 1782.590 37.245 ;
        RECT 1717.000 36.730 1717.260 36.875 ;
        RECT 1734.940 36.730 1735.200 36.875 ;
        RECT 1782.320 36.730 1782.580 36.875 ;
        RECT 2479.220 36.730 2479.480 37.050 ;
        RECT 2479.280 2.400 2479.420 36.730 ;
        RECT 2479.210 0.000 2479.490 2.400 ;
      LAYER via2 ;
        RECT 1690.770 36.920 1691.050 37.200 ;
        RECT 1716.990 36.920 1717.270 37.200 ;
        RECT 1734.930 36.920 1735.210 37.200 ;
        RECT 1782.310 36.920 1782.590 37.200 ;
      LAYER met3 ;
        RECT 1690.745 37.210 1691.075 37.225 ;
        RECT 1716.965 37.210 1717.295 37.225 ;
        RECT 1690.745 36.910 1717.295 37.210 ;
        RECT 1690.745 36.895 1691.075 36.910 ;
        RECT 1716.965 36.895 1717.295 36.910 ;
        RECT 1734.905 37.210 1735.235 37.225 ;
        RECT 1782.285 37.210 1782.615 37.225 ;
        RECT 1734.905 36.910 1782.615 37.210 ;
        RECT 1734.905 36.895 1735.235 36.910 ;
        RECT 1782.285 36.895 1782.615 36.910 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1698.185 37.655 1698.355 39.695 ;
        RECT 1698.185 37.485 1704.795 37.655 ;
        RECT 1789.725 37.145 1790.815 37.315 ;
      LAYER mcon ;
        RECT 1698.185 39.525 1698.355 39.695 ;
        RECT 1704.625 37.485 1704.795 37.655 ;
        RECT 1790.645 37.145 1790.815 37.315 ;
      LAYER met1 ;
        RECT 1671.430 39.680 1671.750 39.740 ;
        RECT 1698.125 39.680 1698.415 39.725 ;
        RECT 1671.430 39.540 1698.415 39.680 ;
        RECT 1671.430 39.480 1671.750 39.540 ;
        RECT 1698.125 39.495 1698.415 39.540 ;
        RECT 1704.565 37.640 1704.855 37.685 ;
        RECT 1704.565 37.500 1705.700 37.640 ;
        RECT 1704.565 37.455 1704.855 37.500 ;
        RECT 1705.560 37.300 1705.700 37.500 ;
        RECT 1789.665 37.300 1789.955 37.345 ;
        RECT 1705.560 37.160 1789.955 37.300 ;
        RECT 1789.665 37.115 1789.955 37.160 ;
        RECT 1790.585 37.300 1790.875 37.345 ;
        RECT 2497.130 37.300 2497.450 37.360 ;
        RECT 1790.585 37.160 2497.450 37.300 ;
        RECT 1790.585 37.115 1790.875 37.160 ;
        RECT 2497.130 37.100 2497.450 37.160 ;
      LAYER via ;
        RECT 1671.460 39.480 1671.720 39.740 ;
        RECT 2497.160 37.100 2497.420 37.360 ;
      LAYER met2 ;
        RECT 1671.520 39.770 1671.660 54.000 ;
        RECT 1671.460 39.450 1671.720 39.770 ;
        RECT 2497.160 37.070 2497.420 37.390 ;
        RECT 2497.220 2.400 2497.360 37.070 ;
        RECT 2497.150 0.000 2497.430 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1706.465 36.975 1706.635 37.655 ;
        RECT 2369.325 37.485 2370.415 37.655 ;
        RECT 1706.005 36.805 1706.635 36.975 ;
      LAYER mcon ;
        RECT 1706.465 37.485 1706.635 37.655 ;
        RECT 2370.245 37.485 2370.415 37.655 ;
      LAYER met1 ;
        RECT 1706.405 37.640 1706.695 37.685 ;
        RECT 2369.265 37.640 2369.555 37.685 ;
        RECT 1706.405 37.500 2369.555 37.640 ;
        RECT 1706.405 37.455 1706.695 37.500 ;
        RECT 2369.265 37.455 2369.555 37.500 ;
        RECT 2370.185 37.640 2370.475 37.685 ;
        RECT 2514.610 37.640 2514.930 37.700 ;
        RECT 2370.185 37.500 2514.930 37.640 ;
        RECT 2370.185 37.455 2370.475 37.500 ;
        RECT 2514.610 37.440 2514.930 37.500 ;
        RECT 1671.890 36.960 1672.210 37.020 ;
        RECT 1705.945 36.960 1706.235 37.005 ;
        RECT 1671.890 36.820 1706.235 36.960 ;
        RECT 1671.890 36.760 1672.210 36.820 ;
        RECT 1705.945 36.775 1706.235 36.820 ;
      LAYER via ;
        RECT 2514.640 37.440 2514.900 37.700 ;
        RECT 1671.920 36.760 1672.180 37.020 ;
      LAYER met2 ;
        RECT 1671.980 37.050 1672.120 54.000 ;
        RECT 2514.640 37.410 2514.900 37.730 ;
        RECT 1671.920 36.730 1672.180 37.050 ;
        RECT 2514.700 2.400 2514.840 37.410 ;
        RECT 2514.630 0.000 2514.910 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1706.390 41.380 1706.710 41.440 ;
        RECT 2532.550 41.380 2532.870 41.440 ;
        RECT 1706.390 41.240 2532.870 41.380 ;
        RECT 1706.390 41.180 1706.710 41.240 ;
        RECT 2532.550 41.180 2532.870 41.240 ;
        RECT 1678.330 37.640 1678.650 37.700 ;
        RECT 1704.090 37.640 1704.410 37.700 ;
        RECT 1678.330 37.500 1704.410 37.640 ;
        RECT 1678.330 37.440 1678.650 37.500 ;
        RECT 1704.090 37.440 1704.410 37.500 ;
      LAYER via ;
        RECT 1706.420 41.180 1706.680 41.440 ;
        RECT 2532.580 41.180 2532.840 41.440 ;
        RECT 1678.360 37.440 1678.620 37.700 ;
        RECT 1704.120 37.440 1704.380 37.700 ;
      LAYER met2 ;
        RECT 1678.420 37.730 1678.560 54.000 ;
        RECT 1706.420 41.325 1706.680 41.470 ;
        RECT 1704.110 40.955 1704.390 41.325 ;
        RECT 1706.410 40.955 1706.690 41.325 ;
        RECT 2532.580 41.150 2532.840 41.470 ;
        RECT 1704.180 37.730 1704.320 40.955 ;
        RECT 1678.360 37.410 1678.620 37.730 ;
        RECT 1704.120 37.410 1704.380 37.730 ;
        RECT 2532.640 2.400 2532.780 41.150 ;
        RECT 2532.570 0.000 2532.850 2.400 ;
      LAYER via2 ;
        RECT 1704.110 41.000 1704.390 41.280 ;
        RECT 1706.410 41.000 1706.690 41.280 ;
      LAYER met3 ;
        RECT 1704.085 41.290 1704.415 41.305 ;
        RECT 1706.385 41.290 1706.715 41.305 ;
        RECT 1704.085 40.990 1706.715 41.290 ;
        RECT 1704.085 40.975 1704.415 40.990 ;
        RECT 1706.385 40.975 1706.715 40.990 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1706.850 40.360 1707.170 40.420 ;
        RECT 2550.490 40.360 2550.810 40.420 ;
        RECT 1706.850 40.220 2550.810 40.360 ;
        RECT 1706.850 40.160 1707.170 40.220 ;
        RECT 2550.490 40.160 2550.810 40.220 ;
        RECT 1677.870 37.300 1678.190 37.360 ;
        RECT 1703.630 37.300 1703.950 37.360 ;
        RECT 1677.870 37.160 1703.950 37.300 ;
        RECT 1677.870 37.100 1678.190 37.160 ;
        RECT 1703.630 37.100 1703.950 37.160 ;
      LAYER via ;
        RECT 1706.880 40.160 1707.140 40.420 ;
        RECT 2550.520 40.160 2550.780 40.420 ;
        RECT 1677.900 37.100 1678.160 37.360 ;
        RECT 1703.660 37.100 1703.920 37.360 ;
      LAYER met2 ;
        RECT 1677.960 37.390 1678.100 54.000 ;
        RECT 1703.650 40.275 1703.930 40.645 ;
        RECT 1706.870 40.275 1707.150 40.645 ;
        RECT 1703.720 37.390 1703.860 40.275 ;
        RECT 1706.880 40.130 1707.140 40.275 ;
        RECT 2550.520 40.130 2550.780 40.450 ;
        RECT 1677.900 37.070 1678.160 37.390 ;
        RECT 1703.660 37.070 1703.920 37.390 ;
        RECT 2550.580 2.400 2550.720 40.130 ;
        RECT 2550.510 0.000 2550.790 2.400 ;
      LAYER via2 ;
        RECT 1703.650 40.320 1703.930 40.600 ;
        RECT 1706.870 40.320 1707.150 40.600 ;
      LAYER met3 ;
        RECT 1703.625 40.610 1703.955 40.625 ;
        RECT 1706.845 40.610 1707.175 40.625 ;
        RECT 1703.625 40.310 1707.175 40.610 ;
        RECT 1703.625 40.295 1703.955 40.310 ;
        RECT 1706.845 40.295 1707.175 40.310 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1706.465 40.205 1706.635 45.815 ;
        RECT 1753.385 39.355 1753.555 45.815 ;
        RECT 1754.305 39.865 1754.935 40.035 ;
        RECT 1754.305 39.355 1754.475 39.865 ;
        RECT 1753.385 39.185 1754.475 39.355 ;
      LAYER mcon ;
        RECT 1706.465 45.645 1706.635 45.815 ;
        RECT 1753.385 45.645 1753.555 45.815 ;
        RECT 1754.765 39.865 1754.935 40.035 ;
      LAYER met1 ;
        RECT 1706.405 45.800 1706.695 45.845 ;
        RECT 1753.325 45.800 1753.615 45.845 ;
        RECT 1706.405 45.660 1753.615 45.800 ;
        RECT 1706.405 45.615 1706.695 45.660 ;
        RECT 1753.325 45.615 1753.615 45.660 ;
        RECT 1684.770 40.360 1685.090 40.420 ;
        RECT 1706.405 40.360 1706.695 40.405 ;
        RECT 1684.770 40.220 1706.695 40.360 ;
        RECT 1684.770 40.160 1685.090 40.220 ;
        RECT 1706.405 40.175 1706.695 40.220 ;
        RECT 1754.705 40.020 1754.995 40.065 ;
        RECT 2568.430 40.020 2568.750 40.080 ;
        RECT 1754.705 39.880 2568.750 40.020 ;
        RECT 1754.705 39.835 1754.995 39.880 ;
        RECT 2568.430 39.820 2568.750 39.880 ;
      LAYER via ;
        RECT 1684.800 40.160 1685.060 40.420 ;
        RECT 2568.460 39.820 2568.720 40.080 ;
      LAYER met2 ;
        RECT 1684.860 40.450 1685.000 54.000 ;
        RECT 1684.800 40.130 1685.060 40.450 ;
        RECT 2568.460 39.790 2568.720 40.110 ;
        RECT 2568.520 2.400 2568.660 39.790 ;
        RECT 2568.450 0.000 2568.730 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1706.005 41.225 1706.175 45.475 ;
        RECT 1753.845 39.525 1754.015 45.475 ;
      LAYER mcon ;
        RECT 1706.005 45.305 1706.175 45.475 ;
        RECT 1753.845 45.305 1754.015 45.475 ;
      LAYER met1 ;
        RECT 1705.945 45.460 1706.235 45.505 ;
        RECT 1753.785 45.460 1754.075 45.505 ;
        RECT 1705.945 45.320 1754.075 45.460 ;
        RECT 1705.945 45.275 1706.235 45.320 ;
        RECT 1753.785 45.275 1754.075 45.320 ;
        RECT 1685.230 41.380 1685.550 41.440 ;
        RECT 1705.945 41.380 1706.235 41.425 ;
        RECT 1685.230 41.240 1706.235 41.380 ;
        RECT 1685.230 41.180 1685.550 41.240 ;
        RECT 1705.945 41.195 1706.235 41.240 ;
        RECT 1753.785 39.680 1754.075 39.725 ;
        RECT 2586.370 39.680 2586.690 39.740 ;
        RECT 1753.785 39.540 2586.690 39.680 ;
        RECT 1753.785 39.495 1754.075 39.540 ;
        RECT 2586.370 39.480 2586.690 39.540 ;
      LAYER via ;
        RECT 1685.260 41.180 1685.520 41.440 ;
        RECT 2586.400 39.480 2586.660 39.740 ;
      LAYER met2 ;
        RECT 1685.320 41.470 1685.460 54.000 ;
        RECT 1685.260 41.150 1685.520 41.470 ;
        RECT 2586.400 39.450 2586.660 39.770 ;
        RECT 2586.460 2.400 2586.600 39.450 ;
        RECT 2586.390 0.000 2586.670 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 819.970 32.200 820.290 32.260 ;
        RECT 1315.850 32.200 1316.170 32.260 ;
        RECT 819.970 32.060 1316.170 32.200 ;
        RECT 819.970 32.000 820.290 32.060 ;
        RECT 1315.850 32.000 1316.170 32.060 ;
      LAYER via ;
        RECT 820.000 32.000 820.260 32.260 ;
        RECT 1315.880 32.000 1316.140 32.260 ;
      LAYER met2 ;
        RECT 1315.940 32.290 1316.080 54.000 ;
        RECT 820.000 31.970 820.260 32.290 ;
        RECT 1315.880 31.970 1316.140 32.290 ;
        RECT 820.060 2.400 820.200 31.970 ;
        RECT 819.990 0.000 820.270 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1691.210 39.340 1691.530 39.400 ;
        RECT 2604.310 39.340 2604.630 39.400 ;
        RECT 1691.210 39.200 2604.630 39.340 ;
        RECT 1691.210 39.140 1691.530 39.200 ;
        RECT 2604.310 39.140 2604.630 39.200 ;
      LAYER via ;
        RECT 1691.240 39.140 1691.500 39.400 ;
        RECT 2604.340 39.140 2604.600 39.400 ;
      LAYER met2 ;
        RECT 1691.300 39.430 1691.440 54.000 ;
        RECT 1691.240 39.110 1691.500 39.430 ;
        RECT 2604.340 39.110 2604.600 39.430 ;
        RECT 2604.400 7.210 2604.540 39.110 ;
        RECT 2603.940 7.070 2604.540 7.210 ;
        RECT 2603.940 2.400 2604.080 7.070 ;
        RECT 2603.870 0.000 2604.150 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2287.905 38.845 2288.075 41.735 ;
      LAYER mcon ;
        RECT 2287.905 41.565 2288.075 41.735 ;
      LAYER met1 ;
        RECT 1806.210 41.720 1806.530 41.780 ;
        RECT 2287.845 41.720 2288.135 41.765 ;
        RECT 1806.210 41.580 2288.135 41.720 ;
        RECT 1806.210 41.520 1806.530 41.580 ;
        RECT 2287.845 41.535 2288.135 41.580 ;
        RECT 1691.670 40.020 1691.990 40.080 ;
        RECT 1754.230 40.020 1754.550 40.080 ;
        RECT 1691.670 39.880 1754.550 40.020 ;
        RECT 1691.670 39.820 1691.990 39.880 ;
        RECT 1754.230 39.820 1754.550 39.880 ;
        RECT 2287.845 39.000 2288.135 39.045 ;
        RECT 2621.790 39.000 2622.110 39.060 ;
        RECT 2287.845 38.860 2622.110 39.000 ;
        RECT 2287.845 38.815 2288.135 38.860 ;
        RECT 2621.790 38.800 2622.110 38.860 ;
      LAYER via ;
        RECT 1806.240 41.520 1806.500 41.780 ;
        RECT 1691.700 39.820 1691.960 40.080 ;
        RECT 1754.260 39.820 1754.520 40.080 ;
        RECT 2621.820 38.800 2622.080 39.060 ;
      LAYER met2 ;
        RECT 1691.760 40.110 1691.900 54.000 ;
        RECT 1806.240 41.490 1806.500 41.810 ;
        RECT 1691.700 39.790 1691.960 40.110 ;
        RECT 1754.260 39.790 1754.520 40.110 ;
        RECT 1754.320 39.285 1754.460 39.790 ;
        RECT 1806.300 39.285 1806.440 41.490 ;
        RECT 1754.250 38.915 1754.530 39.285 ;
        RECT 1806.230 38.915 1806.510 39.285 ;
        RECT 2621.820 38.770 2622.080 39.090 ;
        RECT 2621.880 2.400 2622.020 38.770 ;
        RECT 2621.810 0.000 2622.090 2.400 ;
      LAYER via2 ;
        RECT 1754.250 38.960 1754.530 39.240 ;
        RECT 1806.230 38.960 1806.510 39.240 ;
      LAYER met3 ;
        RECT 1754.225 39.250 1754.555 39.265 ;
        RECT 1806.205 39.250 1806.535 39.265 ;
        RECT 1754.225 38.950 1806.535 39.250 ;
        RECT 1754.225 38.935 1754.555 38.950 ;
        RECT 1806.205 38.935 1806.535 38.950 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2287.445 38.505 2287.615 42.075 ;
      LAYER mcon ;
        RECT 2287.445 41.905 2287.615 42.075 ;
      LAYER met1 ;
        RECT 1780.910 42.060 1781.230 42.120 ;
        RECT 1851.750 42.060 1852.070 42.120 ;
        RECT 1780.910 41.920 1852.070 42.060 ;
        RECT 1780.910 41.860 1781.230 41.920 ;
        RECT 1851.750 41.860 1852.070 41.920 ;
        RECT 1997.110 42.060 1997.430 42.120 ;
        RECT 2045.870 42.060 2046.190 42.120 ;
        RECT 1997.110 41.920 2046.190 42.060 ;
        RECT 1997.110 41.860 1997.430 41.920 ;
        RECT 2045.870 41.860 2046.190 41.920 ;
        RECT 2191.230 42.060 2191.550 42.120 ;
        RECT 2287.385 42.060 2287.675 42.105 ;
        RECT 2191.230 41.920 2287.675 42.060 ;
        RECT 2191.230 41.860 2191.550 41.920 ;
        RECT 2287.385 41.875 2287.675 41.920 ;
        RECT 1698.570 39.680 1698.890 39.740 ;
        RECT 1753.310 39.680 1753.630 39.740 ;
        RECT 1698.570 39.540 1753.630 39.680 ;
        RECT 1698.570 39.480 1698.890 39.540 ;
        RECT 1753.310 39.480 1753.630 39.540 ;
        RECT 2287.385 38.660 2287.675 38.705 ;
        RECT 2639.730 38.660 2640.050 38.720 ;
        RECT 2287.385 38.520 2640.050 38.660 ;
        RECT 2287.385 38.475 2287.675 38.520 ;
        RECT 2639.730 38.460 2640.050 38.520 ;
      LAYER via ;
        RECT 1780.940 41.860 1781.200 42.120 ;
        RECT 1851.780 41.860 1852.040 42.120 ;
        RECT 1997.140 41.860 1997.400 42.120 ;
        RECT 2045.900 41.860 2046.160 42.120 ;
        RECT 2191.260 41.860 2191.520 42.120 ;
        RECT 1698.600 39.480 1698.860 39.740 ;
        RECT 1753.340 39.480 1753.600 39.740 ;
        RECT 2639.760 38.460 2640.020 38.720 ;
      LAYER met2 ;
        RECT 1698.660 39.770 1698.800 54.000 ;
        RECT 1780.940 41.830 1781.200 42.150 ;
        RECT 1851.780 41.830 1852.040 42.150 ;
        RECT 1997.140 41.830 1997.400 42.150 ;
        RECT 2045.900 41.830 2046.160 42.150 ;
        RECT 2191.260 41.830 2191.520 42.150 ;
        RECT 1698.600 39.450 1698.860 39.770 ;
        RECT 1753.340 39.450 1753.600 39.770 ;
        RECT 1753.400 38.605 1753.540 39.450 ;
        RECT 1781.000 38.605 1781.140 41.830 ;
        RECT 1851.840 38.605 1851.980 41.830 ;
        RECT 1997.200 38.605 1997.340 41.830 ;
        RECT 2045.960 38.605 2046.100 41.830 ;
        RECT 2191.320 38.605 2191.460 41.830 ;
        RECT 1753.330 38.235 1753.610 38.605 ;
        RECT 1780.930 38.235 1781.210 38.605 ;
        RECT 1851.770 38.235 1852.050 38.605 ;
        RECT 1997.130 38.235 1997.410 38.605 ;
        RECT 2045.890 38.235 2046.170 38.605 ;
        RECT 2191.250 38.235 2191.530 38.605 ;
        RECT 2639.760 38.430 2640.020 38.750 ;
        RECT 2639.820 2.400 2639.960 38.430 ;
        RECT 2639.750 0.000 2640.030 2.400 ;
      LAYER via2 ;
        RECT 1753.330 38.280 1753.610 38.560 ;
        RECT 1780.930 38.280 1781.210 38.560 ;
        RECT 1851.770 38.280 1852.050 38.560 ;
        RECT 1997.130 38.280 1997.410 38.560 ;
        RECT 2045.890 38.280 2046.170 38.560 ;
        RECT 2191.250 38.280 2191.530 38.560 ;
      LAYER met3 ;
        RECT 1753.305 38.570 1753.635 38.585 ;
        RECT 1780.905 38.570 1781.235 38.585 ;
        RECT 1753.305 38.270 1781.235 38.570 ;
        RECT 1753.305 38.255 1753.635 38.270 ;
        RECT 1780.905 38.255 1781.235 38.270 ;
        RECT 1851.745 38.570 1852.075 38.585 ;
        RECT 1997.105 38.570 1997.435 38.585 ;
        RECT 1851.745 38.270 1997.435 38.570 ;
        RECT 1851.745 38.255 1852.075 38.270 ;
        RECT 1997.105 38.255 1997.435 38.270 ;
        RECT 2045.865 38.570 2046.195 38.585 ;
        RECT 2191.225 38.570 2191.555 38.585 ;
        RECT 2045.865 38.270 2191.555 38.570 ;
        RECT 2045.865 38.255 2046.195 38.270 ;
        RECT 2191.225 38.255 2191.555 38.270 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2657.760 2.400 2657.900 54.000 ;
        RECT 2657.690 0.000 2657.970 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2675.240 2.400 2675.380 54.000 ;
        RECT 2675.170 0.000 2675.450 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2686.650 37.640 2686.970 37.700 ;
        RECT 2693.090 37.640 2693.410 37.700 ;
        RECT 2686.650 37.500 2693.410 37.640 ;
        RECT 2686.650 37.440 2686.970 37.500 ;
        RECT 2693.090 37.440 2693.410 37.500 ;
      LAYER via ;
        RECT 2686.680 37.440 2686.940 37.700 ;
        RECT 2693.120 37.440 2693.380 37.700 ;
      LAYER met2 ;
        RECT 2686.740 37.730 2686.880 54.000 ;
        RECT 2686.680 37.410 2686.940 37.730 ;
        RECT 2693.120 37.410 2693.380 37.730 ;
        RECT 2693.180 2.400 2693.320 37.410 ;
        RECT 2693.110 0.000 2693.390 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2707.425 48.365 2707.595 54.000 ;
      LAYER met1 ;
        RECT 2707.365 48.520 2707.655 48.565 ;
        RECT 2711.030 48.520 2711.350 48.580 ;
        RECT 2707.365 48.380 2711.350 48.520 ;
        RECT 2707.365 48.335 2707.655 48.380 ;
        RECT 2711.030 48.320 2711.350 48.380 ;
      LAYER via ;
        RECT 2711.060 48.320 2711.320 48.580 ;
      LAYER met2 ;
        RECT 2711.060 48.290 2711.320 48.610 ;
        RECT 2711.120 2.400 2711.260 48.290 ;
        RECT 2711.050 0.000 2711.330 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2727.590 48.520 2727.910 48.580 ;
        RECT 2728.970 48.520 2729.290 48.580 ;
        RECT 2727.590 48.380 2729.290 48.520 ;
        RECT 2727.590 48.320 2727.910 48.380 ;
        RECT 2728.970 48.320 2729.290 48.380 ;
      LAYER via ;
        RECT 2727.620 48.320 2727.880 48.580 ;
        RECT 2729.000 48.320 2729.260 48.580 ;
      LAYER met2 ;
        RECT 2727.680 48.610 2727.820 54.000 ;
        RECT 2727.620 48.290 2727.880 48.610 ;
        RECT 2729.000 48.290 2729.260 48.610 ;
        RECT 2729.060 2.400 2729.200 48.290 ;
        RECT 2728.990 0.000 2729.270 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2747.000 2.400 2747.140 54.000 ;
        RECT 2746.930 0.000 2747.210 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2762.625 48.365 2762.795 54.000 ;
      LAYER met1 ;
        RECT 2762.565 48.520 2762.855 48.565 ;
        RECT 2764.390 48.520 2764.710 48.580 ;
        RECT 2762.565 48.380 2764.710 48.520 ;
        RECT 2762.565 48.335 2762.855 48.380 ;
        RECT 2764.390 48.320 2764.710 48.380 ;
      LAYER via ;
        RECT 2764.420 48.320 2764.680 48.580 ;
      LAYER met2 ;
        RECT 2764.420 48.290 2764.680 48.610 ;
        RECT 2764.480 2.400 2764.620 48.290 ;
        RECT 2764.410 0.000 2764.690 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 837.910 33.220 838.230 33.280 ;
        RECT 1322.750 33.220 1323.070 33.280 ;
        RECT 837.910 33.080 1323.070 33.220 ;
        RECT 837.910 33.020 838.230 33.080 ;
        RECT 1322.750 33.020 1323.070 33.080 ;
      LAYER via ;
        RECT 837.940 33.020 838.200 33.280 ;
        RECT 1322.780 33.020 1323.040 33.280 ;
      LAYER met2 ;
        RECT 1322.840 33.310 1322.980 54.000 ;
        RECT 837.940 32.990 838.200 33.310 ;
        RECT 1322.780 32.990 1323.040 33.310 ;
        RECT 838.000 2.400 838.140 32.990 ;
        RECT 837.930 0.000 838.210 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2776.350 37.640 2776.670 37.700 ;
        RECT 2782.330 37.640 2782.650 37.700 ;
        RECT 2776.350 37.500 2782.650 37.640 ;
        RECT 2776.350 37.440 2776.670 37.500 ;
        RECT 2782.330 37.440 2782.650 37.500 ;
      LAYER via ;
        RECT 2776.380 37.440 2776.640 37.700 ;
        RECT 2782.360 37.440 2782.620 37.700 ;
      LAYER met2 ;
        RECT 2776.440 37.730 2776.580 54.000 ;
        RECT 2776.380 37.410 2776.640 37.730 ;
        RECT 2782.360 37.410 2782.620 37.730 ;
        RECT 2782.420 2.400 2782.560 37.410 ;
        RECT 2782.350 0.000 2782.630 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1755.610 47.160 1755.930 47.220 ;
        RECT 2800.270 47.160 2800.590 47.220 ;
        RECT 1755.610 47.020 2800.590 47.160 ;
        RECT 1755.610 46.960 1755.930 47.020 ;
        RECT 2800.270 46.960 2800.590 47.020 ;
        RECT 1733.070 46.820 1733.390 46.880 ;
        RECT 1746.410 46.820 1746.730 46.880 ;
        RECT 1733.070 46.680 1746.730 46.820 ;
        RECT 1733.070 46.620 1733.390 46.680 ;
        RECT 1746.410 46.620 1746.730 46.680 ;
      LAYER via ;
        RECT 1755.640 46.960 1755.900 47.220 ;
        RECT 2800.300 46.960 2800.560 47.220 ;
        RECT 1733.100 46.620 1733.360 46.880 ;
        RECT 1746.440 46.620 1746.700 46.880 ;
      LAYER met2 ;
        RECT 1733.160 46.910 1733.300 54.000 ;
        RECT 1755.640 46.930 1755.900 47.250 ;
        RECT 2800.300 46.930 2800.560 47.250 ;
        RECT 1733.100 46.590 1733.360 46.910 ;
        RECT 1746.440 46.590 1746.700 46.910 ;
        RECT 1746.500 46.085 1746.640 46.590 ;
        RECT 1755.700 46.085 1755.840 46.930 ;
        RECT 1746.430 45.715 1746.710 46.085 ;
        RECT 1755.630 45.715 1755.910 46.085 ;
        RECT 2800.360 2.400 2800.500 46.930 ;
        RECT 2800.290 0.000 2800.570 2.400 ;
      LAYER via2 ;
        RECT 1746.430 45.760 1746.710 46.040 ;
        RECT 1755.630 45.760 1755.910 46.040 ;
      LAYER met3 ;
        RECT 1746.405 46.050 1746.735 46.065 ;
        RECT 1755.605 46.050 1755.935 46.065 ;
        RECT 1746.405 45.750 1755.935 46.050 ;
        RECT 1746.405 45.735 1746.735 45.750 ;
        RECT 1755.605 45.735 1755.935 45.750 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1756.605 44.965 1756.775 54.000 ;
        RECT 1780.065 45.135 1780.235 46.835 ;
        RECT 1778.685 44.965 1780.235 45.135 ;
      LAYER mcon ;
        RECT 1780.065 46.665 1780.235 46.835 ;
      LAYER met1 ;
        RECT 1780.005 46.820 1780.295 46.865 ;
        RECT 2818.210 46.820 2818.530 46.880 ;
        RECT 1780.005 46.680 2818.530 46.820 ;
        RECT 1780.005 46.635 1780.295 46.680 ;
        RECT 2818.210 46.620 2818.530 46.680 ;
        RECT 1756.545 45.120 1756.835 45.165 ;
        RECT 1778.625 45.120 1778.915 45.165 ;
        RECT 1756.545 44.980 1778.915 45.120 ;
        RECT 1756.545 44.935 1756.835 44.980 ;
        RECT 1778.625 44.935 1778.915 44.980 ;
      LAYER via ;
        RECT 2818.240 46.620 2818.500 46.880 ;
      LAYER met2 ;
        RECT 2818.240 46.590 2818.500 46.910 ;
        RECT 2818.300 2.400 2818.440 46.590 ;
        RECT 2818.230 0.000 2818.510 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1755.225 47.005 1755.855 47.175 ;
        RECT 1755.685 45.645 1755.855 47.005 ;
      LAYER met1 ;
        RECT 1754.230 47.160 1754.550 47.220 ;
        RECT 1755.165 47.160 1755.455 47.205 ;
        RECT 1754.230 47.020 1755.455 47.160 ;
        RECT 1754.230 46.960 1754.550 47.020 ;
        RECT 1755.165 46.975 1755.455 47.020 ;
        RECT 1755.625 45.800 1755.915 45.845 ;
        RECT 2836.150 45.800 2836.470 45.860 ;
        RECT 1755.625 45.660 2836.470 45.800 ;
        RECT 1755.625 45.615 1755.915 45.660 ;
        RECT 2836.150 45.600 2836.470 45.660 ;
      LAYER via ;
        RECT 1754.260 46.960 1754.520 47.220 ;
        RECT 2836.180 45.600 2836.440 45.860 ;
      LAYER met2 ;
        RECT 1740.060 47.445 1740.200 54.000 ;
        RECT 1739.990 47.075 1740.270 47.445 ;
        RECT 1754.250 47.075 1754.530 47.445 ;
        RECT 1754.260 46.930 1754.520 47.075 ;
        RECT 2836.180 45.570 2836.440 45.890 ;
        RECT 2836.240 2.400 2836.380 45.570 ;
        RECT 2836.170 0.000 2836.450 2.400 ;
      LAYER via2 ;
        RECT 1739.990 47.120 1740.270 47.400 ;
        RECT 1754.250 47.120 1754.530 47.400 ;
      LAYER met3 ;
        RECT 1739.965 47.410 1740.295 47.425 ;
        RECT 1754.225 47.410 1754.555 47.425 ;
        RECT 1739.965 47.110 1754.555 47.410 ;
        RECT 1739.965 47.095 1740.295 47.110 ;
        RECT 1754.225 47.095 1754.555 47.110 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1754.765 46.665 1754.935 54.000 ;
        RECT 1779.605 45.305 1779.775 46.835 ;
      LAYER mcon ;
        RECT 1779.605 46.665 1779.775 46.835 ;
      LAYER met1 ;
        RECT 1754.705 46.820 1754.995 46.865 ;
        RECT 1779.545 46.820 1779.835 46.865 ;
        RECT 1754.705 46.680 1779.835 46.820 ;
        RECT 1754.705 46.635 1754.995 46.680 ;
        RECT 1779.545 46.635 1779.835 46.680 ;
        RECT 1779.545 45.460 1779.835 45.505 ;
        RECT 2853.630 45.460 2853.950 45.520 ;
        RECT 1779.545 45.320 2853.950 45.460 ;
        RECT 1779.545 45.275 1779.835 45.320 ;
        RECT 2853.630 45.260 2853.950 45.320 ;
      LAYER via ;
        RECT 2853.660 45.260 2853.920 45.520 ;
      LAYER met2 ;
        RECT 2853.660 45.230 2853.920 45.550 ;
        RECT 2853.720 2.400 2853.860 45.230 ;
        RECT 2853.650 0.000 2853.930 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1753.385 47.345 1754.475 47.515 ;
        RECT 1753.385 46.665 1753.555 47.345 ;
        RECT 1754.305 46.495 1754.475 47.345 ;
        RECT 1754.305 46.325 1754.935 46.495 ;
        RECT 1754.765 45.305 1754.935 46.325 ;
      LAYER met1 ;
        RECT 1747.330 46.820 1747.650 46.880 ;
        RECT 1753.325 46.820 1753.615 46.865 ;
        RECT 1747.330 46.680 1753.615 46.820 ;
        RECT 1747.330 46.620 1747.650 46.680 ;
        RECT 1753.325 46.635 1753.615 46.680 ;
        RECT 1754.705 45.460 1754.995 45.505 ;
        RECT 1754.705 45.320 1779.300 45.460 ;
        RECT 1754.705 45.275 1754.995 45.320 ;
        RECT 1779.160 45.120 1779.300 45.320 ;
        RECT 2871.570 45.120 2871.890 45.180 ;
        RECT 1779.160 44.980 2871.890 45.120 ;
        RECT 2871.570 44.920 2871.890 44.980 ;
      LAYER via ;
        RECT 1747.360 46.620 1747.620 46.880 ;
        RECT 2871.600 44.920 2871.860 45.180 ;
      LAYER met2 ;
        RECT 1747.420 46.910 1747.560 54.000 ;
        RECT 1747.360 46.590 1747.620 46.910 ;
        RECT 2871.600 44.890 2871.860 45.210 ;
        RECT 2871.660 2.400 2871.800 44.890 ;
        RECT 2871.590 0.000 2871.870 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1753.845 45.815 1754.015 47.175 ;
        RECT 1753.845 45.645 1754.475 45.815 ;
        RECT 1755.225 44.795 1755.395 45.815 ;
        RECT 1755.225 44.625 1755.855 44.795 ;
      LAYER mcon ;
        RECT 1753.845 47.005 1754.015 47.175 ;
        RECT 1754.305 45.645 1754.475 45.815 ;
        RECT 1755.225 45.645 1755.395 45.815 ;
        RECT 1755.685 44.625 1755.855 44.795 ;
      LAYER met1 ;
        RECT 1746.870 47.160 1747.190 47.220 ;
        RECT 1753.785 47.160 1754.075 47.205 ;
        RECT 1746.870 47.020 1754.075 47.160 ;
        RECT 1746.870 46.960 1747.190 47.020 ;
        RECT 1753.785 46.975 1754.075 47.020 ;
        RECT 1754.245 45.800 1754.535 45.845 ;
        RECT 1755.165 45.800 1755.455 45.845 ;
        RECT 1754.245 45.660 1755.455 45.800 ;
        RECT 1754.245 45.615 1754.535 45.660 ;
        RECT 1755.165 45.615 1755.455 45.660 ;
        RECT 1755.625 44.780 1755.915 44.825 ;
        RECT 2889.510 44.780 2889.830 44.840 ;
        RECT 1755.625 44.640 2889.830 44.780 ;
        RECT 1755.625 44.595 1755.915 44.640 ;
        RECT 2889.510 44.580 2889.830 44.640 ;
      LAYER via ;
        RECT 1746.900 46.960 1747.160 47.220 ;
        RECT 2889.540 44.580 2889.800 44.840 ;
      LAYER met2 ;
        RECT 1746.960 47.250 1747.100 54.000 ;
        RECT 1746.900 46.930 1747.160 47.250 ;
        RECT 2889.540 44.550 2889.800 44.870 ;
        RECT 2889.600 2.400 2889.740 44.550 ;
        RECT 2889.530 0.000 2889.810 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1754.780 44.725 1754.920 54.000 ;
        RECT 1754.710 44.355 1754.990 44.725 ;
        RECT 2907.930 44.355 2908.210 44.725 ;
        RECT 2908.000 7.210 2908.140 44.355 ;
        RECT 2907.540 7.070 2908.140 7.210 ;
        RECT 2907.540 2.400 2907.680 7.070 ;
        RECT 2907.470 0.000 2907.750 2.400 ;
      LAYER via2 ;
        RECT 1754.710 44.400 1754.990 44.680 ;
        RECT 2907.930 44.400 2908.210 44.680 ;
      LAYER met3 ;
        RECT 1754.685 44.690 1755.015 44.705 ;
        RECT 2907.905 44.690 2908.235 44.705 ;
        RECT 1754.685 44.390 2908.235 44.690 ;
        RECT 1754.685 44.375 1755.015 44.390 ;
        RECT 2907.905 44.375 2908.235 44.390 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 855.390 33.560 855.710 33.620 ;
        RECT 1327.810 33.560 1328.130 33.620 ;
        RECT 855.390 33.420 1328.130 33.560 ;
        RECT 855.390 33.360 855.710 33.420 ;
        RECT 1327.810 33.360 1328.130 33.420 ;
      LAYER via ;
        RECT 855.420 33.360 855.680 33.620 ;
        RECT 1327.840 33.360 1328.100 33.620 ;
      LAYER met2 ;
        RECT 1327.900 33.650 1328.040 54.000 ;
        RECT 855.420 33.330 855.680 33.650 ;
        RECT 1327.840 33.330 1328.100 33.650 ;
        RECT 855.480 2.400 855.620 33.330 ;
        RECT 855.410 0.000 855.690 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 873.330 33.900 873.650 33.960 ;
        RECT 1330.110 33.900 1330.430 33.960 ;
        RECT 873.330 33.760 1330.430 33.900 ;
        RECT 873.330 33.700 873.650 33.760 ;
        RECT 1330.110 33.700 1330.430 33.760 ;
      LAYER via ;
        RECT 873.360 33.700 873.620 33.960 ;
        RECT 1330.140 33.700 1330.400 33.960 ;
      LAYER met2 ;
        RECT 1330.200 33.990 1330.340 54.000 ;
        RECT 873.360 33.670 873.620 33.990 ;
        RECT 1330.140 33.670 1330.400 33.990 ;
        RECT 873.420 2.400 873.560 33.670 ;
        RECT 873.350 0.000 873.630 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 891.270 34.240 891.590 34.300 ;
        RECT 1334.710 34.240 1335.030 34.300 ;
        RECT 891.270 34.100 1335.030 34.240 ;
        RECT 891.270 34.040 891.590 34.100 ;
        RECT 1334.710 34.040 1335.030 34.100 ;
      LAYER via ;
        RECT 891.300 34.040 891.560 34.300 ;
        RECT 1334.740 34.040 1335.000 34.300 ;
      LAYER met2 ;
        RECT 1334.800 34.330 1334.940 54.000 ;
        RECT 891.300 34.010 891.560 34.330 ;
        RECT 1334.740 34.010 1335.000 34.330 ;
        RECT 891.360 2.400 891.500 34.010 ;
        RECT 891.290 0.000 891.570 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 909.210 30.500 909.530 30.560 ;
        RECT 1336.550 30.500 1336.870 30.560 ;
        RECT 909.210 30.360 1336.870 30.500 ;
        RECT 909.210 30.300 909.530 30.360 ;
        RECT 1336.550 30.300 1336.870 30.360 ;
      LAYER via ;
        RECT 909.240 30.300 909.500 30.560 ;
        RECT 1336.580 30.300 1336.840 30.560 ;
      LAYER met2 ;
        RECT 1336.640 30.590 1336.780 54.000 ;
        RECT 909.240 30.270 909.500 30.590 ;
        RECT 1336.580 30.270 1336.840 30.590 ;
        RECT 909.300 2.400 909.440 30.270 ;
        RECT 909.230 0.000 909.510 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 926.690 29.480 927.010 29.540 ;
        RECT 1342.070 29.480 1342.390 29.540 ;
        RECT 926.690 29.340 1342.390 29.480 ;
        RECT 926.690 29.280 927.010 29.340 ;
        RECT 1342.070 29.280 1342.390 29.340 ;
      LAYER via ;
        RECT 926.720 29.280 926.980 29.540 ;
        RECT 1342.100 29.280 1342.360 29.540 ;
      LAYER met2 ;
        RECT 1342.160 29.570 1342.300 54.000 ;
        RECT 926.720 29.250 926.980 29.570 ;
        RECT 1342.100 29.250 1342.360 29.570 ;
        RECT 926.780 2.400 926.920 29.250 ;
        RECT 926.710 0.000 926.990 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 944.630 29.140 944.950 29.200 ;
        RECT 1341.610 29.140 1341.930 29.200 ;
        RECT 944.630 29.000 1341.930 29.140 ;
        RECT 944.630 28.940 944.950 29.000 ;
        RECT 1341.610 28.940 1341.930 29.000 ;
      LAYER via ;
        RECT 944.660 28.940 944.920 29.200 ;
        RECT 1341.640 28.940 1341.900 29.200 ;
      LAYER met2 ;
        RECT 1341.700 29.230 1341.840 54.000 ;
        RECT 944.660 28.910 944.920 29.230 ;
        RECT 1341.640 28.910 1341.900 29.230 ;
        RECT 944.720 2.400 944.860 28.910 ;
        RECT 944.650 0.000 944.930 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 962.570 28.800 962.890 28.860 ;
        RECT 1349.430 28.800 1349.750 28.860 ;
        RECT 962.570 28.660 1349.750 28.800 ;
        RECT 962.570 28.600 962.890 28.660 ;
        RECT 1349.430 28.600 1349.750 28.660 ;
      LAYER via ;
        RECT 962.600 28.600 962.860 28.860 ;
        RECT 1349.460 28.600 1349.720 28.860 ;
      LAYER met2 ;
        RECT 1349.520 28.890 1349.660 54.000 ;
        RECT 962.600 28.570 962.860 28.890 ;
        RECT 1349.460 28.570 1349.720 28.890 ;
        RECT 962.660 2.400 962.800 28.570 ;
        RECT 962.590 0.000 962.870 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 980.585 13.005 980.755 28.475 ;
      LAYER mcon ;
        RECT 980.585 28.305 980.755 28.475 ;
      LAYER met1 ;
        RECT 980.525 28.460 980.815 28.505 ;
        RECT 1348.970 28.460 1349.290 28.520 ;
        RECT 980.525 28.320 1349.290 28.460 ;
        RECT 980.525 28.275 980.815 28.320 ;
        RECT 1348.970 28.260 1349.290 28.320 ;
        RECT 980.510 13.160 980.830 13.220 ;
        RECT 980.315 13.020 980.830 13.160 ;
        RECT 980.510 12.960 980.830 13.020 ;
      LAYER via ;
        RECT 1349.000 28.260 1349.260 28.520 ;
        RECT 980.540 12.960 980.800 13.220 ;
      LAYER met2 ;
        RECT 1349.060 28.550 1349.200 54.000 ;
        RECT 1349.000 28.230 1349.260 28.550 ;
        RECT 980.540 12.930 980.800 13.250 ;
        RECT 980.600 2.400 980.740 12.930 ;
        RECT 980.530 0.000 980.810 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 659.430 31.860 659.750 31.920 ;
        RECT 1286.870 31.860 1287.190 31.920 ;
        RECT 659.430 31.720 1287.190 31.860 ;
        RECT 659.430 31.660 659.750 31.720 ;
        RECT 1286.870 31.660 1287.190 31.720 ;
      LAYER via ;
        RECT 659.460 31.660 659.720 31.920 ;
        RECT 1286.900 31.660 1287.160 31.920 ;
      LAYER met2 ;
        RECT 1286.960 31.950 1287.100 54.000 ;
        RECT 659.460 31.630 659.720 31.950 ;
        RECT 1286.900 31.630 1287.160 31.950 ;
        RECT 659.520 2.400 659.660 31.630 ;
        RECT 659.450 0.000 659.730 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 998.450 28.120 998.770 28.180 ;
        RECT 1356.330 28.120 1356.650 28.180 ;
        RECT 998.450 27.980 1356.650 28.120 ;
        RECT 998.450 27.920 998.770 27.980 ;
        RECT 1356.330 27.920 1356.650 27.980 ;
      LAYER via ;
        RECT 998.480 27.920 998.740 28.180 ;
        RECT 1356.360 27.920 1356.620 28.180 ;
      LAYER met2 ;
        RECT 1356.420 28.210 1356.560 54.000 ;
        RECT 998.480 27.890 998.740 28.210 ;
        RECT 1356.360 27.890 1356.620 28.210 ;
        RECT 998.540 2.400 998.680 27.890 ;
        RECT 998.470 0.000 998.750 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1015.930 27.780 1016.250 27.840 ;
        RECT 1355.870 27.780 1356.190 27.840 ;
        RECT 1015.930 27.640 1356.190 27.780 ;
        RECT 1015.930 27.580 1016.250 27.640 ;
        RECT 1355.870 27.580 1356.190 27.640 ;
      LAYER via ;
        RECT 1015.960 27.580 1016.220 27.840 ;
        RECT 1355.900 27.580 1356.160 27.840 ;
      LAYER met2 ;
        RECT 1355.960 27.870 1356.100 54.000 ;
        RECT 1015.960 27.550 1016.220 27.870 ;
        RECT 1355.900 27.550 1356.160 27.870 ;
        RECT 1016.020 2.400 1016.160 27.550 ;
        RECT 1015.950 0.000 1016.230 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1364.225 30.685 1364.395 41.395 ;
      LAYER mcon ;
        RECT 1364.225 41.225 1364.395 41.395 ;
      LAYER met1 ;
        RECT 1364.150 41.380 1364.470 41.440 ;
        RECT 1363.955 41.240 1364.470 41.380 ;
        RECT 1364.150 41.180 1364.470 41.240 ;
        RECT 1079.410 30.840 1079.730 30.900 ;
        RECT 1364.165 30.840 1364.455 30.885 ;
        RECT 1079.410 30.700 1364.455 30.840 ;
        RECT 1079.410 30.640 1079.730 30.700 ;
        RECT 1364.165 30.655 1364.455 30.700 ;
      LAYER via ;
        RECT 1364.180 41.180 1364.440 41.440 ;
        RECT 1079.440 30.640 1079.700 30.900 ;
      LAYER met2 ;
        RECT 1364.240 41.470 1364.380 54.000 ;
        RECT 1364.180 41.150 1364.440 41.470 ;
        RECT 1079.440 30.610 1079.700 30.930 ;
        RECT 1079.500 29.765 1079.640 30.610 ;
        RECT 1033.890 29.395 1034.170 29.765 ;
        RECT 1079.430 29.395 1079.710 29.765 ;
        RECT 1033.960 2.400 1034.100 29.395 ;
        RECT 1033.890 0.000 1034.170 2.400 ;
      LAYER via2 ;
        RECT 1033.890 29.440 1034.170 29.720 ;
        RECT 1079.430 29.440 1079.710 29.720 ;
      LAYER met3 ;
        RECT 1033.865 29.730 1034.195 29.745 ;
        RECT 1079.405 29.730 1079.735 29.745 ;
        RECT 1033.865 29.430 1079.735 29.730 ;
        RECT 1033.865 29.415 1034.195 29.430 ;
        RECT 1079.405 29.415 1079.735 29.430 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1126.330 31.180 1126.650 31.240 ;
        RECT 1363.230 31.180 1363.550 31.240 ;
        RECT 1126.330 31.040 1363.550 31.180 ;
        RECT 1126.330 30.980 1126.650 31.040 ;
        RECT 1363.230 30.980 1363.550 31.040 ;
      LAYER via ;
        RECT 1126.360 30.980 1126.620 31.240 ;
        RECT 1363.260 30.980 1363.520 31.240 ;
      LAYER met2 ;
        RECT 1363.320 31.270 1363.460 54.000 ;
        RECT 1126.360 30.950 1126.620 31.270 ;
        RECT 1363.260 30.950 1363.520 31.270 ;
        RECT 1126.420 29.085 1126.560 30.950 ;
        RECT 1051.830 28.715 1052.110 29.085 ;
        RECT 1126.350 28.715 1126.630 29.085 ;
        RECT 1051.900 2.400 1052.040 28.715 ;
        RECT 1051.830 0.000 1052.110 2.400 ;
      LAYER via2 ;
        RECT 1051.830 28.760 1052.110 29.040 ;
        RECT 1126.350 28.760 1126.630 29.040 ;
      LAYER met3 ;
        RECT 1051.805 29.050 1052.135 29.065 ;
        RECT 1126.325 29.050 1126.655 29.065 ;
        RECT 1051.805 28.750 1126.655 29.050 ;
        RECT 1051.805 28.735 1052.135 28.750 ;
        RECT 1126.325 28.735 1126.655 28.750 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1072.600 48.805 1072.740 54.000 ;
        RECT 1069.770 48.435 1070.050 48.805 ;
        RECT 1072.530 48.435 1072.810 48.805 ;
        RECT 1069.840 2.400 1069.980 48.435 ;
        RECT 1069.770 0.000 1070.050 2.400 ;
      LAYER via2 ;
        RECT 1069.770 48.480 1070.050 48.760 ;
        RECT 1072.530 48.480 1072.810 48.760 ;
      LAYER met3 ;
        RECT 1069.745 48.770 1070.075 48.785 ;
        RECT 1072.505 48.770 1072.835 48.785 ;
        RECT 1069.745 48.470 1072.835 48.770 ;
        RECT 1069.745 48.455 1070.075 48.470 ;
        RECT 1072.505 48.455 1072.835 48.470 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1087.690 19.960 1088.010 20.020 ;
        RECT 1092.290 19.960 1092.610 20.020 ;
        RECT 1087.690 19.820 1092.610 19.960 ;
        RECT 1087.690 19.760 1088.010 19.820 ;
        RECT 1092.290 19.760 1092.610 19.820 ;
      LAYER via ;
        RECT 1087.720 19.760 1087.980 20.020 ;
        RECT 1092.320 19.760 1092.580 20.020 ;
      LAYER met2 ;
        RECT 1092.380 20.050 1092.520 54.000 ;
        RECT 1087.720 19.730 1087.980 20.050 ;
        RECT 1092.320 19.730 1092.580 20.050 ;
        RECT 1087.780 2.400 1087.920 19.730 ;
        RECT 1087.710 0.000 1087.990 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1105.170 2.960 1105.490 3.020 ;
        RECT 1106.090 2.960 1106.410 3.020 ;
        RECT 1105.170 2.820 1106.410 2.960 ;
        RECT 1105.170 2.760 1105.490 2.820 ;
        RECT 1106.090 2.760 1106.410 2.820 ;
      LAYER via ;
        RECT 1105.200 2.760 1105.460 3.020 ;
        RECT 1106.120 2.760 1106.380 3.020 ;
      LAYER met2 ;
        RECT 1106.180 3.050 1106.320 54.000 ;
        RECT 1105.200 2.730 1105.460 3.050 ;
        RECT 1106.120 2.730 1106.380 3.050 ;
        RECT 1105.260 2.400 1105.400 2.730 ;
        RECT 1105.190 0.000 1105.470 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1125.500 48.805 1125.640 54.000 ;
        RECT 1125.430 48.435 1125.710 48.805 ;
        RECT 1126.350 48.435 1126.630 48.805 ;
        RECT 1126.420 39.965 1126.560 48.435 ;
        RECT 1123.130 39.595 1123.410 39.965 ;
        RECT 1126.350 39.595 1126.630 39.965 ;
        RECT 1123.200 2.400 1123.340 39.595 ;
        RECT 1123.130 0.000 1123.410 2.400 ;
      LAYER via2 ;
        RECT 1125.430 48.480 1125.710 48.760 ;
        RECT 1126.350 48.480 1126.630 48.760 ;
        RECT 1123.130 39.640 1123.410 39.920 ;
        RECT 1126.350 39.640 1126.630 39.920 ;
      LAYER met3 ;
        RECT 1125.405 48.770 1125.735 48.785 ;
        RECT 1126.325 48.770 1126.655 48.785 ;
        RECT 1125.405 48.470 1126.655 48.770 ;
        RECT 1125.405 48.455 1125.735 48.470 ;
        RECT 1126.325 48.455 1126.655 48.470 ;
        RECT 1123.105 39.930 1123.435 39.945 ;
        RECT 1126.325 39.930 1126.655 39.945 ;
        RECT 1123.105 39.630 1126.655 39.930 ;
        RECT 1123.105 39.615 1123.435 39.630 ;
        RECT 1126.325 39.615 1126.655 39.630 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1141.050 20.300 1141.370 20.360 ;
        RECT 1147.490 20.300 1147.810 20.360 ;
        RECT 1141.050 20.160 1147.810 20.300 ;
        RECT 1141.050 20.100 1141.370 20.160 ;
        RECT 1147.490 20.100 1147.810 20.160 ;
      LAYER via ;
        RECT 1141.080 20.100 1141.340 20.360 ;
        RECT 1147.520 20.100 1147.780 20.360 ;
      LAYER met2 ;
        RECT 1147.580 20.390 1147.720 54.000 ;
        RECT 1141.080 20.070 1141.340 20.390 ;
        RECT 1147.520 20.070 1147.780 20.390 ;
        RECT 1141.140 2.400 1141.280 20.070 ;
        RECT 1141.070 0.000 1141.350 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1158.990 2.960 1159.310 3.020 ;
        RECT 1159.910 2.960 1160.230 3.020 ;
        RECT 1158.990 2.820 1160.230 2.960 ;
        RECT 1158.990 2.760 1159.310 2.820 ;
        RECT 1159.910 2.760 1160.230 2.820 ;
      LAYER via ;
        RECT 1159.020 2.760 1159.280 3.020 ;
        RECT 1159.940 2.760 1160.200 3.020 ;
      LAYER met2 ;
        RECT 1160.920 48.805 1161.060 54.000 ;
        RECT 1159.470 48.435 1159.750 48.805 ;
        RECT 1160.850 48.435 1161.130 48.805 ;
        RECT 1159.540 24.890 1159.680 48.435 ;
        RECT 1159.540 24.750 1160.140 24.890 ;
        RECT 1160.000 3.050 1160.140 24.750 ;
        RECT 1159.020 2.730 1159.280 3.050 ;
        RECT 1159.940 2.730 1160.200 3.050 ;
        RECT 1159.080 2.400 1159.220 2.730 ;
        RECT 1159.010 0.000 1159.290 2.400 ;
      LAYER via2 ;
        RECT 1159.470 48.480 1159.750 48.760 ;
        RECT 1160.850 48.480 1161.130 48.760 ;
      LAYER met3 ;
        RECT 1159.445 48.770 1159.775 48.785 ;
        RECT 1160.825 48.770 1161.155 48.785 ;
        RECT 1159.445 48.470 1161.155 48.770 ;
        RECT 1159.445 48.455 1159.775 48.470 ;
        RECT 1160.825 48.455 1161.155 48.470 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 676.540 48.805 676.680 54.000 ;
        RECT 676.470 48.435 676.750 48.805 ;
        RECT 677.390 48.435 677.670 48.805 ;
        RECT 677.460 3.130 677.600 48.435 ;
        RECT 677.000 2.990 677.600 3.130 ;
        RECT 677.000 2.400 677.140 2.990 ;
        RECT 676.930 0.000 677.210 2.400 ;
      LAYER via2 ;
        RECT 676.470 48.480 676.750 48.760 ;
        RECT 677.390 48.480 677.670 48.760 ;
      LAYER met3 ;
        RECT 676.445 48.770 676.775 48.785 ;
        RECT 677.365 48.770 677.695 48.785 ;
        RECT 676.445 48.470 677.695 48.770 ;
        RECT 676.445 48.455 676.775 48.470 ;
        RECT 677.365 48.455 677.695 48.470 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1176.470 20.640 1176.790 20.700 ;
        RECT 1181.990 20.640 1182.310 20.700 ;
        RECT 1176.470 20.500 1182.310 20.640 ;
        RECT 1176.470 20.440 1176.790 20.500 ;
        RECT 1181.990 20.440 1182.310 20.500 ;
      LAYER via ;
        RECT 1176.500 20.440 1176.760 20.700 ;
        RECT 1182.020 20.440 1182.280 20.700 ;
      LAYER met2 ;
        RECT 1182.080 20.730 1182.220 54.000 ;
        RECT 1176.500 20.410 1176.760 20.730 ;
        RECT 1182.020 20.410 1182.280 20.730 ;
        RECT 1176.560 2.400 1176.700 20.410 ;
        RECT 1176.490 0.000 1176.770 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1194.410 39.340 1194.730 39.400 ;
        RECT 1397.730 39.340 1398.050 39.400 ;
        RECT 1194.410 39.200 1398.050 39.340 ;
        RECT 1194.410 39.140 1194.730 39.200 ;
        RECT 1397.730 39.140 1398.050 39.200 ;
      LAYER via ;
        RECT 1194.440 39.140 1194.700 39.400 ;
        RECT 1397.760 39.140 1398.020 39.400 ;
      LAYER met2 ;
        RECT 1397.820 39.430 1397.960 54.000 ;
        RECT 1194.440 39.110 1194.700 39.430 ;
        RECT 1397.760 39.110 1398.020 39.430 ;
        RECT 1194.500 2.400 1194.640 39.110 ;
        RECT 1194.430 0.000 1194.710 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1212.350 39.680 1212.670 39.740 ;
        RECT 1399.110 39.680 1399.430 39.740 ;
        RECT 1212.350 39.540 1399.430 39.680 ;
        RECT 1212.350 39.480 1212.670 39.540 ;
        RECT 1399.110 39.480 1399.430 39.540 ;
      LAYER via ;
        RECT 1212.380 39.480 1212.640 39.740 ;
        RECT 1399.140 39.480 1399.400 39.740 ;
      LAYER met2 ;
        RECT 1399.200 39.770 1399.340 54.000 ;
        RECT 1212.380 39.450 1212.640 39.770 ;
        RECT 1399.140 39.450 1399.400 39.770 ;
        RECT 1212.440 2.400 1212.580 39.450 ;
        RECT 1212.370 0.000 1212.650 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1229.830 40.020 1230.150 40.080 ;
        RECT 1404.170 40.020 1404.490 40.080 ;
        RECT 1229.830 39.880 1404.490 40.020 ;
        RECT 1229.830 39.820 1230.150 39.880 ;
        RECT 1404.170 39.820 1404.490 39.880 ;
      LAYER via ;
        RECT 1229.860 39.820 1230.120 40.080 ;
        RECT 1404.200 39.820 1404.460 40.080 ;
      LAYER met2 ;
        RECT 1404.260 40.110 1404.400 54.000 ;
        RECT 1229.860 39.790 1230.120 40.110 ;
        RECT 1404.200 39.790 1404.460 40.110 ;
        RECT 1229.920 20.130 1230.060 39.790 ;
        RECT 1229.920 19.990 1230.520 20.130 ;
        RECT 1230.380 2.400 1230.520 19.990 ;
        RECT 1230.310 0.000 1230.590 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1248.230 40.360 1248.550 40.420 ;
        RECT 1403.710 40.360 1404.030 40.420 ;
        RECT 1248.230 40.220 1404.030 40.360 ;
        RECT 1248.230 40.160 1248.550 40.220 ;
        RECT 1403.710 40.160 1404.030 40.220 ;
      LAYER via ;
        RECT 1248.260 40.160 1248.520 40.420 ;
        RECT 1403.740 40.160 1404.000 40.420 ;
      LAYER met2 ;
        RECT 1403.800 40.450 1403.940 54.000 ;
        RECT 1248.260 40.130 1248.520 40.450 ;
        RECT 1403.740 40.130 1404.000 40.450 ;
        RECT 1248.320 2.400 1248.460 40.130 ;
        RECT 1248.250 0.000 1248.530 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1265.710 15.880 1266.030 15.940 ;
        RECT 1270.770 15.880 1271.090 15.940 ;
        RECT 1265.710 15.740 1271.090 15.880 ;
        RECT 1265.710 15.680 1266.030 15.740 ;
        RECT 1270.770 15.680 1271.090 15.740 ;
      LAYER via ;
        RECT 1265.740 15.680 1266.000 15.940 ;
        RECT 1270.800 15.680 1271.060 15.940 ;
      LAYER met2 ;
        RECT 1271.320 46.650 1271.460 54.000 ;
        RECT 1270.860 46.510 1271.460 46.650 ;
        RECT 1270.860 15.970 1271.000 46.510 ;
        RECT 1265.740 15.650 1266.000 15.970 ;
        RECT 1270.800 15.650 1271.060 15.970 ;
        RECT 1265.800 2.400 1265.940 15.650 ;
        RECT 1265.730 0.000 1266.010 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1283.650 2.960 1283.970 3.020 ;
        RECT 1285.490 2.960 1285.810 3.020 ;
        RECT 1283.650 2.820 1285.810 2.960 ;
        RECT 1283.650 2.760 1283.970 2.820 ;
        RECT 1285.490 2.760 1285.810 2.820 ;
      LAYER via ;
        RECT 1283.680 2.760 1283.940 3.020 ;
        RECT 1285.520 2.760 1285.780 3.020 ;
      LAYER met2 ;
        RECT 1285.580 3.050 1285.720 54.000 ;
        RECT 1283.680 2.730 1283.940 3.050 ;
        RECT 1285.520 2.730 1285.780 3.050 ;
        RECT 1283.740 2.400 1283.880 2.730 ;
        RECT 1283.670 0.000 1283.950 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1301.590 20.640 1301.910 20.700 ;
        RECT 1306.190 20.640 1306.510 20.700 ;
        RECT 1301.590 20.500 1306.510 20.640 ;
        RECT 1301.590 20.440 1301.910 20.500 ;
        RECT 1306.190 20.440 1306.510 20.500 ;
      LAYER via ;
        RECT 1301.620 20.440 1301.880 20.700 ;
        RECT 1306.220 20.440 1306.480 20.700 ;
      LAYER met2 ;
        RECT 1306.280 20.730 1306.420 54.000 ;
        RECT 1301.620 20.410 1301.880 20.730 ;
        RECT 1306.220 20.410 1306.480 20.730 ;
        RECT 1301.680 2.400 1301.820 20.410 ;
        RECT 1301.610 0.000 1301.890 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1319.530 18.600 1319.850 18.660 ;
        RECT 1418.430 18.600 1418.750 18.660 ;
        RECT 1319.530 18.460 1418.750 18.600 ;
        RECT 1319.530 18.400 1319.850 18.460 ;
        RECT 1418.430 18.400 1418.750 18.460 ;
      LAYER via ;
        RECT 1319.560 18.400 1319.820 18.660 ;
        RECT 1418.460 18.400 1418.720 18.660 ;
      LAYER met2 ;
        RECT 1418.520 18.690 1418.660 54.000 ;
        RECT 1319.560 18.370 1319.820 18.690 ;
        RECT 1418.460 18.370 1418.720 18.690 ;
        RECT 1319.620 2.400 1319.760 18.370 ;
        RECT 1319.550 0.000 1319.830 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1337.470 19.960 1337.790 20.020 ;
        RECT 1424.410 19.960 1424.730 20.020 ;
        RECT 1337.470 19.820 1424.730 19.960 ;
        RECT 1337.470 19.760 1337.790 19.820 ;
        RECT 1424.410 19.760 1424.730 19.820 ;
      LAYER via ;
        RECT 1337.500 19.760 1337.760 20.020 ;
        RECT 1424.440 19.760 1424.700 20.020 ;
      LAYER met2 ;
        RECT 1424.500 20.050 1424.640 54.000 ;
        RECT 1337.500 19.730 1337.760 20.050 ;
        RECT 1424.440 19.730 1424.700 20.050 ;
        RECT 1337.560 2.400 1337.700 19.730 ;
        RECT 1337.490 0.000 1337.770 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 694.850 18.260 695.170 18.320 ;
        RECT 698.990 18.260 699.310 18.320 ;
        RECT 694.850 18.120 699.310 18.260 ;
        RECT 694.850 18.060 695.170 18.120 ;
        RECT 698.990 18.060 699.310 18.120 ;
      LAYER via ;
        RECT 694.880 18.060 695.140 18.320 ;
        RECT 699.020 18.060 699.280 18.320 ;
      LAYER met2 ;
        RECT 699.080 18.350 699.220 54.000 ;
        RECT 694.880 18.030 695.140 18.350 ;
        RECT 699.020 18.030 699.280 18.350 ;
        RECT 694.940 2.400 695.080 18.030 ;
        RECT 694.870 0.000 695.150 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1354.950 15.880 1355.270 15.940 ;
        RECT 1354.950 15.740 1390.600 15.880 ;
        RECT 1354.950 15.680 1355.270 15.740 ;
        RECT 1390.460 15.540 1390.600 15.740 ;
        RECT 1427.630 15.540 1427.950 15.600 ;
        RECT 1390.460 15.400 1427.950 15.540 ;
        RECT 1427.630 15.340 1427.950 15.400 ;
      LAYER via ;
        RECT 1354.980 15.680 1355.240 15.940 ;
        RECT 1427.660 15.340 1427.920 15.600 ;
      LAYER met2 ;
        RECT 1354.980 15.650 1355.240 15.970 ;
        RECT 1355.040 2.400 1355.180 15.650 ;
        RECT 1427.720 15.630 1427.860 54.000 ;
        RECT 1427.660 15.310 1427.920 15.630 ;
        RECT 1354.970 0.000 1355.250 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1372.890 14.860 1373.210 14.920 ;
        RECT 1433.150 14.860 1433.470 14.920 ;
        RECT 1372.890 14.720 1433.470 14.860 ;
        RECT 1372.890 14.660 1373.210 14.720 ;
        RECT 1433.150 14.660 1433.470 14.720 ;
      LAYER via ;
        RECT 1372.920 14.660 1373.180 14.920 ;
        RECT 1433.180 14.660 1433.440 14.920 ;
      LAYER met2 ;
        RECT 1433.240 14.950 1433.380 54.000 ;
        RECT 1372.920 14.630 1373.180 14.950 ;
        RECT 1433.180 14.630 1433.440 14.950 ;
        RECT 1372.980 2.400 1373.120 14.630 ;
        RECT 1372.910 0.000 1373.190 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1390.830 15.880 1391.150 15.940 ;
        RECT 1434.070 15.880 1434.390 15.940 ;
        RECT 1390.830 15.740 1434.390 15.880 ;
        RECT 1390.830 15.680 1391.150 15.740 ;
        RECT 1434.070 15.680 1434.390 15.740 ;
      LAYER via ;
        RECT 1390.860 15.680 1391.120 15.940 ;
        RECT 1434.100 15.680 1434.360 15.940 ;
      LAYER met2 ;
        RECT 1434.160 15.970 1434.300 54.000 ;
        RECT 1390.860 15.650 1391.120 15.970 ;
        RECT 1434.100 15.650 1434.360 15.970 ;
        RECT 1390.920 2.400 1391.060 15.650 ;
        RECT 1390.850 0.000 1391.130 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1408.770 14.180 1409.090 14.240 ;
        RECT 1440.970 14.180 1441.290 14.240 ;
        RECT 1408.770 14.040 1441.290 14.180 ;
        RECT 1408.770 13.980 1409.090 14.040 ;
        RECT 1440.970 13.980 1441.290 14.040 ;
      LAYER via ;
        RECT 1408.800 13.980 1409.060 14.240 ;
        RECT 1441.000 13.980 1441.260 14.240 ;
      LAYER met2 ;
        RECT 1441.060 14.270 1441.200 54.000 ;
        RECT 1408.800 13.950 1409.060 14.270 ;
        RECT 1441.000 13.950 1441.260 14.270 ;
        RECT 1408.860 2.400 1409.000 13.950 ;
        RECT 1408.790 0.000 1409.070 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1426.250 18.260 1426.570 18.320 ;
        RECT 1448.330 18.260 1448.650 18.320 ;
        RECT 1426.250 18.120 1448.650 18.260 ;
        RECT 1426.250 18.060 1426.570 18.120 ;
        RECT 1448.330 18.060 1448.650 18.120 ;
      LAYER via ;
        RECT 1426.280 18.060 1426.540 18.320 ;
        RECT 1448.360 18.060 1448.620 18.320 ;
      LAYER met2 ;
        RECT 1448.420 18.350 1448.560 54.000 ;
        RECT 1426.280 18.030 1426.540 18.350 ;
        RECT 1448.360 18.030 1448.620 18.350 ;
        RECT 1426.340 2.400 1426.480 18.030 ;
        RECT 1426.270 0.000 1426.550 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1444.190 20.640 1444.510 20.700 ;
        RECT 1446.950 20.640 1447.270 20.700 ;
        RECT 1444.190 20.500 1447.270 20.640 ;
        RECT 1444.190 20.440 1444.510 20.500 ;
        RECT 1446.950 20.440 1447.270 20.500 ;
      LAYER via ;
        RECT 1444.220 20.440 1444.480 20.700 ;
        RECT 1446.980 20.440 1447.240 20.700 ;
      LAYER met2 ;
        RECT 1447.040 20.730 1447.180 54.000 ;
        RECT 1444.220 20.410 1444.480 20.730 ;
        RECT 1446.980 20.410 1447.240 20.730 ;
        RECT 1444.280 2.400 1444.420 20.410 ;
        RECT 1444.210 0.000 1444.490 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1457.530 20.640 1457.850 20.700 ;
        RECT 1462.130 20.640 1462.450 20.700 ;
        RECT 1457.530 20.500 1462.450 20.640 ;
        RECT 1457.530 20.440 1457.850 20.500 ;
        RECT 1462.130 20.440 1462.450 20.500 ;
      LAYER via ;
        RECT 1457.560 20.440 1457.820 20.700 ;
        RECT 1462.160 20.440 1462.420 20.700 ;
      LAYER met2 ;
        RECT 1457.620 20.730 1457.760 54.000 ;
        RECT 1457.560 20.410 1457.820 20.730 ;
        RECT 1462.160 20.410 1462.420 20.730 ;
        RECT 1462.220 2.400 1462.360 20.410 ;
        RECT 1462.150 0.000 1462.430 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1461.670 15.540 1461.990 15.600 ;
        RECT 1480.070 15.540 1480.390 15.600 ;
        RECT 1461.670 15.400 1480.390 15.540 ;
        RECT 1461.670 15.340 1461.990 15.400 ;
        RECT 1480.070 15.340 1480.390 15.400 ;
      LAYER via ;
        RECT 1461.700 15.340 1461.960 15.600 ;
        RECT 1480.100 15.340 1480.360 15.600 ;
      LAYER met2 ;
        RECT 1461.760 15.630 1461.900 54.000 ;
        RECT 1461.700 15.310 1461.960 15.630 ;
        RECT 1480.100 15.310 1480.360 15.630 ;
        RECT 1480.160 2.400 1480.300 15.310 ;
        RECT 1480.090 0.000 1480.370 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1464.430 18.600 1464.750 18.660 ;
        RECT 1498.010 18.600 1498.330 18.660 ;
        RECT 1464.430 18.460 1498.330 18.600 ;
        RECT 1464.430 18.400 1464.750 18.460 ;
        RECT 1498.010 18.400 1498.330 18.460 ;
      LAYER via ;
        RECT 1464.460 18.400 1464.720 18.660 ;
        RECT 1498.040 18.400 1498.300 18.660 ;
      LAYER met2 ;
        RECT 1464.520 18.690 1464.660 54.000 ;
        RECT 1464.460 18.370 1464.720 18.690 ;
        RECT 1498.040 18.370 1498.300 18.690 ;
        RECT 1498.100 2.400 1498.240 18.370 ;
        RECT 1498.030 0.000 1498.310 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1493.025 14.025 1493.195 16.915 ;
      LAYER mcon ;
        RECT 1493.025 16.745 1493.195 16.915 ;
      LAYER met1 ;
        RECT 1492.965 16.900 1493.255 16.945 ;
        RECT 1515.490 16.900 1515.810 16.960 ;
        RECT 1492.965 16.760 1515.810 16.900 ;
        RECT 1492.965 16.715 1493.255 16.760 ;
        RECT 1515.490 16.700 1515.810 16.760 ;
        RECT 1469.030 14.180 1469.350 14.240 ;
        RECT 1492.965 14.180 1493.255 14.225 ;
        RECT 1469.030 14.040 1493.255 14.180 ;
        RECT 1469.030 13.980 1469.350 14.040 ;
        RECT 1492.965 13.995 1493.255 14.040 ;
      LAYER via ;
        RECT 1515.520 16.700 1515.780 16.960 ;
        RECT 1469.060 13.980 1469.320 14.240 ;
      LAYER met2 ;
        RECT 1469.120 14.270 1469.260 54.000 ;
        RECT 1515.520 16.670 1515.780 16.990 ;
        RECT 1469.060 13.950 1469.320 14.270 ;
        RECT 1515.580 2.400 1515.720 16.670 ;
        RECT 1515.510 0.000 1515.790 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 712.420 17.580 712.560 54.000 ;
        RECT 712.420 17.440 713.020 17.580 ;
        RECT 712.880 2.400 713.020 17.440 ;
        RECT 712.810 0.000 713.090 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1470.870 15.200 1471.190 15.260 ;
        RECT 1470.870 15.060 1510.200 15.200 ;
        RECT 1470.870 15.000 1471.190 15.060 ;
        RECT 1510.060 14.520 1510.200 15.060 ;
        RECT 1533.430 14.520 1533.750 14.580 ;
        RECT 1510.060 14.380 1533.750 14.520 ;
        RECT 1533.430 14.320 1533.750 14.380 ;
      LAYER via ;
        RECT 1470.900 15.000 1471.160 15.260 ;
        RECT 1533.460 14.320 1533.720 14.580 ;
      LAYER met2 ;
        RECT 1470.960 15.290 1471.100 54.000 ;
        RECT 1470.900 14.970 1471.160 15.290 ;
        RECT 1533.460 14.290 1533.720 14.610 ;
        RECT 1533.520 2.400 1533.660 14.290 ;
        RECT 1533.450 0.000 1533.730 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1505.445 15.725 1505.615 17.255 ;
      LAYER mcon ;
        RECT 1505.445 17.085 1505.615 17.255 ;
      LAYER met1 ;
        RECT 1505.385 17.240 1505.675 17.285 ;
        RECT 1551.370 17.240 1551.690 17.300 ;
        RECT 1505.385 17.100 1551.690 17.240 ;
        RECT 1505.385 17.055 1505.675 17.100 ;
        RECT 1551.370 17.040 1551.690 17.100 ;
        RECT 1470.410 15.880 1470.730 15.940 ;
        RECT 1505.385 15.880 1505.675 15.925 ;
        RECT 1470.410 15.740 1505.675 15.880 ;
        RECT 1470.410 15.680 1470.730 15.740 ;
        RECT 1505.385 15.695 1505.675 15.740 ;
      LAYER via ;
        RECT 1551.400 17.040 1551.660 17.300 ;
        RECT 1470.440 15.680 1470.700 15.940 ;
      LAYER met2 ;
        RECT 1470.500 15.970 1470.640 54.000 ;
        RECT 1551.400 17.010 1551.660 17.330 ;
        RECT 1470.440 15.650 1470.700 15.970 ;
        RECT 1551.460 2.400 1551.600 17.010 ;
        RECT 1551.390 0.000 1551.670 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1478.690 18.260 1479.010 18.320 ;
        RECT 1569.310 18.260 1569.630 18.320 ;
        RECT 1478.690 18.120 1569.630 18.260 ;
        RECT 1478.690 18.060 1479.010 18.120 ;
        RECT 1569.310 18.060 1569.630 18.120 ;
      LAYER via ;
        RECT 1478.720 18.060 1478.980 18.320 ;
        RECT 1569.340 18.060 1569.600 18.320 ;
      LAYER met2 ;
        RECT 1478.780 18.350 1478.920 54.000 ;
        RECT 1478.720 18.030 1478.980 18.350 ;
        RECT 1569.340 18.030 1569.600 18.350 ;
        RECT 1569.400 2.400 1569.540 18.030 ;
        RECT 1569.330 0.000 1569.610 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1513.265 25.415 1513.435 26.435 ;
        RECT 1512.805 25.245 1513.435 25.415 ;
      LAYER mcon ;
        RECT 1513.265 26.265 1513.435 26.435 ;
      LAYER met1 ;
        RECT 1513.205 26.420 1513.495 26.465 ;
        RECT 1562.870 26.420 1563.190 26.480 ;
        RECT 1513.205 26.280 1563.190 26.420 ;
        RECT 1513.205 26.235 1513.495 26.280 ;
        RECT 1562.870 26.220 1563.190 26.280 ;
        RECT 1478.230 25.400 1478.550 25.460 ;
        RECT 1512.745 25.400 1513.035 25.445 ;
        RECT 1478.230 25.260 1513.035 25.400 ;
        RECT 1478.230 25.200 1478.550 25.260 ;
        RECT 1512.745 25.215 1513.035 25.260 ;
      LAYER via ;
        RECT 1562.900 26.220 1563.160 26.480 ;
        RECT 1478.260 25.200 1478.520 25.460 ;
      LAYER met2 ;
        RECT 1478.320 25.490 1478.460 54.000 ;
        RECT 1562.900 26.365 1563.160 26.510 ;
        RECT 1562.890 25.995 1563.170 26.365 ;
        RECT 1587.270 25.995 1587.550 26.365 ;
        RECT 1478.260 25.170 1478.520 25.490 ;
        RECT 1587.340 2.400 1587.480 25.995 ;
        RECT 1587.270 0.000 1587.550 2.400 ;
      LAYER via2 ;
        RECT 1562.890 26.040 1563.170 26.320 ;
        RECT 1587.270 26.040 1587.550 26.320 ;
      LAYER met3 ;
        RECT 1562.865 26.330 1563.195 26.345 ;
        RECT 1587.245 26.330 1587.575 26.345 ;
        RECT 1562.865 26.030 1587.575 26.330 ;
        RECT 1562.865 26.015 1563.195 26.030 ;
        RECT 1587.245 26.015 1587.575 26.030 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1562.025 24.735 1562.195 26.095 ;
        RECT 1562.025 24.565 1563.115 24.735 ;
        RECT 1562.945 20.145 1563.115 24.565 ;
      LAYER mcon ;
        RECT 1562.025 25.925 1562.195 26.095 ;
      LAYER met1 ;
        RECT 1483.750 26.080 1484.070 26.140 ;
        RECT 1561.965 26.080 1562.255 26.125 ;
        RECT 1483.750 25.940 1562.255 26.080 ;
        RECT 1483.750 25.880 1484.070 25.940 ;
        RECT 1561.965 25.895 1562.255 25.940 ;
        RECT 1562.885 20.300 1563.175 20.345 ;
        RECT 1604.730 20.300 1605.050 20.360 ;
        RECT 1562.885 20.160 1605.050 20.300 ;
        RECT 1562.885 20.115 1563.175 20.160 ;
        RECT 1604.730 20.100 1605.050 20.160 ;
      LAYER via ;
        RECT 1483.780 25.880 1484.040 26.140 ;
        RECT 1604.760 20.100 1605.020 20.360 ;
      LAYER met2 ;
        RECT 1483.840 26.170 1483.980 54.000 ;
        RECT 1483.780 25.850 1484.040 26.170 ;
        RECT 1604.760 20.070 1605.020 20.390 ;
        RECT 1604.820 2.400 1604.960 20.070 ;
        RECT 1604.750 0.000 1605.030 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1505.905 20.145 1506.075 25.755 ;
      LAYER mcon ;
        RECT 1505.905 25.585 1506.075 25.755 ;
      LAYER met1 ;
        RECT 1484.210 25.740 1484.530 25.800 ;
        RECT 1505.845 25.740 1506.135 25.785 ;
        RECT 1484.210 25.600 1506.135 25.740 ;
        RECT 1484.210 25.540 1484.530 25.600 ;
        RECT 1505.845 25.555 1506.135 25.600 ;
        RECT 1513.190 21.320 1513.510 21.380 ;
        RECT 1622.670 21.320 1622.990 21.380 ;
        RECT 1513.190 21.180 1622.990 21.320 ;
        RECT 1513.190 21.120 1513.510 21.180 ;
        RECT 1622.670 21.120 1622.990 21.180 ;
        RECT 1505.845 20.300 1506.135 20.345 ;
        RECT 1512.730 20.300 1513.050 20.360 ;
        RECT 1505.845 20.160 1513.050 20.300 ;
        RECT 1505.845 20.115 1506.135 20.160 ;
        RECT 1512.730 20.100 1513.050 20.160 ;
      LAYER via ;
        RECT 1484.240 25.540 1484.500 25.800 ;
        RECT 1513.220 21.120 1513.480 21.380 ;
        RECT 1622.700 21.120 1622.960 21.380 ;
        RECT 1512.760 20.100 1513.020 20.360 ;
      LAYER met2 ;
        RECT 1484.300 25.830 1484.440 54.000 ;
        RECT 1484.240 25.510 1484.500 25.830 ;
        RECT 1513.220 21.090 1513.480 21.410 ;
        RECT 1622.700 21.090 1622.960 21.410 ;
        RECT 1512.760 20.300 1513.020 20.390 ;
        RECT 1513.280 20.300 1513.420 21.090 ;
        RECT 1512.760 20.160 1513.420 20.300 ;
        RECT 1512.760 20.070 1513.020 20.160 ;
        RECT 1622.760 2.400 1622.900 21.090 ;
        RECT 1622.690 0.000 1622.970 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1492.030 22.680 1492.350 22.740 ;
        RECT 1512.730 22.680 1513.050 22.740 ;
        RECT 1492.030 22.540 1513.050 22.680 ;
        RECT 1492.030 22.480 1492.350 22.540 ;
        RECT 1512.730 22.480 1513.050 22.540 ;
        RECT 1515.490 22.680 1515.810 22.740 ;
        RECT 1640.610 22.680 1640.930 22.740 ;
        RECT 1515.490 22.540 1640.930 22.680 ;
        RECT 1515.490 22.480 1515.810 22.540 ;
        RECT 1640.610 22.480 1640.930 22.540 ;
      LAYER via ;
        RECT 1492.060 22.480 1492.320 22.740 ;
        RECT 1512.760 22.480 1513.020 22.740 ;
        RECT 1515.520 22.480 1515.780 22.740 ;
        RECT 1640.640 22.480 1640.900 22.740 ;
      LAYER met2 ;
        RECT 1492.120 22.770 1492.260 54.000 ;
        RECT 1492.060 22.450 1492.320 22.770 ;
        RECT 1512.750 22.595 1513.030 22.965 ;
        RECT 1515.510 22.595 1515.790 22.965 ;
        RECT 1512.760 22.450 1513.020 22.595 ;
        RECT 1515.520 22.450 1515.780 22.595 ;
        RECT 1640.640 22.450 1640.900 22.770 ;
        RECT 1640.700 2.400 1640.840 22.450 ;
        RECT 1640.630 0.000 1640.910 2.400 ;
      LAYER via2 ;
        RECT 1512.750 22.640 1513.030 22.920 ;
        RECT 1515.510 22.640 1515.790 22.920 ;
      LAYER met3 ;
        RECT 1512.725 22.930 1513.055 22.945 ;
        RECT 1515.485 22.930 1515.815 22.945 ;
        RECT 1512.725 22.630 1515.815 22.930 ;
        RECT 1512.725 22.615 1513.055 22.630 ;
        RECT 1515.485 22.615 1515.815 22.630 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1513.265 21.335 1513.435 22.695 ;
        RECT 1512.805 21.165 1513.435 21.335 ;
      LAYER mcon ;
        RECT 1513.265 22.525 1513.435 22.695 ;
      LAYER met1 ;
        RECT 1561.030 25.400 1561.350 25.460 ;
        RECT 1658.550 25.400 1658.870 25.460 ;
        RECT 1561.030 25.260 1658.870 25.400 ;
        RECT 1561.030 25.200 1561.350 25.260 ;
        RECT 1658.550 25.200 1658.870 25.260 ;
        RECT 1513.205 22.680 1513.495 22.725 ;
        RECT 1514.110 22.680 1514.430 22.740 ;
        RECT 1513.205 22.540 1514.430 22.680 ;
        RECT 1513.205 22.495 1513.495 22.540 ;
        RECT 1514.110 22.480 1514.430 22.540 ;
        RECT 1491.110 21.320 1491.430 21.380 ;
        RECT 1512.745 21.320 1513.035 21.365 ;
        RECT 1491.110 21.180 1513.035 21.320 ;
        RECT 1491.110 21.120 1491.430 21.180 ;
        RECT 1512.745 21.135 1513.035 21.180 ;
      LAYER via ;
        RECT 1561.060 25.200 1561.320 25.460 ;
        RECT 1658.580 25.200 1658.840 25.460 ;
        RECT 1514.140 22.480 1514.400 22.740 ;
        RECT 1491.140 21.120 1491.400 21.380 ;
      LAYER met2 ;
        RECT 1491.200 21.410 1491.340 54.000 ;
        RECT 1561.060 25.170 1561.320 25.490 ;
        RECT 1658.580 25.170 1658.840 25.490 ;
        RECT 1561.120 25.005 1561.260 25.170 ;
        RECT 1514.130 24.635 1514.410 25.005 ;
        RECT 1561.050 24.635 1561.330 25.005 ;
        RECT 1514.200 22.770 1514.340 24.635 ;
        RECT 1514.140 22.450 1514.400 22.770 ;
        RECT 1491.140 21.090 1491.400 21.410 ;
        RECT 1658.640 2.400 1658.780 25.170 ;
        RECT 1658.570 0.000 1658.850 2.400 ;
      LAYER via2 ;
        RECT 1514.130 24.680 1514.410 24.960 ;
        RECT 1561.050 24.680 1561.330 24.960 ;
      LAYER met3 ;
        RECT 1514.105 24.970 1514.435 24.985 ;
        RECT 1561.025 24.970 1561.355 24.985 ;
        RECT 1514.105 24.670 1561.355 24.970 ;
        RECT 1514.105 24.655 1514.435 24.670 ;
        RECT 1561.025 24.655 1561.355 24.670 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1538.105 23.205 1538.275 25.075 ;
      LAYER mcon ;
        RECT 1538.105 24.905 1538.275 25.075 ;
      LAYER met1 ;
        RECT 1538.045 25.060 1538.335 25.105 ;
        RECT 1676.030 25.060 1676.350 25.120 ;
        RECT 1538.045 24.920 1676.350 25.060 ;
        RECT 1538.045 24.875 1538.335 24.920 ;
        RECT 1676.030 24.860 1676.350 24.920 ;
        RECT 1499.390 23.360 1499.710 23.420 ;
        RECT 1538.045 23.360 1538.335 23.405 ;
        RECT 1499.390 23.220 1538.335 23.360 ;
        RECT 1499.390 23.160 1499.710 23.220 ;
        RECT 1538.045 23.175 1538.335 23.220 ;
      LAYER via ;
        RECT 1676.060 24.860 1676.320 25.120 ;
        RECT 1499.420 23.160 1499.680 23.420 ;
      LAYER met2 ;
        RECT 1499.480 23.450 1499.620 54.000 ;
        RECT 1676.060 24.830 1676.320 25.150 ;
        RECT 1499.420 23.130 1499.680 23.450 ;
        RECT 1676.120 2.400 1676.260 24.830 ;
        RECT 1676.050 0.000 1676.330 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1562.485 20.145 1562.655 23.715 ;
      LAYER mcon ;
        RECT 1562.485 23.545 1562.655 23.715 ;
      LAYER met1 ;
        RECT 1506.290 25.740 1506.610 25.800 ;
        RECT 1513.650 25.740 1513.970 25.800 ;
        RECT 1506.290 25.600 1513.970 25.740 ;
        RECT 1506.290 25.540 1506.610 25.600 ;
        RECT 1513.650 25.540 1513.970 25.600 ;
        RECT 1562.425 23.700 1562.715 23.745 ;
        RECT 1693.970 23.700 1694.290 23.760 ;
        RECT 1562.425 23.560 1694.290 23.700 ;
        RECT 1562.425 23.515 1562.715 23.560 ;
        RECT 1693.970 23.500 1694.290 23.560 ;
        RECT 1513.650 20.300 1513.970 20.360 ;
        RECT 1562.425 20.300 1562.715 20.345 ;
        RECT 1513.650 20.160 1562.715 20.300 ;
        RECT 1513.650 20.100 1513.970 20.160 ;
        RECT 1562.425 20.115 1562.715 20.160 ;
      LAYER via ;
        RECT 1506.320 25.540 1506.580 25.800 ;
        RECT 1513.680 25.540 1513.940 25.800 ;
        RECT 1694.000 23.500 1694.260 23.760 ;
        RECT 1513.680 20.100 1513.940 20.360 ;
      LAYER met2 ;
        RECT 1506.380 25.830 1506.520 54.000 ;
        RECT 1506.320 25.510 1506.580 25.830 ;
        RECT 1513.680 25.510 1513.940 25.830 ;
        RECT 1513.740 20.390 1513.880 25.510 ;
        RECT 1694.000 23.470 1694.260 23.790 ;
        RECT 1513.680 20.070 1513.940 20.390 ;
        RECT 1694.060 2.400 1694.200 23.470 ;
        RECT 1693.990 0.000 1694.270 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 730.730 37.640 731.050 37.700 ;
        RECT 1301.590 37.640 1301.910 37.700 ;
        RECT 730.730 37.500 1301.910 37.640 ;
        RECT 730.730 37.440 731.050 37.500 ;
        RECT 1301.590 37.440 1301.910 37.500 ;
      LAYER via ;
        RECT 730.760 37.440 731.020 37.700 ;
        RECT 1301.620 37.440 1301.880 37.700 ;
      LAYER met2 ;
        RECT 1301.680 37.730 1301.820 54.000 ;
        RECT 730.760 37.410 731.020 37.730 ;
        RECT 1301.620 37.410 1301.880 37.730 ;
        RECT 730.820 2.400 730.960 37.410 ;
        RECT 730.750 0.000 731.030 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1513.725 25.585 1514.355 25.755 ;
        RECT 1537.185 25.585 1538.735 25.755 ;
        RECT 1513.725 23.885 1513.895 25.585 ;
        RECT 1538.565 23.205 1538.735 25.585 ;
        RECT 1561.565 23.375 1561.735 26.775 ;
        RECT 1662.305 25.585 1662.475 26.435 ;
        RECT 1561.105 23.205 1561.735 23.375 ;
      LAYER mcon ;
        RECT 1561.565 26.605 1561.735 26.775 ;
        RECT 1514.185 25.585 1514.355 25.755 ;
        RECT 1662.305 26.265 1662.475 26.435 ;
      LAYER met1 ;
        RECT 1561.505 26.760 1561.795 26.805 ;
        RECT 1561.505 26.620 1586.100 26.760 ;
        RECT 1561.505 26.575 1561.795 26.620 ;
        RECT 1585.960 26.420 1586.100 26.620 ;
        RECT 1662.245 26.420 1662.535 26.465 ;
        RECT 1585.960 26.280 1662.535 26.420 ;
        RECT 1662.245 26.235 1662.535 26.280 ;
        RECT 1514.125 25.740 1514.415 25.785 ;
        RECT 1537.125 25.740 1537.415 25.785 ;
        RECT 1514.125 25.600 1537.415 25.740 ;
        RECT 1514.125 25.555 1514.415 25.600 ;
        RECT 1537.125 25.555 1537.415 25.600 ;
        RECT 1662.245 25.740 1662.535 25.785 ;
        RECT 1711.910 25.740 1712.230 25.800 ;
        RECT 1662.245 25.600 1712.230 25.740 ;
        RECT 1662.245 25.555 1662.535 25.600 ;
        RECT 1711.910 25.540 1712.230 25.600 ;
        RECT 1505.830 24.040 1506.150 24.100 ;
        RECT 1513.665 24.040 1513.955 24.085 ;
        RECT 1505.830 23.900 1513.955 24.040 ;
        RECT 1505.830 23.840 1506.150 23.900 ;
        RECT 1513.665 23.855 1513.955 23.900 ;
        RECT 1538.505 23.360 1538.795 23.405 ;
        RECT 1561.045 23.360 1561.335 23.405 ;
        RECT 1538.505 23.220 1561.335 23.360 ;
        RECT 1538.505 23.175 1538.795 23.220 ;
        RECT 1561.045 23.175 1561.335 23.220 ;
      LAYER via ;
        RECT 1711.940 25.540 1712.200 25.800 ;
        RECT 1505.860 23.840 1506.120 24.100 ;
      LAYER met2 ;
        RECT 1505.920 24.130 1506.060 54.000 ;
        RECT 1711.940 25.510 1712.200 25.830 ;
        RECT 1505.860 23.810 1506.120 24.130 ;
        RECT 1712.000 2.400 1712.140 25.510 ;
        RECT 1711.930 0.000 1712.210 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1560.645 25.245 1560.815 28.475 ;
        RECT 1562.485 25.925 1562.655 28.475 ;
      LAYER mcon ;
        RECT 1560.645 28.305 1560.815 28.475 ;
        RECT 1562.485 28.305 1562.655 28.475 ;
      LAYER met1 ;
        RECT 1560.585 28.460 1560.875 28.505 ;
        RECT 1562.425 28.460 1562.715 28.505 ;
        RECT 1560.585 28.320 1562.715 28.460 ;
        RECT 1560.585 28.275 1560.875 28.320 ;
        RECT 1562.425 28.275 1562.715 28.320 ;
        RECT 1562.425 26.080 1562.715 26.125 ;
        RECT 1729.850 26.080 1730.170 26.140 ;
        RECT 1562.425 25.940 1730.170 26.080 ;
        RECT 1562.425 25.895 1562.715 25.940 ;
        RECT 1729.850 25.880 1730.170 25.940 ;
        RECT 1513.190 25.400 1513.510 25.460 ;
        RECT 1560.585 25.400 1560.875 25.445 ;
        RECT 1513.190 25.260 1560.875 25.400 ;
        RECT 1513.190 25.200 1513.510 25.260 ;
        RECT 1560.585 25.215 1560.875 25.260 ;
      LAYER via ;
        RECT 1729.880 25.880 1730.140 26.140 ;
        RECT 1513.220 25.200 1513.480 25.460 ;
      LAYER met2 ;
        RECT 1513.280 25.490 1513.420 54.000 ;
        RECT 1729.880 25.850 1730.140 26.170 ;
        RECT 1513.220 25.170 1513.480 25.490 ;
        RECT 1729.940 2.400 1730.080 25.850 ;
        RECT 1729.870 0.000 1730.150 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1608.945 31.025 1609.115 34.595 ;
      LAYER mcon ;
        RECT 1608.945 34.425 1609.115 34.595 ;
      LAYER met1 ;
        RECT 1608.885 34.580 1609.175 34.625 ;
        RECT 1611.170 34.580 1611.490 34.640 ;
        RECT 1608.885 34.440 1611.490 34.580 ;
        RECT 1608.885 34.395 1609.175 34.440 ;
        RECT 1611.170 34.380 1611.490 34.440 ;
        RECT 1512.270 31.180 1512.590 31.240 ;
        RECT 1608.885 31.180 1609.175 31.225 ;
        RECT 1512.270 31.040 1609.175 31.180 ;
        RECT 1512.270 30.980 1512.590 31.040 ;
        RECT 1608.885 30.995 1609.175 31.040 ;
      LAYER via ;
        RECT 1611.200 34.380 1611.460 34.640 ;
        RECT 1512.300 30.980 1512.560 31.240 ;
      LAYER met2 ;
        RECT 1512.360 31.270 1512.500 54.000 ;
        RECT 1611.200 34.350 1611.460 34.670 ;
        RECT 1611.260 31.805 1611.400 34.350 ;
        RECT 1611.190 31.435 1611.470 31.805 ;
        RECT 1747.810 31.435 1748.090 31.805 ;
        RECT 1512.300 30.950 1512.560 31.270 ;
        RECT 1747.880 2.400 1748.020 31.435 ;
        RECT 1747.810 0.000 1748.090 2.400 ;
      LAYER via2 ;
        RECT 1611.190 31.480 1611.470 31.760 ;
        RECT 1747.810 31.480 1748.090 31.760 ;
      LAYER met3 ;
        RECT 1611.165 31.770 1611.495 31.785 ;
        RECT 1747.785 31.770 1748.115 31.785 ;
        RECT 1611.165 31.470 1748.115 31.770 ;
        RECT 1611.165 31.455 1611.495 31.470 ;
        RECT 1747.785 31.455 1748.115 31.470 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1519.630 44.780 1519.950 44.840 ;
        RECT 1755.150 44.780 1755.470 44.840 ;
        RECT 1519.630 44.640 1755.470 44.780 ;
        RECT 1519.630 44.580 1519.950 44.640 ;
        RECT 1755.150 44.580 1755.470 44.640 ;
        RECT 1755.610 41.720 1755.930 41.780 ;
        RECT 1765.270 41.720 1765.590 41.780 ;
        RECT 1755.610 41.580 1765.590 41.720 ;
        RECT 1755.610 41.520 1755.930 41.580 ;
        RECT 1765.270 41.520 1765.590 41.580 ;
      LAYER via ;
        RECT 1519.660 44.580 1519.920 44.840 ;
        RECT 1755.180 44.580 1755.440 44.840 ;
        RECT 1755.640 41.520 1755.900 41.780 ;
        RECT 1765.300 41.520 1765.560 41.780 ;
      LAYER met2 ;
        RECT 1519.720 44.870 1519.860 54.000 ;
        RECT 1519.660 44.550 1519.920 44.870 ;
        RECT 1755.180 44.610 1755.440 44.870 ;
        RECT 1755.180 44.550 1755.840 44.610 ;
        RECT 1755.240 44.470 1755.840 44.550 ;
        RECT 1755.700 41.810 1755.840 44.470 ;
        RECT 1755.640 41.490 1755.900 41.810 ;
        RECT 1765.300 41.490 1765.560 41.810 ;
        RECT 1765.360 2.400 1765.500 41.490 ;
        RECT 1765.290 0.000 1765.570 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1518.710 45.120 1519.030 45.180 ;
        RECT 1756.070 45.120 1756.390 45.180 ;
        RECT 1518.710 44.980 1756.390 45.120 ;
        RECT 1518.710 44.920 1519.030 44.980 ;
        RECT 1756.070 44.920 1756.390 44.980 ;
      LAYER via ;
        RECT 1518.740 44.920 1519.000 45.180 ;
        RECT 1756.100 44.920 1756.360 45.180 ;
      LAYER met2 ;
        RECT 1518.800 45.210 1518.940 54.000 ;
        RECT 1518.740 44.890 1519.000 45.210 ;
        RECT 1756.090 45.035 1756.370 45.405 ;
        RECT 1783.230 45.035 1783.510 45.405 ;
        RECT 1756.100 44.890 1756.360 45.035 ;
        RECT 1783.300 2.400 1783.440 45.035 ;
        RECT 1783.230 0.000 1783.510 2.400 ;
      LAYER via2 ;
        RECT 1756.090 45.080 1756.370 45.360 ;
        RECT 1783.230 45.080 1783.510 45.360 ;
      LAYER met3 ;
        RECT 1756.065 45.370 1756.395 45.385 ;
        RECT 1783.205 45.370 1783.535 45.385 ;
        RECT 1756.065 45.070 1783.535 45.370 ;
        RECT 1756.065 45.055 1756.395 45.070 ;
        RECT 1783.205 45.055 1783.535 45.070 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1526.530 41.720 1526.850 41.780 ;
        RECT 1755.150 41.720 1755.470 41.780 ;
        RECT 1526.530 41.580 1755.470 41.720 ;
        RECT 1526.530 41.520 1526.850 41.580 ;
        RECT 1755.150 41.520 1755.470 41.580 ;
      LAYER via ;
        RECT 1526.560 41.520 1526.820 41.780 ;
        RECT 1755.180 41.520 1755.440 41.780 ;
      LAYER met2 ;
        RECT 1526.620 41.810 1526.760 54.000 ;
        RECT 1526.560 41.490 1526.820 41.810 ;
        RECT 1755.170 41.635 1755.450 42.005 ;
        RECT 1801.170 41.635 1801.450 42.005 ;
        RECT 1755.180 41.490 1755.440 41.635 ;
        RECT 1801.240 2.400 1801.380 41.635 ;
        RECT 1801.170 0.000 1801.450 2.400 ;
      LAYER via2 ;
        RECT 1755.170 41.680 1755.450 41.960 ;
        RECT 1801.170 41.680 1801.450 41.960 ;
      LAYER met3 ;
        RECT 1755.145 41.970 1755.475 41.985 ;
        RECT 1801.145 41.970 1801.475 41.985 ;
        RECT 1755.145 41.670 1801.475 41.970 ;
        RECT 1755.145 41.655 1755.475 41.670 ;
        RECT 1801.145 41.655 1801.475 41.670 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1777.765 42.245 1778.855 42.415 ;
        RECT 1777.765 41.905 1777.935 42.245 ;
      LAYER mcon ;
        RECT 1778.685 42.245 1778.855 42.415 ;
      LAYER met1 ;
        RECT 1525.150 48.520 1525.470 48.580 ;
        RECT 1525.610 48.520 1525.930 48.580 ;
        RECT 1525.150 48.380 1525.930 48.520 ;
        RECT 1525.150 48.320 1525.470 48.380 ;
        RECT 1525.610 48.320 1525.930 48.380 ;
        RECT 1778.625 42.400 1778.915 42.445 ;
        RECT 1819.090 42.400 1819.410 42.460 ;
        RECT 1778.625 42.260 1819.410 42.400 ;
        RECT 1778.625 42.215 1778.915 42.260 ;
        RECT 1819.090 42.200 1819.410 42.260 ;
        RECT 1525.150 42.060 1525.470 42.120 ;
        RECT 1777.705 42.060 1777.995 42.105 ;
        RECT 1525.150 41.920 1777.995 42.060 ;
        RECT 1525.150 41.860 1525.470 41.920 ;
        RECT 1777.705 41.875 1777.995 41.920 ;
      LAYER via ;
        RECT 1525.180 48.320 1525.440 48.580 ;
        RECT 1525.640 48.320 1525.900 48.580 ;
        RECT 1819.120 42.200 1819.380 42.460 ;
        RECT 1525.180 41.860 1525.440 42.120 ;
      LAYER met2 ;
        RECT 1525.700 48.610 1525.840 54.000 ;
        RECT 1525.180 48.290 1525.440 48.610 ;
        RECT 1525.640 48.290 1525.900 48.610 ;
        RECT 1525.240 42.150 1525.380 48.290 ;
        RECT 1819.120 42.170 1819.380 42.490 ;
        RECT 1525.180 41.830 1525.440 42.150 ;
        RECT 1819.180 2.400 1819.320 42.170 ;
        RECT 1819.110 0.000 1819.390 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1533.430 42.400 1533.750 42.460 ;
        RECT 1819.550 42.400 1819.870 42.460 ;
        RECT 1837.030 42.400 1837.350 42.460 ;
        RECT 1533.430 42.260 1778.380 42.400 ;
        RECT 1533.430 42.200 1533.750 42.260 ;
        RECT 1778.240 41.720 1778.380 42.260 ;
        RECT 1819.550 42.260 1837.350 42.400 ;
        RECT 1819.550 42.200 1819.870 42.260 ;
        RECT 1837.030 42.200 1837.350 42.260 ;
        RECT 1805.750 41.720 1806.070 41.780 ;
        RECT 1778.240 41.580 1806.070 41.720 ;
        RECT 1805.750 41.520 1806.070 41.580 ;
      LAYER via ;
        RECT 1533.460 42.200 1533.720 42.460 ;
        RECT 1819.580 42.200 1819.840 42.460 ;
        RECT 1837.060 42.200 1837.320 42.460 ;
        RECT 1805.780 41.520 1806.040 41.780 ;
      LAYER met2 ;
        RECT 1533.520 42.490 1533.660 54.000 ;
        RECT 1533.460 42.170 1533.720 42.490 ;
        RECT 1819.580 42.170 1819.840 42.490 ;
        RECT 1837.060 42.170 1837.320 42.490 ;
        RECT 1819.640 42.005 1819.780 42.170 ;
        RECT 1805.770 41.635 1806.050 42.005 ;
        RECT 1819.570 41.635 1819.850 42.005 ;
        RECT 1805.780 41.490 1806.040 41.635 ;
        RECT 1837.120 2.400 1837.260 42.170 ;
        RECT 1837.050 0.000 1837.330 2.400 ;
      LAYER via2 ;
        RECT 1805.770 41.680 1806.050 41.960 ;
        RECT 1819.570 41.680 1819.850 41.960 ;
      LAYER met3 ;
        RECT 1805.745 41.970 1806.075 41.985 ;
        RECT 1819.545 41.970 1819.875 41.985 ;
        RECT 1805.745 41.670 1819.875 41.970 ;
        RECT 1805.745 41.655 1806.075 41.670 ;
        RECT 1819.545 41.655 1819.875 41.670 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1532.050 42.740 1532.370 42.800 ;
        RECT 1854.050 42.740 1854.370 42.800 ;
        RECT 1532.050 42.600 1854.370 42.740 ;
        RECT 1532.050 42.540 1532.370 42.600 ;
        RECT 1854.050 42.540 1854.370 42.600 ;
      LAYER via ;
        RECT 1532.080 42.540 1532.340 42.800 ;
        RECT 1854.080 42.540 1854.340 42.800 ;
      LAYER met2 ;
        RECT 1532.140 42.830 1532.280 54.000 ;
        RECT 1532.080 42.510 1532.340 42.830 ;
        RECT 1854.080 42.510 1854.340 42.830 ;
        RECT 1854.140 24.890 1854.280 42.510 ;
        RECT 1854.140 24.750 1854.740 24.890 ;
        RECT 1854.600 2.400 1854.740 24.750 ;
        RECT 1854.530 0.000 1854.810 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1539.870 43.080 1540.190 43.140 ;
        RECT 1872.910 43.080 1873.230 43.140 ;
        RECT 1539.870 42.940 1873.230 43.080 ;
        RECT 1539.870 42.880 1540.190 42.940 ;
        RECT 1872.910 42.880 1873.230 42.940 ;
      LAYER via ;
        RECT 1539.900 42.880 1540.160 43.140 ;
        RECT 1872.940 42.880 1873.200 43.140 ;
      LAYER met2 ;
        RECT 1539.960 43.170 1540.100 54.000 ;
        RECT 1539.900 42.850 1540.160 43.170 ;
        RECT 1872.940 42.850 1873.200 43.170 ;
        RECT 1873.000 41.210 1873.140 42.850 ;
        RECT 1872.540 41.070 1873.140 41.210 ;
        RECT 1872.540 2.400 1872.680 41.070 ;
        RECT 1872.470 0.000 1872.750 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 748.670 37.300 748.990 37.360 ;
        RECT 1300.210 37.300 1300.530 37.360 ;
        RECT 748.670 37.160 1300.530 37.300 ;
        RECT 748.670 37.100 748.990 37.160 ;
        RECT 1300.210 37.100 1300.530 37.160 ;
      LAYER via ;
        RECT 748.700 37.100 748.960 37.360 ;
        RECT 1300.240 37.100 1300.500 37.360 ;
      LAYER met2 ;
        RECT 1300.300 37.390 1300.440 54.000 ;
        RECT 748.700 37.070 748.960 37.390 ;
        RECT 1300.240 37.070 1300.500 37.390 ;
        RECT 748.760 2.400 748.900 37.070 ;
        RECT 748.690 0.000 748.970 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1540.330 44.100 1540.650 44.160 ;
        RECT 1890.390 44.100 1890.710 44.160 ;
        RECT 1540.330 43.960 1890.710 44.100 ;
        RECT 1540.330 43.900 1540.650 43.960 ;
        RECT 1890.390 43.900 1890.710 43.960 ;
      LAYER via ;
        RECT 1540.360 43.900 1540.620 44.160 ;
        RECT 1890.420 43.900 1890.680 44.160 ;
      LAYER met2 ;
        RECT 1540.420 44.190 1540.560 54.000 ;
        RECT 1540.360 43.870 1540.620 44.190 ;
        RECT 1890.420 43.870 1890.680 44.190 ;
        RECT 1890.480 2.400 1890.620 43.870 ;
        RECT 1890.410 0.000 1890.690 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1546.310 44.440 1546.630 44.500 ;
        RECT 1908.330 44.440 1908.650 44.500 ;
        RECT 1546.310 44.300 1908.650 44.440 ;
        RECT 1546.310 44.240 1546.630 44.300 ;
        RECT 1908.330 44.240 1908.650 44.300 ;
      LAYER via ;
        RECT 1546.340 44.240 1546.600 44.500 ;
        RECT 1908.360 44.240 1908.620 44.500 ;
      LAYER met2 ;
        RECT 1546.400 44.530 1546.540 54.000 ;
        RECT 1546.340 44.210 1546.600 44.530 ;
        RECT 1908.360 44.210 1908.620 44.530 ;
        RECT 1908.420 2.400 1908.560 44.210 ;
        RECT 1908.350 0.000 1908.630 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1545.850 48.180 1546.170 48.240 ;
        RECT 1925.810 48.180 1926.130 48.240 ;
        RECT 1545.850 48.040 1926.130 48.180 ;
        RECT 1545.850 47.980 1546.170 48.040 ;
        RECT 1925.810 47.980 1926.130 48.040 ;
      LAYER via ;
        RECT 1545.880 47.980 1546.140 48.240 ;
        RECT 1925.840 47.980 1926.100 48.240 ;
      LAYER met2 ;
        RECT 1545.940 48.270 1546.080 54.000 ;
        RECT 1545.880 47.950 1546.140 48.270 ;
        RECT 1925.840 47.950 1926.100 48.270 ;
        RECT 1925.900 2.400 1926.040 47.950 ;
        RECT 1925.830 0.000 1926.110 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1553.210 47.840 1553.530 47.900 ;
        RECT 1943.750 47.840 1944.070 47.900 ;
        RECT 1553.210 47.700 1944.070 47.840 ;
        RECT 1553.210 47.640 1553.530 47.700 ;
        RECT 1943.750 47.640 1944.070 47.700 ;
      LAYER via ;
        RECT 1553.240 47.640 1553.500 47.900 ;
        RECT 1943.780 47.640 1944.040 47.900 ;
      LAYER met2 ;
        RECT 1553.300 47.930 1553.440 54.000 ;
        RECT 1553.240 47.610 1553.500 47.930 ;
        RECT 1943.780 47.610 1944.040 47.930 ;
        RECT 1943.840 2.400 1943.980 47.610 ;
        RECT 1943.770 0.000 1944.050 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1560.110 47.500 1560.430 47.560 ;
        RECT 1961.690 47.500 1962.010 47.560 ;
        RECT 1560.110 47.360 1962.010 47.500 ;
        RECT 1560.110 47.300 1560.430 47.360 ;
        RECT 1961.690 47.300 1962.010 47.360 ;
      LAYER via ;
        RECT 1560.140 47.300 1560.400 47.560 ;
        RECT 1961.720 47.300 1961.980 47.560 ;
      LAYER met2 ;
        RECT 1560.200 47.590 1560.340 54.000 ;
        RECT 1560.140 47.270 1560.400 47.590 ;
        RECT 1961.720 47.270 1961.980 47.590 ;
        RECT 1961.780 2.400 1961.920 47.270 ;
        RECT 1961.710 0.000 1961.990 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1975.950 2.960 1976.270 3.020 ;
        RECT 1979.630 2.960 1979.950 3.020 ;
        RECT 1975.950 2.820 1979.950 2.960 ;
        RECT 1975.950 2.760 1976.270 2.820 ;
        RECT 1979.630 2.760 1979.950 2.820 ;
      LAYER via ;
        RECT 1975.980 2.760 1976.240 3.020 ;
        RECT 1979.660 2.760 1979.920 3.020 ;
      LAYER met2 ;
        RECT 1976.040 3.050 1976.180 54.000 ;
        RECT 1975.980 2.730 1976.240 3.050 ;
        RECT 1979.660 2.730 1979.920 3.050 ;
        RECT 1979.720 2.400 1979.860 2.730 ;
        RECT 1979.650 0.000 1979.930 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1996.740 3.130 1996.880 54.000 ;
        RECT 1996.740 2.990 1997.800 3.130 ;
        RECT 1997.660 2.400 1997.800 2.990 ;
        RECT 1997.590 0.000 1997.870 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2010.450 2.960 2010.770 3.020 ;
        RECT 2015.050 2.960 2015.370 3.020 ;
        RECT 2010.450 2.820 2015.370 2.960 ;
        RECT 2010.450 2.760 2010.770 2.820 ;
        RECT 2015.050 2.760 2015.370 2.820 ;
      LAYER via ;
        RECT 2010.480 2.760 2010.740 3.020 ;
        RECT 2015.080 2.760 2015.340 3.020 ;
      LAYER met2 ;
        RECT 2010.540 3.050 2010.680 54.000 ;
        RECT 2010.480 2.730 2010.740 3.050 ;
        RECT 2015.080 2.730 2015.340 3.050 ;
        RECT 2015.140 2.400 2015.280 2.730 ;
        RECT 2015.070 0.000 2015.350 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2031.150 2.960 2031.470 3.020 ;
        RECT 2032.990 2.960 2033.310 3.020 ;
        RECT 2031.150 2.820 2033.310 2.960 ;
        RECT 2031.150 2.760 2031.470 2.820 ;
        RECT 2032.990 2.760 2033.310 2.820 ;
      LAYER via ;
        RECT 2031.180 2.760 2031.440 3.020 ;
        RECT 2033.020 2.760 2033.280 3.020 ;
      LAYER met2 ;
        RECT 2031.240 3.050 2031.380 54.000 ;
        RECT 2031.180 2.730 2031.440 3.050 ;
        RECT 2033.020 2.730 2033.280 3.050 ;
        RECT 2033.080 2.400 2033.220 2.730 ;
        RECT 2033.010 0.000 2033.290 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2051.020 2.400 2051.160 54.000 ;
        RECT 2050.950 0.000 2051.230 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 766.150 36.960 766.470 37.020 ;
        RECT 1308.950 36.960 1309.270 37.020 ;
        RECT 766.150 36.820 1309.270 36.960 ;
        RECT 766.150 36.760 766.470 36.820 ;
        RECT 1308.950 36.760 1309.270 36.820 ;
      LAYER via ;
        RECT 766.180 36.760 766.440 37.020 ;
        RECT 1308.980 36.760 1309.240 37.020 ;
      LAYER met2 ;
        RECT 1309.040 37.050 1309.180 54.000 ;
        RECT 766.180 36.730 766.440 37.050 ;
        RECT 1308.980 36.730 1309.240 37.050 ;
        RECT 766.240 2.400 766.380 36.730 ;
        RECT 766.170 0.000 766.450 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2066.200 48.805 2066.340 54.000 ;
        RECT 2066.130 48.435 2066.410 48.805 ;
        RECT 2068.890 48.435 2069.170 48.805 ;
        RECT 2068.960 2.400 2069.100 48.435 ;
        RECT 2068.890 0.000 2069.170 2.400 ;
      LAYER via2 ;
        RECT 2066.130 48.480 2066.410 48.760 ;
        RECT 2068.890 48.480 2069.170 48.760 ;
      LAYER met3 ;
        RECT 2066.105 48.770 2066.435 48.785 ;
        RECT 2068.865 48.770 2069.195 48.785 ;
        RECT 2066.105 48.470 2069.195 48.770 ;
        RECT 2066.105 48.455 2066.435 48.470 ;
        RECT 2068.865 48.455 2069.195 48.470 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2086.900 2.400 2087.040 54.000 ;
        RECT 2086.830 0.000 2087.110 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2104.365 2.805 2104.535 14.195 ;
      LAYER mcon ;
        RECT 2104.365 14.025 2104.535 14.195 ;
      LAYER met1 ;
        RECT 2100.150 14.180 2100.470 14.240 ;
        RECT 2104.305 14.180 2104.595 14.225 ;
        RECT 2100.150 14.040 2104.595 14.180 ;
        RECT 2100.150 13.980 2100.470 14.040 ;
        RECT 2104.305 13.995 2104.595 14.040 ;
        RECT 2104.290 2.960 2104.610 3.020 ;
        RECT 2104.095 2.820 2104.610 2.960 ;
        RECT 2104.290 2.760 2104.610 2.820 ;
      LAYER via ;
        RECT 2100.180 13.980 2100.440 14.240 ;
        RECT 2104.320 2.760 2104.580 3.020 ;
      LAYER met2 ;
        RECT 2100.240 14.270 2100.380 54.000 ;
        RECT 2100.180 13.950 2100.440 14.270 ;
        RECT 2104.320 2.730 2104.580 3.050 ;
        RECT 2104.380 2.400 2104.520 2.730 ;
        RECT 2104.310 0.000 2104.590 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1587.710 52.600 1588.030 52.660 ;
        RECT 2044.950 52.600 2045.270 52.660 ;
        RECT 1587.710 52.460 2045.270 52.600 ;
        RECT 1587.710 52.400 1588.030 52.460 ;
        RECT 2044.950 52.400 2045.270 52.460 ;
        RECT 2120.850 2.960 2121.170 3.020 ;
        RECT 2122.230 2.960 2122.550 3.020 ;
        RECT 2120.850 2.820 2122.550 2.960 ;
        RECT 2120.850 2.760 2121.170 2.820 ;
        RECT 2122.230 2.760 2122.550 2.820 ;
      LAYER via ;
        RECT 1587.740 52.400 1588.000 52.660 ;
        RECT 2044.980 52.400 2045.240 52.660 ;
        RECT 2120.880 2.760 2121.140 3.020 ;
        RECT 2122.260 2.760 2122.520 3.020 ;
      LAYER met2 ;
        RECT 1587.800 52.690 1587.940 54.000 ;
        RECT 1587.740 52.370 1588.000 52.690 ;
        RECT 2044.970 52.515 2045.250 52.885 ;
        RECT 2120.870 52.515 2121.150 52.885 ;
        RECT 2044.980 52.370 2045.240 52.515 ;
        RECT 2120.940 3.050 2121.080 52.515 ;
        RECT 2120.880 2.730 2121.140 3.050 ;
        RECT 2122.260 2.730 2122.520 3.050 ;
        RECT 2122.320 2.400 2122.460 2.730 ;
        RECT 2122.250 0.000 2122.530 2.400 ;
      LAYER via2 ;
        RECT 2044.970 52.560 2045.250 52.840 ;
        RECT 2120.870 52.560 2121.150 52.840 ;
      LAYER met3 ;
        RECT 2044.945 52.850 2045.275 52.865 ;
        RECT 2120.845 52.850 2121.175 52.865 ;
        RECT 2044.945 52.550 2121.175 52.850 ;
        RECT 2044.945 52.535 2045.275 52.550 ;
        RECT 2120.845 52.535 2121.175 52.550 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2093.325 52.615 2093.495 52.955 ;
        RECT 2093.325 52.445 2093.955 52.615 ;
        RECT 2093.785 47.685 2093.955 52.445 ;
      LAYER mcon ;
        RECT 2093.325 52.785 2093.495 52.955 ;
      LAYER met1 ;
        RECT 1594.150 52.940 1594.470 53.000 ;
        RECT 2093.265 52.940 2093.555 52.985 ;
        RECT 1594.150 52.800 2093.555 52.940 ;
        RECT 1594.150 52.740 1594.470 52.800 ;
        RECT 2093.265 52.755 2093.555 52.800 ;
        RECT 2093.725 47.840 2094.015 47.885 ;
        RECT 2134.650 47.840 2134.970 47.900 ;
        RECT 2093.725 47.700 2134.970 47.840 ;
        RECT 2093.725 47.655 2094.015 47.700 ;
        RECT 2134.650 47.640 2134.970 47.700 ;
        RECT 2134.650 2.960 2134.970 3.020 ;
        RECT 2140.170 2.960 2140.490 3.020 ;
        RECT 2134.650 2.820 2140.490 2.960 ;
        RECT 2134.650 2.760 2134.970 2.820 ;
        RECT 2140.170 2.760 2140.490 2.820 ;
      LAYER via ;
        RECT 1594.180 52.740 1594.440 53.000 ;
        RECT 2134.680 47.640 2134.940 47.900 ;
        RECT 2134.680 2.760 2134.940 3.020 ;
        RECT 2140.200 2.760 2140.460 3.020 ;
      LAYER met2 ;
        RECT 1594.240 53.030 1594.380 54.000 ;
        RECT 1594.180 52.710 1594.440 53.030 ;
        RECT 2134.680 47.610 2134.940 47.930 ;
        RECT 2134.740 3.050 2134.880 47.610 ;
        RECT 2134.680 2.730 2134.940 3.050 ;
        RECT 2140.200 2.730 2140.460 3.050 ;
        RECT 2140.260 2.400 2140.400 2.730 ;
        RECT 2140.190 0.000 2140.470 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2093.325 48.025 2093.495 52.275 ;
      LAYER mcon ;
        RECT 2093.325 52.105 2093.495 52.275 ;
      LAYER met1 ;
        RECT 1593.230 52.260 1593.550 52.320 ;
        RECT 2093.265 52.260 2093.555 52.305 ;
        RECT 1593.230 52.120 2093.555 52.260 ;
        RECT 1593.230 52.060 1593.550 52.120 ;
        RECT 2093.265 52.075 2093.555 52.120 ;
        RECT 2093.265 48.180 2093.555 48.225 ;
        RECT 2155.350 48.180 2155.670 48.240 ;
        RECT 2093.265 48.040 2155.670 48.180 ;
        RECT 2093.265 47.995 2093.555 48.040 ;
        RECT 2155.350 47.980 2155.670 48.040 ;
        RECT 2155.350 2.960 2155.670 3.020 ;
        RECT 2158.110 2.960 2158.430 3.020 ;
        RECT 2155.350 2.820 2158.430 2.960 ;
        RECT 2155.350 2.760 2155.670 2.820 ;
        RECT 2158.110 2.760 2158.430 2.820 ;
      LAYER via ;
        RECT 1593.260 52.060 1593.520 52.320 ;
        RECT 2155.380 47.980 2155.640 48.240 ;
        RECT 2155.380 2.760 2155.640 3.020 ;
        RECT 2158.140 2.760 2158.400 3.020 ;
      LAYER met2 ;
        RECT 1593.320 52.350 1593.460 54.000 ;
        RECT 1593.260 52.030 1593.520 52.350 ;
        RECT 2155.380 47.950 2155.640 48.270 ;
        RECT 2155.440 3.050 2155.580 47.950 ;
        RECT 2155.380 2.730 2155.640 3.050 ;
        RECT 2158.140 2.730 2158.400 3.050 ;
        RECT 2158.200 2.400 2158.340 2.730 ;
        RECT 2158.130 0.000 2158.410 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2141.625 47.345 2141.795 48.535 ;
      LAYER mcon ;
        RECT 2141.625 48.365 2141.795 48.535 ;
      LAYER met1 ;
        RECT 1600.590 48.520 1600.910 48.580 ;
        RECT 2141.565 48.520 2141.855 48.565 ;
        RECT 2175.590 48.520 2175.910 48.580 ;
        RECT 1600.590 48.380 2141.855 48.520 ;
        RECT 1600.590 48.320 1600.910 48.380 ;
        RECT 2141.565 48.335 2141.855 48.380 ;
        RECT 2156.360 48.380 2175.910 48.520 ;
        RECT 2141.565 47.500 2141.855 47.545 ;
        RECT 2156.360 47.500 2156.500 48.380 ;
        RECT 2175.590 48.320 2175.910 48.380 ;
        RECT 2141.565 47.360 2156.500 47.500 ;
        RECT 2141.565 47.315 2141.855 47.360 ;
      LAYER via ;
        RECT 1600.620 48.320 1600.880 48.580 ;
        RECT 2175.620 48.320 2175.880 48.580 ;
      LAYER met2 ;
        RECT 1600.680 48.610 1600.820 54.000 ;
        RECT 1600.620 48.290 1600.880 48.610 ;
        RECT 2175.620 48.290 2175.880 48.610 ;
        RECT 2175.680 2.400 2175.820 48.290 ;
        RECT 2175.610 0.000 2175.890 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1601.050 49.540 1601.370 49.600 ;
        RECT 2189.850 49.540 2190.170 49.600 ;
        RECT 1601.050 49.400 2190.170 49.540 ;
        RECT 1601.050 49.340 1601.370 49.400 ;
        RECT 2189.850 49.340 2190.170 49.400 ;
      LAYER via ;
        RECT 1601.080 49.340 1601.340 49.600 ;
        RECT 2189.880 49.340 2190.140 49.600 ;
      LAYER met2 ;
        RECT 1601.140 49.630 1601.280 54.000 ;
        RECT 1601.080 49.310 1601.340 49.630 ;
        RECT 2189.880 49.310 2190.140 49.630 ;
        RECT 2189.940 3.130 2190.080 49.310 ;
        RECT 2189.940 2.990 2193.300 3.130 ;
        RECT 2193.160 2.960 2193.300 2.990 ;
        RECT 2193.160 2.820 2193.760 2.960 ;
        RECT 2193.620 2.400 2193.760 2.820 ;
        RECT 2193.550 0.000 2193.830 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1608.870 49.880 1609.190 49.940 ;
        RECT 2210.550 49.880 2210.870 49.940 ;
        RECT 1608.870 49.740 2210.870 49.880 ;
        RECT 1608.870 49.680 1609.190 49.740 ;
        RECT 2210.550 49.680 2210.870 49.740 ;
        RECT 2210.550 2.960 2210.870 3.020 ;
        RECT 2211.470 2.960 2211.790 3.020 ;
        RECT 2210.550 2.820 2211.790 2.960 ;
        RECT 2210.550 2.760 2210.870 2.820 ;
        RECT 2211.470 2.760 2211.790 2.820 ;
      LAYER via ;
        RECT 1608.900 49.680 1609.160 49.940 ;
        RECT 2210.580 49.680 2210.840 49.940 ;
        RECT 2210.580 2.760 2210.840 3.020 ;
        RECT 2211.500 2.760 2211.760 3.020 ;
      LAYER met2 ;
        RECT 1608.960 49.970 1609.100 54.000 ;
        RECT 1608.900 49.650 1609.160 49.970 ;
        RECT 2210.580 49.650 2210.840 49.970 ;
        RECT 2210.640 3.050 2210.780 49.650 ;
        RECT 2210.580 2.730 2210.840 3.050 ;
        RECT 2211.500 2.730 2211.760 3.050 ;
        RECT 2211.560 2.400 2211.700 2.730 ;
        RECT 2211.490 0.000 2211.770 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1615.310 53.620 1615.630 53.680 ;
        RECT 1641.990 53.620 1642.310 53.680 ;
        RECT 1615.310 53.480 1642.310 53.620 ;
        RECT 1615.310 53.420 1615.630 53.480 ;
        RECT 1641.990 53.420 1642.310 53.480 ;
        RECT 1658.090 50.220 1658.410 50.280 ;
        RECT 2224.350 50.220 2224.670 50.280 ;
        RECT 1658.090 50.080 2224.670 50.220 ;
        RECT 1658.090 50.020 1658.410 50.080 ;
        RECT 2224.350 50.020 2224.670 50.080 ;
        RECT 2224.350 2.960 2224.670 3.020 ;
        RECT 2229.410 2.960 2229.730 3.020 ;
        RECT 2224.350 2.820 2229.730 2.960 ;
        RECT 2224.350 2.760 2224.670 2.820 ;
        RECT 2229.410 2.760 2229.730 2.820 ;
      LAYER via ;
        RECT 1615.340 53.420 1615.600 53.680 ;
        RECT 1642.020 53.420 1642.280 53.680 ;
        RECT 1658.120 50.020 1658.380 50.280 ;
        RECT 2224.380 50.020 2224.640 50.280 ;
        RECT 2224.380 2.760 2224.640 3.020 ;
        RECT 2229.440 2.760 2229.700 3.020 ;
      LAYER met2 ;
        RECT 1615.400 53.710 1615.540 54.000 ;
        RECT 1615.340 53.390 1615.600 53.710 ;
        RECT 1642.020 53.390 1642.280 53.710 ;
        RECT 1642.080 50.165 1642.220 53.390 ;
        RECT 1658.120 50.165 1658.380 50.310 ;
        RECT 1642.010 49.795 1642.290 50.165 ;
        RECT 1658.110 49.795 1658.390 50.165 ;
        RECT 2224.380 49.990 2224.640 50.310 ;
        RECT 2224.440 3.050 2224.580 49.990 ;
        RECT 2224.380 2.730 2224.640 3.050 ;
        RECT 2229.440 2.730 2229.700 3.050 ;
        RECT 2229.500 2.400 2229.640 2.730 ;
        RECT 2229.430 0.000 2229.710 2.400 ;
      LAYER via2 ;
        RECT 1642.010 49.840 1642.290 50.120 ;
        RECT 1658.110 49.840 1658.390 50.120 ;
      LAYER met3 ;
        RECT 1641.985 50.130 1642.315 50.145 ;
        RECT 1658.085 50.130 1658.415 50.145 ;
        RECT 1641.985 49.830 1658.415 50.130 ;
        RECT 1641.985 49.815 1642.315 49.830 ;
        RECT 1658.085 49.815 1658.415 49.830 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 784.090 36.620 784.410 36.680 ;
        RECT 1308.490 36.620 1308.810 36.680 ;
        RECT 784.090 36.480 1308.810 36.620 ;
        RECT 784.090 36.420 784.410 36.480 ;
        RECT 1308.490 36.420 1308.810 36.480 ;
      LAYER via ;
        RECT 784.120 36.420 784.380 36.680 ;
        RECT 1308.520 36.420 1308.780 36.680 ;
      LAYER met2 ;
        RECT 1308.580 36.710 1308.720 54.000 ;
        RECT 784.120 36.390 784.380 36.710 ;
        RECT 1308.520 36.390 1308.780 36.710 ;
        RECT 784.180 2.400 784.320 36.390 ;
        RECT 784.110 0.000 784.390 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1656.710 50.560 1657.030 50.620 ;
        RECT 2245.050 50.560 2245.370 50.620 ;
        RECT 1656.710 50.420 2245.370 50.560 ;
        RECT 1656.710 50.360 1657.030 50.420 ;
        RECT 2245.050 50.360 2245.370 50.420 ;
        RECT 2245.050 2.960 2245.370 3.020 ;
        RECT 2247.350 2.960 2247.670 3.020 ;
        RECT 2245.050 2.820 2247.670 2.960 ;
        RECT 2245.050 2.760 2245.370 2.820 ;
        RECT 2247.350 2.760 2247.670 2.820 ;
      LAYER via ;
        RECT 1656.740 50.360 1657.000 50.620 ;
        RECT 2245.080 50.360 2245.340 50.620 ;
        RECT 2245.080 2.760 2245.340 3.020 ;
        RECT 2247.380 2.760 2247.640 3.020 ;
      LAYER met2 ;
        RECT 1656.800 50.650 1656.940 54.000 ;
        RECT 1656.740 50.330 1657.000 50.650 ;
        RECT 2245.080 50.330 2245.340 50.650 ;
        RECT 2245.140 3.050 2245.280 50.330 ;
        RECT 2245.080 2.730 2245.340 3.050 ;
        RECT 2247.380 2.730 2247.640 3.050 ;
        RECT 2247.440 2.400 2247.580 2.730 ;
        RECT 2247.370 0.000 2247.650 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1622.210 53.280 1622.530 53.340 ;
        RECT 1649.350 53.280 1649.670 53.340 ;
        RECT 1622.210 53.140 1649.670 53.280 ;
        RECT 1622.210 53.080 1622.530 53.140 ;
        RECT 1649.350 53.080 1649.670 53.140 ;
        RECT 1658.090 50.900 1658.410 50.960 ;
        RECT 2259.310 50.900 2259.630 50.960 ;
        RECT 1658.090 50.760 2259.630 50.900 ;
        RECT 1658.090 50.700 1658.410 50.760 ;
        RECT 2259.310 50.700 2259.630 50.760 ;
        RECT 2259.310 2.960 2259.630 3.020 ;
        RECT 2264.830 2.960 2265.150 3.020 ;
        RECT 2259.310 2.820 2265.150 2.960 ;
        RECT 2259.310 2.760 2259.630 2.820 ;
        RECT 2264.830 2.760 2265.150 2.820 ;
      LAYER via ;
        RECT 1622.240 53.080 1622.500 53.340 ;
        RECT 1649.380 53.080 1649.640 53.340 ;
        RECT 1658.120 50.700 1658.380 50.960 ;
        RECT 2259.340 50.700 2259.600 50.960 ;
        RECT 2259.340 2.760 2259.600 3.020 ;
        RECT 2264.860 2.760 2265.120 3.020 ;
      LAYER met2 ;
        RECT 1622.300 53.370 1622.440 54.000 ;
        RECT 1622.240 53.050 1622.500 53.370 ;
        RECT 1649.380 53.050 1649.640 53.370 ;
        RECT 1649.440 52.885 1649.580 53.050 ;
        RECT 1649.370 52.515 1649.650 52.885 ;
        RECT 1658.110 52.515 1658.390 52.885 ;
        RECT 1658.180 50.990 1658.320 52.515 ;
        RECT 1658.120 50.670 1658.380 50.990 ;
        RECT 2259.340 50.670 2259.600 50.990 ;
        RECT 2259.400 3.050 2259.540 50.670 ;
        RECT 2259.340 2.730 2259.600 3.050 ;
        RECT 2264.860 2.730 2265.120 3.050 ;
        RECT 2264.920 2.400 2265.060 2.730 ;
        RECT 2264.850 0.000 2265.130 2.400 ;
      LAYER via2 ;
        RECT 1649.370 52.560 1649.650 52.840 ;
        RECT 1658.110 52.560 1658.390 52.840 ;
      LAYER met3 ;
        RECT 1649.345 52.850 1649.675 52.865 ;
        RECT 1658.085 52.850 1658.415 52.865 ;
        RECT 1649.345 52.550 1658.415 52.850 ;
        RECT 1649.345 52.535 1649.675 52.550 ;
        RECT 1658.085 52.535 1658.415 52.550 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1657.705 50.575 1657.875 50.915 ;
        RECT 1657.245 50.405 1657.875 50.575 ;
        RECT 1657.245 50.235 1657.415 50.405 ;
        RECT 1655.865 50.065 1657.415 50.235 ;
      LAYER mcon ;
        RECT 1657.705 50.745 1657.875 50.915 ;
      LAYER met1 ;
        RECT 2279.550 51.240 2279.870 51.300 ;
        RECT 1657.720 51.100 2279.870 51.240 ;
        RECT 1657.720 50.945 1657.860 51.100 ;
        RECT 2279.550 51.040 2279.870 51.100 ;
        RECT 1657.645 50.715 1657.935 50.945 ;
        RECT 1622.670 50.220 1622.990 50.280 ;
        RECT 1655.805 50.220 1656.095 50.265 ;
        RECT 1622.670 50.080 1656.095 50.220 ;
        RECT 1622.670 50.020 1622.990 50.080 ;
        RECT 1655.805 50.035 1656.095 50.080 ;
      LAYER via ;
        RECT 2279.580 51.040 2279.840 51.300 ;
        RECT 1622.700 50.020 1622.960 50.280 ;
      LAYER met2 ;
        RECT 1622.760 50.310 1622.900 54.000 ;
        RECT 2279.580 51.010 2279.840 51.330 ;
        RECT 1622.700 49.990 1622.960 50.310 ;
        RECT 2279.640 3.130 2279.780 51.010 ;
        RECT 2279.640 2.990 2282.540 3.130 ;
        RECT 2282.400 2.960 2282.540 2.990 ;
        RECT 2282.400 2.820 2283.000 2.960 ;
        RECT 2282.860 2.400 2283.000 2.820 ;
        RECT 2282.790 0.000 2283.070 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1657.245 50.745 1657.415 54.000 ;
      LAYER met1 ;
        RECT 1629.110 50.900 1629.430 50.960 ;
        RECT 1657.185 50.900 1657.475 50.945 ;
        RECT 1629.110 50.760 1657.475 50.900 ;
        RECT 1629.110 50.700 1629.430 50.760 ;
        RECT 1657.185 50.715 1657.475 50.760 ;
      LAYER via ;
        RECT 1629.140 50.700 1629.400 50.960 ;
      LAYER met2 ;
        RECT 1629.200 50.990 1629.340 54.000 ;
        RECT 1629.140 50.670 1629.400 50.990 ;
        RECT 2300.800 2.400 2300.940 54.000 ;
        RECT 2300.730 0.000 2301.010 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1658.165 50.235 1658.335 53.975 ;
        RECT 1657.705 50.065 1658.335 50.235 ;
      LAYER mcon ;
        RECT 1658.165 53.805 1658.335 53.975 ;
      LAYER met1 ;
        RECT 1658.105 53.960 1658.395 54.000 ;
        RECT 2314.050 53.960 2314.370 54.000 ;
        RECT 1658.105 53.820 2314.370 53.960 ;
        RECT 1658.105 53.775 1658.395 53.820 ;
        RECT 2314.050 53.760 2314.370 53.820 ;
        RECT 1629.570 50.560 1629.890 50.620 ;
        RECT 1629.570 50.420 1656.480 50.560 ;
        RECT 1629.570 50.360 1629.890 50.420 ;
        RECT 1656.340 50.220 1656.480 50.420 ;
        RECT 1657.645 50.220 1657.935 50.265 ;
        RECT 1656.340 50.080 1657.935 50.220 ;
        RECT 1657.645 50.035 1657.935 50.080 ;
        RECT 2314.050 2.960 2314.370 3.020 ;
        RECT 2318.650 2.960 2318.970 3.020 ;
        RECT 2314.050 2.820 2318.970 2.960 ;
        RECT 2314.050 2.760 2314.370 2.820 ;
        RECT 2318.650 2.760 2318.970 2.820 ;
      LAYER via ;
        RECT 2314.080 53.760 2314.340 54.000 ;
        RECT 1629.600 50.360 1629.860 50.620 ;
        RECT 2314.080 2.760 2314.340 3.020 ;
        RECT 2318.680 2.760 2318.940 3.020 ;
      LAYER met2 ;
        RECT 1629.660 50.650 1629.800 54.000 ;
        RECT 2314.080 53.730 2314.340 54.000 ;
        RECT 1629.600 50.330 1629.860 50.650 ;
        RECT 2314.140 3.050 2314.280 53.730 ;
        RECT 2314.080 2.730 2314.340 3.050 ;
        RECT 2318.680 2.730 2318.940 3.050 ;
        RECT 2318.740 2.400 2318.880 2.730 ;
        RECT 2318.670 0.000 2318.950 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1657.705 53.805 1657.875 54.000 ;
        RECT 1706.465 53.465 1706.635 54.000 ;
      LAYER met1 ;
        RECT 1636.010 53.960 1636.330 54.000 ;
        RECT 1657.645 53.960 1657.935 54.000 ;
        RECT 1636.010 53.820 1657.935 53.960 ;
        RECT 1636.010 53.760 1636.330 53.820 ;
        RECT 1657.645 53.775 1657.935 53.820 ;
        RECT 1706.405 53.620 1706.695 53.665 ;
        RECT 2334.750 53.620 2335.070 53.680 ;
        RECT 1706.405 53.480 2335.070 53.620 ;
        RECT 1706.405 53.435 1706.695 53.480 ;
        RECT 2334.750 53.420 2335.070 53.480 ;
        RECT 2334.750 2.960 2335.070 3.020 ;
        RECT 2336.590 2.960 2336.910 3.020 ;
        RECT 2334.750 2.820 2336.910 2.960 ;
        RECT 2334.750 2.760 2335.070 2.820 ;
        RECT 2336.590 2.760 2336.910 2.820 ;
      LAYER via ;
        RECT 1636.040 53.760 1636.300 54.000 ;
        RECT 2334.780 53.420 2335.040 53.680 ;
        RECT 2334.780 2.760 2335.040 3.020 ;
        RECT 2336.620 2.760 2336.880 3.020 ;
      LAYER met2 ;
        RECT 1636.040 53.730 1636.300 54.000 ;
        RECT 2334.780 53.390 2335.040 53.710 ;
        RECT 2334.840 3.050 2334.980 53.390 ;
        RECT 2334.780 2.730 2335.040 3.050 ;
        RECT 2336.620 2.730 2336.880 3.050 ;
        RECT 2336.680 2.400 2336.820 2.730 ;
        RECT 2336.610 0.000 2336.890 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1656.325 51.085 1656.495 54.000 ;
        RECT 1706.005 53.125 1706.175 54.000 ;
      LAYER met1 ;
        RECT 1705.945 53.280 1706.235 53.325 ;
        RECT 2348.550 53.280 2348.870 53.340 ;
        RECT 1705.945 53.140 2348.870 53.280 ;
        RECT 1705.945 53.095 1706.235 53.140 ;
        RECT 2348.550 53.080 2348.870 53.140 ;
        RECT 1635.550 51.240 1635.870 51.300 ;
        RECT 1656.265 51.240 1656.555 51.285 ;
        RECT 1635.550 51.100 1656.555 51.240 ;
        RECT 1635.550 51.040 1635.870 51.100 ;
        RECT 1656.265 51.055 1656.555 51.100 ;
        RECT 2348.550 2.960 2348.870 3.020 ;
        RECT 2354.070 2.960 2354.390 3.020 ;
        RECT 2348.550 2.820 2354.390 2.960 ;
        RECT 2348.550 2.760 2348.870 2.820 ;
        RECT 2354.070 2.760 2354.390 2.820 ;
      LAYER via ;
        RECT 2348.580 53.080 2348.840 53.340 ;
        RECT 1635.580 51.040 1635.840 51.300 ;
        RECT 2348.580 2.760 2348.840 3.020 ;
        RECT 2354.100 2.760 2354.360 3.020 ;
      LAYER met2 ;
        RECT 1635.640 51.330 1635.780 54.000 ;
        RECT 2348.580 53.050 2348.840 53.370 ;
        RECT 1635.580 51.010 1635.840 51.330 ;
        RECT 2348.640 3.050 2348.780 53.050 ;
        RECT 2348.580 2.730 2348.840 3.050 ;
        RECT 2354.100 2.730 2354.360 3.050 ;
        RECT 2354.160 2.400 2354.300 2.730 ;
        RECT 2354.090 0.000 2354.370 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1705.545 53.125 1705.715 54.000 ;
        RECT 2092.865 52.445 2093.035 54.000 ;
      LAYER met1 ;
        RECT 1642.450 53.620 1642.770 53.680 ;
        RECT 1642.450 53.480 1659.240 53.620 ;
        RECT 1642.450 53.420 1642.770 53.480 ;
        RECT 1659.100 53.280 1659.240 53.480 ;
        RECT 1705.485 53.280 1705.775 53.325 ;
        RECT 1659.100 53.140 1705.775 53.280 ;
        RECT 1705.485 53.095 1705.775 53.140 ;
        RECT 2372.010 52.940 2372.330 53.000 ;
        RECT 2117.260 52.800 2372.330 52.940 ;
        RECT 2092.805 52.600 2093.095 52.645 ;
        RECT 2117.260 52.600 2117.400 52.800 ;
        RECT 2372.010 52.740 2372.330 52.800 ;
        RECT 2092.805 52.460 2117.400 52.600 ;
        RECT 2092.805 52.415 2093.095 52.460 ;
      LAYER via ;
        RECT 1642.480 53.420 1642.740 53.680 ;
        RECT 2372.040 52.740 2372.300 53.000 ;
      LAYER met2 ;
        RECT 1642.540 53.710 1642.680 54.000 ;
        RECT 1642.480 53.390 1642.740 53.710 ;
        RECT 2372.040 52.710 2372.300 53.030 ;
        RECT 2372.100 2.400 2372.240 52.710 ;
        RECT 2372.030 0.000 2372.310 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1659.545 53.465 1659.715 54.000 ;
        RECT 1704.625 53.465 1704.795 54.000 ;
        RECT 2045.485 52.445 2045.655 54.000 ;
        RECT 2092.405 52.445 2092.575 54.000 ;
        RECT 2093.785 52.785 2093.955 54.000 ;
        RECT 2116.785 52.615 2116.955 52.955 ;
        RECT 2116.785 52.445 2117.875 52.615 ;
      LAYER mcon ;
        RECT 2116.785 52.785 2116.955 52.955 ;
        RECT 2117.705 52.445 2117.875 52.615 ;
      LAYER met1 ;
        RECT 1659.485 53.620 1659.775 53.665 ;
        RECT 1704.565 53.620 1704.855 53.665 ;
        RECT 1659.485 53.480 1704.855 53.620 ;
        RECT 1659.485 53.435 1659.775 53.480 ;
        RECT 1704.565 53.435 1704.855 53.480 ;
        RECT 2093.725 52.940 2094.015 52.985 ;
        RECT 2116.725 52.940 2117.015 52.985 ;
        RECT 2093.725 52.800 2117.015 52.940 ;
        RECT 2093.725 52.755 2094.015 52.800 ;
        RECT 2116.725 52.755 2117.015 52.800 ;
        RECT 2045.425 52.600 2045.715 52.645 ;
        RECT 2092.345 52.600 2092.635 52.645 ;
        RECT 2045.425 52.460 2092.635 52.600 ;
        RECT 2045.425 52.415 2045.715 52.460 ;
        RECT 2092.345 52.415 2092.635 52.460 ;
        RECT 2117.645 52.600 2117.935 52.645 ;
        RECT 2389.950 52.600 2390.270 52.660 ;
        RECT 2117.645 52.460 2390.270 52.600 ;
        RECT 2117.645 52.415 2117.935 52.460 ;
        RECT 2389.950 52.400 2390.270 52.460 ;
      LAYER via ;
        RECT 2389.980 52.400 2390.240 52.660 ;
      LAYER met2 ;
        RECT 2389.980 52.370 2390.240 52.690 ;
        RECT 2390.040 2.400 2390.180 52.370 ;
        RECT 2389.970 0.000 2390.250 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1658.625 53.125 1658.795 54.000 ;
      LAYER met1 ;
        RECT 1649.810 53.280 1650.130 53.340 ;
        RECT 1658.565 53.280 1658.855 53.325 ;
        RECT 1649.810 53.140 1658.855 53.280 ;
        RECT 1649.810 53.080 1650.130 53.140 ;
        RECT 1658.565 53.095 1658.855 53.140 ;
        RECT 2093.710 52.260 2094.030 52.320 ;
        RECT 2407.890 52.260 2408.210 52.320 ;
        RECT 2093.710 52.120 2408.210 52.260 ;
        RECT 2093.710 52.060 2094.030 52.120 ;
        RECT 2407.890 52.060 2408.210 52.120 ;
      LAYER via ;
        RECT 1649.840 53.080 1650.100 53.340 ;
        RECT 2093.740 52.060 2094.000 52.320 ;
        RECT 2407.920 52.060 2408.180 52.320 ;
      LAYER met2 ;
        RECT 1649.900 53.370 1650.040 54.000 ;
        RECT 1649.840 53.050 1650.100 53.370 ;
        RECT 1707.400 52.205 1707.540 54.000 ;
        RECT 2093.740 52.205 2094.000 52.350 ;
        RECT 1707.330 51.835 1707.610 52.205 ;
        RECT 2093.730 51.835 2094.010 52.205 ;
        RECT 2407.920 52.030 2408.180 52.350 ;
        RECT 2407.980 2.400 2408.120 52.030 ;
        RECT 2407.910 0.000 2408.190 2.400 ;
      LAYER via2 ;
        RECT 1707.330 51.880 1707.610 52.160 ;
        RECT 2093.730 51.880 2094.010 52.160 ;
      LAYER met3 ;
        RECT 1707.305 52.170 1707.635 52.185 ;
        RECT 2093.705 52.170 2094.035 52.185 ;
        RECT 1707.305 51.870 2094.035 52.170 ;
        RECT 1707.305 51.855 1707.635 51.870 ;
        RECT 2093.705 51.855 2094.035 51.870 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 802.030 36.280 802.350 36.340 ;
        RECT 1316.310 36.280 1316.630 36.340 ;
        RECT 802.030 36.140 1316.630 36.280 ;
        RECT 802.030 36.080 802.350 36.140 ;
        RECT 1316.310 36.080 1316.630 36.140 ;
      LAYER via ;
        RECT 802.060 36.080 802.320 36.340 ;
        RECT 1316.340 36.080 1316.600 36.340 ;
      LAYER met2 ;
        RECT 1316.400 36.370 1316.540 54.000 ;
        RECT 802.060 36.050 802.320 36.370 ;
        RECT 1316.340 36.050 1316.600 36.370 ;
        RECT 802.120 2.400 802.260 36.050 ;
        RECT 802.050 0.000 802.330 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 647.470 41.380 647.790 41.440 ;
        RECT 1280.430 41.380 1280.750 41.440 ;
        RECT 647.470 41.240 1280.750 41.380 ;
        RECT 647.470 41.180 647.790 41.240 ;
        RECT 1280.430 41.180 1280.750 41.240 ;
      LAYER via ;
        RECT 647.500 41.180 647.760 41.440 ;
        RECT 1280.460 41.180 1280.720 41.440 ;
      LAYER met2 ;
        RECT 1280.520 41.470 1280.660 54.000 ;
        RECT 647.500 41.150 647.760 41.470 ;
        RECT 1280.460 41.150 1280.720 41.470 ;
        RECT 647.560 2.400 647.700 41.150 ;
        RECT 647.490 0.000 647.770 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1656.340 51.525 1656.480 54.000 ;
        RECT 1656.270 51.155 1656.550 51.525 ;
        RECT 2432.290 51.155 2432.570 51.525 ;
        RECT 2432.360 35.090 2432.500 51.155 ;
        RECT 2431.440 34.950 2432.500 35.090 ;
        RECT 2431.440 2.400 2431.580 34.950 ;
        RECT 2431.370 0.000 2431.650 2.400 ;
      LAYER via2 ;
        RECT 1656.270 51.200 1656.550 51.480 ;
        RECT 2432.290 51.200 2432.570 51.480 ;
      LAYER met3 ;
        RECT 1656.245 51.490 1656.575 51.505 ;
        RECT 2432.265 51.490 2432.595 51.505 ;
        RECT 1656.245 51.190 2432.595 51.490 ;
        RECT 1656.245 51.175 1656.575 51.190 ;
        RECT 2432.265 51.175 2432.595 51.190 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2449.380 2.400 2449.520 54.000 ;
        RECT 2449.310 0.000 2449.590 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2465.940 3.130 2466.080 54.000 ;
        RECT 2465.940 2.990 2467.000 3.130 ;
        RECT 2466.860 2.960 2467.000 2.990 ;
        RECT 2466.860 2.820 2467.460 2.960 ;
        RECT 2467.320 2.400 2467.460 2.820 ;
        RECT 2467.250 0.000 2467.530 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2479.650 2.960 2479.970 3.020 ;
        RECT 2485.170 2.960 2485.490 3.020 ;
        RECT 2479.650 2.820 2485.490 2.960 ;
        RECT 2479.650 2.760 2479.970 2.820 ;
        RECT 2485.170 2.760 2485.490 2.820 ;
      LAYER via ;
        RECT 2479.680 2.760 2479.940 3.020 ;
        RECT 2485.200 2.760 2485.460 3.020 ;
      LAYER met2 ;
        RECT 2479.740 3.050 2479.880 54.000 ;
        RECT 2479.680 2.730 2479.940 3.050 ;
        RECT 2485.200 2.730 2485.460 3.050 ;
        RECT 2485.260 2.400 2485.400 2.730 ;
        RECT 2485.190 0.000 2485.470 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2500.350 2.960 2500.670 3.020 ;
        RECT 2503.110 2.960 2503.430 3.020 ;
        RECT 2500.350 2.820 2503.430 2.960 ;
        RECT 2500.350 2.760 2500.670 2.820 ;
        RECT 2503.110 2.760 2503.430 2.820 ;
      LAYER via ;
        RECT 2500.380 2.760 2500.640 3.020 ;
        RECT 2503.140 2.760 2503.400 3.020 ;
      LAYER met2 ;
        RECT 2500.440 3.050 2500.580 54.000 ;
        RECT 2500.380 2.730 2500.640 3.050 ;
        RECT 2503.140 2.730 2503.400 3.050 ;
        RECT 2503.200 2.400 2503.340 2.730 ;
        RECT 2503.130 0.000 2503.410 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2520.680 2.400 2520.820 54.000 ;
        RECT 2520.610 0.000 2520.890 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2534.850 2.960 2535.170 3.020 ;
        RECT 2538.530 2.960 2538.850 3.020 ;
        RECT 2534.850 2.820 2538.850 2.960 ;
        RECT 2534.850 2.760 2535.170 2.820 ;
        RECT 2538.530 2.760 2538.850 2.820 ;
      LAYER via ;
        RECT 2534.880 2.760 2535.140 3.020 ;
        RECT 2538.560 2.760 2538.820 3.020 ;
      LAYER met2 ;
        RECT 2534.940 3.050 2535.080 54.000 ;
        RECT 2534.880 2.730 2535.140 3.050 ;
        RECT 2538.560 2.730 2538.820 3.050 ;
        RECT 2538.620 2.400 2538.760 2.730 ;
        RECT 2538.550 0.000 2538.830 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2556.560 2.400 2556.700 54.000 ;
        RECT 2556.490 0.000 2556.770 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2574.500 2.400 2574.640 54.000 ;
        RECT 2574.430 0.000 2574.710 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2591.980 2.400 2592.120 54.000 ;
        RECT 2591.910 0.000 2592.190 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 825.950 35.940 826.270 36.000 ;
        RECT 1321.370 35.940 1321.690 36.000 ;
        RECT 825.950 35.800 1321.690 35.940 ;
        RECT 825.950 35.740 826.270 35.800 ;
        RECT 1321.370 35.740 1321.690 35.800 ;
      LAYER via ;
        RECT 825.980 35.740 826.240 36.000 ;
        RECT 1321.400 35.740 1321.660 36.000 ;
      LAYER met2 ;
        RECT 1321.460 36.030 1321.600 54.000 ;
        RECT 825.980 35.710 826.240 36.030 ;
        RECT 1321.400 35.710 1321.660 36.030 ;
        RECT 826.040 2.400 826.180 35.710 ;
        RECT 825.970 0.000 826.250 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2603.850 37.640 2604.170 37.700 ;
        RECT 2609.830 37.640 2610.150 37.700 ;
        RECT 2603.850 37.500 2610.150 37.640 ;
        RECT 2603.850 37.440 2604.170 37.500 ;
        RECT 2609.830 37.440 2610.150 37.500 ;
      LAYER via ;
        RECT 2603.880 37.440 2604.140 37.700 ;
        RECT 2609.860 37.440 2610.120 37.700 ;
      LAYER met2 ;
        RECT 2603.940 37.730 2604.080 54.000 ;
        RECT 2603.880 37.410 2604.140 37.730 ;
        RECT 2609.860 37.410 2610.120 37.730 ;
        RECT 2609.920 2.400 2610.060 37.410 ;
        RECT 2609.850 0.000 2610.130 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2627.860 2.400 2628.000 54.000 ;
        RECT 2627.790 0.000 2628.070 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2645.325 48.365 2645.495 54.000 ;
      LAYER met1 ;
        RECT 2645.265 48.520 2645.555 48.565 ;
        RECT 2645.710 48.520 2646.030 48.580 ;
        RECT 2645.265 48.380 2646.030 48.520 ;
        RECT 2645.265 48.335 2645.555 48.380 ;
        RECT 2645.710 48.320 2646.030 48.380 ;
        RECT 2645.710 2.960 2646.030 3.020 ;
        RECT 2646.170 2.960 2646.490 3.020 ;
        RECT 2645.710 2.820 2646.490 2.960 ;
        RECT 2645.710 2.760 2646.030 2.820 ;
        RECT 2646.170 2.760 2646.490 2.820 ;
      LAYER via ;
        RECT 2645.740 48.320 2646.000 48.580 ;
        RECT 2645.740 2.760 2646.000 3.020 ;
        RECT 2646.200 2.760 2646.460 3.020 ;
      LAYER met2 ;
        RECT 2645.740 48.290 2646.000 48.610 ;
        RECT 2645.800 48.010 2645.940 48.290 ;
        RECT 2645.800 47.870 2646.400 48.010 ;
        RECT 2646.260 3.050 2646.400 47.870 ;
        RECT 2645.740 2.730 2646.000 3.050 ;
        RECT 2646.200 2.730 2646.460 3.050 ;
        RECT 2645.800 2.400 2645.940 2.730 ;
        RECT 2645.730 0.000 2646.010 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2663.740 2.400 2663.880 54.000 ;
        RECT 2663.670 0.000 2663.950 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2679.825 48.365 2679.995 54.000 ;
      LAYER met1 ;
        RECT 2679.765 48.520 2680.055 48.565 ;
        RECT 2681.130 48.520 2681.450 48.580 ;
        RECT 2679.765 48.380 2681.450 48.520 ;
        RECT 2679.765 48.335 2680.055 48.380 ;
        RECT 2681.130 48.320 2681.450 48.380 ;
      LAYER via ;
        RECT 2681.160 48.320 2681.420 48.580 ;
      LAYER met2 ;
        RECT 2681.160 48.290 2681.420 48.610 ;
        RECT 2681.220 2.400 2681.360 48.290 ;
        RECT 2681.150 0.000 2681.430 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2699.160 2.400 2699.300 54.000 ;
        RECT 2699.090 0.000 2699.370 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2717.100 2.400 2717.240 54.000 ;
        RECT 2717.030 0.000 2717.310 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2735.040 2.400 2735.180 54.000 ;
        RECT 2734.970 0.000 2735.250 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2752.980 2.400 2753.120 54.000 ;
        RECT 2752.910 0.000 2753.190 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2770.460 2.400 2770.600 54.000 ;
        RECT 2770.390 0.000 2770.670 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 843.430 34.920 843.750 34.980 ;
        RECT 1320.910 34.920 1321.230 34.980 ;
        RECT 843.430 34.780 1321.230 34.920 ;
        RECT 843.430 34.720 843.750 34.780 ;
        RECT 1320.910 34.720 1321.230 34.780 ;
      LAYER via ;
        RECT 843.460 34.720 843.720 34.980 ;
        RECT 1320.940 34.720 1321.200 34.980 ;
      LAYER met2 ;
        RECT 1321.000 35.010 1321.140 54.000 ;
        RECT 843.460 34.690 843.720 35.010 ;
        RECT 1320.940 34.690 1321.200 35.010 ;
        RECT 843.520 2.400 843.660 34.690 ;
        RECT 843.450 0.000 843.730 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2788.400 2.400 2788.540 54.000 ;
        RECT 2788.330 0.000 2788.610 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2804.025 48.365 2804.195 54.000 ;
      LAYER met1 ;
        RECT 2803.965 48.520 2804.255 48.565 ;
        RECT 2806.250 48.520 2806.570 48.580 ;
        RECT 2803.965 48.380 2806.570 48.520 ;
        RECT 2803.965 48.335 2804.255 48.380 ;
        RECT 2806.250 48.320 2806.570 48.380 ;
      LAYER via ;
        RECT 2806.280 48.320 2806.540 48.580 ;
      LAYER met2 ;
        RECT 2806.280 48.290 2806.540 48.610 ;
        RECT 2806.340 2.400 2806.480 48.290 ;
        RECT 2806.270 0.000 2806.550 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2817.750 37.640 2818.070 37.700 ;
        RECT 2824.190 37.640 2824.510 37.700 ;
        RECT 2817.750 37.500 2824.510 37.640 ;
        RECT 2817.750 37.440 2818.070 37.500 ;
        RECT 2824.190 37.440 2824.510 37.500 ;
      LAYER via ;
        RECT 2817.780 37.440 2818.040 37.700 ;
        RECT 2824.220 37.440 2824.480 37.700 ;
      LAYER met2 ;
        RECT 2817.840 37.730 2817.980 54.000 ;
        RECT 2817.780 37.410 2818.040 37.730 ;
        RECT 2824.220 37.410 2824.480 37.730 ;
        RECT 2824.280 2.400 2824.420 37.410 ;
        RECT 2824.210 0.000 2824.490 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2841.760 2.400 2841.900 54.000 ;
        RECT 2841.690 0.000 2841.970 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2859.225 48.365 2859.395 54.000 ;
      LAYER met1 ;
        RECT 2859.165 48.520 2859.455 48.565 ;
        RECT 2859.610 48.520 2859.930 48.580 ;
        RECT 2859.165 48.380 2859.930 48.520 ;
        RECT 2859.165 48.335 2859.455 48.380 ;
        RECT 2859.610 48.320 2859.930 48.380 ;
      LAYER via ;
        RECT 2859.640 48.320 2859.900 48.580 ;
      LAYER met2 ;
        RECT 2859.640 48.290 2859.900 48.610 ;
        RECT 2859.700 2.400 2859.840 48.290 ;
        RECT 2859.630 0.000 2859.910 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2872.950 1307.540 2873.270 1307.600 ;
        RECT 2870.580 1307.400 2873.270 1307.540 ;
        RECT 2872.950 1307.340 2873.270 1307.400 ;
        RECT 2872.950 62.120 2873.270 62.180 ;
        RECT 2877.550 62.120 2877.870 62.180 ;
        RECT 2872.950 61.980 2877.870 62.120 ;
        RECT 2872.950 61.920 2873.270 61.980 ;
        RECT 2877.550 61.920 2877.870 61.980 ;
      LAYER via ;
        RECT 2872.980 1307.340 2873.240 1307.600 ;
        RECT 2872.980 61.920 2873.240 62.180 ;
        RECT 2877.580 61.920 2877.840 62.180 ;
      LAYER met2 ;
        RECT 2872.980 1307.310 2873.240 1307.630 ;
        RECT 2873.040 62.210 2873.180 1307.310 ;
        RECT 2872.980 61.890 2873.240 62.210 ;
        RECT 2877.580 61.890 2877.840 62.210 ;
        RECT 2877.640 2.400 2877.780 61.890 ;
        RECT 2877.570 0.000 2877.850 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2889.970 1418.040 2890.290 1418.100 ;
        RECT 2870.580 1417.900 2890.290 1418.040 ;
        RECT 2889.970 1417.840 2890.290 1417.900 ;
        RECT 2889.970 20.640 2890.290 20.700 ;
        RECT 2895.490 20.640 2895.810 20.700 ;
        RECT 2889.970 20.500 2895.810 20.640 ;
        RECT 2889.970 20.440 2890.290 20.500 ;
        RECT 2895.490 20.440 2895.810 20.500 ;
      LAYER via ;
        RECT 2890.000 1417.840 2890.260 1418.100 ;
        RECT 2890.000 20.440 2890.260 20.700 ;
        RECT 2895.520 20.440 2895.780 20.700 ;
      LAYER met2 ;
        RECT 2890.000 1417.810 2890.260 1418.130 ;
        RECT 2890.060 20.730 2890.200 1417.810 ;
        RECT 2890.000 20.410 2890.260 20.730 ;
        RECT 2895.520 20.410 2895.780 20.730 ;
        RECT 2895.580 2.400 2895.720 20.410 ;
        RECT 2895.510 0.000 2895.790 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2907.450 1266.060 2907.770 1266.120 ;
        RECT 2870.580 1265.920 2907.770 1266.060 ;
        RECT 2907.450 1265.860 2907.770 1265.920 ;
        RECT 2907.450 37.640 2907.770 37.700 ;
        RECT 2913.430 37.640 2913.750 37.700 ;
        RECT 2907.450 37.500 2913.750 37.640 ;
        RECT 2907.450 37.440 2907.770 37.500 ;
        RECT 2913.430 37.440 2913.750 37.500 ;
      LAYER via ;
        RECT 2907.480 1265.860 2907.740 1266.120 ;
        RECT 2907.480 37.440 2907.740 37.700 ;
        RECT 2913.460 37.440 2913.720 37.700 ;
      LAYER met2 ;
        RECT 2907.480 1265.830 2907.740 1266.150 ;
        RECT 2907.540 37.730 2907.680 1265.830 ;
        RECT 2907.480 37.410 2907.740 37.730 ;
        RECT 2913.460 37.410 2913.720 37.730 ;
        RECT 2913.520 2.400 2913.660 37.410 ;
        RECT 2913.450 0.000 2913.730 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 861.370 34.580 861.690 34.640 ;
        RECT 1328.730 34.580 1329.050 34.640 ;
        RECT 861.370 34.440 1329.050 34.580 ;
        RECT 861.370 34.380 861.690 34.440 ;
        RECT 1328.730 34.380 1329.050 34.440 ;
      LAYER via ;
        RECT 861.400 34.380 861.660 34.640 ;
        RECT 1328.760 34.380 1329.020 34.640 ;
      LAYER met2 ;
        RECT 1328.820 34.670 1328.960 54.000 ;
        RECT 861.400 34.350 861.660 34.670 ;
        RECT 1328.760 34.350 1329.020 34.670 ;
        RECT 861.460 2.400 861.600 34.350 ;
        RECT 861.390 0.000 861.670 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 885.825 29.325 885.995 41.735 ;
        RECT 975.065 38.505 975.235 41.735 ;
      LAYER mcon ;
        RECT 885.825 41.565 885.995 41.735 ;
        RECT 975.065 41.565 975.235 41.735 ;
      LAYER met1 ;
        RECT 885.765 41.720 886.055 41.765 ;
        RECT 975.005 41.720 975.295 41.765 ;
        RECT 885.765 41.580 975.295 41.720 ;
        RECT 885.765 41.535 886.055 41.580 ;
        RECT 975.005 41.535 975.295 41.580 ;
        RECT 975.005 38.660 975.295 38.705 ;
        RECT 1328.270 38.660 1328.590 38.720 ;
        RECT 975.005 38.520 1328.590 38.660 ;
        RECT 975.005 38.475 975.295 38.520 ;
        RECT 1328.270 38.460 1328.590 38.520 ;
        RECT 879.310 29.480 879.630 29.540 ;
        RECT 885.765 29.480 886.055 29.525 ;
        RECT 879.310 29.340 886.055 29.480 ;
        RECT 879.310 29.280 879.630 29.340 ;
        RECT 885.765 29.295 886.055 29.340 ;
      LAYER via ;
        RECT 1328.300 38.460 1328.560 38.720 ;
        RECT 879.340 29.280 879.600 29.540 ;
      LAYER met2 ;
        RECT 1328.360 38.750 1328.500 54.000 ;
        RECT 1328.300 38.430 1328.560 38.750 ;
        RECT 879.340 29.250 879.600 29.570 ;
        RECT 879.400 2.400 879.540 29.250 ;
        RECT 879.330 0.000 879.610 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 933.665 28.985 933.835 39.015 ;
      LAYER mcon ;
        RECT 933.665 38.845 933.835 39.015 ;
      LAYER met1 ;
        RECT 933.605 39.000 933.895 39.045 ;
        RECT 1335.170 39.000 1335.490 39.060 ;
        RECT 933.605 38.860 1335.490 39.000 ;
        RECT 933.605 38.815 933.895 38.860 ;
        RECT 1335.170 38.800 1335.490 38.860 ;
        RECT 897.250 29.140 897.570 29.200 ;
        RECT 933.605 29.140 933.895 29.185 ;
        RECT 897.250 29.000 933.895 29.140 ;
        RECT 897.250 28.940 897.570 29.000 ;
        RECT 933.605 28.955 933.895 29.000 ;
      LAYER via ;
        RECT 1335.200 38.800 1335.460 39.060 ;
        RECT 897.280 28.940 897.540 29.200 ;
      LAYER met2 ;
        RECT 1335.260 39.090 1335.400 54.000 ;
        RECT 1335.200 38.770 1335.460 39.090 ;
        RECT 897.280 28.910 897.540 29.230 ;
        RECT 897.340 2.400 897.480 28.910 ;
        RECT 897.270 0.000 897.550 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 915.190 2.960 915.510 3.020 ;
        RECT 919.790 2.960 920.110 3.020 ;
        RECT 915.190 2.820 920.110 2.960 ;
        RECT 915.190 2.760 915.510 2.820 ;
        RECT 919.790 2.760 920.110 2.820 ;
      LAYER via ;
        RECT 915.220 2.760 915.480 3.020 ;
        RECT 919.820 2.760 920.080 3.020 ;
      LAYER met2 ;
        RECT 919.880 3.050 920.020 54.000 ;
        RECT 915.220 2.730 915.480 3.050 ;
        RECT 919.820 2.730 920.080 3.050 ;
        RECT 915.280 2.400 915.420 2.730 ;
        RECT 915.210 0.000 915.490 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 933.680 3.130 933.820 54.000 ;
        RECT 933.220 2.990 933.820 3.130 ;
        RECT 933.220 2.960 933.360 2.990 ;
        RECT 932.760 2.820 933.360 2.960 ;
        RECT 932.760 2.400 932.900 2.820 ;
        RECT 932.690 0.000 932.970 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 950.610 2.960 950.930 3.020 ;
        RECT 951.990 2.960 952.310 3.020 ;
        RECT 950.610 2.820 952.310 2.960 ;
        RECT 950.610 2.760 950.930 2.820 ;
        RECT 951.990 2.760 952.310 2.820 ;
      LAYER via ;
        RECT 950.640 2.760 950.900 3.020 ;
        RECT 952.020 2.760 952.280 3.020 ;
      LAYER met2 ;
        RECT 952.080 48.805 952.220 54.000 ;
        RECT 952.010 48.435 952.290 48.805 ;
        RECT 952.930 48.435 953.210 48.805 ;
        RECT 953.000 48.010 953.140 48.435 ;
        RECT 952.080 47.870 953.140 48.010 ;
        RECT 952.080 3.050 952.220 47.870 ;
        RECT 950.640 2.730 950.900 3.050 ;
        RECT 952.020 2.730 952.280 3.050 ;
        RECT 950.700 2.400 950.840 2.730 ;
        RECT 950.630 0.000 950.910 2.400 ;
      LAYER via2 ;
        RECT 952.010 48.480 952.290 48.760 ;
        RECT 952.930 48.480 953.210 48.760 ;
      LAYER met3 ;
        RECT 951.985 48.770 952.315 48.785 ;
        RECT 952.905 48.770 953.235 48.785 ;
        RECT 951.985 48.470 953.235 48.770 ;
        RECT 951.985 48.455 952.315 48.470 ;
        RECT 952.905 48.455 953.235 48.470 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 968.550 38.660 968.870 38.720 ;
        RECT 974.530 38.660 974.850 38.720 ;
        RECT 968.550 38.520 974.850 38.660 ;
        RECT 968.550 38.460 968.870 38.520 ;
        RECT 974.530 38.460 974.850 38.520 ;
      LAYER via ;
        RECT 968.580 38.460 968.840 38.720 ;
        RECT 974.560 38.460 974.820 38.720 ;
      LAYER met2 ;
        RECT 974.620 38.750 974.760 54.000 ;
        RECT 968.580 38.430 968.840 38.750 ;
        RECT 974.560 38.430 974.820 38.750 ;
        RECT 968.640 2.400 968.780 38.430 ;
        RECT 968.570 0.000 968.850 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 986.490 2.960 986.810 3.020 ;
        RECT 988.790 2.960 989.110 3.020 ;
        RECT 986.490 2.820 989.110 2.960 ;
        RECT 986.490 2.760 986.810 2.820 ;
        RECT 988.790 2.760 989.110 2.820 ;
      LAYER via ;
        RECT 986.520 2.760 986.780 3.020 ;
        RECT 988.820 2.760 989.080 3.020 ;
      LAYER met2 ;
        RECT 988.880 3.050 989.020 54.000 ;
        RECT 986.520 2.730 986.780 3.050 ;
        RECT 988.820 2.730 989.080 3.050 ;
        RECT 986.580 2.400 986.720 2.730 ;
        RECT 986.510 0.000 986.790 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 665.410 19.960 665.730 20.020 ;
        RECT 670.930 19.960 671.250 20.020 ;
        RECT 665.410 19.820 671.250 19.960 ;
        RECT 665.410 19.760 665.730 19.820 ;
        RECT 670.930 19.760 671.250 19.820 ;
      LAYER via ;
        RECT 665.440 19.760 665.700 20.020 ;
        RECT 670.960 19.760 671.220 20.020 ;
      LAYER met2 ;
        RECT 671.020 20.050 671.160 54.000 ;
        RECT 665.440 19.730 665.700 20.050 ;
        RECT 670.960 19.730 671.220 20.050 ;
        RECT 665.500 2.400 665.640 19.730 ;
        RECT 665.430 0.000 665.710 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1004.430 2.960 1004.750 3.020 ;
        RECT 1009.490 2.960 1009.810 3.020 ;
        RECT 1004.430 2.820 1009.810 2.960 ;
        RECT 1004.430 2.760 1004.750 2.820 ;
        RECT 1009.490 2.760 1009.810 2.820 ;
      LAYER via ;
        RECT 1004.460 2.760 1004.720 3.020 ;
        RECT 1009.520 2.760 1009.780 3.020 ;
      LAYER met2 ;
        RECT 1009.580 3.050 1009.720 54.000 ;
        RECT 1004.460 2.730 1004.720 3.050 ;
        RECT 1009.520 2.730 1009.780 3.050 ;
        RECT 1004.520 2.400 1004.660 2.730 ;
        RECT 1004.450 0.000 1004.730 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1023.380 3.130 1023.520 54.000 ;
        RECT 1022.000 2.990 1023.520 3.130 ;
        RECT 1022.000 2.400 1022.140 2.990 ;
        RECT 1021.930 0.000 1022.210 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1039.850 43.080 1040.170 43.140 ;
        RECT 1363.690 43.080 1364.010 43.140 ;
        RECT 1039.850 42.940 1364.010 43.080 ;
        RECT 1039.850 42.880 1040.170 42.940 ;
        RECT 1363.690 42.880 1364.010 42.940 ;
      LAYER via ;
        RECT 1039.880 42.880 1040.140 43.140 ;
        RECT 1363.720 42.880 1363.980 43.140 ;
      LAYER met2 ;
        RECT 1363.780 43.170 1363.920 54.000 ;
        RECT 1039.880 42.850 1040.140 43.170 ;
        RECT 1363.720 42.850 1363.980 43.170 ;
        RECT 1039.940 2.400 1040.080 42.850 ;
        RECT 1039.870 0.000 1040.150 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1057.790 42.740 1058.110 42.800 ;
        RECT 1369.670 42.740 1369.990 42.800 ;
        RECT 1057.790 42.600 1369.990 42.740 ;
        RECT 1057.790 42.540 1058.110 42.600 ;
        RECT 1369.670 42.540 1369.990 42.600 ;
      LAYER via ;
        RECT 1057.820 42.540 1058.080 42.800 ;
        RECT 1369.700 42.540 1369.960 42.800 ;
      LAYER met2 ;
        RECT 1369.760 42.830 1369.900 54.000 ;
        RECT 1057.820 42.510 1058.080 42.830 ;
        RECT 1369.700 42.510 1369.960 42.830 ;
        RECT 1057.880 2.400 1058.020 42.510 ;
        RECT 1057.810 0.000 1058.090 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1371.970 42.400 1372.290 42.460 ;
        RECT 1093.300 42.260 1372.290 42.400 ;
        RECT 1075.730 42.060 1076.050 42.120 ;
        RECT 1093.300 42.060 1093.440 42.260 ;
        RECT 1371.970 42.200 1372.290 42.260 ;
        RECT 1075.730 41.920 1093.440 42.060 ;
        RECT 1075.730 41.860 1076.050 41.920 ;
      LAYER via ;
        RECT 1075.760 41.860 1076.020 42.120 ;
        RECT 1372.000 42.200 1372.260 42.460 ;
      LAYER met2 ;
        RECT 1372.060 42.490 1372.200 54.000 ;
        RECT 1372.000 42.170 1372.260 42.490 ;
        RECT 1075.760 41.830 1076.020 42.150 ;
        RECT 1075.820 2.400 1075.960 41.830 ;
        RECT 1075.750 0.000 1076.030 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1125.945 41.905 1127.035 42.075 ;
        RECT 1125.945 41.565 1126.115 41.905 ;
      LAYER mcon ;
        RECT 1126.865 41.905 1127.035 42.075 ;
      LAYER met1 ;
        RECT 1126.805 42.060 1127.095 42.105 ;
        RECT 1376.570 42.060 1376.890 42.120 ;
        RECT 1126.805 41.920 1376.890 42.060 ;
        RECT 1126.805 41.875 1127.095 41.920 ;
        RECT 1376.570 41.860 1376.890 41.920 ;
        RECT 1092.750 41.720 1093.070 41.780 ;
        RECT 1125.885 41.720 1126.175 41.765 ;
        RECT 1092.750 41.580 1126.175 41.720 ;
        RECT 1092.750 41.520 1093.070 41.580 ;
        RECT 1125.885 41.535 1126.175 41.580 ;
      LAYER via ;
        RECT 1376.600 41.860 1376.860 42.120 ;
        RECT 1092.780 41.520 1093.040 41.780 ;
      LAYER met2 ;
        RECT 1376.660 42.150 1376.800 54.000 ;
        RECT 1376.600 41.830 1376.860 42.150 ;
        RECT 1092.780 41.490 1093.040 41.810 ;
        RECT 1092.840 14.010 1092.980 41.490 ;
        RECT 1092.840 13.870 1093.440 14.010 ;
        RECT 1093.300 2.400 1093.440 13.870 ;
        RECT 1093.230 0.000 1093.510 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1112.530 42.060 1112.850 42.120 ;
        RECT 1112.530 41.920 1126.560 42.060 ;
        RECT 1112.530 41.860 1112.850 41.920 ;
        RECT 1126.420 41.720 1126.560 41.920 ;
        RECT 1377.030 41.720 1377.350 41.780 ;
        RECT 1126.420 41.580 1377.350 41.720 ;
        RECT 1377.030 41.520 1377.350 41.580 ;
      LAYER via ;
        RECT 1112.560 41.860 1112.820 42.120 ;
        RECT 1377.060 41.520 1377.320 41.780 ;
      LAYER met2 ;
        RECT 1112.560 41.830 1112.820 42.150 ;
        RECT 1112.620 3.130 1112.760 41.830 ;
        RECT 1377.120 41.810 1377.260 54.000 ;
        RECT 1377.060 41.490 1377.320 41.810 ;
        RECT 1111.240 2.990 1112.760 3.130 ;
        RECT 1111.240 2.400 1111.380 2.990 ;
        RECT 1111.170 0.000 1111.450 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.090 44.780 1175.410 44.840 ;
        RECT 1383.470 44.780 1383.790 44.840 ;
        RECT 1175.090 44.640 1383.790 44.780 ;
        RECT 1175.090 44.580 1175.410 44.640 ;
        RECT 1383.470 44.580 1383.790 44.640 ;
      LAYER via ;
        RECT 1175.120 44.580 1175.380 44.840 ;
        RECT 1383.500 44.580 1383.760 44.840 ;
      LAYER met2 ;
        RECT 1383.560 44.870 1383.700 54.000 ;
        RECT 1175.120 44.550 1175.380 44.870 ;
        RECT 1383.500 44.550 1383.760 44.870 ;
        RECT 1175.180 44.045 1175.320 44.550 ;
        RECT 1129.110 43.675 1129.390 44.045 ;
        RECT 1175.110 43.675 1175.390 44.045 ;
        RECT 1129.180 2.400 1129.320 43.675 ;
        RECT 1129.110 0.000 1129.390 2.400 ;
      LAYER via2 ;
        RECT 1129.110 43.720 1129.390 44.000 ;
        RECT 1175.110 43.720 1175.390 44.000 ;
      LAYER met3 ;
        RECT 1129.085 44.010 1129.415 44.025 ;
        RECT 1175.085 44.010 1175.415 44.025 ;
        RECT 1129.085 43.710 1175.415 44.010 ;
        RECT 1129.085 43.695 1129.415 43.710 ;
        RECT 1175.085 43.695 1175.415 43.710 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1174.630 45.120 1174.950 45.180 ;
        RECT 1383.930 45.120 1384.250 45.180 ;
        RECT 1174.630 44.980 1384.250 45.120 ;
        RECT 1174.630 44.920 1174.950 44.980 ;
        RECT 1383.930 44.920 1384.250 44.980 ;
      LAYER via ;
        RECT 1174.660 44.920 1174.920 45.180 ;
        RECT 1383.960 44.920 1384.220 45.180 ;
      LAYER met2 ;
        RECT 1384.020 45.210 1384.160 54.000 ;
        RECT 1174.660 44.890 1174.920 45.210 ;
        RECT 1383.960 44.890 1384.220 45.210 ;
        RECT 1174.720 44.725 1174.860 44.890 ;
        RECT 1147.050 44.355 1147.330 44.725 ;
        RECT 1174.650 44.355 1174.930 44.725 ;
        RECT 1147.120 2.400 1147.260 44.355 ;
        RECT 1147.050 0.000 1147.330 2.400 ;
      LAYER via2 ;
        RECT 1147.050 44.400 1147.330 44.680 ;
        RECT 1174.650 44.400 1174.930 44.680 ;
      LAYER met3 ;
        RECT 1147.025 44.690 1147.355 44.705 ;
        RECT 1174.625 44.690 1174.955 44.705 ;
        RECT 1147.025 44.390 1174.955 44.690 ;
        RECT 1147.025 44.375 1147.355 44.390 ;
        RECT 1174.625 44.375 1174.955 44.390 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1390.830 45.460 1391.150 45.520 ;
        RECT 1174.260 45.320 1391.150 45.460 ;
        RECT 1164.970 44.780 1165.290 44.840 ;
        RECT 1174.260 44.780 1174.400 45.320 ;
        RECT 1390.830 45.260 1391.150 45.320 ;
        RECT 1164.970 44.640 1174.400 44.780 ;
        RECT 1164.970 44.580 1165.290 44.640 ;
      LAYER via ;
        RECT 1165.000 44.580 1165.260 44.840 ;
        RECT 1390.860 45.260 1391.120 45.520 ;
      LAYER met2 ;
        RECT 1390.920 45.550 1391.060 54.000 ;
        RECT 1390.860 45.230 1391.120 45.550 ;
        RECT 1165.000 44.550 1165.260 44.870 ;
        RECT 1165.060 2.400 1165.200 44.550 ;
        RECT 1164.990 0.000 1165.270 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1272.685 48.025 1272.855 50.575 ;
      LAYER mcon ;
        RECT 1272.685 50.405 1272.855 50.575 ;
      LAYER met1 ;
        RECT 1223.850 50.560 1224.170 50.620 ;
        RECT 1272.625 50.560 1272.915 50.605 ;
        RECT 1223.850 50.420 1272.915 50.560 ;
        RECT 1223.850 50.360 1224.170 50.420 ;
        RECT 1272.625 50.375 1272.915 50.420 ;
        RECT 1272.625 48.180 1272.915 48.225 ;
        RECT 1287.330 48.180 1287.650 48.240 ;
        RECT 1272.625 48.040 1287.650 48.180 ;
        RECT 1272.625 47.995 1272.915 48.040 ;
        RECT 1287.330 47.980 1287.650 48.040 ;
        RECT 682.890 45.800 683.210 45.860 ;
        RECT 1223.850 45.800 1224.170 45.860 ;
        RECT 682.890 45.660 1224.170 45.800 ;
        RECT 682.890 45.600 683.210 45.660 ;
        RECT 1223.850 45.600 1224.170 45.660 ;
      LAYER via ;
        RECT 1223.880 50.360 1224.140 50.620 ;
        RECT 1287.360 47.980 1287.620 48.240 ;
        RECT 682.920 45.600 683.180 45.860 ;
        RECT 1223.880 45.600 1224.140 45.860 ;
      LAYER met2 ;
        RECT 1223.880 50.330 1224.140 50.650 ;
        RECT 1223.940 45.890 1224.080 50.330 ;
        RECT 1287.420 48.270 1287.560 54.000 ;
        RECT 1287.360 47.950 1287.620 48.270 ;
        RECT 682.920 45.570 683.180 45.890 ;
        RECT 1223.880 45.570 1224.140 45.890 ;
        RECT 682.980 2.400 683.120 45.570 ;
        RECT 682.910 0.000 683.190 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1224.310 45.800 1224.630 45.860 ;
        RECT 1271.230 45.800 1271.550 45.860 ;
        RECT 1224.310 45.660 1271.550 45.800 ;
        RECT 1224.310 45.600 1224.630 45.660 ;
        RECT 1271.230 45.600 1271.550 45.660 ;
        RECT 1272.610 45.800 1272.930 45.860 ;
        RECT 1390.370 45.800 1390.690 45.860 ;
        RECT 1272.610 45.660 1390.690 45.800 ;
        RECT 1272.610 45.600 1272.930 45.660 ;
        RECT 1390.370 45.600 1390.690 45.660 ;
        RECT 1182.450 20.640 1182.770 20.700 ;
        RECT 1188.890 20.640 1189.210 20.700 ;
        RECT 1182.450 20.500 1189.210 20.640 ;
        RECT 1182.450 20.440 1182.770 20.500 ;
        RECT 1188.890 20.440 1189.210 20.500 ;
      LAYER via ;
        RECT 1224.340 45.600 1224.600 45.860 ;
        RECT 1271.260 45.600 1271.520 45.860 ;
        RECT 1272.640 45.600 1272.900 45.860 ;
        RECT 1390.400 45.600 1390.660 45.860 ;
        RECT 1182.480 20.440 1182.740 20.700 ;
        RECT 1188.920 20.440 1189.180 20.700 ;
      LAYER met2 ;
        RECT 1188.910 45.715 1189.190 46.085 ;
        RECT 1224.330 45.715 1224.610 46.085 ;
        RECT 1271.250 45.715 1271.530 46.085 ;
        RECT 1272.630 45.715 1272.910 46.085 ;
        RECT 1390.460 45.890 1390.600 54.000 ;
        RECT 1188.980 20.730 1189.120 45.715 ;
        RECT 1224.340 45.570 1224.600 45.715 ;
        RECT 1271.260 45.570 1271.520 45.715 ;
        RECT 1272.640 45.570 1272.900 45.715 ;
        RECT 1390.400 45.570 1390.660 45.890 ;
        RECT 1182.480 20.410 1182.740 20.730 ;
        RECT 1188.920 20.410 1189.180 20.730 ;
        RECT 1182.540 2.400 1182.680 20.410 ;
        RECT 1182.470 0.000 1182.750 2.400 ;
      LAYER via2 ;
        RECT 1188.910 45.760 1189.190 46.040 ;
        RECT 1224.330 45.760 1224.610 46.040 ;
        RECT 1271.250 45.760 1271.530 46.040 ;
        RECT 1272.630 45.760 1272.910 46.040 ;
      LAYER met3 ;
        RECT 1188.885 46.050 1189.215 46.065 ;
        RECT 1224.305 46.050 1224.635 46.065 ;
        RECT 1188.885 45.750 1224.635 46.050 ;
        RECT 1188.885 45.735 1189.215 45.750 ;
        RECT 1224.305 45.735 1224.635 45.750 ;
        RECT 1271.225 46.050 1271.555 46.065 ;
        RECT 1272.605 46.050 1272.935 46.065 ;
        RECT 1271.225 45.750 1272.935 46.050 ;
        RECT 1271.225 45.735 1271.555 45.750 ;
        RECT 1272.605 45.735 1272.935 45.750 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1224.310 46.820 1224.630 46.880 ;
        RECT 1398.190 46.820 1398.510 46.880 ;
        RECT 1224.310 46.680 1398.510 46.820 ;
        RECT 1224.310 46.620 1224.630 46.680 ;
        RECT 1398.190 46.620 1398.510 46.680 ;
      LAYER via ;
        RECT 1224.340 46.620 1224.600 46.880 ;
        RECT 1398.220 46.620 1398.480 46.880 ;
      LAYER met2 ;
        RECT 1398.280 46.910 1398.420 54.000 ;
        RECT 1224.340 46.765 1224.600 46.910 ;
        RECT 1200.410 46.395 1200.690 46.765 ;
        RECT 1224.330 46.395 1224.610 46.765 ;
        RECT 1398.220 46.590 1398.480 46.910 ;
        RECT 1200.480 2.400 1200.620 46.395 ;
        RECT 1200.410 0.000 1200.690 2.400 ;
      LAYER via2 ;
        RECT 1200.410 46.440 1200.690 46.720 ;
        RECT 1224.330 46.440 1224.610 46.720 ;
      LAYER met3 ;
        RECT 1200.385 46.730 1200.715 46.745 ;
        RECT 1224.305 46.730 1224.635 46.745 ;
        RECT 1200.385 46.430 1224.635 46.730 ;
        RECT 1200.385 46.415 1200.715 46.430 ;
        RECT 1224.305 46.415 1224.635 46.430 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1344.445 14.025 1344.615 17.935 ;
      LAYER mcon ;
        RECT 1344.445 17.765 1344.615 17.935 ;
      LAYER met1 ;
        RECT 1218.330 18.260 1218.650 18.320 ;
        RECT 1218.330 18.120 1236.040 18.260 ;
        RECT 1218.330 18.060 1218.650 18.120 ;
        RECT 1235.900 17.920 1236.040 18.120 ;
        RECT 1344.385 17.920 1344.675 17.965 ;
        RECT 1235.900 17.780 1344.675 17.920 ;
        RECT 1344.385 17.735 1344.675 17.780 ;
        RECT 1344.385 14.180 1344.675 14.225 ;
        RECT 1396.350 14.180 1396.670 14.240 ;
        RECT 1344.385 14.040 1396.670 14.180 ;
        RECT 1344.385 13.995 1344.675 14.040 ;
        RECT 1396.350 13.980 1396.670 14.040 ;
      LAYER via ;
        RECT 1218.360 18.060 1218.620 18.320 ;
        RECT 1396.380 13.980 1396.640 14.240 ;
      LAYER met2 ;
        RECT 1218.360 18.030 1218.620 18.350 ;
        RECT 1218.420 2.400 1218.560 18.030 ;
        RECT 1396.440 14.270 1396.580 54.000 ;
        RECT 1396.380 13.950 1396.640 14.270 ;
        RECT 1218.350 0.000 1218.630 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1236.270 18.260 1236.590 18.320 ;
        RECT 1236.270 18.120 1393.360 18.260 ;
        RECT 1236.270 18.060 1236.590 18.120 ;
        RECT 1393.220 17.920 1393.360 18.120 ;
        RECT 1405.090 17.920 1405.410 17.980 ;
        RECT 1393.220 17.780 1405.410 17.920 ;
        RECT 1405.090 17.720 1405.410 17.780 ;
      LAYER via ;
        RECT 1236.300 18.060 1236.560 18.320 ;
        RECT 1405.120 17.720 1405.380 17.980 ;
      LAYER met2 ;
        RECT 1236.300 18.030 1236.560 18.350 ;
        RECT 1236.360 2.400 1236.500 18.030 ;
        RECT 1405.180 18.010 1405.320 54.000 ;
        RECT 1405.120 17.690 1405.380 18.010 ;
        RECT 1236.290 0.000 1236.570 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1254.210 15.200 1254.530 15.260 ;
        RECT 1257.890 15.200 1258.210 15.260 ;
        RECT 1254.210 15.060 1258.210 15.200 ;
        RECT 1254.210 15.000 1254.530 15.060 ;
        RECT 1257.890 15.000 1258.210 15.060 ;
      LAYER via ;
        RECT 1254.240 15.000 1254.500 15.260 ;
        RECT 1257.920 15.000 1258.180 15.260 ;
      LAYER met2 ;
        RECT 1257.980 15.290 1258.120 54.000 ;
        RECT 1254.240 14.970 1254.500 15.290 ;
        RECT 1257.920 14.970 1258.180 15.290 ;
        RECT 1254.300 2.400 1254.440 14.970 ;
        RECT 1254.230 0.000 1254.510 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1271.780 2.400 1271.920 54.000 ;
        RECT 1271.710 0.000 1271.990 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1393.205 17.255 1393.375 17.595 ;
        RECT 1378.485 15.045 1378.655 17.255 ;
        RECT 1392.285 17.085 1393.375 17.255 ;
        RECT 1392.285 15.045 1392.455 17.085 ;
      LAYER mcon ;
        RECT 1393.205 17.425 1393.375 17.595 ;
        RECT 1378.485 17.085 1378.655 17.255 ;
      LAYER met1 ;
        RECT 1393.145 17.580 1393.435 17.625 ;
        RECT 1411.530 17.580 1411.850 17.640 ;
        RECT 1393.145 17.440 1411.850 17.580 ;
        RECT 1393.145 17.395 1393.435 17.440 ;
        RECT 1411.530 17.380 1411.850 17.440 ;
        RECT 1378.425 17.240 1378.715 17.285 ;
        RECT 1313.640 17.100 1378.715 17.240 ;
        RECT 1289.630 16.900 1289.950 16.960 ;
        RECT 1313.640 16.900 1313.780 17.100 ;
        RECT 1378.425 17.055 1378.715 17.100 ;
        RECT 1289.630 16.760 1313.780 16.900 ;
        RECT 1289.630 16.700 1289.950 16.760 ;
        RECT 1378.425 15.200 1378.715 15.245 ;
        RECT 1392.225 15.200 1392.515 15.245 ;
        RECT 1378.425 15.060 1392.515 15.200 ;
        RECT 1378.425 15.015 1378.715 15.060 ;
        RECT 1392.225 15.015 1392.515 15.060 ;
      LAYER via ;
        RECT 1411.560 17.380 1411.820 17.640 ;
        RECT 1289.660 16.700 1289.920 16.960 ;
      LAYER met2 ;
        RECT 1411.620 17.670 1411.760 54.000 ;
        RECT 1411.560 17.350 1411.820 17.670 ;
        RECT 1289.660 16.670 1289.920 16.990 ;
        RECT 1289.720 2.400 1289.860 16.670 ;
        RECT 1289.650 0.000 1289.930 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1307.570 17.240 1307.890 17.300 ;
        RECT 1313.090 17.240 1313.410 17.300 ;
        RECT 1307.570 17.100 1313.410 17.240 ;
        RECT 1307.570 17.040 1307.890 17.100 ;
        RECT 1313.090 17.040 1313.410 17.100 ;
      LAYER via ;
        RECT 1307.600 17.040 1307.860 17.300 ;
        RECT 1313.120 17.040 1313.380 17.300 ;
      LAYER met2 ;
        RECT 1313.180 17.330 1313.320 54.000 ;
        RECT 1307.600 17.010 1307.860 17.330 ;
        RECT 1313.120 17.010 1313.380 17.330 ;
        RECT 1307.660 2.400 1307.800 17.010 ;
        RECT 1307.590 0.000 1307.870 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1393.665 17.935 1393.835 18.275 ;
        RECT 1392.745 17.765 1393.835 17.935 ;
        RECT 1392.745 17.425 1392.915 17.765 ;
      LAYER mcon ;
        RECT 1393.665 18.105 1393.835 18.275 ;
      LAYER met1 ;
        RECT 1393.605 18.260 1393.895 18.305 ;
        RECT 1425.790 18.260 1426.110 18.320 ;
        RECT 1393.605 18.120 1426.110 18.260 ;
        RECT 1393.605 18.075 1393.895 18.120 ;
        RECT 1425.790 18.060 1426.110 18.120 ;
        RECT 1325.510 17.580 1325.830 17.640 ;
        RECT 1392.685 17.580 1392.975 17.625 ;
        RECT 1325.510 17.440 1392.975 17.580 ;
        RECT 1325.510 17.380 1325.830 17.440 ;
        RECT 1392.685 17.395 1392.975 17.440 ;
      LAYER via ;
        RECT 1425.820 18.060 1426.080 18.320 ;
        RECT 1325.540 17.380 1325.800 17.640 ;
      LAYER met2 ;
        RECT 1425.880 18.350 1426.020 54.000 ;
        RECT 1425.820 18.030 1426.080 18.350 ;
        RECT 1325.540 17.350 1325.800 17.670 ;
        RECT 1325.600 2.400 1325.740 17.350 ;
        RECT 1325.530 0.000 1325.810 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1419.885 19.635 1420.055 20.315 ;
        RECT 1419.885 19.465 1420.975 19.635 ;
      LAYER mcon ;
        RECT 1419.885 20.145 1420.055 20.315 ;
        RECT 1420.805 19.465 1420.975 19.635 ;
      LAYER met1 ;
        RECT 1425.330 48.520 1425.650 48.580 ;
        RECT 1426.250 48.520 1426.570 48.580 ;
        RECT 1425.330 48.380 1426.570 48.520 ;
        RECT 1425.330 48.320 1425.650 48.380 ;
        RECT 1426.250 48.320 1426.570 48.380 ;
        RECT 1342.990 20.300 1343.310 20.360 ;
        RECT 1419.825 20.300 1420.115 20.345 ;
        RECT 1342.990 20.160 1420.115 20.300 ;
        RECT 1342.990 20.100 1343.310 20.160 ;
        RECT 1419.825 20.115 1420.115 20.160 ;
        RECT 1420.745 19.620 1421.035 19.665 ;
        RECT 1426.250 19.620 1426.570 19.680 ;
        RECT 1420.745 19.480 1426.570 19.620 ;
        RECT 1420.745 19.435 1421.035 19.480 ;
        RECT 1426.250 19.420 1426.570 19.480 ;
      LAYER via ;
        RECT 1425.360 48.320 1425.620 48.580 ;
        RECT 1426.280 48.320 1426.540 48.580 ;
        RECT 1343.020 20.100 1343.280 20.360 ;
        RECT 1426.280 19.420 1426.540 19.680 ;
      LAYER met2 ;
        RECT 1425.420 48.610 1425.560 54.000 ;
        RECT 1425.360 48.290 1425.620 48.610 ;
        RECT 1426.280 48.290 1426.540 48.610 ;
        RECT 1343.020 20.070 1343.280 20.390 ;
        RECT 1343.080 2.400 1343.220 20.070 ;
        RECT 1426.340 19.710 1426.480 48.290 ;
        RECT 1426.280 19.390 1426.540 19.710 ;
        RECT 1343.010 0.000 1343.290 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1224.385 46.835 1224.555 47.515 ;
        RECT 740.465 44.965 740.635 46.835 ;
        RECT 1223.925 46.665 1224.555 46.835 ;
      LAYER mcon ;
        RECT 1224.385 47.345 1224.555 47.515 ;
        RECT 740.465 46.665 740.635 46.835 ;
      LAYER met1 ;
        RECT 1224.325 47.500 1224.615 47.545 ;
        RECT 1295.150 47.500 1295.470 47.560 ;
        RECT 1224.325 47.360 1295.470 47.500 ;
        RECT 1224.325 47.315 1224.615 47.360 ;
        RECT 1295.150 47.300 1295.470 47.360 ;
        RECT 740.405 46.820 740.695 46.865 ;
        RECT 1223.865 46.820 1224.155 46.865 ;
        RECT 740.405 46.680 1224.155 46.820 ;
        RECT 740.405 46.635 740.695 46.680 ;
        RECT 1223.865 46.635 1224.155 46.680 ;
        RECT 700.830 45.120 701.150 45.180 ;
        RECT 740.405 45.120 740.695 45.165 ;
        RECT 700.830 44.980 740.695 45.120 ;
        RECT 700.830 44.920 701.150 44.980 ;
        RECT 740.405 44.935 740.695 44.980 ;
      LAYER via ;
        RECT 1295.180 47.300 1295.440 47.560 ;
        RECT 700.860 44.920 701.120 45.180 ;
      LAYER met2 ;
        RECT 1295.240 47.590 1295.380 54.000 ;
        RECT 1295.180 47.270 1295.440 47.590 ;
        RECT 700.860 44.890 701.120 45.210 ;
        RECT 700.920 2.400 701.060 44.890 ;
        RECT 700.850 0.000 701.130 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1392.745 15.045 1392.915 16.915 ;
      LAYER mcon ;
        RECT 1392.745 16.745 1392.915 16.915 ;
      LAYER met1 ;
        RECT 1360.930 16.900 1361.250 16.960 ;
        RECT 1392.685 16.900 1392.975 16.945 ;
        RECT 1360.930 16.760 1392.975 16.900 ;
        RECT 1360.930 16.700 1361.250 16.760 ;
        RECT 1392.685 16.715 1392.975 16.760 ;
        RECT 1392.685 15.200 1392.975 15.245 ;
        RECT 1431.770 15.200 1432.090 15.260 ;
        RECT 1392.685 15.060 1432.090 15.200 ;
        RECT 1392.685 15.015 1392.975 15.060 ;
        RECT 1431.770 15.000 1432.090 15.060 ;
      LAYER via ;
        RECT 1360.960 16.700 1361.220 16.960 ;
        RECT 1431.800 15.000 1432.060 15.260 ;
      LAYER met2 ;
        RECT 1360.960 16.670 1361.220 16.990 ;
        RECT 1361.020 2.400 1361.160 16.670 ;
        RECT 1431.860 15.290 1432.000 54.000 ;
        RECT 1431.800 14.970 1432.060 15.290 ;
        RECT 1360.950 0.000 1361.230 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1378.870 17.240 1379.190 17.300 ;
        RECT 1378.870 17.100 1393.360 17.240 ;
        RECT 1378.870 17.040 1379.190 17.100 ;
        RECT 1393.220 16.900 1393.360 17.100 ;
        RECT 1433.610 16.900 1433.930 16.960 ;
        RECT 1393.220 16.760 1433.930 16.900 ;
        RECT 1433.610 16.700 1433.930 16.760 ;
      LAYER via ;
        RECT 1378.900 17.040 1379.160 17.300 ;
        RECT 1433.640 16.700 1433.900 16.960 ;
      LAYER met2 ;
        RECT 1378.900 17.010 1379.160 17.330 ;
        RECT 1378.960 2.400 1379.100 17.010 ;
        RECT 1433.700 16.990 1433.840 54.000 ;
        RECT 1433.640 16.670 1433.900 16.990 ;
        RECT 1378.890 0.000 1379.170 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1400.490 17.240 1400.810 17.300 ;
        RECT 1440.510 17.240 1440.830 17.300 ;
        RECT 1400.490 17.100 1440.830 17.240 ;
        RECT 1400.490 17.040 1400.810 17.100 ;
        RECT 1440.510 17.040 1440.830 17.100 ;
      LAYER via ;
        RECT 1400.520 17.040 1400.780 17.300 ;
        RECT 1440.540 17.040 1440.800 17.300 ;
      LAYER met2 ;
        RECT 1440.600 17.330 1440.740 54.000 ;
        RECT 1400.520 17.010 1400.780 17.330 ;
        RECT 1440.540 17.010 1440.800 17.330 ;
        RECT 1400.580 9.250 1400.720 17.010 ;
        RECT 1396.900 9.110 1400.720 9.250 ;
        RECT 1396.900 2.400 1397.040 9.110 ;
        RECT 1396.830 0.000 1397.110 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1414.750 17.920 1415.070 17.980 ;
        RECT 1439.590 17.920 1439.910 17.980 ;
        RECT 1414.750 17.780 1439.910 17.920 ;
        RECT 1414.750 17.720 1415.070 17.780 ;
        RECT 1439.590 17.720 1439.910 17.780 ;
      LAYER via ;
        RECT 1414.780 17.720 1415.040 17.980 ;
        RECT 1439.620 17.720 1439.880 17.980 ;
      LAYER met2 ;
        RECT 1439.680 18.010 1439.820 54.000 ;
        RECT 1414.780 17.690 1415.040 18.010 ;
        RECT 1439.620 17.690 1439.880 18.010 ;
        RECT 1414.840 2.400 1414.980 17.690 ;
        RECT 1414.770 0.000 1415.050 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1432.230 19.960 1432.550 20.020 ;
        RECT 1445.570 19.960 1445.890 20.020 ;
        RECT 1432.230 19.820 1445.890 19.960 ;
        RECT 1432.230 19.760 1432.550 19.820 ;
        RECT 1445.570 19.760 1445.890 19.820 ;
      LAYER via ;
        RECT 1432.260 19.760 1432.520 20.020 ;
        RECT 1445.600 19.760 1445.860 20.020 ;
      LAYER met2 ;
        RECT 1445.660 20.050 1445.800 54.000 ;
        RECT 1432.260 19.730 1432.520 20.050 ;
        RECT 1445.600 19.730 1445.860 20.050 ;
        RECT 1432.320 2.400 1432.460 19.730 ;
        RECT 1432.250 0.000 1432.530 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1447.870 20.640 1448.190 20.700 ;
        RECT 1450.170 20.640 1450.490 20.700 ;
        RECT 1447.870 20.500 1450.490 20.640 ;
        RECT 1447.870 20.440 1448.190 20.500 ;
        RECT 1450.170 20.440 1450.490 20.500 ;
      LAYER via ;
        RECT 1447.900 20.440 1448.160 20.700 ;
        RECT 1450.200 20.440 1450.460 20.700 ;
      LAYER met2 ;
        RECT 1447.960 20.730 1448.100 54.000 ;
        RECT 1447.900 20.410 1448.160 20.730 ;
        RECT 1450.200 20.410 1450.460 20.730 ;
        RECT 1450.260 2.400 1450.400 20.410 ;
        RECT 1450.190 0.000 1450.470 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1457.070 17.240 1457.390 17.300 ;
        RECT 1468.110 17.240 1468.430 17.300 ;
        RECT 1457.070 17.100 1468.430 17.240 ;
        RECT 1457.070 17.040 1457.390 17.100 ;
        RECT 1468.110 17.040 1468.430 17.100 ;
      LAYER via ;
        RECT 1457.100 17.040 1457.360 17.300 ;
        RECT 1468.140 17.040 1468.400 17.300 ;
      LAYER met2 ;
        RECT 1457.160 17.330 1457.300 54.000 ;
        RECT 1457.100 17.010 1457.360 17.330 ;
        RECT 1468.140 17.010 1468.400 17.330 ;
        RECT 1468.200 2.400 1468.340 17.010 ;
        RECT 1468.130 0.000 1468.410 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1469.490 20.640 1469.810 20.700 ;
        RECT 1486.050 20.640 1486.370 20.700 ;
        RECT 1469.490 20.500 1486.370 20.640 ;
        RECT 1469.490 20.440 1469.810 20.500 ;
        RECT 1486.050 20.440 1486.370 20.500 ;
      LAYER via ;
        RECT 1469.520 20.440 1469.780 20.700 ;
        RECT 1486.080 20.440 1486.340 20.700 ;
      LAYER met2 ;
        RECT 1469.580 20.730 1469.720 54.000 ;
        RECT 1469.520 20.410 1469.780 20.730 ;
        RECT 1486.080 20.410 1486.340 20.730 ;
        RECT 1486.140 2.400 1486.280 20.410 ;
        RECT 1486.070 0.000 1486.350 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1463.510 17.580 1463.830 17.640 ;
        RECT 1503.990 17.580 1504.310 17.640 ;
        RECT 1463.510 17.440 1504.310 17.580 ;
        RECT 1463.510 17.380 1463.830 17.440 ;
        RECT 1503.990 17.380 1504.310 17.440 ;
      LAYER via ;
        RECT 1463.540 17.380 1463.800 17.640 ;
        RECT 1504.020 17.380 1504.280 17.640 ;
      LAYER met2 ;
        RECT 1463.600 17.670 1463.740 54.000 ;
        RECT 1463.540 17.350 1463.800 17.670 ;
        RECT 1504.020 17.350 1504.280 17.670 ;
        RECT 1504.080 2.400 1504.220 17.350 ;
        RECT 1504.010 0.000 1504.290 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1492.565 16.745 1492.735 19.635 ;
      LAYER mcon ;
        RECT 1492.565 19.465 1492.735 19.635 ;
      LAYER met1 ;
        RECT 1521.470 19.960 1521.790 20.020 ;
        RECT 1512.820 19.820 1521.790 19.960 ;
        RECT 1492.505 19.620 1492.795 19.665 ;
        RECT 1512.820 19.620 1512.960 19.820 ;
        RECT 1521.470 19.760 1521.790 19.820 ;
        RECT 1492.505 19.480 1512.960 19.620 ;
        RECT 1492.505 19.435 1492.795 19.480 ;
        RECT 1468.570 16.900 1468.890 16.960 ;
        RECT 1492.505 16.900 1492.795 16.945 ;
        RECT 1468.570 16.760 1492.795 16.900 ;
        RECT 1468.570 16.700 1468.890 16.760 ;
        RECT 1492.505 16.715 1492.795 16.760 ;
      LAYER via ;
        RECT 1521.500 19.760 1521.760 20.020 ;
        RECT 1468.600 16.700 1468.860 16.960 ;
      LAYER met2 ;
        RECT 1468.660 16.990 1468.800 54.000 ;
        RECT 1521.500 19.730 1521.760 20.050 ;
        RECT 1468.600 16.670 1468.860 16.990 ;
        RECT 1521.560 2.400 1521.700 19.730 ;
        RECT 1521.490 0.000 1521.770 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1296.070 47.160 1296.390 47.220 ;
        RECT 740.020 47.020 1296.390 47.160 ;
        RECT 718.770 46.820 719.090 46.880 ;
        RECT 740.020 46.820 740.160 47.020 ;
        RECT 1296.070 46.960 1296.390 47.020 ;
        RECT 718.770 46.680 740.160 46.820 ;
        RECT 718.770 46.620 719.090 46.680 ;
      LAYER via ;
        RECT 718.800 46.620 719.060 46.880 ;
        RECT 1296.100 46.960 1296.360 47.220 ;
      LAYER met2 ;
        RECT 1296.160 47.250 1296.300 54.000 ;
        RECT 1296.100 46.930 1296.360 47.250 ;
        RECT 718.800 46.590 719.060 46.910 ;
        RECT 718.860 2.400 719.000 46.590 ;
        RECT 718.790 0.000 719.070 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1504.985 17.085 1505.155 17.935 ;
      LAYER mcon ;
        RECT 1504.985 17.765 1505.155 17.935 ;
      LAYER met1 ;
        RECT 1504.925 17.920 1505.215 17.965 ;
        RECT 1539.410 17.920 1539.730 17.980 ;
        RECT 1504.925 17.780 1539.730 17.920 ;
        RECT 1504.925 17.735 1505.215 17.780 ;
        RECT 1539.410 17.720 1539.730 17.780 ;
        RECT 1471.790 17.240 1472.110 17.300 ;
        RECT 1504.925 17.240 1505.215 17.285 ;
        RECT 1471.790 17.100 1505.215 17.240 ;
        RECT 1471.790 17.040 1472.110 17.100 ;
        RECT 1504.925 17.055 1505.215 17.100 ;
      LAYER via ;
        RECT 1539.440 17.720 1539.700 17.980 ;
        RECT 1471.820 17.040 1472.080 17.300 ;
      LAYER met2 ;
        RECT 1471.880 17.330 1472.020 54.000 ;
        RECT 1539.440 17.690 1539.700 18.010 ;
        RECT 1471.820 17.010 1472.080 17.330 ;
        RECT 1539.500 2.400 1539.640 17.690 ;
        RECT 1539.430 0.000 1539.710 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1498.545 18.445 1498.715 20.315 ;
      LAYER mcon ;
        RECT 1498.545 20.145 1498.715 20.315 ;
      LAYER met1 ;
        RECT 1471.330 20.300 1471.650 20.360 ;
        RECT 1498.485 20.300 1498.775 20.345 ;
        RECT 1471.330 20.160 1498.775 20.300 ;
        RECT 1471.330 20.100 1471.650 20.160 ;
        RECT 1498.485 20.115 1498.775 20.160 ;
        RECT 1498.485 18.600 1498.775 18.645 ;
        RECT 1557.350 18.600 1557.670 18.660 ;
        RECT 1498.485 18.460 1557.670 18.600 ;
        RECT 1498.485 18.415 1498.775 18.460 ;
        RECT 1557.350 18.400 1557.670 18.460 ;
      LAYER via ;
        RECT 1471.360 20.100 1471.620 20.360 ;
        RECT 1557.380 18.400 1557.640 18.660 ;
      LAYER met2 ;
        RECT 1471.420 20.390 1471.560 54.000 ;
        RECT 1471.360 20.070 1471.620 20.390 ;
        RECT 1557.380 18.370 1557.640 18.690 ;
        RECT 1557.440 2.400 1557.580 18.370 ;
        RECT 1557.370 0.000 1557.650 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1570.780 14.180 1570.920 54.000 ;
        RECT 1570.780 14.040 1575.520 14.180 ;
        RECT 1575.380 2.400 1575.520 14.040 ;
        RECT 1575.310 0.000 1575.590 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1485.590 17.920 1485.910 17.980 ;
        RECT 1485.590 17.780 1504.680 17.920 ;
        RECT 1485.590 17.720 1485.910 17.780 ;
        RECT 1504.540 17.580 1504.680 17.780 ;
        RECT 1592.770 17.580 1593.090 17.640 ;
        RECT 1504.540 17.440 1593.090 17.580 ;
        RECT 1592.770 17.380 1593.090 17.440 ;
      LAYER via ;
        RECT 1485.620 17.720 1485.880 17.980 ;
        RECT 1592.800 17.380 1593.060 17.640 ;
      LAYER met2 ;
        RECT 1485.680 18.010 1485.820 54.000 ;
        RECT 1485.620 17.690 1485.880 18.010 ;
        RECT 1592.800 17.350 1593.060 17.670 ;
        RECT 1592.860 2.400 1593.000 17.350 ;
        RECT 1592.790 0.000 1593.070 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1610.340 3.130 1610.480 54.000 ;
        RECT 1610.340 2.990 1610.940 3.130 ;
        RECT 1610.800 2.400 1610.940 2.990 ;
        RECT 1610.730 0.000 1611.010 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1624.050 2.960 1624.370 3.020 ;
        RECT 1628.650 2.960 1628.970 3.020 ;
        RECT 1624.050 2.820 1628.970 2.960 ;
        RECT 1624.050 2.760 1624.370 2.820 ;
        RECT 1628.650 2.760 1628.970 2.820 ;
      LAYER via ;
        RECT 1624.080 2.760 1624.340 3.020 ;
        RECT 1628.680 2.760 1628.940 3.020 ;
      LAYER met2 ;
        RECT 1624.140 3.050 1624.280 54.000 ;
        RECT 1624.080 2.730 1624.340 3.050 ;
        RECT 1628.680 2.730 1628.940 3.050 ;
        RECT 1628.740 2.400 1628.880 2.730 ;
        RECT 1628.670 0.000 1628.950 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1644.840 14.010 1644.980 54.000 ;
        RECT 1644.840 13.870 1646.360 14.010 ;
        RECT 1646.220 13.330 1646.360 13.870 ;
        RECT 1646.220 13.190 1646.820 13.330 ;
        RECT 1646.680 2.400 1646.820 13.190 ;
        RECT 1646.610 0.000 1646.890 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1658.550 37.640 1658.870 37.700 ;
        RECT 1664.530 37.640 1664.850 37.700 ;
        RECT 1658.550 37.500 1664.850 37.640 ;
        RECT 1658.550 37.440 1658.870 37.500 ;
        RECT 1664.530 37.440 1664.850 37.500 ;
      LAYER via ;
        RECT 1658.580 37.440 1658.840 37.700 ;
        RECT 1664.560 37.440 1664.820 37.700 ;
      LAYER met2 ;
        RECT 1658.640 37.730 1658.780 54.000 ;
        RECT 1658.580 37.410 1658.840 37.730 ;
        RECT 1664.560 37.410 1664.820 37.730 ;
        RECT 1664.620 2.400 1664.760 37.410 ;
        RECT 1664.550 0.000 1664.830 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1680.720 24.210 1680.860 54.000 ;
        RECT 1680.720 24.070 1682.240 24.210 ;
        RECT 1682.100 2.400 1682.240 24.070 ;
        RECT 1682.030 0.000 1682.310 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1700.040 2.400 1700.180 54.000 ;
        RECT 1699.970 0.000 1700.250 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1224.845 47.855 1225.015 48.535 ;
        RECT 1223.925 47.685 1225.015 47.855 ;
        RECT 1223.925 47.345 1224.095 47.685 ;
        RECT 1271.765 45.645 1271.935 48.535 ;
      LAYER mcon ;
        RECT 1224.845 48.365 1225.015 48.535 ;
        RECT 1271.765 48.365 1271.935 48.535 ;
      LAYER met1 ;
        RECT 1224.785 48.520 1225.075 48.565 ;
        RECT 1271.705 48.520 1271.995 48.565 ;
        RECT 1224.785 48.380 1271.995 48.520 ;
        RECT 1224.785 48.335 1225.075 48.380 ;
        RECT 1271.705 48.335 1271.995 48.380 ;
        RECT 736.710 47.500 737.030 47.560 ;
        RECT 1223.865 47.500 1224.155 47.545 ;
        RECT 736.710 47.360 1224.155 47.500 ;
        RECT 736.710 47.300 737.030 47.360 ;
        RECT 1223.865 47.315 1224.155 47.360 ;
        RECT 1271.705 45.800 1271.995 45.845 ;
        RECT 1272.150 45.800 1272.470 45.860 ;
        RECT 1271.705 45.660 1272.470 45.800 ;
        RECT 1271.705 45.615 1271.995 45.660 ;
        RECT 1272.150 45.600 1272.470 45.660 ;
        RECT 1274.450 44.100 1274.770 44.160 ;
        RECT 1302.050 44.100 1302.370 44.160 ;
        RECT 1274.450 43.960 1302.370 44.100 ;
        RECT 1274.450 43.900 1274.770 43.960 ;
        RECT 1302.050 43.900 1302.370 43.960 ;
      LAYER via ;
        RECT 736.740 47.300 737.000 47.560 ;
        RECT 1272.180 45.600 1272.440 45.860 ;
        RECT 1274.480 43.900 1274.740 44.160 ;
        RECT 1302.080 43.900 1302.340 44.160 ;
      LAYER met2 ;
        RECT 736.740 47.270 737.000 47.590 ;
        RECT 736.800 2.400 736.940 47.270 ;
        RECT 1272.180 45.570 1272.440 45.890 ;
        RECT 1272.240 44.725 1272.380 45.570 ;
        RECT 1272.170 44.355 1272.450 44.725 ;
        RECT 1274.470 44.355 1274.750 44.725 ;
        RECT 1274.540 44.190 1274.680 44.355 ;
        RECT 1302.140 44.190 1302.280 54.000 ;
        RECT 1274.480 43.870 1274.740 44.190 ;
        RECT 1302.080 43.870 1302.340 44.190 ;
        RECT 736.730 0.000 737.010 2.400 ;
      LAYER via2 ;
        RECT 1272.170 44.400 1272.450 44.680 ;
        RECT 1274.470 44.400 1274.750 44.680 ;
      LAYER met3 ;
        RECT 1272.145 44.690 1272.475 44.705 ;
        RECT 1274.445 44.690 1274.775 44.705 ;
        RECT 1272.145 44.390 1274.775 44.690 ;
        RECT 1272.145 44.375 1272.475 44.390 ;
        RECT 1274.445 44.375 1274.775 44.390 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1713.840 25.570 1713.980 54.000 ;
        RECT 1713.840 25.430 1718.120 25.570 ;
        RECT 1717.980 2.400 1718.120 25.430 ;
        RECT 1717.910 0.000 1718.190 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1735.460 48.805 1735.600 54.000 ;
        RECT 1734.470 48.435 1734.750 48.805 ;
        RECT 1735.390 48.435 1735.670 48.805 ;
        RECT 1734.540 14.010 1734.680 48.435 ;
        RECT 1734.540 13.870 1735.600 14.010 ;
        RECT 1735.460 13.330 1735.600 13.870 ;
        RECT 1735.460 13.190 1736.060 13.330 ;
        RECT 1735.920 2.400 1736.060 13.190 ;
        RECT 1735.850 0.000 1736.130 2.400 ;
      LAYER via2 ;
        RECT 1734.470 48.480 1734.750 48.760 ;
        RECT 1735.390 48.480 1735.670 48.760 ;
      LAYER met3 ;
        RECT 1734.445 48.770 1734.775 48.785 ;
        RECT 1735.365 48.770 1735.695 48.785 ;
        RECT 1734.445 48.470 1735.695 48.770 ;
        RECT 1734.445 48.455 1734.775 48.470 ;
        RECT 1735.365 48.455 1735.695 48.470 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1748.250 12.140 1748.570 12.200 ;
        RECT 1753.770 12.140 1754.090 12.200 ;
        RECT 1748.250 12.000 1754.090 12.140 ;
        RECT 1748.250 11.940 1748.570 12.000 ;
        RECT 1753.770 11.940 1754.090 12.000 ;
      LAYER via ;
        RECT 1748.280 11.940 1748.540 12.200 ;
        RECT 1753.800 11.940 1754.060 12.200 ;
      LAYER met2 ;
        RECT 1748.340 12.230 1748.480 54.000 ;
        RECT 1748.280 11.910 1748.540 12.230 ;
        RECT 1753.800 11.910 1754.060 12.230 ;
        RECT 1753.860 2.400 1754.000 11.910 ;
        RECT 1753.790 0.000 1754.070 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1768.950 5.680 1769.270 5.740 ;
        RECT 1771.250 5.680 1771.570 5.740 ;
        RECT 1768.950 5.540 1771.570 5.680 ;
        RECT 1768.950 5.480 1769.270 5.540 ;
        RECT 1771.250 5.480 1771.570 5.540 ;
      LAYER via ;
        RECT 1768.980 5.480 1769.240 5.740 ;
        RECT 1771.280 5.480 1771.540 5.740 ;
      LAYER met2 ;
        RECT 1769.040 5.770 1769.180 54.000 ;
        RECT 1768.980 5.450 1769.240 5.770 ;
        RECT 1771.280 5.450 1771.540 5.770 ;
        RECT 1771.340 2.400 1771.480 5.450 ;
        RECT 1771.270 0.000 1771.550 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1782.750 7.040 1783.070 7.100 ;
        RECT 1789.190 7.040 1789.510 7.100 ;
        RECT 1782.750 6.900 1789.510 7.040 ;
        RECT 1782.750 6.840 1783.070 6.900 ;
        RECT 1789.190 6.840 1789.510 6.900 ;
      LAYER via ;
        RECT 1782.780 6.840 1783.040 7.100 ;
        RECT 1789.220 6.840 1789.480 7.100 ;
      LAYER met2 ;
        RECT 1782.840 7.130 1782.980 54.000 ;
        RECT 1782.780 6.810 1783.040 7.130 ;
        RECT 1789.220 6.810 1789.480 7.130 ;
        RECT 1789.280 2.400 1789.420 6.810 ;
        RECT 1789.210 0.000 1789.490 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1803.450 13.160 1803.770 13.220 ;
        RECT 1807.130 13.160 1807.450 13.220 ;
        RECT 1803.450 13.020 1807.450 13.160 ;
        RECT 1803.450 12.960 1803.770 13.020 ;
        RECT 1807.130 12.960 1807.450 13.020 ;
      LAYER via ;
        RECT 1803.480 12.960 1803.740 13.220 ;
        RECT 1807.160 12.960 1807.420 13.220 ;
      LAYER met2 ;
        RECT 1803.540 13.250 1803.680 54.000 ;
        RECT 1803.480 12.930 1803.740 13.250 ;
        RECT 1807.160 12.930 1807.420 13.250 ;
        RECT 1807.220 2.400 1807.360 12.930 ;
        RECT 1807.150 0.000 1807.430 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1824.240 37.810 1824.380 54.000 ;
        RECT 1824.240 37.670 1825.300 37.810 ;
        RECT 1825.160 2.400 1825.300 37.670 ;
        RECT 1825.090 0.000 1825.370 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1842.180 20.810 1842.320 54.000 ;
        RECT 1842.180 20.670 1842.780 20.810 ;
        RECT 1842.640 2.400 1842.780 20.670 ;
        RECT 1842.570 0.000 1842.850 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1860.120 12.650 1860.260 54.000 ;
        RECT 1860.120 12.510 1860.720 12.650 ;
        RECT 1860.580 2.400 1860.720 12.510 ;
        RECT 1860.510 0.000 1860.790 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1872.450 42.060 1872.770 42.120 ;
        RECT 1878.430 42.060 1878.750 42.120 ;
        RECT 1872.450 41.920 1878.750 42.060 ;
        RECT 1872.450 41.860 1872.770 41.920 ;
        RECT 1878.430 41.860 1878.750 41.920 ;
      LAYER via ;
        RECT 1872.480 41.860 1872.740 42.120 ;
        RECT 1878.460 41.860 1878.720 42.120 ;
      LAYER met2 ;
        RECT 1872.540 42.150 1872.680 54.000 ;
        RECT 1872.480 41.830 1872.740 42.150 ;
        RECT 1878.460 41.830 1878.720 42.150 ;
        RECT 1878.520 2.400 1878.660 41.830 ;
        RECT 1878.450 0.000 1878.730 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 754.650 47.840 754.970 47.900 ;
        RECT 1308.030 47.840 1308.350 47.900 ;
        RECT 754.650 47.700 1308.350 47.840 ;
        RECT 754.650 47.640 754.970 47.700 ;
        RECT 1308.030 47.640 1308.350 47.700 ;
      LAYER via ;
        RECT 754.680 47.640 754.940 47.900 ;
        RECT 1308.060 47.640 1308.320 47.900 ;
      LAYER met2 ;
        RECT 1308.120 47.930 1308.260 54.000 ;
        RECT 754.680 47.610 754.940 47.930 ;
        RECT 1308.060 47.610 1308.320 47.930 ;
        RECT 754.740 2.400 754.880 47.610 ;
        RECT 754.670 0.000 754.950 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1893.150 2.960 1893.470 3.020 ;
        RECT 1896.370 2.960 1896.690 3.020 ;
        RECT 1893.150 2.820 1896.690 2.960 ;
        RECT 1893.150 2.760 1893.470 2.820 ;
        RECT 1896.370 2.760 1896.690 2.820 ;
      LAYER via ;
        RECT 1893.180 2.760 1893.440 3.020 ;
        RECT 1896.400 2.760 1896.660 3.020 ;
      LAYER met2 ;
        RECT 1893.240 3.050 1893.380 54.000 ;
        RECT 1893.180 2.730 1893.440 3.050 ;
        RECT 1896.400 2.730 1896.660 3.050 ;
        RECT 1896.460 2.400 1896.600 2.730 ;
        RECT 1896.390 0.000 1896.670 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1852.285 15.555 1852.455 17.935 ;
        RECT 1852.285 15.385 1873.155 15.555 ;
        RECT 1872.985 13.005 1873.155 15.385 ;
      LAYER mcon ;
        RECT 1852.285 17.765 1852.455 17.935 ;
      LAYER met1 ;
        RECT 1547.690 17.920 1548.010 17.980 ;
        RECT 1852.225 17.920 1852.515 17.965 ;
        RECT 1547.690 17.780 1852.515 17.920 ;
        RECT 1547.690 17.720 1548.010 17.780 ;
        RECT 1852.225 17.735 1852.515 17.780 ;
        RECT 1872.925 13.160 1873.215 13.205 ;
        RECT 1914.310 13.160 1914.630 13.220 ;
        RECT 1872.925 13.020 1914.630 13.160 ;
        RECT 1872.925 12.975 1873.215 13.020 ;
        RECT 1914.310 12.960 1914.630 13.020 ;
      LAYER via ;
        RECT 1547.720 17.720 1547.980 17.980 ;
        RECT 1914.340 12.960 1914.600 13.220 ;
      LAYER met2 ;
        RECT 1547.780 18.010 1547.920 54.000 ;
        RECT 1547.720 17.690 1547.980 18.010 ;
        RECT 1914.340 12.930 1914.600 13.250 ;
        RECT 1914.400 2.400 1914.540 12.930 ;
        RECT 1914.330 0.000 1914.610 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1930.040 48.805 1930.180 54.000 ;
        RECT 1929.970 48.435 1930.250 48.805 ;
        RECT 1931.810 48.435 1932.090 48.805 ;
        RECT 1931.880 2.400 1932.020 48.435 ;
        RECT 1931.810 0.000 1932.090 2.400 ;
      LAYER via2 ;
        RECT 1929.970 48.480 1930.250 48.760 ;
        RECT 1931.810 48.480 1932.090 48.760 ;
      LAYER met3 ;
        RECT 1929.945 48.770 1930.275 48.785 ;
        RECT 1931.785 48.770 1932.115 48.785 ;
        RECT 1929.945 48.470 1932.115 48.770 ;
        RECT 1929.945 48.455 1930.275 48.470 ;
        RECT 1931.785 48.455 1932.115 48.470 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1554.590 17.240 1554.910 17.300 ;
        RECT 1949.730 17.240 1950.050 17.300 ;
        RECT 1554.590 17.100 1950.050 17.240 ;
        RECT 1554.590 17.040 1554.910 17.100 ;
        RECT 1949.730 17.040 1950.050 17.100 ;
      LAYER via ;
        RECT 1554.620 17.040 1554.880 17.300 ;
        RECT 1949.760 17.040 1950.020 17.300 ;
      LAYER met2 ;
        RECT 1554.680 17.330 1554.820 54.000 ;
        RECT 1554.620 17.010 1554.880 17.330 ;
        RECT 1949.760 17.010 1950.020 17.330 ;
        RECT 1949.820 2.400 1949.960 17.010 ;
        RECT 1949.750 0.000 1950.030 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1967.760 2.400 1967.900 54.000 ;
        RECT 1967.690 0.000 1967.970 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1559.650 14.180 1559.970 14.240 ;
        RECT 1823.230 14.180 1823.550 14.240 ;
        RECT 1559.650 14.040 1823.550 14.180 ;
        RECT 1559.650 13.980 1559.970 14.040 ;
        RECT 1823.230 13.980 1823.550 14.040 ;
        RECT 1825.530 14.180 1825.850 14.240 ;
        RECT 1985.610 14.180 1985.930 14.240 ;
        RECT 1825.530 14.040 1985.930 14.180 ;
        RECT 1825.530 13.980 1825.850 14.040 ;
        RECT 1985.610 13.980 1985.930 14.040 ;
      LAYER via ;
        RECT 1559.680 13.980 1559.940 14.240 ;
        RECT 1823.260 13.980 1823.520 14.240 ;
        RECT 1825.560 13.980 1825.820 14.240 ;
        RECT 1985.640 13.980 1985.900 14.240 ;
      LAYER met2 ;
        RECT 1561.580 28.970 1561.720 54.000 ;
        RECT 1559.740 28.830 1561.720 28.970 ;
        RECT 1559.740 14.270 1559.880 28.830 ;
        RECT 1559.680 13.950 1559.940 14.270 ;
        RECT 1823.260 14.125 1823.520 14.270 ;
        RECT 1825.560 14.125 1825.820 14.270 ;
        RECT 1823.250 13.755 1823.530 14.125 ;
        RECT 1825.550 13.755 1825.830 14.125 ;
        RECT 1985.640 13.950 1985.900 14.270 ;
        RECT 1985.700 2.400 1985.840 13.950 ;
        RECT 1985.630 0.000 1985.910 2.400 ;
      LAYER via2 ;
        RECT 1823.250 13.800 1823.530 14.080 ;
        RECT 1825.550 13.800 1825.830 14.080 ;
      LAYER met3 ;
        RECT 1823.225 14.090 1823.555 14.105 ;
        RECT 1825.525 14.090 1825.855 14.105 ;
        RECT 1823.225 13.790 1825.855 14.090 ;
        RECT 1823.225 13.775 1823.555 13.790 ;
        RECT 1825.525 13.775 1825.855 13.790 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2003.640 2.400 2003.780 54.000 ;
        RECT 2003.570 0.000 2003.850 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1568.390 14.520 1568.710 14.580 ;
        RECT 1568.390 14.380 2008.840 14.520 ;
        RECT 1568.390 14.320 1568.710 14.380 ;
        RECT 2008.700 14.180 2008.840 14.380 ;
        RECT 2021.030 14.180 2021.350 14.240 ;
        RECT 2008.700 14.040 2021.350 14.180 ;
        RECT 2021.030 13.980 2021.350 14.040 ;
      LAYER via ;
        RECT 1568.420 14.320 1568.680 14.580 ;
        RECT 2021.060 13.980 2021.320 14.240 ;
      LAYER met2 ;
        RECT 1568.480 14.610 1568.620 54.000 ;
        RECT 1568.420 14.290 1568.680 14.610 ;
        RECT 2021.060 13.950 2021.320 14.270 ;
        RECT 2021.120 2.400 2021.260 13.950 ;
        RECT 2021.050 0.000 2021.330 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2038.140 3.130 2038.280 54.000 ;
        RECT 2038.140 2.990 2039.200 3.130 ;
        RECT 2039.060 2.400 2039.200 2.990 ;
        RECT 2038.990 0.000 2039.270 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1775.465 15.045 1777.015 15.215 ;
        RECT 1775.465 14.705 1775.635 15.045 ;
        RECT 1776.845 14.705 1777.015 15.045 ;
      LAYER met1 ;
        RECT 1575.290 14.860 1575.610 14.920 ;
        RECT 1775.405 14.860 1775.695 14.905 ;
        RECT 1575.290 14.720 1775.695 14.860 ;
        RECT 1575.290 14.660 1575.610 14.720 ;
        RECT 1775.405 14.675 1775.695 14.720 ;
        RECT 1776.785 14.860 1777.075 14.905 ;
        RECT 1776.785 14.720 2020.800 14.860 ;
        RECT 1776.785 14.675 1777.075 14.720 ;
        RECT 2020.660 14.520 2020.800 14.720 ;
        RECT 2056.910 14.520 2057.230 14.580 ;
        RECT 2020.660 14.380 2057.230 14.520 ;
        RECT 2056.910 14.320 2057.230 14.380 ;
      LAYER via ;
        RECT 1575.320 14.660 1575.580 14.920 ;
        RECT 2056.940 14.320 2057.200 14.580 ;
      LAYER met2 ;
        RECT 1575.380 14.950 1575.520 54.000 ;
        RECT 1575.320 14.630 1575.580 14.950 ;
        RECT 2056.940 14.290 2057.200 14.610 ;
        RECT 2057.000 2.400 2057.140 14.290 ;
        RECT 2056.930 0.000 2057.210 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 812.685 42.585 812.855 48.195 ;
        RECT 1273.605 44.285 1273.775 48.535 ;
      LAYER mcon ;
        RECT 1273.605 48.365 1273.775 48.535 ;
        RECT 812.685 48.025 812.855 48.195 ;
      LAYER met1 ;
        RECT 1273.545 48.520 1273.835 48.565 ;
        RECT 1272.240 48.380 1273.835 48.520 ;
        RECT 812.625 48.180 812.915 48.225 ;
        RECT 847.570 48.180 847.890 48.240 ;
        RECT 812.625 48.040 847.890 48.180 ;
        RECT 812.625 47.995 812.915 48.040 ;
        RECT 847.570 47.980 847.890 48.040 ;
        RECT 850.790 48.180 851.110 48.240 ;
        RECT 1272.240 48.180 1272.380 48.380 ;
        RECT 1273.545 48.335 1273.835 48.380 ;
        RECT 850.790 48.040 1272.380 48.180 ;
        RECT 850.790 47.980 851.110 48.040 ;
        RECT 1273.545 44.440 1273.835 44.485 ;
        RECT 1309.410 44.440 1309.730 44.500 ;
        RECT 1273.545 44.300 1309.730 44.440 ;
        RECT 1273.545 44.255 1273.835 44.300 ;
        RECT 1309.410 44.240 1309.730 44.300 ;
        RECT 772.130 42.740 772.450 42.800 ;
        RECT 812.625 42.740 812.915 42.785 ;
        RECT 772.130 42.600 812.915 42.740 ;
        RECT 772.130 42.540 772.450 42.600 ;
        RECT 812.625 42.555 812.915 42.600 ;
      LAYER via ;
        RECT 847.600 47.980 847.860 48.240 ;
        RECT 850.820 47.980 851.080 48.240 ;
        RECT 1309.440 44.240 1309.700 44.500 ;
        RECT 772.160 42.540 772.420 42.800 ;
      LAYER met2 ;
        RECT 847.600 47.950 847.860 48.270 ;
        RECT 850.820 47.950 851.080 48.270 ;
        RECT 847.660 47.445 847.800 47.950 ;
        RECT 850.880 47.445 851.020 47.950 ;
        RECT 847.590 47.075 847.870 47.445 ;
        RECT 850.810 47.075 851.090 47.445 ;
        RECT 1309.500 44.530 1309.640 54.000 ;
        RECT 1309.440 44.210 1309.700 44.530 ;
        RECT 772.160 42.510 772.420 42.830 ;
        RECT 772.220 2.400 772.360 42.510 ;
        RECT 772.150 0.000 772.430 2.400 ;
      LAYER via2 ;
        RECT 847.590 47.120 847.870 47.400 ;
        RECT 850.810 47.120 851.090 47.400 ;
      LAYER met3 ;
        RECT 847.565 47.410 847.895 47.425 ;
        RECT 850.785 47.410 851.115 47.425 ;
        RECT 847.565 47.110 851.115 47.410 ;
        RECT 847.565 47.095 847.895 47.110 ;
        RECT 850.785 47.095 851.115 47.110 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2074.940 2.400 2075.080 54.000 ;
        RECT 2074.870 0.000 2075.150 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1582.190 15.200 1582.510 15.260 ;
        RECT 2092.330 15.200 2092.650 15.260 ;
        RECT 1582.190 15.060 2092.650 15.200 ;
        RECT 1582.190 15.000 1582.510 15.060 ;
        RECT 2092.330 15.000 2092.650 15.060 ;
      LAYER via ;
        RECT 1582.220 15.000 1582.480 15.260 ;
        RECT 2092.360 15.000 2092.620 15.260 ;
      LAYER met2 ;
        RECT 1582.280 15.290 1582.420 54.000 ;
        RECT 1582.220 14.970 1582.480 15.290 ;
        RECT 2092.360 14.970 2092.620 15.290 ;
        RECT 2092.420 2.400 2092.560 14.970 ;
        RECT 2092.350 0.000 2092.630 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1589.090 15.540 1589.410 15.600 ;
        RECT 2110.270 15.540 2110.590 15.600 ;
        RECT 1589.090 15.400 2110.590 15.540 ;
        RECT 1589.090 15.340 1589.410 15.400 ;
        RECT 2110.270 15.340 2110.590 15.400 ;
      LAYER via ;
        RECT 1589.120 15.340 1589.380 15.600 ;
        RECT 2110.300 15.340 2110.560 15.600 ;
      LAYER met2 ;
        RECT 1589.180 15.630 1589.320 54.000 ;
        RECT 1589.120 15.310 1589.380 15.630 ;
        RECT 2110.300 15.310 2110.560 15.630 ;
        RECT 2110.360 2.400 2110.500 15.310 ;
        RECT 2110.290 0.000 2110.570 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1595.990 15.880 1596.310 15.940 ;
        RECT 2128.210 15.880 2128.530 15.940 ;
        RECT 1595.990 15.740 2128.530 15.880 ;
        RECT 1595.990 15.680 1596.310 15.740 ;
        RECT 2128.210 15.680 2128.530 15.740 ;
      LAYER via ;
        RECT 1596.020 15.680 1596.280 15.940 ;
        RECT 2128.240 15.680 2128.500 15.940 ;
      LAYER met2 ;
        RECT 1596.080 15.970 1596.220 54.000 ;
        RECT 1596.020 15.650 1596.280 15.970 ;
        RECT 2128.240 15.650 2128.500 15.970 ;
        RECT 2128.300 2.400 2128.440 15.650 ;
        RECT 2128.230 0.000 2128.510 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1595.530 16.900 1595.850 16.960 ;
        RECT 2146.150 16.900 2146.470 16.960 ;
        RECT 1595.530 16.760 2146.470 16.900 ;
        RECT 1595.530 16.700 1595.850 16.760 ;
        RECT 2146.150 16.700 2146.470 16.760 ;
      LAYER via ;
        RECT 1595.560 16.700 1595.820 16.960 ;
        RECT 2146.180 16.700 2146.440 16.960 ;
      LAYER met2 ;
        RECT 1595.620 16.990 1595.760 54.000 ;
        RECT 1595.560 16.670 1595.820 16.990 ;
        RECT 2146.180 16.670 2146.440 16.990 ;
        RECT 2146.240 2.400 2146.380 16.670 ;
        RECT 2146.170 0.000 2146.450 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1614.465 19.465 1614.635 20.655 ;
        RECT 2093.785 15.045 2093.955 20.655 ;
      LAYER mcon ;
        RECT 1614.465 20.485 1614.635 20.655 ;
        RECT 2093.785 20.485 2093.955 20.655 ;
      LAYER met1 ;
        RECT 1614.405 20.640 1614.695 20.685 ;
        RECT 2093.725 20.640 2094.015 20.685 ;
        RECT 1614.405 20.500 2094.015 20.640 ;
        RECT 1614.405 20.455 1614.695 20.500 ;
        RECT 2093.725 20.455 2094.015 20.500 ;
        RECT 1602.430 19.620 1602.750 19.680 ;
        RECT 1614.405 19.620 1614.695 19.665 ;
        RECT 1602.430 19.480 1614.695 19.620 ;
        RECT 1602.430 19.420 1602.750 19.480 ;
        RECT 1614.405 19.435 1614.695 19.480 ;
        RECT 2164.090 15.540 2164.410 15.600 ;
        RECT 2111.280 15.400 2164.410 15.540 ;
        RECT 2093.725 15.200 2094.015 15.245 ;
        RECT 2111.280 15.200 2111.420 15.400 ;
        RECT 2164.090 15.340 2164.410 15.400 ;
        RECT 2093.725 15.060 2111.420 15.200 ;
        RECT 2093.725 15.015 2094.015 15.060 ;
      LAYER via ;
        RECT 1602.460 19.420 1602.720 19.680 ;
        RECT 2164.120 15.340 2164.380 15.600 ;
      LAYER met2 ;
        RECT 1602.520 19.710 1602.660 54.000 ;
        RECT 1602.460 19.390 1602.720 19.710 ;
        RECT 2164.120 15.310 2164.380 15.630 ;
        RECT 2164.180 2.400 2164.320 15.310 ;
        RECT 2164.110 0.000 2164.390 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1602.890 20.640 1603.210 20.700 ;
        RECT 1602.890 20.500 1614.160 20.640 ;
        RECT 1602.890 20.440 1603.210 20.500 ;
        RECT 1614.020 20.300 1614.160 20.500 ;
        RECT 2181.570 20.300 2181.890 20.360 ;
        RECT 1614.020 20.160 2181.890 20.300 ;
        RECT 2181.570 20.100 2181.890 20.160 ;
      LAYER via ;
        RECT 1602.920 20.440 1603.180 20.700 ;
        RECT 2181.600 20.100 2181.860 20.360 ;
      LAYER met2 ;
        RECT 1602.980 20.730 1603.120 54.000 ;
        RECT 1602.920 20.410 1603.180 20.730 ;
        RECT 2181.600 20.070 2181.860 20.390 ;
        RECT 2181.660 2.400 2181.800 20.070 ;
        RECT 2181.590 0.000 2181.870 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1609.330 19.960 1609.650 20.020 ;
        RECT 2199.510 19.960 2199.830 20.020 ;
        RECT 1609.330 19.820 2199.830 19.960 ;
        RECT 1609.330 19.760 1609.650 19.820 ;
        RECT 2199.510 19.760 2199.830 19.820 ;
      LAYER via ;
        RECT 1609.360 19.760 1609.620 20.020 ;
        RECT 2199.540 19.760 2199.800 20.020 ;
      LAYER met2 ;
        RECT 1609.880 41.210 1610.020 54.000 ;
        RECT 1609.420 41.070 1610.020 41.210 ;
        RECT 1609.420 20.050 1609.560 41.070 ;
        RECT 1609.360 19.730 1609.620 20.050 ;
        RECT 2199.540 19.730 2199.800 20.050 ;
        RECT 2199.600 2.400 2199.740 19.730 ;
        RECT 2199.530 0.000 2199.810 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1630.105 17.425 1630.275 19.635 ;
      LAYER mcon ;
        RECT 1630.105 19.465 1630.275 19.635 ;
      LAYER met1 ;
        RECT 1630.045 19.620 1630.335 19.665 ;
        RECT 2217.450 19.620 2217.770 19.680 ;
        RECT 1630.045 19.480 2217.770 19.620 ;
        RECT 1630.045 19.435 1630.335 19.480 ;
        RECT 2217.450 19.420 2217.770 19.480 ;
        RECT 1608.870 17.580 1609.190 17.640 ;
        RECT 1630.045 17.580 1630.335 17.625 ;
        RECT 1608.870 17.440 1630.335 17.580 ;
        RECT 1608.870 17.380 1609.190 17.440 ;
        RECT 1630.045 17.395 1630.335 17.440 ;
      LAYER via ;
        RECT 2217.480 19.420 2217.740 19.680 ;
        RECT 1608.900 17.380 1609.160 17.640 ;
      LAYER met2 ;
        RECT 1609.420 41.890 1609.560 54.000 ;
        RECT 1608.960 41.750 1609.560 41.890 ;
        RECT 1608.960 17.670 1609.100 41.750 ;
        RECT 2217.480 19.390 2217.740 19.710 ;
        RECT 1608.900 17.350 1609.160 17.670 ;
        RECT 2217.540 2.400 2217.680 19.390 ;
        RECT 2217.470 0.000 2217.750 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1620.905 19.465 1621.075 20.995 ;
        RECT 1658.165 18.445 1658.335 20.995 ;
      LAYER mcon ;
        RECT 1620.905 20.825 1621.075 20.995 ;
        RECT 1658.165 20.825 1658.335 20.995 ;
      LAYER met1 ;
        RECT 1620.845 20.980 1621.135 21.025 ;
        RECT 1658.105 20.980 1658.395 21.025 ;
        RECT 1620.845 20.840 1658.395 20.980 ;
        RECT 1620.845 20.795 1621.135 20.840 ;
        RECT 1658.105 20.795 1658.395 20.840 ;
        RECT 1614.850 19.620 1615.170 19.680 ;
        RECT 1620.845 19.620 1621.135 19.665 ;
        RECT 1614.850 19.480 1621.135 19.620 ;
        RECT 1614.850 19.420 1615.170 19.480 ;
        RECT 1620.845 19.435 1621.135 19.480 ;
        RECT 1658.105 18.600 1658.395 18.645 ;
        RECT 2235.390 18.600 2235.710 18.660 ;
        RECT 1658.105 18.460 2235.710 18.600 ;
        RECT 1658.105 18.415 1658.395 18.460 ;
        RECT 2235.390 18.400 2235.710 18.460 ;
      LAYER via ;
        RECT 1614.880 19.420 1615.140 19.680 ;
        RECT 2235.420 18.400 2235.680 18.660 ;
      LAYER met2 ;
        RECT 1614.480 40.530 1614.620 54.000 ;
        RECT 1614.480 40.390 1615.080 40.530 ;
        RECT 1614.940 19.710 1615.080 40.390 ;
        RECT 1614.880 19.390 1615.140 19.710 ;
        RECT 2235.420 18.370 2235.680 18.690 ;
        RECT 2235.480 2.400 2235.620 18.370 ;
        RECT 2235.410 0.000 2235.690 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 814.525 42.925 814.695 44.455 ;
        RECT 1274.065 43.945 1274.235 48.535 ;
      LAYER mcon ;
        RECT 1274.065 48.365 1274.235 48.535 ;
        RECT 814.525 44.285 814.695 44.455 ;
      LAYER met1 ;
        RECT 1274.005 48.520 1274.295 48.565 ;
        RECT 1274.005 48.380 1288.020 48.520 ;
        RECT 1274.005 48.335 1274.295 48.380 ;
        RECT 1287.880 48.180 1288.020 48.380 ;
        RECT 1314.010 48.180 1314.330 48.240 ;
        RECT 1287.880 48.040 1314.330 48.180 ;
        RECT 1314.010 47.980 1314.330 48.040 ;
        RECT 814.465 44.440 814.755 44.485 ;
        RECT 814.465 44.300 1272.840 44.440 ;
        RECT 814.465 44.255 814.755 44.300 ;
        RECT 1272.700 44.100 1272.840 44.300 ;
        RECT 1274.005 44.100 1274.295 44.145 ;
        RECT 1272.700 43.960 1274.295 44.100 ;
        RECT 1274.005 43.915 1274.295 43.960 ;
        RECT 790.070 43.080 790.390 43.140 ;
        RECT 814.465 43.080 814.755 43.125 ;
        RECT 790.070 42.940 814.755 43.080 ;
        RECT 790.070 42.880 790.390 42.940 ;
        RECT 814.465 42.895 814.755 42.940 ;
      LAYER via ;
        RECT 1314.040 47.980 1314.300 48.240 ;
        RECT 790.100 42.880 790.360 43.140 ;
      LAYER met2 ;
        RECT 1314.100 48.270 1314.240 54.000 ;
        RECT 1314.040 47.950 1314.300 48.270 ;
        RECT 790.100 42.850 790.360 43.170 ;
        RECT 790.160 2.400 790.300 42.850 ;
        RECT 790.090 0.000 790.370 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1616.230 18.260 1616.550 18.320 ;
        RECT 2253.330 18.260 2253.650 18.320 ;
        RECT 1616.230 18.120 2253.650 18.260 ;
        RECT 1616.230 18.060 1616.550 18.120 ;
        RECT 2253.330 18.060 2253.650 18.120 ;
      LAYER via ;
        RECT 1616.260 18.060 1616.520 18.320 ;
        RECT 2253.360 18.060 2253.620 18.320 ;
      LAYER met2 ;
        RECT 1616.320 18.350 1616.460 54.000 ;
        RECT 1616.260 18.030 1616.520 18.350 ;
        RECT 2253.360 18.030 2253.620 18.350 ;
        RECT 2253.420 2.400 2253.560 18.030 ;
        RECT 2253.350 0.000 2253.630 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1629.645 19.805 1631.655 19.975 ;
        RECT 1629.645 19.465 1629.815 19.805 ;
        RECT 1631.485 17.425 1631.655 19.805 ;
        RECT 1706.925 17.425 1707.095 22.695 ;
        RECT 1728.085 12.665 1728.255 22.695 ;
        RECT 1776.385 13.005 1776.555 14.875 ;
        RECT 1803.525 14.195 1803.695 17.595 ;
        RECT 1851.825 14.195 1851.995 17.595 ;
        RECT 1803.525 14.025 1823.475 14.195 ;
        RECT 1823.305 13.005 1823.475 14.025 ;
        RECT 1824.685 13.005 1824.855 14.195 ;
        RECT 1851.825 14.025 1871.775 14.195 ;
        RECT 1871.605 13.005 1871.775 14.025 ;
        RECT 1920.365 12.665 1920.535 17.935 ;
      LAYER mcon ;
        RECT 1706.925 22.525 1707.095 22.695 ;
        RECT 1728.085 22.525 1728.255 22.695 ;
        RECT 1920.365 17.765 1920.535 17.935 ;
        RECT 1803.525 17.425 1803.695 17.595 ;
        RECT 1776.385 14.705 1776.555 14.875 ;
        RECT 1851.825 17.425 1851.995 17.595 ;
        RECT 1824.685 14.025 1824.855 14.195 ;
      LAYER met1 ;
        RECT 1706.865 22.680 1707.155 22.725 ;
        RECT 1728.025 22.680 1728.315 22.725 ;
        RECT 1706.865 22.540 1728.315 22.680 ;
        RECT 1706.865 22.495 1707.155 22.540 ;
        RECT 1728.025 22.495 1728.315 22.540 ;
        RECT 1621.290 19.620 1621.610 19.680 ;
        RECT 1629.585 19.620 1629.875 19.665 ;
        RECT 1621.290 19.480 1629.875 19.620 ;
        RECT 1621.290 19.420 1621.610 19.480 ;
        RECT 1629.585 19.435 1629.875 19.480 ;
        RECT 1920.305 17.920 1920.595 17.965 ;
        RECT 2270.810 17.920 2271.130 17.980 ;
        RECT 1920.305 17.780 2271.130 17.920 ;
        RECT 1920.305 17.735 1920.595 17.780 ;
        RECT 2270.810 17.720 2271.130 17.780 ;
        RECT 1631.425 17.580 1631.715 17.625 ;
        RECT 1706.865 17.580 1707.155 17.625 ;
        RECT 1631.425 17.440 1707.155 17.580 ;
        RECT 1631.425 17.395 1631.715 17.440 ;
        RECT 1706.865 17.395 1707.155 17.440 ;
        RECT 1802.990 17.580 1803.310 17.640 ;
        RECT 1803.465 17.580 1803.755 17.625 ;
        RECT 1802.990 17.440 1803.755 17.580 ;
        RECT 1802.990 17.380 1803.310 17.440 ;
        RECT 1803.465 17.395 1803.755 17.440 ;
        RECT 1851.290 17.580 1851.610 17.640 ;
        RECT 1851.765 17.580 1852.055 17.625 ;
        RECT 1851.290 17.440 1852.055 17.580 ;
        RECT 1851.290 17.380 1851.610 17.440 ;
        RECT 1851.765 17.395 1852.055 17.440 ;
        RECT 1776.310 14.860 1776.630 14.920 ;
        RECT 1776.115 14.720 1776.630 14.860 ;
        RECT 1776.310 14.660 1776.630 14.720 ;
        RECT 1824.610 14.180 1824.930 14.240 ;
        RECT 1824.610 14.040 1825.125 14.180 ;
        RECT 1824.610 13.980 1824.930 14.040 ;
        RECT 1776.325 13.160 1776.615 13.205 ;
        RECT 1736.840 13.020 1776.615 13.160 ;
        RECT 1728.025 12.820 1728.315 12.865 ;
        RECT 1736.840 12.820 1736.980 13.020 ;
        RECT 1776.325 12.975 1776.615 13.020 ;
        RECT 1823.245 13.160 1823.535 13.205 ;
        RECT 1824.625 13.160 1824.915 13.205 ;
        RECT 1823.245 13.020 1824.915 13.160 ;
        RECT 1823.245 12.975 1823.535 13.020 ;
        RECT 1824.625 12.975 1824.915 13.020 ;
        RECT 1871.545 13.160 1871.835 13.205 ;
        RECT 1871.545 13.020 1872.680 13.160 ;
        RECT 1871.545 12.975 1871.835 13.020 ;
        RECT 1728.025 12.680 1736.980 12.820 ;
        RECT 1872.540 12.820 1872.680 13.020 ;
        RECT 1920.305 12.820 1920.595 12.865 ;
        RECT 1872.540 12.680 1920.595 12.820 ;
        RECT 1728.025 12.635 1728.315 12.680 ;
        RECT 1920.305 12.635 1920.595 12.680 ;
      LAYER via ;
        RECT 1621.320 19.420 1621.580 19.680 ;
        RECT 2270.840 17.720 2271.100 17.980 ;
        RECT 1803.020 17.380 1803.280 17.640 ;
        RECT 1851.320 17.380 1851.580 17.640 ;
        RECT 1776.340 14.660 1776.600 14.920 ;
        RECT 1824.640 13.980 1824.900 14.240 ;
      LAYER met2 ;
        RECT 1621.380 19.710 1621.520 54.000 ;
        RECT 1621.320 19.390 1621.580 19.710 ;
        RECT 2270.840 17.690 2271.100 18.010 ;
        RECT 1803.020 17.350 1803.280 17.670 ;
        RECT 1851.320 17.525 1851.580 17.670 ;
        RECT 1776.340 14.805 1776.600 14.950 ;
        RECT 1803.080 14.805 1803.220 17.350 ;
        RECT 1824.630 17.155 1824.910 17.525 ;
        RECT 1851.310 17.155 1851.590 17.525 ;
        RECT 1776.330 14.435 1776.610 14.805 ;
        RECT 1803.010 14.435 1803.290 14.805 ;
        RECT 1824.700 14.270 1824.840 17.155 ;
        RECT 1824.640 13.950 1824.900 14.270 ;
        RECT 2270.900 2.400 2271.040 17.690 ;
        RECT 2270.830 0.000 2271.110 2.400 ;
      LAYER via2 ;
        RECT 1824.630 17.200 1824.910 17.480 ;
        RECT 1851.310 17.200 1851.590 17.480 ;
        RECT 1776.330 14.480 1776.610 14.760 ;
        RECT 1803.010 14.480 1803.290 14.760 ;
      LAYER met3 ;
        RECT 1824.605 17.490 1824.935 17.505 ;
        RECT 1851.285 17.490 1851.615 17.505 ;
        RECT 1824.605 17.190 1851.615 17.490 ;
        RECT 1824.605 17.175 1824.935 17.190 ;
        RECT 1851.285 17.175 1851.615 17.190 ;
        RECT 1776.305 14.770 1776.635 14.785 ;
        RECT 1802.985 14.770 1803.315 14.785 ;
        RECT 1776.305 14.470 1803.315 14.770 ;
        RECT 1776.305 14.455 1776.635 14.470 ;
        RECT 1802.985 14.455 1803.315 14.470 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1657.705 18.445 1657.875 21.335 ;
        RECT 1753.845 12.665 1754.015 17.595 ;
        RECT 1823.765 12.665 1823.935 14.195 ;
      LAYER mcon ;
        RECT 1657.705 21.165 1657.875 21.335 ;
        RECT 1753.845 17.425 1754.015 17.595 ;
        RECT 1823.765 14.025 1823.935 14.195 ;
      LAYER met1 ;
        RECT 1657.645 21.320 1657.935 21.365 ;
        RECT 1683.390 21.320 1683.710 21.380 ;
        RECT 1657.645 21.180 1683.710 21.320 ;
        RECT 1657.645 21.135 1657.935 21.180 ;
        RECT 1683.390 21.120 1683.710 21.180 ;
        RECT 1623.130 18.600 1623.450 18.660 ;
        RECT 1657.645 18.600 1657.935 18.645 ;
        RECT 1623.130 18.460 1657.935 18.600 ;
        RECT 1623.130 18.400 1623.450 18.460 ;
        RECT 1657.645 18.415 1657.935 18.460 ;
        RECT 1707.310 17.580 1707.630 17.640 ;
        RECT 1753.785 17.580 1754.075 17.625 ;
        RECT 1707.310 17.440 1754.075 17.580 ;
        RECT 1707.310 17.380 1707.630 17.440 ;
        RECT 1753.785 17.395 1754.075 17.440 ;
        RECT 1852.670 17.580 1852.990 17.640 ;
        RECT 2288.750 17.580 2289.070 17.640 ;
        RECT 1852.670 17.440 2289.070 17.580 ;
        RECT 1852.670 17.380 1852.990 17.440 ;
        RECT 2288.750 17.380 2289.070 17.440 ;
        RECT 1823.690 14.180 1824.010 14.240 ;
        RECT 1823.690 14.040 1824.205 14.180 ;
        RECT 1823.690 13.980 1824.010 14.040 ;
        RECT 1753.785 12.820 1754.075 12.865 ;
        RECT 1823.705 12.820 1823.995 12.865 ;
        RECT 1753.785 12.680 1823.995 12.820 ;
        RECT 1753.785 12.635 1754.075 12.680 ;
        RECT 1823.705 12.635 1823.995 12.680 ;
      LAYER via ;
        RECT 1683.420 21.120 1683.680 21.380 ;
        RECT 1623.160 18.400 1623.420 18.660 ;
        RECT 1707.340 17.380 1707.600 17.640 ;
        RECT 1852.700 17.380 1852.960 17.640 ;
        RECT 2288.780 17.380 2289.040 17.640 ;
        RECT 1823.720 13.980 1823.980 14.240 ;
      LAYER met2 ;
        RECT 1623.220 18.690 1623.360 54.000 ;
        RECT 1683.420 21.090 1683.680 21.410 ;
        RECT 1623.160 18.370 1623.420 18.690 ;
        RECT 1683.480 17.525 1683.620 21.090 ;
        RECT 1707.340 17.525 1707.600 17.670 ;
        RECT 1683.410 17.155 1683.690 17.525 ;
        RECT 1707.330 17.155 1707.610 17.525 ;
        RECT 1852.700 17.350 1852.960 17.670 ;
        RECT 2288.780 17.350 2289.040 17.670 ;
        RECT 1852.760 15.485 1852.900 17.350 ;
        RECT 1852.690 15.115 1852.970 15.485 ;
        RECT 1823.710 14.435 1823.990 14.805 ;
        RECT 1823.780 14.270 1823.920 14.435 ;
        RECT 1823.720 13.950 1823.980 14.270 ;
        RECT 2288.840 2.400 2288.980 17.350 ;
        RECT 2288.770 0.000 2289.050 2.400 ;
      LAYER via2 ;
        RECT 1683.410 17.200 1683.690 17.480 ;
        RECT 1707.330 17.200 1707.610 17.480 ;
        RECT 1852.690 15.160 1852.970 15.440 ;
        RECT 1823.710 14.480 1823.990 14.760 ;
      LAYER met3 ;
        RECT 1683.385 17.490 1683.715 17.505 ;
        RECT 1707.305 17.490 1707.635 17.505 ;
        RECT 1683.385 17.190 1707.635 17.490 ;
        RECT 1683.385 17.175 1683.715 17.190 ;
        RECT 1707.305 17.175 1707.635 17.190 ;
        RECT 1852.665 15.450 1852.995 15.465 ;
        RECT 1828.070 15.150 1852.995 15.450 ;
        RECT 1823.685 14.770 1824.015 14.785 ;
        RECT 1828.070 14.770 1828.370 15.150 ;
        RECT 1852.665 15.135 1852.995 15.150 ;
        RECT 1823.685 14.470 1828.370 14.770 ;
        RECT 1823.685 14.455 1824.015 14.470 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1631.025 13.005 1631.195 17.595 ;
        RECT 1919.905 13.005 1920.075 17.935 ;
        RECT 1950.265 13.005 1950.435 17.255 ;
      LAYER mcon ;
        RECT 1919.905 17.765 1920.075 17.935 ;
        RECT 1631.025 17.425 1631.195 17.595 ;
        RECT 1950.265 17.085 1950.435 17.255 ;
      LAYER met1 ;
        RECT 1853.130 17.920 1853.450 17.980 ;
        RECT 1919.845 17.920 1920.135 17.965 ;
        RECT 1853.130 17.780 1920.135 17.920 ;
        RECT 1853.130 17.720 1853.450 17.780 ;
        RECT 1919.845 17.735 1920.135 17.780 ;
        RECT 1630.490 17.580 1630.810 17.640 ;
        RECT 1630.965 17.580 1631.255 17.625 ;
        RECT 1630.490 17.440 1631.255 17.580 ;
        RECT 1630.490 17.380 1630.810 17.440 ;
        RECT 1630.965 17.395 1631.255 17.440 ;
        RECT 1755.610 17.580 1755.930 17.640 ;
        RECT 1802.530 17.580 1802.850 17.640 ;
        RECT 1755.610 17.440 1802.850 17.580 ;
        RECT 1755.610 17.380 1755.930 17.440 ;
        RECT 1802.530 17.380 1802.850 17.440 ;
        RECT 1803.910 17.580 1804.230 17.640 ;
        RECT 1850.830 17.580 1851.150 17.640 ;
        RECT 1803.910 17.440 1851.150 17.580 ;
        RECT 1803.910 17.380 1804.230 17.440 ;
        RECT 1850.830 17.380 1851.150 17.440 ;
        RECT 1950.205 17.240 1950.495 17.285 ;
        RECT 2306.690 17.240 2307.010 17.300 ;
        RECT 1950.205 17.100 2307.010 17.240 ;
        RECT 1950.205 17.055 1950.495 17.100 ;
        RECT 2306.690 17.040 2307.010 17.100 ;
        RECT 1630.965 13.160 1631.255 13.205 ;
        RECT 1731.690 13.160 1732.010 13.220 ;
        RECT 1630.965 13.020 1732.010 13.160 ;
        RECT 1630.965 12.975 1631.255 13.020 ;
        RECT 1731.690 12.960 1732.010 13.020 ;
        RECT 1919.845 13.160 1920.135 13.205 ;
        RECT 1950.205 13.160 1950.495 13.205 ;
        RECT 1919.845 13.020 1950.495 13.160 ;
        RECT 1919.845 12.975 1920.135 13.020 ;
        RECT 1950.205 12.975 1950.495 13.020 ;
      LAYER via ;
        RECT 1853.160 17.720 1853.420 17.980 ;
        RECT 1630.520 17.380 1630.780 17.640 ;
        RECT 1755.640 17.380 1755.900 17.640 ;
        RECT 1802.560 17.380 1802.820 17.640 ;
        RECT 1803.940 17.380 1804.200 17.640 ;
        RECT 1850.860 17.380 1851.120 17.640 ;
        RECT 2306.720 17.040 2306.980 17.300 ;
        RECT 1731.720 12.960 1731.980 13.220 ;
      LAYER met2 ;
        RECT 1630.580 17.670 1630.720 54.000 ;
        RECT 1853.160 17.690 1853.420 18.010 ;
        RECT 1630.520 17.350 1630.780 17.670 ;
        RECT 1755.640 17.350 1755.900 17.670 ;
        RECT 1802.560 17.350 1802.820 17.670 ;
        RECT 1803.940 17.350 1804.200 17.670 ;
        RECT 1850.860 17.350 1851.120 17.670 ;
        RECT 1755.700 16.165 1755.840 17.350 ;
        RECT 1802.620 16.165 1802.760 17.350 ;
        RECT 1804.000 16.165 1804.140 17.350 ;
        RECT 1850.920 16.165 1851.060 17.350 ;
        RECT 1853.220 16.165 1853.360 17.690 ;
        RECT 2306.720 17.010 2306.980 17.330 ;
        RECT 1731.710 15.795 1731.990 16.165 ;
        RECT 1755.630 15.795 1755.910 16.165 ;
        RECT 1802.550 15.795 1802.830 16.165 ;
        RECT 1803.930 15.795 1804.210 16.165 ;
        RECT 1850.850 15.795 1851.130 16.165 ;
        RECT 1853.150 15.795 1853.430 16.165 ;
        RECT 1731.780 13.250 1731.920 15.795 ;
        RECT 1731.720 12.930 1731.980 13.250 ;
        RECT 2306.780 2.400 2306.920 17.010 ;
        RECT 2306.710 0.000 2306.990 2.400 ;
      LAYER via2 ;
        RECT 1731.710 15.840 1731.990 16.120 ;
        RECT 1755.630 15.840 1755.910 16.120 ;
        RECT 1802.550 15.840 1802.830 16.120 ;
        RECT 1803.930 15.840 1804.210 16.120 ;
        RECT 1850.850 15.840 1851.130 16.120 ;
        RECT 1853.150 15.840 1853.430 16.120 ;
      LAYER met3 ;
        RECT 1731.685 16.130 1732.015 16.145 ;
        RECT 1755.605 16.130 1755.935 16.145 ;
        RECT 1731.685 15.830 1755.935 16.130 ;
        RECT 1731.685 15.815 1732.015 15.830 ;
        RECT 1755.605 15.815 1755.935 15.830 ;
        RECT 1802.525 16.130 1802.855 16.145 ;
        RECT 1803.905 16.130 1804.235 16.145 ;
        RECT 1802.525 15.830 1804.235 16.130 ;
        RECT 1802.525 15.815 1802.855 15.830 ;
        RECT 1803.905 15.815 1804.235 15.830 ;
        RECT 1850.825 16.130 1851.155 16.145 ;
        RECT 1853.125 16.130 1853.455 16.145 ;
        RECT 1850.825 15.830 1853.455 16.130 ;
        RECT 1850.825 15.815 1851.155 15.830 ;
        RECT 1853.125 15.815 1853.455 15.830 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1630.120 20.245 1630.260 54.000 ;
        RECT 1630.050 19.875 1630.330 20.245 ;
        RECT 2324.650 19.875 2324.930 20.245 ;
        RECT 2324.720 2.400 2324.860 19.875 ;
        RECT 2324.650 0.000 2324.930 2.400 ;
      LAYER via2 ;
        RECT 1630.050 19.920 1630.330 20.200 ;
        RECT 2324.650 19.920 2324.930 20.200 ;
      LAYER met3 ;
        RECT 1630.025 20.210 1630.355 20.225 ;
        RECT 2324.625 20.210 2324.955 20.225 ;
        RECT 1630.025 19.910 2324.955 20.210 ;
        RECT 1630.025 19.895 1630.355 19.910 ;
        RECT 2324.625 19.895 2324.955 19.910 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1637.020 19.565 1637.160 54.000 ;
        RECT 1636.950 19.195 1637.230 19.565 ;
        RECT 2342.130 19.195 2342.410 19.565 ;
        RECT 2342.200 2.400 2342.340 19.195 ;
        RECT 2342.130 0.000 2342.410 2.400 ;
      LAYER via2 ;
        RECT 1636.950 19.240 1637.230 19.520 ;
        RECT 2342.130 19.240 2342.410 19.520 ;
      LAYER met3 ;
        RECT 1636.925 19.530 1637.255 19.545 ;
        RECT 2342.105 19.530 2342.435 19.545 ;
        RECT 1636.925 19.230 2342.435 19.530 ;
        RECT 1636.925 19.215 1637.255 19.230 ;
        RECT 2342.105 19.215 2342.435 19.230 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1637.480 18.885 1637.620 54.000 ;
        RECT 1637.410 18.515 1637.690 18.885 ;
        RECT 2360.070 18.515 2360.350 18.885 ;
        RECT 2360.140 2.400 2360.280 18.515 ;
        RECT 2360.070 0.000 2360.350 2.400 ;
      LAYER via2 ;
        RECT 1637.410 18.560 1637.690 18.840 ;
        RECT 2360.070 18.560 2360.350 18.840 ;
      LAYER met3 ;
        RECT 1637.385 18.850 1637.715 18.865 ;
        RECT 2360.045 18.850 2360.375 18.865 ;
        RECT 1637.385 18.550 2360.375 18.850 ;
        RECT 1637.385 18.535 1637.715 18.550 ;
        RECT 2360.045 18.535 2360.375 18.550 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1643.920 18.205 1644.060 54.000 ;
        RECT 1643.850 17.835 1644.130 18.205 ;
        RECT 2378.010 17.835 2378.290 18.205 ;
        RECT 2378.080 2.400 2378.220 17.835 ;
        RECT 2378.010 0.000 2378.290 2.400 ;
      LAYER via2 ;
        RECT 1643.850 17.880 1644.130 18.160 ;
        RECT 2378.010 17.880 2378.290 18.160 ;
      LAYER met3 ;
        RECT 1643.825 18.170 1644.155 18.185 ;
        RECT 1739.710 18.170 1740.090 18.180 ;
        RECT 1643.825 17.870 1740.090 18.170 ;
        RECT 1643.825 17.855 1644.155 17.870 ;
        RECT 1739.710 17.860 1740.090 17.870 ;
        RECT 1742.470 18.170 1742.850 18.180 ;
        RECT 2377.985 18.170 2378.315 18.185 ;
        RECT 1742.470 17.870 2378.315 18.170 ;
        RECT 1742.470 17.860 1742.850 17.870 ;
        RECT 2377.985 17.855 2378.315 17.870 ;
      LAYER via3 ;
        RECT 1739.740 17.860 1740.060 18.180 ;
        RECT 1742.500 17.860 1742.820 18.180 ;
      LAYER met4 ;
        RECT 1739.750 18.550 1742.810 18.850 ;
        RECT 1739.750 18.185 1740.050 18.550 ;
        RECT 1742.510 18.185 1742.810 18.550 ;
        RECT 1739.735 17.855 1740.065 18.185 ;
        RECT 1742.495 17.855 1742.825 18.185 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1644.380 17.525 1644.520 54.000 ;
        RECT 1644.310 17.155 1644.590 17.525 ;
        RECT 1875.690 17.155 1875.970 17.525 ;
        RECT 2167.790 17.155 2168.070 17.525 ;
        RECT 2168.710 17.155 2168.990 17.525 ;
        RECT 2395.950 17.155 2396.230 17.525 ;
        RECT 1692.610 16.730 1692.890 16.845 ;
        RECT 1691.760 16.590 1692.890 16.730 ;
        RECT 1691.760 16.165 1691.900 16.590 ;
        RECT 1692.610 16.475 1692.890 16.590 ;
        RECT 1826.470 16.475 1826.750 16.845 ;
        RECT 1691.690 15.795 1691.970 16.165 ;
        RECT 1826.540 14.690 1826.680 16.475 ;
        RECT 1875.760 14.805 1875.900 17.155 ;
        RECT 2167.860 16.900 2168.000 17.155 ;
        RECT 2168.780 16.900 2168.920 17.155 ;
        RECT 2167.860 16.760 2168.920 16.900 ;
        RECT 1828.770 14.690 1829.050 14.805 ;
        RECT 1826.540 14.550 1829.050 14.690 ;
        RECT 1828.770 14.435 1829.050 14.550 ;
        RECT 1875.690 14.435 1875.970 14.805 ;
        RECT 2396.020 2.400 2396.160 17.155 ;
        RECT 2395.950 0.000 2396.230 2.400 ;
      LAYER via2 ;
        RECT 1644.310 17.200 1644.590 17.480 ;
        RECT 1875.690 17.200 1875.970 17.480 ;
        RECT 2167.790 17.200 2168.070 17.480 ;
        RECT 2168.710 17.200 2168.990 17.480 ;
        RECT 2395.950 17.200 2396.230 17.480 ;
        RECT 1692.610 16.520 1692.890 16.800 ;
        RECT 1826.470 16.520 1826.750 16.800 ;
        RECT 1691.690 15.840 1691.970 16.120 ;
        RECT 1828.770 14.480 1829.050 14.760 ;
        RECT 1875.690 14.480 1875.970 14.760 ;
      LAYER met3 ;
        RECT 1644.285 17.490 1644.615 17.505 ;
        RECT 1740.900 17.490 1742.120 17.660 ;
        RECT 1875.665 17.490 1875.995 17.505 ;
        RECT 2167.765 17.490 2168.095 17.505 ;
        RECT 1644.285 17.190 1668.290 17.490 ;
        RECT 1644.285 17.175 1644.615 17.190 ;
        RECT 1667.990 16.130 1668.290 17.190 ;
        RECT 1716.750 17.360 1813.650 17.490 ;
        RECT 1716.750 17.190 1741.200 17.360 ;
        RECT 1741.820 17.190 1813.650 17.360 ;
        RECT 1692.585 16.810 1692.915 16.825 ;
        RECT 1716.750 16.810 1717.050 17.190 ;
        RECT 1692.585 16.510 1717.050 16.810 ;
        RECT 1813.350 16.810 1813.650 17.190 ;
        RECT 1875.665 17.190 2168.095 17.490 ;
        RECT 1875.665 17.175 1875.995 17.190 ;
        RECT 2167.765 17.175 2168.095 17.190 ;
        RECT 2168.685 17.490 2169.015 17.505 ;
        RECT 2395.925 17.490 2396.255 17.505 ;
        RECT 2168.685 17.190 2396.255 17.490 ;
        RECT 2168.685 17.175 2169.015 17.190 ;
        RECT 2395.925 17.175 2396.255 17.190 ;
        RECT 1826.445 16.810 1826.775 16.825 ;
        RECT 1813.350 16.510 1826.775 16.810 ;
        RECT 1692.585 16.495 1692.915 16.510 ;
        RECT 1826.445 16.495 1826.775 16.510 ;
        RECT 1691.665 16.130 1691.995 16.145 ;
        RECT 1667.990 15.830 1691.995 16.130 ;
        RECT 1691.665 15.815 1691.995 15.830 ;
        RECT 1828.745 14.770 1829.075 14.785 ;
        RECT 1875.665 14.770 1875.995 14.785 ;
        RECT 1828.745 14.470 1875.995 14.770 ;
        RECT 1828.745 14.455 1829.075 14.470 ;
        RECT 1875.665 14.455 1875.995 14.470 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2169.150 16.900 2169.470 16.960 ;
        RECT 2258.390 16.900 2258.710 16.960 ;
        RECT 2169.150 16.760 2258.710 16.900 ;
        RECT 2169.150 16.700 2169.470 16.760 ;
        RECT 2258.390 16.700 2258.710 16.760 ;
        RECT 2332.910 16.900 2333.230 16.960 ;
        RECT 2403.290 16.900 2403.610 16.960 ;
        RECT 2332.910 16.760 2403.610 16.900 ;
        RECT 2332.910 16.700 2333.230 16.760 ;
        RECT 2403.290 16.700 2403.610 16.760 ;
        RECT 2034.370 14.860 2034.690 14.920 ;
        RECT 2058.290 14.860 2058.610 14.920 ;
        RECT 2034.370 14.720 2058.610 14.860 ;
        RECT 2034.370 14.660 2034.690 14.720 ;
        RECT 2058.290 14.660 2058.610 14.720 ;
        RECT 2073.010 14.860 2073.330 14.920 ;
        RECT 2120.390 14.860 2120.710 14.920 ;
        RECT 2073.010 14.720 2120.710 14.860 ;
        RECT 2073.010 14.660 2073.330 14.720 ;
        RECT 2120.390 14.660 2120.710 14.720 ;
      LAYER via ;
        RECT 2169.180 16.700 2169.440 16.960 ;
        RECT 2258.420 16.700 2258.680 16.960 ;
        RECT 2332.940 16.700 2333.200 16.960 ;
        RECT 2403.320 16.700 2403.580 16.960 ;
        RECT 2034.400 14.660 2034.660 14.920 ;
        RECT 2058.320 14.660 2058.580 14.920 ;
        RECT 2073.040 14.660 2073.300 14.920 ;
        RECT 2120.420 14.660 2120.680 14.920 ;
      LAYER met2 ;
        RECT 1648.980 53.990 1649.580 54.000 ;
        RECT 1648.980 14.805 1649.120 53.990 ;
        RECT 2072.640 17.270 2073.240 17.410 ;
        RECT 2072.640 16.845 2072.780 17.270 ;
        RECT 1731.250 16.475 1731.530 16.845 ;
        RECT 1878.910 16.730 1879.190 16.845 ;
        RECT 1879.830 16.730 1880.110 16.845 ;
        RECT 1878.910 16.590 1880.110 16.730 ;
        RECT 1878.910 16.475 1879.190 16.590 ;
        RECT 1879.830 16.475 1880.110 16.590 ;
        RECT 1962.170 16.475 1962.450 16.845 ;
        RECT 2058.310 16.475 2058.590 16.845 ;
        RECT 2072.570 16.475 2072.850 16.845 ;
        RECT 1731.320 14.805 1731.460 16.475 ;
        RECT 1962.240 14.805 1962.380 16.475 ;
        RECT 2010.010 15.795 2010.290 16.165 ;
        RECT 2034.390 15.795 2034.670 16.165 ;
        RECT 2010.080 14.805 2010.220 15.795 ;
        RECT 2034.460 14.950 2034.600 15.795 ;
        RECT 2058.380 14.950 2058.520 16.475 ;
        RECT 2073.100 14.950 2073.240 17.270 ;
        RECT 2169.180 16.845 2169.440 16.990 ;
        RECT 2169.170 16.475 2169.450 16.845 ;
        RECT 2258.420 16.670 2258.680 16.990 ;
        RECT 2332.940 16.670 2333.200 16.990 ;
        RECT 2403.320 16.670 2403.580 16.990 ;
        RECT 2258.480 16.165 2258.620 16.670 ;
        RECT 2333.000 16.165 2333.140 16.670 ;
        RECT 2403.380 16.165 2403.520 16.670 ;
        RECT 2120.410 15.795 2120.690 16.165 ;
        RECT 2258.410 15.795 2258.690 16.165 ;
        RECT 2313.610 15.795 2313.890 16.165 ;
        RECT 2332.930 15.795 2333.210 16.165 ;
        RECT 2403.310 15.795 2403.590 16.165 ;
        RECT 2413.890 15.795 2414.170 16.165 ;
        RECT 2120.480 14.950 2120.620 15.795 ;
        RECT 2313.680 15.485 2313.820 15.795 ;
        RECT 2313.610 15.115 2313.890 15.485 ;
        RECT 1648.910 14.435 1649.190 14.805 ;
        RECT 1731.250 14.435 1731.530 14.805 ;
        RECT 1962.170 14.435 1962.450 14.805 ;
        RECT 2010.010 14.435 2010.290 14.805 ;
        RECT 2034.400 14.630 2034.660 14.950 ;
        RECT 2058.320 14.630 2058.580 14.950 ;
        RECT 2073.040 14.630 2073.300 14.950 ;
        RECT 2120.420 14.630 2120.680 14.950 ;
        RECT 2413.960 2.400 2414.100 15.795 ;
        RECT 2413.890 0.000 2414.170 2.400 ;
      LAYER via2 ;
        RECT 1731.250 16.520 1731.530 16.800 ;
        RECT 1878.910 16.520 1879.190 16.800 ;
        RECT 1879.830 16.520 1880.110 16.800 ;
        RECT 1962.170 16.520 1962.450 16.800 ;
        RECT 2058.310 16.520 2058.590 16.800 ;
        RECT 2072.570 16.520 2072.850 16.800 ;
        RECT 2010.010 15.840 2010.290 16.120 ;
        RECT 2034.390 15.840 2034.670 16.120 ;
        RECT 2169.170 16.520 2169.450 16.800 ;
        RECT 2120.410 15.840 2120.690 16.120 ;
        RECT 2258.410 15.840 2258.690 16.120 ;
        RECT 2313.610 15.840 2313.890 16.120 ;
        RECT 2332.930 15.840 2333.210 16.120 ;
        RECT 2403.310 15.840 2403.590 16.120 ;
        RECT 2413.890 15.840 2414.170 16.120 ;
        RECT 2313.610 15.160 2313.890 15.440 ;
        RECT 1648.910 14.480 1649.190 14.760 ;
        RECT 1731.250 14.480 1731.530 14.760 ;
        RECT 1962.170 14.480 1962.450 14.760 ;
        RECT 2010.010 14.480 2010.290 14.760 ;
      LAYER met3 ;
        RECT 1731.225 16.810 1731.555 16.825 ;
        RECT 1878.885 16.810 1879.215 16.825 ;
        RECT 1731.225 16.510 1779.610 16.810 ;
        RECT 1731.225 16.495 1731.555 16.510 ;
        RECT 1779.310 15.450 1779.610 16.510 ;
        RECT 1827.150 16.510 1879.215 16.810 ;
        RECT 1827.150 15.450 1827.450 16.510 ;
        RECT 1878.885 16.495 1879.215 16.510 ;
        RECT 1879.805 16.810 1880.135 16.825 ;
        RECT 1962.145 16.810 1962.475 16.825 ;
        RECT 1879.805 16.510 1962.475 16.810 ;
        RECT 1879.805 16.495 1880.135 16.510 ;
        RECT 1962.145 16.495 1962.475 16.510 ;
        RECT 2058.285 16.810 2058.615 16.825 ;
        RECT 2072.545 16.810 2072.875 16.825 ;
        RECT 2169.145 16.810 2169.475 16.825 ;
        RECT 2058.285 16.510 2072.875 16.810 ;
        RECT 2058.285 16.495 2058.615 16.510 ;
        RECT 2072.545 16.495 2072.875 16.510 ;
        RECT 2168.470 16.510 2169.475 16.810 ;
        RECT 2009.985 16.130 2010.315 16.145 ;
        RECT 2034.365 16.130 2034.695 16.145 ;
        RECT 2009.985 15.830 2034.695 16.130 ;
        RECT 2009.985 15.815 2010.315 15.830 ;
        RECT 2034.365 15.815 2034.695 15.830 ;
        RECT 2120.385 16.130 2120.715 16.145 ;
        RECT 2120.385 15.830 2140.250 16.130 ;
        RECT 2120.385 15.815 2120.715 15.830 ;
        RECT 1779.310 15.150 1827.450 15.450 ;
        RECT 2139.950 15.450 2140.250 15.830 ;
        RECT 2168.470 15.450 2168.770 16.510 ;
        RECT 2169.145 16.495 2169.475 16.510 ;
        RECT 2258.385 16.130 2258.715 16.145 ;
        RECT 2313.585 16.130 2313.915 16.145 ;
        RECT 2332.905 16.130 2333.235 16.145 ;
        RECT 2258.385 15.830 2266.290 16.130 ;
        RECT 2258.385 15.815 2258.715 15.830 ;
        RECT 2139.950 15.150 2168.770 15.450 ;
        RECT 2265.990 15.450 2266.290 15.830 ;
        RECT 2313.585 15.830 2333.235 16.130 ;
        RECT 2313.585 15.815 2313.915 15.830 ;
        RECT 2332.905 15.815 2333.235 15.830 ;
        RECT 2403.285 16.130 2403.615 16.145 ;
        RECT 2413.865 16.130 2414.195 16.145 ;
        RECT 2403.285 15.830 2414.195 16.130 ;
        RECT 2403.285 15.815 2403.615 15.830 ;
        RECT 2413.865 15.815 2414.195 15.830 ;
        RECT 2313.585 15.450 2313.915 15.465 ;
        RECT 2265.990 15.150 2313.915 15.450 ;
        RECT 2313.585 15.135 2313.915 15.150 ;
        RECT 1648.885 14.770 1649.215 14.785 ;
        RECT 1731.225 14.770 1731.555 14.785 ;
        RECT 1648.885 14.470 1731.555 14.770 ;
        RECT 1648.885 14.455 1649.215 14.470 ;
        RECT 1731.225 14.455 1731.555 14.470 ;
        RECT 1962.145 14.770 1962.475 14.785 ;
        RECT 2009.985 14.770 2010.315 14.785 ;
        RECT 1962.145 14.470 2010.315 14.770 ;
        RECT 1962.145 14.455 1962.475 14.470 ;
        RECT 2009.985 14.455 2010.315 14.470 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1273.145 44.115 1273.315 49.555 ;
        RECT 1295.685 47.345 1295.855 49.555 ;
        RECT 1272.225 43.945 1273.315 44.115 ;
      LAYER mcon ;
        RECT 1273.145 49.385 1273.315 49.555 ;
        RECT 1295.685 49.385 1295.855 49.555 ;
      LAYER met1 ;
        RECT 1273.085 49.540 1273.375 49.585 ;
        RECT 1295.625 49.540 1295.915 49.585 ;
        RECT 1273.085 49.400 1295.915 49.540 ;
        RECT 1273.085 49.355 1273.375 49.400 ;
        RECT 1295.625 49.355 1295.915 49.400 ;
        RECT 1295.625 47.500 1295.915 47.545 ;
        RECT 1314.470 47.500 1314.790 47.560 ;
        RECT 1295.625 47.360 1314.790 47.500 ;
        RECT 1295.625 47.315 1295.915 47.360 ;
        RECT 1314.470 47.300 1314.790 47.360 ;
        RECT 808.010 44.440 808.330 44.500 ;
        RECT 808.010 44.300 814.220 44.440 ;
        RECT 808.010 44.240 808.330 44.300 ;
        RECT 814.080 44.100 814.220 44.300 ;
        RECT 1272.165 44.100 1272.455 44.145 ;
        RECT 814.080 43.960 1272.455 44.100 ;
        RECT 1272.165 43.915 1272.455 43.960 ;
      LAYER via ;
        RECT 1314.500 47.300 1314.760 47.560 ;
        RECT 808.040 44.240 808.300 44.500 ;
      LAYER met2 ;
        RECT 1314.560 47.590 1314.700 54.000 ;
        RECT 1314.500 47.270 1314.760 47.590 ;
        RECT 808.040 44.210 808.300 44.530 ;
        RECT 808.100 2.400 808.240 44.210 ;
        RECT 808.030 0.000 808.310 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2919.430 0.000 2919.710 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1103.405 23.885 1103.575 25.415 ;
        RECT 1137.905 25.075 1138.075 25.415 ;
        RECT 1137.905 24.905 1138.995 25.075 ;
      LAYER mcon ;
        RECT 1103.405 25.245 1103.575 25.415 ;
        RECT 1137.905 25.245 1138.075 25.415 ;
        RECT 1138.825 24.905 1138.995 25.075 ;
      LAYER met1 ;
        RECT 1103.345 25.400 1103.635 25.445 ;
        RECT 1137.845 25.400 1138.135 25.445 ;
        RECT 1103.345 25.260 1138.135 25.400 ;
        RECT 1103.345 25.215 1103.635 25.260 ;
        RECT 1137.845 25.215 1138.135 25.260 ;
        RECT 1138.765 25.060 1139.055 25.105 ;
        RECT 1148.410 25.060 1148.730 25.120 ;
        RECT 1138.765 24.920 1148.730 25.060 ;
        RECT 1138.765 24.875 1139.055 24.920 ;
        RECT 1148.410 24.860 1148.730 24.920 ;
        RECT 5.310 24.040 5.630 24.100 ;
        RECT 1103.345 24.040 1103.635 24.085 ;
        RECT 5.310 23.900 1103.635 24.040 ;
        RECT 5.310 23.840 5.630 23.900 ;
        RECT 1103.345 23.855 1103.635 23.900 ;
      LAYER via ;
        RECT 1148.440 24.860 1148.700 25.120 ;
        RECT 5.340 23.840 5.600 24.100 ;
      LAYER met2 ;
        RECT 1148.500 25.150 1148.640 54.000 ;
        RECT 1148.440 24.830 1148.700 25.150 ;
        RECT 5.340 23.810 5.600 24.130 ;
        RECT 5.400 2.400 5.540 23.810 ;
        RECT 5.330 0.000 5.610 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1146.645 25.585 1147.735 25.755 ;
        RECT 1146.645 25.245 1146.815 25.585 ;
        RECT 1147.565 25.075 1147.735 25.585 ;
        RECT 1147.565 24.905 1149.115 25.075 ;
      LAYER mcon ;
        RECT 1148.945 24.905 1149.115 25.075 ;
      LAYER met1 ;
        RECT 10.830 25.400 11.150 25.460 ;
        RECT 1146.585 25.400 1146.875 25.445 ;
        RECT 10.830 25.260 1103.100 25.400 ;
        RECT 10.830 25.200 11.150 25.260 ;
        RECT 1102.960 25.060 1103.100 25.260 ;
        RECT 1138.380 25.260 1146.875 25.400 ;
        RECT 1138.380 25.060 1138.520 25.260 ;
        RECT 1146.585 25.215 1146.875 25.260 ;
        RECT 1102.960 24.920 1138.520 25.060 ;
        RECT 1148.885 25.060 1149.175 25.105 ;
        RECT 1150.710 25.060 1151.030 25.120 ;
        RECT 1148.885 24.920 1151.030 25.060 ;
        RECT 1148.885 24.875 1149.175 24.920 ;
        RECT 1150.710 24.860 1151.030 24.920 ;
      LAYER via ;
        RECT 10.860 25.200 11.120 25.460 ;
        RECT 1150.740 24.860 1151.000 25.120 ;
      LAYER met2 ;
        RECT 10.860 25.170 11.120 25.490 ;
        RECT 10.920 2.400 11.060 25.170 ;
        RECT 1150.800 25.150 1150.940 54.000 ;
        RECT 1150.740 24.830 1151.000 25.150 ;
        RECT 10.850 0.000 11.130 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1102.485 23.715 1102.655 25.075 ;
        RECT 1103.865 23.715 1104.035 24.055 ;
        RECT 1102.485 23.545 1104.035 23.715 ;
      LAYER mcon ;
        RECT 1102.485 24.905 1102.655 25.075 ;
        RECT 1103.865 23.885 1104.035 24.055 ;
      LAYER met1 ;
        RECT 16.810 25.060 17.130 25.120 ;
        RECT 1102.425 25.060 1102.715 25.105 ;
        RECT 16.810 24.920 1102.715 25.060 ;
        RECT 16.810 24.860 17.130 24.920 ;
        RECT 1102.425 24.875 1102.715 24.920 ;
        RECT 1103.805 24.040 1104.095 24.085 ;
        RECT 1126.330 24.040 1126.650 24.100 ;
        RECT 1103.805 23.900 1126.650 24.040 ;
        RECT 1103.805 23.855 1104.095 23.900 ;
        RECT 1126.330 23.840 1126.650 23.900 ;
      LAYER via ;
        RECT 16.840 24.860 17.100 25.120 ;
        RECT 1126.360 23.840 1126.620 24.100 ;
      LAYER met2 ;
        RECT 1158.160 27.045 1158.300 54.000 ;
        RECT 1158.090 26.675 1158.370 27.045 ;
        RECT 1126.350 25.995 1126.630 26.365 ;
        RECT 16.840 24.830 17.100 25.150 ;
        RECT 16.900 2.400 17.040 24.830 ;
        RECT 1126.420 24.130 1126.560 25.995 ;
        RECT 1126.360 23.810 1126.620 24.130 ;
        RECT 16.830 0.000 17.110 2.400 ;
      LAYER via2 ;
        RECT 1158.090 26.720 1158.370 27.000 ;
        RECT 1126.350 26.040 1126.630 26.320 ;
      LAYER met3 ;
        RECT 1158.065 27.010 1158.395 27.025 ;
        RECT 1127.950 26.710 1158.395 27.010 ;
        RECT 1126.325 26.330 1126.655 26.345 ;
        RECT 1127.950 26.330 1128.250 26.710 ;
        RECT 1158.065 26.695 1158.395 26.710 ;
        RECT 1126.325 26.030 1128.250 26.330 ;
        RECT 1126.325 26.015 1126.655 26.030 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 40.730 25.740 41.050 25.800 ;
        RECT 1134.610 25.740 1134.930 25.800 ;
        RECT 40.730 25.600 1134.930 25.740 ;
        RECT 40.730 25.540 41.050 25.600 ;
        RECT 1134.610 25.540 1134.930 25.600 ;
      LAYER via ;
        RECT 40.760 25.540 41.020 25.800 ;
        RECT 1134.640 25.540 1134.900 25.800 ;
      LAYER met2 ;
        RECT 1155.400 26.365 1155.540 54.000 ;
        RECT 1134.630 25.995 1134.910 26.365 ;
        RECT 1155.330 25.995 1155.610 26.365 ;
        RECT 1134.700 25.830 1134.840 25.995 ;
        RECT 40.760 25.510 41.020 25.830 ;
        RECT 1134.640 25.510 1134.900 25.830 ;
        RECT 40.820 2.400 40.960 25.510 ;
        RECT 40.750 0.000 41.030 2.400 ;
      LAYER via2 ;
        RECT 1134.630 26.040 1134.910 26.320 ;
        RECT 1155.330 26.040 1155.610 26.320 ;
      LAYER met3 ;
        RECT 1134.605 26.330 1134.935 26.345 ;
        RECT 1155.305 26.330 1155.635 26.345 ;
        RECT 1134.605 26.030 1155.635 26.330 ;
        RECT 1134.605 26.015 1134.935 26.030 ;
        RECT 1155.305 26.015 1155.635 26.030 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.260 31.125 1197.400 54.000 ;
        RECT 243.150 30.755 243.430 31.125 ;
        RECT 1197.190 30.755 1197.470 31.125 ;
        RECT 243.220 2.400 243.360 30.755 ;
        RECT 243.150 0.000 243.430 2.400 ;
      LAYER via2 ;
        RECT 243.150 30.800 243.430 31.080 ;
        RECT 1197.190 30.800 1197.470 31.080 ;
      LAYER met3 ;
        RECT 243.125 31.090 243.455 31.105 ;
        RECT 1197.165 31.090 1197.495 31.105 ;
        RECT 243.125 30.790 1197.495 31.090 ;
        RECT 243.125 30.775 243.455 30.790 ;
        RECT 1197.165 30.775 1197.495 30.790 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1079.485 30.855 1079.655 31.535 ;
        RECT 1079.025 30.685 1079.655 30.855 ;
      LAYER mcon ;
        RECT 1079.485 31.365 1079.655 31.535 ;
      LAYER met1 ;
        RECT 1079.425 31.520 1079.715 31.565 ;
        RECT 1175.550 31.520 1175.870 31.580 ;
        RECT 1079.425 31.380 1175.870 31.520 ;
        RECT 1079.425 31.335 1079.715 31.380 ;
        RECT 1175.550 31.320 1175.870 31.380 ;
        RECT 260.610 30.840 260.930 30.900 ;
        RECT 1078.965 30.840 1079.255 30.885 ;
        RECT 260.610 30.700 1079.255 30.840 ;
        RECT 260.610 30.640 260.930 30.700 ;
        RECT 1078.965 30.655 1079.255 30.700 ;
      LAYER via ;
        RECT 1175.580 31.320 1175.840 31.580 ;
        RECT 260.640 30.640 260.900 30.900 ;
      LAYER met2 ;
        RECT 1205.080 33.165 1205.220 54.000 ;
        RECT 1175.570 32.795 1175.850 33.165 ;
        RECT 1205.010 32.795 1205.290 33.165 ;
        RECT 1175.640 31.610 1175.780 32.795 ;
        RECT 1175.580 31.290 1175.840 31.610 ;
        RECT 260.640 30.610 260.900 30.930 ;
        RECT 260.700 2.400 260.840 30.610 ;
        RECT 260.630 0.000 260.910 2.400 ;
      LAYER via2 ;
        RECT 1175.570 32.840 1175.850 33.120 ;
        RECT 1205.010 32.840 1205.290 33.120 ;
      LAYER met3 ;
        RECT 1175.545 33.130 1175.875 33.145 ;
        RECT 1204.985 33.130 1205.315 33.145 ;
        RECT 1175.545 32.830 1205.315 33.130 ;
        RECT 1175.545 32.815 1175.875 32.830 ;
        RECT 1204.985 32.815 1205.315 32.830 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 278.550 31.180 278.870 31.240 ;
        RECT 1125.870 31.180 1126.190 31.240 ;
        RECT 278.550 31.040 1126.190 31.180 ;
        RECT 278.550 30.980 278.870 31.040 ;
        RECT 1125.870 30.980 1126.190 31.040 ;
      LAYER via ;
        RECT 278.580 30.980 278.840 31.240 ;
        RECT 1125.900 30.980 1126.160 31.240 ;
      LAYER met2 ;
        RECT 1204.160 31.805 1204.300 54.000 ;
        RECT 1125.890 31.435 1126.170 31.805 ;
        RECT 1204.090 31.435 1204.370 31.805 ;
        RECT 1125.960 31.270 1126.100 31.435 ;
        RECT 278.580 30.950 278.840 31.270 ;
        RECT 1125.900 30.950 1126.160 31.270 ;
        RECT 278.640 2.400 278.780 30.950 ;
        RECT 278.570 0.000 278.850 2.400 ;
      LAYER via2 ;
        RECT 1125.890 31.480 1126.170 31.760 ;
        RECT 1204.090 31.480 1204.370 31.760 ;
      LAYER met3 ;
        RECT 1125.865 31.770 1126.195 31.785 ;
        RECT 1204.065 31.770 1204.395 31.785 ;
        RECT 1125.865 31.470 1204.395 31.770 ;
        RECT 1125.865 31.455 1126.195 31.470 ;
        RECT 1204.065 31.455 1204.395 31.470 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 296.490 31.520 296.810 31.580 ;
        RECT 1078.950 31.520 1079.270 31.580 ;
        RECT 296.490 31.380 1079.270 31.520 ;
        RECT 296.490 31.320 296.810 31.380 ;
        RECT 1078.950 31.320 1079.270 31.380 ;
      LAYER via ;
        RECT 296.520 31.320 296.780 31.580 ;
        RECT 1078.980 31.320 1079.240 31.580 ;
      LAYER met2 ;
        RECT 1211.060 32.485 1211.200 54.000 ;
        RECT 1127.270 32.115 1127.550 32.485 ;
        RECT 1210.990 32.115 1211.270 32.485 ;
        RECT 296.520 31.290 296.780 31.610 ;
        RECT 1078.980 31.290 1079.240 31.610 ;
        RECT 296.580 2.400 296.720 31.290 ;
        RECT 1079.040 30.445 1079.180 31.290 ;
        RECT 1078.970 30.075 1079.250 30.445 ;
        RECT 1127.340 29.765 1127.480 32.115 ;
        RECT 1127.270 29.395 1127.550 29.765 ;
        RECT 296.510 0.000 296.790 2.400 ;
      LAYER via2 ;
        RECT 1127.270 32.160 1127.550 32.440 ;
        RECT 1210.990 32.160 1211.270 32.440 ;
        RECT 1078.970 30.120 1079.250 30.400 ;
        RECT 1127.270 29.440 1127.550 29.720 ;
      LAYER met3 ;
        RECT 1127.245 32.450 1127.575 32.465 ;
        RECT 1210.965 32.450 1211.295 32.465 ;
        RECT 1127.245 32.150 1211.295 32.450 ;
        RECT 1127.245 32.135 1127.575 32.150 ;
        RECT 1210.965 32.135 1211.295 32.150 ;
        RECT 1078.945 30.410 1079.275 30.425 ;
        RECT 1078.945 30.110 1085.010 30.410 ;
        RECT 1078.945 30.095 1079.275 30.110 ;
        RECT 1084.710 29.730 1085.010 30.110 ;
        RECT 1127.245 29.730 1127.575 29.745 ;
        RECT 1084.710 29.430 1127.575 29.730 ;
        RECT 1127.245 29.415 1127.575 29.430 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 314.430 39.680 314.750 39.740 ;
        RECT 1211.890 39.680 1212.210 39.740 ;
        RECT 314.430 39.540 1212.210 39.680 ;
        RECT 314.430 39.480 314.750 39.540 ;
        RECT 1211.890 39.480 1212.210 39.540 ;
      LAYER via ;
        RECT 314.460 39.480 314.720 39.740 ;
        RECT 1211.920 39.480 1212.180 39.740 ;
      LAYER met2 ;
        RECT 1212.440 40.530 1212.580 54.000 ;
        RECT 1211.980 40.390 1212.580 40.530 ;
        RECT 1211.980 39.770 1212.120 40.390 ;
        RECT 314.460 39.450 314.720 39.770 ;
        RECT 1211.920 39.450 1212.180 39.770 ;
        RECT 314.520 2.400 314.660 39.450 ;
        RECT 314.450 0.000 314.730 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 332.370 40.020 332.690 40.080 ;
        RECT 1217.870 40.020 1218.190 40.080 ;
        RECT 332.370 39.880 1218.190 40.020 ;
        RECT 332.370 39.820 332.690 39.880 ;
        RECT 1217.870 39.820 1218.190 39.880 ;
      LAYER via ;
        RECT 332.400 39.820 332.660 40.080 ;
        RECT 1217.900 39.820 1218.160 40.080 ;
      LAYER met2 ;
        RECT 1217.960 40.110 1218.100 54.000 ;
        RECT 332.400 39.790 332.660 40.110 ;
        RECT 1217.900 39.790 1218.160 40.110 ;
        RECT 332.460 2.400 332.600 39.790 ;
        RECT 332.390 0.000 332.670 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 349.850 40.360 350.170 40.420 ;
        RECT 1220.170 40.360 1220.490 40.420 ;
        RECT 349.850 40.220 1220.490 40.360 ;
        RECT 349.850 40.160 350.170 40.220 ;
        RECT 1220.170 40.160 1220.490 40.220 ;
      LAYER via ;
        RECT 349.880 40.160 350.140 40.420 ;
        RECT 1220.200 40.160 1220.460 40.420 ;
      LAYER met2 ;
        RECT 1220.260 40.450 1220.400 54.000 ;
        RECT 349.880 40.130 350.140 40.450 ;
        RECT 1220.200 40.130 1220.460 40.450 ;
        RECT 349.940 2.400 350.080 40.130 ;
        RECT 349.870 0.000 350.150 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 367.880 2.400 368.020 54.000 ;
        RECT 367.810 0.000 368.090 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 385.730 15.540 386.050 15.600 ;
        RECT 388.490 15.540 388.810 15.600 ;
        RECT 385.730 15.400 388.810 15.540 ;
        RECT 385.730 15.340 386.050 15.400 ;
        RECT 388.490 15.340 388.810 15.400 ;
      LAYER via ;
        RECT 385.760 15.340 386.020 15.600 ;
        RECT 388.520 15.340 388.780 15.600 ;
      LAYER met2 ;
        RECT 388.580 15.630 388.720 54.000 ;
        RECT 385.760 15.310 386.020 15.630 ;
        RECT 388.520 15.310 388.780 15.630 ;
        RECT 385.820 2.400 385.960 15.310 ;
        RECT 385.750 0.000 386.030 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 403.670 15.540 403.990 15.600 ;
        RECT 409.190 15.540 409.510 15.600 ;
        RECT 403.670 15.400 409.510 15.540 ;
        RECT 403.670 15.340 403.990 15.400 ;
        RECT 409.190 15.340 409.510 15.400 ;
      LAYER via ;
        RECT 403.700 15.340 403.960 15.600 ;
        RECT 409.220 15.340 409.480 15.600 ;
      LAYER met2 ;
        RECT 409.280 15.630 409.420 54.000 ;
        RECT 403.700 15.310 403.960 15.630 ;
        RECT 409.220 15.310 409.480 15.630 ;
        RECT 403.760 2.400 403.900 15.310 ;
        RECT 403.690 0.000 403.970 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 933.205 38.845 933.375 42.075 ;
        RECT 981.965 39.185 982.135 42.075 ;
      LAYER mcon ;
        RECT 933.205 41.905 933.375 42.075 ;
        RECT 981.965 41.905 982.135 42.075 ;
      LAYER met1 ;
        RECT 933.145 42.060 933.435 42.105 ;
        RECT 981.905 42.060 982.195 42.105 ;
        RECT 933.145 41.920 982.195 42.060 ;
        RECT 933.145 41.875 933.435 41.920 ;
        RECT 981.905 41.875 982.195 41.920 ;
        RECT 981.905 39.340 982.195 39.385 ;
        RECT 1078.950 39.340 1079.270 39.400 ;
        RECT 981.905 39.200 1079.270 39.340 ;
        RECT 981.905 39.155 982.195 39.200 ;
        RECT 1078.950 39.140 1079.270 39.200 ;
        RECT 1156.690 39.340 1157.010 39.400 ;
        RECT 1162.670 39.340 1162.990 39.400 ;
        RECT 1156.690 39.200 1162.990 39.340 ;
        RECT 1156.690 39.140 1157.010 39.200 ;
        RECT 1162.670 39.140 1162.990 39.200 ;
        RECT 64.650 39.000 64.970 39.060 ;
        RECT 933.145 39.000 933.435 39.045 ;
        RECT 64.650 38.860 933.435 39.000 ;
        RECT 64.650 38.800 64.970 38.860 ;
        RECT 933.145 38.815 933.435 38.860 ;
      LAYER via ;
        RECT 1078.980 39.140 1079.240 39.400 ;
        RECT 1156.720 39.140 1156.980 39.400 ;
        RECT 1162.700 39.140 1162.960 39.400 ;
        RECT 64.680 38.800 64.940 39.060 ;
      LAYER met2 ;
        RECT 1078.970 39.595 1079.250 39.965 ;
        RECT 1079.040 39.430 1079.180 39.595 ;
        RECT 1162.760 39.430 1162.900 54.000 ;
        RECT 1078.980 39.110 1079.240 39.430 ;
        RECT 1156.720 39.285 1156.980 39.430 ;
        RECT 64.680 38.770 64.940 39.090 ;
        RECT 1156.710 38.915 1156.990 39.285 ;
        RECT 1162.700 39.110 1162.960 39.430 ;
        RECT 64.740 2.400 64.880 38.770 ;
        RECT 64.670 0.000 64.950 2.400 ;
      LAYER via2 ;
        RECT 1078.970 39.640 1079.250 39.920 ;
        RECT 1156.710 38.960 1156.990 39.240 ;
      LAYER met3 ;
        RECT 1078.945 39.930 1079.275 39.945 ;
        RECT 1078.945 39.630 1082.250 39.930 ;
        RECT 1078.945 39.615 1079.275 39.630 ;
        RECT 1081.950 39.250 1082.250 39.630 ;
        RECT 1156.685 39.250 1157.015 39.265 ;
        RECT 1081.950 38.950 1157.015 39.250 ;
        RECT 1156.685 38.935 1157.015 38.950 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 423.080 16.730 423.220 54.000 ;
        RECT 421.700 16.590 423.220 16.730 ;
        RECT 421.700 2.400 421.840 16.590 ;
        RECT 421.630 0.000 421.910 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 439.090 15.200 439.410 15.260 ;
        RECT 443.690 15.200 444.010 15.260 ;
        RECT 439.090 15.060 444.010 15.200 ;
        RECT 439.090 15.000 439.410 15.060 ;
        RECT 443.690 15.000 444.010 15.060 ;
      LAYER via ;
        RECT 439.120 15.000 439.380 15.260 ;
        RECT 443.720 15.000 443.980 15.260 ;
      LAYER met2 ;
        RECT 443.780 15.290 443.920 54.000 ;
        RECT 439.120 14.970 439.380 15.290 ;
        RECT 443.720 14.970 443.980 15.290 ;
        RECT 439.180 2.400 439.320 14.970 ;
        RECT 439.110 0.000 439.390 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 457.565 48.365 457.735 54.000 ;
      LAYER met1 ;
        RECT 457.490 48.520 457.810 48.580 ;
        RECT 457.295 48.380 457.810 48.520 ;
        RECT 457.490 48.320 457.810 48.380 ;
      LAYER via ;
        RECT 457.520 48.320 457.780 48.580 ;
      LAYER met2 ;
        RECT 457.520 48.290 457.780 48.610 ;
        RECT 457.580 24.210 457.720 48.290 ;
        RECT 457.120 24.070 457.720 24.210 ;
        RECT 457.120 2.400 457.260 24.070 ;
        RECT 457.050 0.000 457.330 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 474.970 17.580 475.290 17.640 ;
        RECT 478.190 17.580 478.510 17.640 ;
        RECT 474.970 17.440 478.510 17.580 ;
        RECT 474.970 17.380 475.290 17.440 ;
        RECT 478.190 17.380 478.510 17.440 ;
      LAYER via ;
        RECT 475.000 17.380 475.260 17.640 ;
        RECT 478.220 17.380 478.480 17.640 ;
      LAYER met2 ;
        RECT 478.280 17.670 478.420 54.000 ;
        RECT 475.000 17.350 475.260 17.670 ;
        RECT 478.220 17.350 478.480 17.670 ;
        RECT 475.060 2.400 475.200 17.350 ;
        RECT 474.990 0.000 475.270 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 492.910 17.580 493.230 17.640 ;
        RECT 498.890 17.580 499.210 17.640 ;
        RECT 492.910 17.440 499.210 17.580 ;
        RECT 492.910 17.380 493.230 17.440 ;
        RECT 498.890 17.380 499.210 17.440 ;
      LAYER via ;
        RECT 492.940 17.380 493.200 17.640 ;
        RECT 498.920 17.380 499.180 17.640 ;
      LAYER met2 ;
        RECT 498.980 17.670 499.120 54.000 ;
        RECT 492.940 17.350 493.200 17.670 ;
        RECT 498.920 17.350 499.180 17.670 ;
        RECT 493.000 2.400 493.140 17.350 ;
        RECT 492.930 0.000 493.210 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 512.690 50.220 513.010 50.280 ;
        RECT 1251.910 50.220 1252.230 50.280 ;
        RECT 512.690 50.080 1252.230 50.220 ;
        RECT 512.690 50.020 513.010 50.080 ;
        RECT 1251.910 50.020 1252.230 50.080 ;
        RECT 510.390 15.200 510.710 15.260 ;
        RECT 512.690 15.200 513.010 15.260 ;
        RECT 510.390 15.060 513.010 15.200 ;
        RECT 510.390 15.000 510.710 15.060 ;
        RECT 512.690 15.000 513.010 15.060 ;
      LAYER via ;
        RECT 512.720 50.020 512.980 50.280 ;
        RECT 1251.940 50.020 1252.200 50.280 ;
        RECT 510.420 15.000 510.680 15.260 ;
        RECT 512.720 15.000 512.980 15.260 ;
      LAYER met2 ;
        RECT 1252.000 50.310 1252.140 54.000 ;
        RECT 512.720 49.990 512.980 50.310 ;
        RECT 1251.940 49.990 1252.200 50.310 ;
        RECT 512.780 15.290 512.920 49.990 ;
        RECT 510.420 14.970 510.680 15.290 ;
        RECT 512.720 14.970 512.980 15.290 ;
        RECT 510.480 2.400 510.620 14.970 ;
        RECT 510.410 0.000 510.690 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 533.390 49.880 533.710 49.940 ;
        RECT 1261.570 49.880 1261.890 49.940 ;
        RECT 533.390 49.740 1261.890 49.880 ;
        RECT 533.390 49.680 533.710 49.740 ;
        RECT 1261.570 49.680 1261.890 49.740 ;
        RECT 528.330 14.860 528.650 14.920 ;
        RECT 533.390 14.860 533.710 14.920 ;
        RECT 528.330 14.720 533.710 14.860 ;
        RECT 528.330 14.660 528.650 14.720 ;
        RECT 533.390 14.660 533.710 14.720 ;
      LAYER via ;
        RECT 533.420 49.680 533.680 49.940 ;
        RECT 1261.600 49.680 1261.860 49.940 ;
        RECT 528.360 14.660 528.620 14.920 ;
        RECT 533.420 14.660 533.680 14.920 ;
      LAYER met2 ;
        RECT 1261.660 49.970 1261.800 54.000 ;
        RECT 533.420 49.650 533.680 49.970 ;
        RECT 1261.600 49.650 1261.860 49.970 ;
        RECT 533.480 14.950 533.620 49.650 ;
        RECT 528.360 14.630 528.620 14.950 ;
        RECT 533.420 14.630 533.680 14.950 ;
        RECT 528.420 2.400 528.560 14.630 ;
        RECT 528.350 0.000 528.630 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 547.190 49.540 547.510 49.600 ;
        RECT 1259.270 49.540 1259.590 49.600 ;
        RECT 547.190 49.400 1259.590 49.540 ;
        RECT 547.190 49.340 547.510 49.400 ;
        RECT 1259.270 49.340 1259.590 49.400 ;
      LAYER via ;
        RECT 547.220 49.340 547.480 49.600 ;
        RECT 1259.300 49.340 1259.560 49.600 ;
      LAYER met2 ;
        RECT 1259.360 49.630 1259.500 54.000 ;
        RECT 547.220 49.310 547.480 49.630 ;
        RECT 1259.300 49.310 1259.560 49.630 ;
        RECT 547.280 17.410 547.420 49.310 ;
        RECT 546.360 17.270 547.420 17.410 ;
        RECT 546.360 2.400 546.500 17.270 ;
        RECT 546.290 0.000 546.570 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1224.385 48.365 1224.555 50.915 ;
      LAYER mcon ;
        RECT 1224.385 50.745 1224.555 50.915 ;
      LAYER met1 ;
        RECT 1224.325 50.900 1224.615 50.945 ;
        RECT 1267.550 50.900 1267.870 50.960 ;
        RECT 1224.325 50.760 1267.870 50.900 ;
        RECT 1224.325 50.715 1224.615 50.760 ;
        RECT 1267.550 50.700 1267.870 50.760 ;
        RECT 567.890 48.520 568.210 48.580 ;
        RECT 1224.325 48.520 1224.615 48.565 ;
        RECT 567.890 48.380 1224.615 48.520 ;
        RECT 567.890 48.320 568.210 48.380 ;
        RECT 1224.325 48.335 1224.615 48.380 ;
        RECT 564.210 14.180 564.530 14.240 ;
        RECT 566.510 14.180 566.830 14.240 ;
        RECT 564.210 14.040 566.830 14.180 ;
        RECT 564.210 13.980 564.530 14.040 ;
        RECT 566.510 13.980 566.830 14.040 ;
      LAYER via ;
        RECT 1267.580 50.700 1267.840 50.960 ;
        RECT 567.920 48.320 568.180 48.580 ;
        RECT 564.240 13.980 564.500 14.240 ;
        RECT 566.540 13.980 566.800 14.240 ;
      LAYER met2 ;
        RECT 1267.640 50.990 1267.780 54.000 ;
        RECT 1267.580 50.670 1267.840 50.990 ;
        RECT 567.920 48.290 568.180 48.610 ;
        RECT 564.240 13.950 564.500 14.270 ;
        RECT 566.540 14.010 566.800 14.270 ;
        RECT 567.980 14.010 568.120 48.290 ;
        RECT 566.540 13.950 568.120 14.010 ;
        RECT 564.300 2.400 564.440 13.950 ;
        RECT 566.600 13.870 568.120 13.950 ;
        RECT 564.230 0.000 564.510 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 669.165 52.105 669.335 54.000 ;
      LAYER met1 ;
        RECT 669.105 52.260 669.395 52.305 ;
        RECT 1265.710 52.260 1266.030 52.320 ;
        RECT 669.105 52.120 1266.030 52.260 ;
        RECT 669.105 52.075 669.395 52.120 ;
        RECT 1265.710 52.060 1266.030 52.120 ;
        RECT 582.150 17.580 582.470 17.640 ;
        RECT 587.210 17.580 587.530 17.640 ;
        RECT 582.150 17.440 587.530 17.580 ;
        RECT 582.150 17.380 582.470 17.440 ;
        RECT 587.210 17.380 587.530 17.440 ;
      LAYER via ;
        RECT 1265.740 52.060 1266.000 52.320 ;
        RECT 582.180 17.380 582.440 17.640 ;
        RECT 587.240 17.380 587.500 17.640 ;
      LAYER met2 ;
        RECT 588.220 18.090 588.360 54.000 ;
        RECT 1265.800 52.350 1265.940 54.000 ;
        RECT 1265.740 52.030 1266.000 52.350 ;
        RECT 587.300 17.950 588.360 18.090 ;
        RECT 587.300 17.670 587.440 17.950 ;
        RECT 582.180 17.350 582.440 17.670 ;
        RECT 587.240 17.350 587.500 17.670 ;
        RECT 582.240 2.400 582.380 17.350 ;
        RECT 582.170 0.000 582.450 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 88.570 39.340 88.890 39.400 ;
        RECT 981.430 39.340 981.750 39.400 ;
        RECT 88.570 39.200 981.750 39.340 ;
        RECT 88.570 39.140 88.890 39.200 ;
        RECT 981.430 39.140 981.750 39.200 ;
        RECT 1126.790 39.340 1127.110 39.400 ;
        RECT 1127.250 39.340 1127.570 39.400 ;
        RECT 1126.790 39.200 1127.570 39.340 ;
        RECT 1126.790 39.140 1127.110 39.200 ;
        RECT 1127.250 39.140 1127.570 39.200 ;
      LAYER via ;
        RECT 88.600 39.140 88.860 39.400 ;
        RECT 981.460 39.140 981.720 39.400 ;
        RECT 1126.820 39.140 1127.080 39.400 ;
        RECT 1127.280 39.140 1127.540 39.400 ;
      LAYER met2 ;
        RECT 1170.120 39.965 1170.260 54.000 ;
        RECT 1127.270 39.595 1127.550 39.965 ;
        RECT 1170.050 39.595 1170.330 39.965 ;
        RECT 1127.340 39.430 1127.480 39.595 ;
        RECT 88.600 39.110 88.860 39.430 ;
        RECT 981.460 39.285 981.720 39.430 ;
        RECT 88.660 2.400 88.800 39.110 ;
        RECT 981.450 38.915 981.730 39.285 ;
        RECT 1126.820 39.110 1127.080 39.430 ;
        RECT 1127.280 39.110 1127.540 39.430 ;
        RECT 1126.880 37.925 1127.020 39.110 ;
        RECT 1126.810 37.555 1127.090 37.925 ;
        RECT 88.590 0.000 88.870 2.400 ;
      LAYER via2 ;
        RECT 1127.270 39.640 1127.550 39.920 ;
        RECT 1170.050 39.640 1170.330 39.920 ;
        RECT 981.450 38.960 981.730 39.240 ;
        RECT 1126.810 37.600 1127.090 37.880 ;
      LAYER met3 ;
        RECT 1127.245 39.930 1127.575 39.945 ;
        RECT 1170.025 39.930 1170.355 39.945 ;
        RECT 1127.245 39.630 1170.355 39.930 ;
        RECT 1127.245 39.615 1127.575 39.630 ;
        RECT 1170.025 39.615 1170.355 39.630 ;
        RECT 981.425 39.250 981.755 39.265 ;
        RECT 981.425 38.950 1080.410 39.250 ;
        RECT 981.425 38.935 981.755 38.950 ;
        RECT 1080.110 37.890 1080.410 38.950 ;
        RECT 1126.785 37.890 1127.115 37.905 ;
        RECT 1080.110 37.590 1127.115 37.890 ;
        RECT 1126.785 37.575 1127.115 37.590 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 617.570 52.940 617.890 53.000 ;
        RECT 1274.910 52.940 1275.230 53.000 ;
        RECT 617.570 52.800 1275.230 52.940 ;
        RECT 617.570 52.740 617.890 52.800 ;
        RECT 1274.910 52.740 1275.230 52.800 ;
        RECT 599.630 17.580 599.950 17.640 ;
        RECT 602.390 17.580 602.710 17.640 ;
        RECT 599.630 17.440 602.710 17.580 ;
        RECT 599.630 17.380 599.950 17.440 ;
        RECT 602.390 17.380 602.710 17.440 ;
      LAYER via ;
        RECT 617.600 52.740 617.860 53.000 ;
        RECT 1274.940 52.740 1275.200 53.000 ;
        RECT 599.660 17.380 599.920 17.640 ;
        RECT 602.420 17.380 602.680 17.640 ;
      LAYER met2 ;
        RECT 1275.000 53.030 1275.140 54.000 ;
        RECT 617.600 52.885 617.860 53.030 ;
        RECT 602.410 52.515 602.690 52.885 ;
        RECT 617.590 52.515 617.870 52.885 ;
        RECT 1274.940 52.710 1275.200 53.030 ;
        RECT 602.480 17.670 602.620 52.515 ;
        RECT 599.660 17.350 599.920 17.670 ;
        RECT 602.420 17.350 602.680 17.670 ;
        RECT 599.720 2.400 599.860 17.350 ;
        RECT 599.650 0.000 599.930 2.400 ;
      LAYER via2 ;
        RECT 602.410 52.560 602.690 52.840 ;
        RECT 617.590 52.560 617.870 52.840 ;
      LAYER met3 ;
        RECT 602.385 52.850 602.715 52.865 ;
        RECT 617.565 52.850 617.895 52.865 ;
        RECT 602.385 52.550 617.895 52.850 ;
        RECT 602.385 52.535 602.715 52.550 ;
        RECT 617.565 52.535 617.895 52.550 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 692.090 52.600 692.410 52.660 ;
        RECT 1273.070 52.600 1273.390 52.660 ;
        RECT 692.090 52.460 1273.390 52.600 ;
        RECT 692.090 52.400 692.410 52.460 ;
        RECT 1273.070 52.400 1273.390 52.460 ;
        RECT 623.090 48.180 623.410 48.240 ;
        RECT 691.170 48.180 691.490 48.240 ;
        RECT 623.090 48.040 691.490 48.180 ;
        RECT 623.090 47.980 623.410 48.040 ;
        RECT 691.170 47.980 691.490 48.040 ;
        RECT 617.570 17.580 617.890 17.640 ;
        RECT 623.090 17.580 623.410 17.640 ;
        RECT 617.570 17.440 623.410 17.580 ;
        RECT 617.570 17.380 617.890 17.440 ;
        RECT 623.090 17.380 623.410 17.440 ;
      LAYER via ;
        RECT 692.120 52.400 692.380 52.660 ;
        RECT 1273.100 52.400 1273.360 52.660 ;
        RECT 623.120 47.980 623.380 48.240 ;
        RECT 691.200 47.980 691.460 48.240 ;
        RECT 617.600 17.380 617.860 17.640 ;
        RECT 623.120 17.380 623.380 17.640 ;
      LAYER met2 ;
        RECT 1273.160 52.690 1273.300 54.000 ;
        RECT 692.120 52.370 692.380 52.690 ;
        RECT 1273.100 52.370 1273.360 52.690 ;
        RECT 692.180 49.370 692.320 52.370 ;
        RECT 691.260 49.230 692.320 49.370 ;
        RECT 691.260 48.270 691.400 49.230 ;
        RECT 623.120 47.950 623.380 48.270 ;
        RECT 691.200 47.950 691.460 48.270 ;
        RECT 623.180 17.670 623.320 47.950 ;
        RECT 617.600 17.350 617.860 17.670 ;
        RECT 623.120 17.350 623.380 17.670 ;
        RECT 617.660 2.400 617.800 17.350 ;
        RECT 617.590 0.000 617.870 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 157.645 44.285 157.815 45.135 ;
        RECT 182.025 44.965 182.195 45.815 ;
        RECT 213.305 44.285 213.475 45.815 ;
        RECT 271.265 44.285 271.435 45.815 ;
        RECT 326.925 44.965 327.095 45.815 ;
        RECT 375.225 44.965 375.395 45.815 ;
        RECT 406.045 44.285 406.215 45.815 ;
        RECT 429.505 44.285 430.135 44.455 ;
        RECT 464.465 44.285 464.635 45.815 ;
        RECT 520.125 44.965 520.295 45.815 ;
        RECT 568.425 44.965 568.595 45.815 ;
        RECT 581.305 44.965 581.475 45.815 ;
        RECT 700.445 44.455 700.615 45.135 ;
        RECT 700.445 44.285 701.535 44.455 ;
        RECT 813.145 43.945 813.315 45.135 ;
        RECT 861.445 42.925 861.615 45.135 ;
        RECT 909.745 42.925 909.915 45.135 ;
        RECT 958.045 42.925 958.215 45.135 ;
        RECT 1006.345 42.925 1006.515 45.135 ;
        RECT 1054.645 41.565 1054.815 45.135 ;
        RECT 1079.485 41.565 1079.655 45.135 ;
      LAYER mcon ;
        RECT 182.025 45.645 182.195 45.815 ;
        RECT 157.645 44.965 157.815 45.135 ;
        RECT 213.305 45.645 213.475 45.815 ;
        RECT 271.265 45.645 271.435 45.815 ;
        RECT 326.925 45.645 327.095 45.815 ;
        RECT 375.225 45.645 375.395 45.815 ;
        RECT 406.045 45.645 406.215 45.815 ;
        RECT 464.465 45.645 464.635 45.815 ;
        RECT 520.125 45.645 520.295 45.815 ;
        RECT 568.425 45.645 568.595 45.815 ;
        RECT 581.305 45.645 581.475 45.815 ;
        RECT 700.445 44.965 700.615 45.135 ;
        RECT 429.965 44.285 430.135 44.455 ;
        RECT 813.145 44.965 813.315 45.135 ;
        RECT 701.365 44.285 701.535 44.455 ;
        RECT 861.445 44.965 861.615 45.135 ;
        RECT 909.745 44.965 909.915 45.135 ;
        RECT 958.045 44.965 958.215 45.135 ;
        RECT 1006.345 44.965 1006.515 45.135 ;
        RECT 1054.645 44.965 1054.815 45.135 ;
        RECT 1079.485 44.965 1079.655 45.135 ;
      LAYER met1 ;
        RECT 181.965 45.800 182.255 45.845 ;
        RECT 213.245 45.800 213.535 45.845 ;
        RECT 181.965 45.660 213.535 45.800 ;
        RECT 181.965 45.615 182.255 45.660 ;
        RECT 213.245 45.615 213.535 45.660 ;
        RECT 271.205 45.800 271.495 45.845 ;
        RECT 326.865 45.800 327.155 45.845 ;
        RECT 271.205 45.660 327.155 45.800 ;
        RECT 271.205 45.615 271.495 45.660 ;
        RECT 326.865 45.615 327.155 45.660 ;
        RECT 375.165 45.800 375.455 45.845 ;
        RECT 405.985 45.800 406.275 45.845 ;
        RECT 375.165 45.660 406.275 45.800 ;
        RECT 375.165 45.615 375.455 45.660 ;
        RECT 405.985 45.615 406.275 45.660 ;
        RECT 464.405 45.800 464.695 45.845 ;
        RECT 520.065 45.800 520.355 45.845 ;
        RECT 464.405 45.660 520.355 45.800 ;
        RECT 464.405 45.615 464.695 45.660 ;
        RECT 520.065 45.615 520.355 45.660 ;
        RECT 568.365 45.800 568.655 45.845 ;
        RECT 581.245 45.800 581.535 45.845 ;
        RECT 568.365 45.660 581.535 45.800 ;
        RECT 568.365 45.615 568.655 45.660 ;
        RECT 581.245 45.615 581.535 45.660 ;
        RECT 157.585 45.120 157.875 45.165 ;
        RECT 181.965 45.120 182.255 45.165 ;
        RECT 157.585 44.980 182.255 45.120 ;
        RECT 157.585 44.935 157.875 44.980 ;
        RECT 181.965 44.935 182.255 44.980 ;
        RECT 326.865 45.120 327.155 45.165 ;
        RECT 375.165 45.120 375.455 45.165 ;
        RECT 326.865 44.980 375.455 45.120 ;
        RECT 326.865 44.935 327.155 44.980 ;
        RECT 375.165 44.935 375.455 44.980 ;
        RECT 520.065 45.120 520.355 45.165 ;
        RECT 568.365 45.120 568.655 45.165 ;
        RECT 520.065 44.980 568.655 45.120 ;
        RECT 520.065 44.935 520.355 44.980 ;
        RECT 568.365 44.935 568.655 44.980 ;
        RECT 581.245 45.120 581.535 45.165 ;
        RECT 700.385 45.120 700.675 45.165 ;
        RECT 581.245 44.980 700.675 45.120 ;
        RECT 581.245 44.935 581.535 44.980 ;
        RECT 700.385 44.935 700.675 44.980 ;
        RECT 813.085 45.120 813.375 45.165 ;
        RECT 861.385 45.120 861.675 45.165 ;
        RECT 813.085 44.980 861.675 45.120 ;
        RECT 813.085 44.935 813.375 44.980 ;
        RECT 861.385 44.935 861.675 44.980 ;
        RECT 909.685 45.120 909.975 45.165 ;
        RECT 957.985 45.120 958.275 45.165 ;
        RECT 909.685 44.980 958.275 45.120 ;
        RECT 909.685 44.935 909.975 44.980 ;
        RECT 957.985 44.935 958.275 44.980 ;
        RECT 1006.285 45.120 1006.575 45.165 ;
        RECT 1054.585 45.120 1054.875 45.165 ;
        RECT 1006.285 44.980 1054.875 45.120 ;
        RECT 1006.285 44.935 1006.575 44.980 ;
        RECT 1054.585 44.935 1054.875 44.980 ;
        RECT 1079.425 45.120 1079.715 45.165 ;
        RECT 1169.110 45.120 1169.430 45.180 ;
        RECT 1079.425 44.980 1169.430 45.120 ;
        RECT 1079.425 44.935 1079.715 44.980 ;
        RECT 1169.110 44.920 1169.430 44.980 ;
        RECT 112.030 44.440 112.350 44.500 ;
        RECT 157.585 44.440 157.875 44.485 ;
        RECT 112.030 44.300 157.875 44.440 ;
        RECT 112.030 44.240 112.350 44.300 ;
        RECT 157.585 44.255 157.875 44.300 ;
        RECT 213.245 44.440 213.535 44.485 ;
        RECT 271.205 44.440 271.495 44.485 ;
        RECT 213.245 44.300 271.495 44.440 ;
        RECT 213.245 44.255 213.535 44.300 ;
        RECT 271.205 44.255 271.495 44.300 ;
        RECT 405.985 44.440 406.275 44.485 ;
        RECT 429.445 44.440 429.735 44.485 ;
        RECT 405.985 44.300 429.735 44.440 ;
        RECT 405.985 44.255 406.275 44.300 ;
        RECT 429.445 44.255 429.735 44.300 ;
        RECT 429.905 44.440 430.195 44.485 ;
        RECT 464.405 44.440 464.695 44.485 ;
        RECT 429.905 44.300 464.695 44.440 ;
        RECT 429.905 44.255 430.195 44.300 ;
        RECT 464.405 44.255 464.695 44.300 ;
        RECT 701.305 44.440 701.595 44.485 ;
        RECT 701.305 44.300 741.080 44.440 ;
        RECT 701.305 44.255 701.595 44.300 ;
        RECT 740.940 44.100 741.080 44.300 ;
        RECT 813.085 44.100 813.375 44.145 ;
        RECT 740.940 43.960 813.375 44.100 ;
        RECT 813.085 43.915 813.375 43.960 ;
        RECT 861.385 43.080 861.675 43.125 ;
        RECT 909.685 43.080 909.975 43.125 ;
        RECT 861.385 42.940 909.975 43.080 ;
        RECT 861.385 42.895 861.675 42.940 ;
        RECT 909.685 42.895 909.975 42.940 ;
        RECT 957.985 43.080 958.275 43.125 ;
        RECT 1006.285 43.080 1006.575 43.125 ;
        RECT 957.985 42.940 1006.575 43.080 ;
        RECT 957.985 42.895 958.275 42.940 ;
        RECT 1006.285 42.895 1006.575 42.940 ;
        RECT 1054.585 41.720 1054.875 41.765 ;
        RECT 1079.425 41.720 1079.715 41.765 ;
        RECT 1054.585 41.580 1079.715 41.720 ;
        RECT 1054.585 41.535 1054.875 41.580 ;
        RECT 1079.425 41.535 1079.715 41.580 ;
      LAYER via ;
        RECT 1169.140 44.920 1169.400 45.180 ;
        RECT 112.060 44.240 112.320 44.500 ;
      LAYER met2 ;
        RECT 1169.200 45.210 1169.340 54.000 ;
        RECT 1169.140 44.890 1169.400 45.210 ;
        RECT 112.060 44.210 112.320 44.530 ;
        RECT 112.120 2.400 112.260 44.210 ;
        RECT 112.050 0.000 112.330 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1173.785 45.305 1173.955 54.000 ;
      LAYER met1 ;
        RECT 135.950 45.460 136.270 45.520 ;
        RECT 1173.725 45.460 1174.015 45.505 ;
        RECT 135.950 45.320 1174.015 45.460 ;
        RECT 135.950 45.260 136.270 45.320 ;
        RECT 1173.725 45.275 1174.015 45.320 ;
      LAYER via ;
        RECT 135.980 45.260 136.240 45.520 ;
      LAYER met2 ;
        RECT 135.980 45.230 136.240 45.550 ;
        RECT 136.040 2.400 136.180 45.230 ;
        RECT 135.970 0.000 136.250 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1183.000 51.525 1183.140 54.000 ;
        RECT 153.450 51.155 153.730 51.525 ;
        RECT 1182.930 51.155 1183.210 51.525 ;
        RECT 153.520 17.410 153.660 51.155 ;
        RECT 153.520 17.270 154.120 17.410 ;
        RECT 153.980 2.400 154.120 17.270 ;
        RECT 153.910 0.000 154.190 2.400 ;
      LAYER via2 ;
        RECT 153.450 51.200 153.730 51.480 ;
        RECT 1182.930 51.200 1183.210 51.480 ;
      LAYER met3 ;
        RECT 153.425 51.490 153.755 51.505 ;
        RECT 1182.905 51.490 1183.235 51.505 ;
        RECT 153.425 51.190 1183.235 51.490 ;
        RECT 153.425 51.175 153.755 51.190 ;
        RECT 1182.905 51.175 1183.235 51.190 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 668.245 52.105 668.415 54.000 ;
      LAYER met1 ;
        RECT 174.590 52.260 174.910 52.320 ;
        RECT 668.185 52.260 668.475 52.305 ;
        RECT 174.590 52.120 668.475 52.260 ;
        RECT 174.590 52.060 174.910 52.120 ;
        RECT 668.185 52.075 668.475 52.120 ;
        RECT 171.830 17.580 172.150 17.640 ;
        RECT 174.590 17.580 174.910 17.640 ;
        RECT 171.830 17.440 174.910 17.580 ;
        RECT 171.830 17.380 172.150 17.440 ;
        RECT 174.590 17.380 174.910 17.440 ;
      LAYER via ;
        RECT 174.620 52.060 174.880 52.320 ;
        RECT 171.860 17.380 172.120 17.640 ;
        RECT 174.620 17.380 174.880 17.640 ;
      LAYER met2 ;
        RECT 174.620 52.030 174.880 52.350 ;
        RECT 174.680 17.670 174.820 52.030 ;
        RECT 171.860 17.350 172.120 17.670 ;
        RECT 174.620 17.350 174.880 17.670 ;
        RECT 171.920 2.400 172.060 17.350 ;
        RECT 171.850 0.000 172.130 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 616.725 52.445 616.895 54.000 ;
        RECT 644.785 53.805 644.955 54.000 ;
        RECT 861.905 53.295 862.075 53.635 ;
        RECT 884.445 53.465 884.615 54.000 ;
        RECT 860.985 53.125 862.075 53.295 ;
        RECT 1150.785 53.125 1150.955 53.975 ;
      LAYER mcon ;
        RECT 861.905 53.465 862.075 53.635 ;
        RECT 1150.785 53.805 1150.955 53.975 ;
      LAYER met1 ;
        RECT 644.725 53.960 645.015 54.000 ;
        RECT 739.010 53.960 739.330 54.000 ;
        RECT 644.725 53.820 739.330 53.960 ;
        RECT 644.725 53.775 645.015 53.820 ;
        RECT 739.010 53.760 739.330 53.820 ;
        RECT 742.230 53.960 742.550 54.000 ;
        RECT 765.230 53.960 765.550 54.000 ;
        RECT 742.230 53.820 765.550 53.960 ;
        RECT 742.230 53.760 742.550 53.820 ;
        RECT 765.230 53.760 765.550 53.820 ;
        RECT 935.430 53.960 935.750 54.000 ;
        RECT 958.430 53.960 958.750 54.000 ;
        RECT 935.430 53.820 958.750 53.960 ;
        RECT 935.430 53.760 935.750 53.820 ;
        RECT 958.430 53.760 958.750 53.820 ;
        RECT 1150.725 53.960 1151.015 54.000 ;
        RECT 1173.250 53.960 1173.570 54.000 ;
        RECT 1150.725 53.820 1173.570 53.960 ;
        RECT 1150.725 53.775 1151.015 53.820 ;
        RECT 1173.250 53.760 1173.570 53.820 ;
        RECT 861.845 53.620 862.135 53.665 ;
        RECT 884.385 53.620 884.675 53.665 ;
        RECT 861.845 53.480 884.675 53.620 ;
        RECT 861.845 53.435 862.135 53.480 ;
        RECT 884.385 53.435 884.675 53.480 ;
        RECT 765.230 53.280 765.550 53.340 ;
        RECT 860.925 53.280 861.215 53.325 ;
        RECT 765.230 53.140 861.215 53.280 ;
        RECT 765.230 53.080 765.550 53.140 ;
        RECT 860.925 53.095 861.215 53.140 ;
        RECT 958.430 53.280 958.750 53.340 ;
        RECT 1150.725 53.280 1151.015 53.325 ;
        RECT 958.430 53.140 1151.015 53.280 ;
        RECT 958.430 53.080 958.750 53.140 ;
        RECT 1150.725 53.095 1151.015 53.140 ;
        RECT 1176.930 53.280 1177.250 53.340 ;
        RECT 1191.190 53.280 1191.510 53.340 ;
        RECT 1176.930 53.140 1191.510 53.280 ;
        RECT 1176.930 53.080 1177.250 53.140 ;
        RECT 1191.190 53.080 1191.510 53.140 ;
        RECT 195.290 52.600 195.610 52.660 ;
        RECT 616.665 52.600 616.955 52.645 ;
        RECT 195.290 52.460 616.955 52.600 ;
        RECT 195.290 52.400 195.610 52.460 ;
        RECT 616.665 52.415 616.955 52.460 ;
        RECT 189.310 17.920 189.630 17.980 ;
        RECT 195.290 17.920 195.610 17.980 ;
        RECT 189.310 17.780 195.610 17.920 ;
        RECT 189.310 17.720 189.630 17.780 ;
        RECT 195.290 17.720 195.610 17.780 ;
      LAYER via ;
        RECT 739.040 53.760 739.300 54.000 ;
        RECT 742.260 53.760 742.520 54.000 ;
        RECT 765.260 53.760 765.520 54.000 ;
        RECT 935.460 53.760 935.720 54.000 ;
        RECT 958.460 53.760 958.720 54.000 ;
        RECT 1173.280 53.760 1173.540 54.000 ;
        RECT 765.260 53.080 765.520 53.340 ;
        RECT 958.460 53.080 958.720 53.340 ;
        RECT 1176.960 53.080 1177.220 53.340 ;
        RECT 1191.220 53.080 1191.480 53.340 ;
        RECT 195.320 52.400 195.580 52.660 ;
        RECT 189.340 17.720 189.600 17.980 ;
        RECT 195.320 17.720 195.580 17.980 ;
      LAYER met2 ;
        RECT 739.040 53.730 739.300 54.000 ;
        RECT 742.260 53.730 742.520 54.000 ;
        RECT 765.260 53.730 765.520 54.000 ;
        RECT 739.100 52.885 739.240 53.730 ;
        RECT 742.320 52.885 742.460 53.730 ;
        RECT 765.320 53.370 765.460 53.730 ;
        RECT 765.260 53.050 765.520 53.370 ;
        RECT 886.300 52.885 886.440 54.000 ;
        RECT 935.460 53.730 935.720 54.000 ;
        RECT 958.460 53.730 958.720 54.000 ;
        RECT 1173.280 53.730 1173.540 54.000 ;
        RECT 935.520 52.885 935.660 53.730 ;
        RECT 958.520 53.370 958.660 53.730 ;
        RECT 958.460 53.050 958.720 53.370 ;
        RECT 1173.340 52.885 1173.480 53.730 ;
        RECT 1191.280 53.370 1191.420 54.000 ;
        RECT 1176.960 53.050 1177.220 53.370 ;
        RECT 1191.220 53.050 1191.480 53.370 ;
        RECT 1177.020 52.885 1177.160 53.050 ;
        RECT 195.320 52.370 195.580 52.690 ;
        RECT 739.030 52.515 739.310 52.885 ;
        RECT 742.250 52.515 742.530 52.885 ;
        RECT 886.230 52.515 886.510 52.885 ;
        RECT 935.450 52.515 935.730 52.885 ;
        RECT 1173.270 52.515 1173.550 52.885 ;
        RECT 1176.950 52.515 1177.230 52.885 ;
        RECT 195.380 18.010 195.520 52.370 ;
        RECT 189.340 17.690 189.600 18.010 ;
        RECT 195.320 17.690 195.580 18.010 ;
        RECT 189.400 2.400 189.540 17.690 ;
        RECT 189.330 0.000 189.610 2.400 ;
      LAYER via2 ;
        RECT 739.030 52.560 739.310 52.840 ;
        RECT 742.250 52.560 742.530 52.840 ;
        RECT 886.230 52.560 886.510 52.840 ;
        RECT 935.450 52.560 935.730 52.840 ;
        RECT 1173.270 52.560 1173.550 52.840 ;
        RECT 1176.950 52.560 1177.230 52.840 ;
      LAYER met3 ;
        RECT 739.005 52.850 739.335 52.865 ;
        RECT 742.225 52.850 742.555 52.865 ;
        RECT 739.005 52.550 742.555 52.850 ;
        RECT 739.005 52.535 739.335 52.550 ;
        RECT 742.225 52.535 742.555 52.550 ;
        RECT 886.205 52.850 886.535 52.865 ;
        RECT 935.425 52.850 935.755 52.865 ;
        RECT 886.205 52.550 935.755 52.850 ;
        RECT 886.205 52.535 886.535 52.550 ;
        RECT 935.425 52.535 935.755 52.550 ;
        RECT 1173.245 52.850 1173.575 52.865 ;
        RECT 1176.925 52.850 1177.255 52.865 ;
        RECT 1173.245 52.550 1177.255 52.850 ;
        RECT 1173.245 52.535 1173.575 52.550 ;
        RECT 1176.925 52.535 1177.255 52.550 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 739.545 53.465 739.715 54.000 ;
        RECT 741.845 53.465 742.015 54.000 ;
        RECT 764.385 53.805 765.935 53.975 ;
        RECT 883.525 53.805 883.695 54.000 ;
        RECT 764.385 53.465 764.555 53.805 ;
        RECT 935.045 53.465 935.215 54.000 ;
        RECT 957.585 53.805 959.135 53.975 ;
        RECT 1150.325 53.805 1150.495 54.000 ;
        RECT 957.585 53.465 957.755 53.805 ;
        RECT 1151.705 53.465 1151.875 54.000 ;
        RECT 1177.465 53.805 1177.635 54.000 ;
        RECT 668.705 52.445 668.875 53.295 ;
      LAYER mcon ;
        RECT 765.765 53.805 765.935 53.975 ;
        RECT 958.965 53.805 959.135 53.975 ;
        RECT 668.705 53.125 668.875 53.295 ;
      LAYER met1 ;
        RECT 765.705 53.960 765.995 54.000 ;
        RECT 883.465 53.960 883.755 54.000 ;
        RECT 765.705 53.820 883.755 53.960 ;
        RECT 765.705 53.775 765.995 53.820 ;
        RECT 883.465 53.775 883.755 53.820 ;
        RECT 958.905 53.960 959.195 54.000 ;
        RECT 1150.265 53.960 1150.555 54.000 ;
        RECT 958.905 53.820 1150.555 53.960 ;
        RECT 958.905 53.775 959.195 53.820 ;
        RECT 1150.265 53.775 1150.555 53.820 ;
        RECT 1177.405 53.960 1177.695 54.000 ;
        RECT 1190.730 53.960 1191.050 54.000 ;
        RECT 1177.405 53.820 1191.050 53.960 ;
        RECT 1177.405 53.775 1177.695 53.820 ;
        RECT 1190.730 53.760 1191.050 53.820 ;
        RECT 739.485 53.620 739.775 53.665 ;
        RECT 717.020 53.480 739.775 53.620 ;
        RECT 668.645 53.280 668.935 53.325 ;
        RECT 717.020 53.280 717.160 53.480 ;
        RECT 739.485 53.435 739.775 53.480 ;
        RECT 741.785 53.620 742.075 53.665 ;
        RECT 764.325 53.620 764.615 53.665 ;
        RECT 741.785 53.480 764.615 53.620 ;
        RECT 741.785 53.435 742.075 53.480 ;
        RECT 764.325 53.435 764.615 53.480 ;
        RECT 934.985 53.620 935.275 53.665 ;
        RECT 957.525 53.620 957.815 53.665 ;
        RECT 934.985 53.480 957.815 53.620 ;
        RECT 934.985 53.435 935.275 53.480 ;
        RECT 957.525 53.435 957.815 53.480 ;
        RECT 1151.645 53.620 1151.935 53.665 ;
        RECT 1174.170 53.620 1174.490 53.680 ;
        RECT 1151.645 53.480 1174.490 53.620 ;
        RECT 1151.645 53.435 1151.935 53.480 ;
        RECT 1174.170 53.420 1174.490 53.480 ;
        RECT 668.645 53.140 717.160 53.280 ;
        RECT 668.645 53.095 668.935 53.140 ;
        RECT 209.090 52.940 209.410 53.000 ;
        RECT 209.090 52.800 617.340 52.940 ;
        RECT 209.090 52.740 209.410 52.800 ;
        RECT 617.200 52.600 617.340 52.800 ;
        RECT 668.645 52.600 668.935 52.645 ;
        RECT 617.200 52.460 668.935 52.600 ;
        RECT 668.645 52.415 668.935 52.460 ;
      LAYER via ;
        RECT 1190.760 53.760 1191.020 54.000 ;
        RECT 1174.200 53.420 1174.460 53.680 ;
        RECT 209.120 52.740 209.380 53.000 ;
      LAYER met2 ;
        RECT 1174.260 53.710 1174.400 54.000 ;
        RECT 1190.760 53.730 1191.020 54.000 ;
        RECT 1174.200 53.390 1174.460 53.710 ;
        RECT 209.120 52.710 209.380 53.030 ;
        RECT 209.180 16.730 209.320 52.710 ;
        RECT 207.340 16.590 209.320 16.730 ;
        RECT 207.340 2.400 207.480 16.590 ;
        RECT 207.270 0.000 207.550 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 716.545 53.465 717.635 53.635 ;
        RECT 717.465 53.125 717.635 53.465 ;
      LAYER met1 ;
        RECT 716.485 53.620 716.775 53.665 ;
        RECT 1196.250 53.620 1196.570 53.680 ;
        RECT 668.260 53.480 716.775 53.620 ;
        RECT 229.790 53.280 230.110 53.340 ;
        RECT 668.260 53.280 668.400 53.480 ;
        RECT 716.485 53.435 716.775 53.480 ;
        RECT 764.860 53.480 861.600 53.620 ;
        RECT 229.790 53.140 668.400 53.280 ;
        RECT 717.405 53.280 717.695 53.325 ;
        RECT 764.860 53.280 765.000 53.480 ;
        RECT 717.405 53.140 765.000 53.280 ;
        RECT 861.460 53.280 861.600 53.480 ;
        RECT 958.060 53.480 1151.400 53.620 ;
        RECT 958.060 53.280 958.200 53.480 ;
        RECT 861.460 53.140 958.200 53.280 ;
        RECT 1151.260 53.280 1151.400 53.480 ;
        RECT 1176.100 53.480 1196.570 53.620 ;
        RECT 1176.100 53.280 1176.240 53.480 ;
        RECT 1196.250 53.420 1196.570 53.480 ;
        RECT 1151.260 53.140 1176.240 53.280 ;
        RECT 229.790 53.080 230.110 53.140 ;
        RECT 717.405 53.095 717.695 53.140 ;
        RECT 225.190 16.900 225.510 16.960 ;
        RECT 229.790 16.900 230.110 16.960 ;
        RECT 225.190 16.760 230.110 16.900 ;
        RECT 225.190 16.700 225.510 16.760 ;
        RECT 229.790 16.700 230.110 16.760 ;
      LAYER via ;
        RECT 229.820 53.080 230.080 53.340 ;
        RECT 1196.280 53.420 1196.540 53.680 ;
        RECT 225.220 16.700 225.480 16.960 ;
        RECT 229.820 16.700 230.080 16.960 ;
      LAYER met2 ;
        RECT 1196.340 53.710 1196.480 54.000 ;
        RECT 1196.280 53.390 1196.540 53.710 ;
        RECT 229.820 53.050 230.080 53.370 ;
        RECT 229.880 16.990 230.020 53.050 ;
        RECT 225.220 16.670 225.480 16.990 ;
        RECT 229.820 16.670 230.080 16.990 ;
        RECT 225.280 2.400 225.420 16.670 ;
        RECT 225.210 0.000 225.490 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1079.410 39.340 1079.730 39.400 ;
        RECT 1126.330 39.340 1126.650 39.400 ;
        RECT 1079.410 39.200 1126.650 39.340 ;
        RECT 1079.410 39.140 1079.730 39.200 ;
        RECT 1126.330 39.140 1126.650 39.200 ;
        RECT 1127.710 39.340 1128.030 39.400 ;
        RECT 1156.230 39.340 1156.550 39.400 ;
        RECT 1127.710 39.200 1156.550 39.340 ;
        RECT 1127.710 39.140 1128.030 39.200 ;
        RECT 1156.230 39.140 1156.550 39.200 ;
        RECT 22.790 38.660 23.110 38.720 ;
        RECT 968.090 38.660 968.410 38.720 ;
        RECT 22.790 38.520 968.410 38.660 ;
        RECT 22.790 38.460 23.110 38.520 ;
        RECT 968.090 38.460 968.410 38.520 ;
      LAYER via ;
        RECT 1079.440 39.140 1079.700 39.400 ;
        RECT 1126.360 39.140 1126.620 39.400 ;
        RECT 1127.740 39.140 1128.000 39.400 ;
        RECT 1156.260 39.140 1156.520 39.400 ;
        RECT 22.820 38.460 23.080 38.720 ;
        RECT 968.120 38.460 968.380 38.720 ;
      LAYER met2 ;
        RECT 1156.320 39.430 1156.460 54.000 ;
        RECT 1079.440 39.110 1079.700 39.430 ;
        RECT 1126.360 39.110 1126.620 39.430 ;
        RECT 1127.740 39.110 1128.000 39.430 ;
        RECT 1156.260 39.110 1156.520 39.430 ;
        RECT 22.820 38.430 23.080 38.750 ;
        RECT 968.120 38.605 968.380 38.750 ;
        RECT 1079.500 38.605 1079.640 39.110 ;
        RECT 1126.420 38.605 1126.560 39.110 ;
        RECT 1127.800 38.605 1127.940 39.110 ;
        RECT 22.880 2.400 23.020 38.430 ;
        RECT 968.110 38.235 968.390 38.605 ;
        RECT 1079.430 38.235 1079.710 38.605 ;
        RECT 1126.350 38.235 1126.630 38.605 ;
        RECT 1127.730 38.235 1128.010 38.605 ;
        RECT 22.810 0.000 23.090 2.400 ;
      LAYER via2 ;
        RECT 968.110 38.280 968.390 38.560 ;
        RECT 1079.430 38.280 1079.710 38.560 ;
        RECT 1126.350 38.280 1126.630 38.560 ;
        RECT 1127.730 38.280 1128.010 38.560 ;
      LAYER met3 ;
        RECT 968.085 38.570 968.415 38.585 ;
        RECT 1079.405 38.570 1079.735 38.585 ;
        RECT 968.085 38.270 1079.735 38.570 ;
        RECT 968.085 38.255 968.415 38.270 ;
        RECT 1079.405 38.255 1079.735 38.270 ;
        RECT 1126.325 38.570 1126.655 38.585 ;
        RECT 1127.705 38.570 1128.035 38.585 ;
        RECT 1126.325 38.270 1128.035 38.570 ;
        RECT 1126.325 38.255 1126.655 38.270 ;
        RECT 1127.705 38.255 1128.035 38.270 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 92.325 44.625 92.495 45.815 ;
        RECT 140.165 44.625 140.335 45.815 ;
        RECT 428.585 44.965 430.135 45.135 ;
        RECT 188.925 42.925 189.095 44.795 ;
        RECT 236.765 42.925 236.935 44.795 ;
        RECT 285.525 43.945 285.695 44.795 ;
        RECT 333.365 43.945 333.535 44.795 ;
        RECT 340.725 43.945 340.895 44.795 ;
        RECT 428.585 43.945 428.755 44.965 ;
        RECT 575.325 42.925 575.495 44.795 ;
        RECT 623.165 42.925 623.335 44.795 ;
        RECT 671.925 43.945 672.095 44.795 ;
        RECT 692.625 44.115 692.795 44.795 ;
        RECT 692.165 43.945 692.795 44.115 ;
      LAYER mcon ;
        RECT 92.325 45.645 92.495 45.815 ;
        RECT 140.165 45.645 140.335 45.815 ;
        RECT 429.965 44.965 430.135 45.135 ;
        RECT 188.925 44.625 189.095 44.795 ;
        RECT 236.765 44.625 236.935 44.795 ;
        RECT 285.525 44.625 285.695 44.795 ;
        RECT 333.365 44.625 333.535 44.795 ;
        RECT 340.725 44.625 340.895 44.795 ;
        RECT 575.325 44.625 575.495 44.795 ;
        RECT 623.165 44.625 623.335 44.795 ;
        RECT 671.925 44.625 672.095 44.795 ;
        RECT 692.625 44.625 692.795 44.795 ;
      LAYER met1 ;
        RECT 92.265 45.800 92.555 45.845 ;
        RECT 140.105 45.800 140.395 45.845 ;
        RECT 92.265 45.660 140.395 45.800 ;
        RECT 92.265 45.615 92.555 45.660 ;
        RECT 140.105 45.615 140.395 45.660 ;
        RECT 429.905 44.935 430.195 45.165 ;
        RECT 46.710 44.780 47.030 44.840 ;
        RECT 92.265 44.780 92.555 44.825 ;
        RECT 46.710 44.640 92.555 44.780 ;
        RECT 46.710 44.580 47.030 44.640 ;
        RECT 92.265 44.595 92.555 44.640 ;
        RECT 140.105 44.780 140.395 44.825 ;
        RECT 188.865 44.780 189.155 44.825 ;
        RECT 140.105 44.640 189.155 44.780 ;
        RECT 140.105 44.595 140.395 44.640 ;
        RECT 188.865 44.595 189.155 44.640 ;
        RECT 236.705 44.780 236.995 44.825 ;
        RECT 285.465 44.780 285.755 44.825 ;
        RECT 236.705 44.640 285.755 44.780 ;
        RECT 236.705 44.595 236.995 44.640 ;
        RECT 285.465 44.595 285.755 44.640 ;
        RECT 333.305 44.780 333.595 44.825 ;
        RECT 340.665 44.780 340.955 44.825 ;
        RECT 333.305 44.640 340.955 44.780 ;
        RECT 429.980 44.780 430.120 44.935 ;
        RECT 575.265 44.780 575.555 44.825 ;
        RECT 429.980 44.640 575.555 44.780 ;
        RECT 333.305 44.595 333.595 44.640 ;
        RECT 340.665 44.595 340.955 44.640 ;
        RECT 575.265 44.595 575.555 44.640 ;
        RECT 623.105 44.780 623.395 44.825 ;
        RECT 671.865 44.780 672.155 44.825 ;
        RECT 623.105 44.640 672.155 44.780 ;
        RECT 623.105 44.595 623.395 44.640 ;
        RECT 671.865 44.595 672.155 44.640 ;
        RECT 692.565 44.780 692.855 44.825 ;
        RECT 1156.690 44.780 1157.010 44.840 ;
        RECT 692.565 44.640 1157.010 44.780 ;
        RECT 692.565 44.595 692.855 44.640 ;
        RECT 1156.690 44.580 1157.010 44.640 ;
        RECT 285.465 44.100 285.755 44.145 ;
        RECT 333.305 44.100 333.595 44.145 ;
        RECT 285.465 43.960 333.595 44.100 ;
        RECT 285.465 43.915 285.755 43.960 ;
        RECT 333.305 43.915 333.595 43.960 ;
        RECT 340.665 44.100 340.955 44.145 ;
        RECT 428.525 44.100 428.815 44.145 ;
        RECT 340.665 43.960 428.815 44.100 ;
        RECT 340.665 43.915 340.955 43.960 ;
        RECT 428.525 43.915 428.815 43.960 ;
        RECT 671.865 44.100 672.155 44.145 ;
        RECT 692.105 44.100 692.395 44.145 ;
        RECT 671.865 43.960 692.395 44.100 ;
        RECT 671.865 43.915 672.155 43.960 ;
        RECT 692.105 43.915 692.395 43.960 ;
        RECT 188.865 43.080 189.155 43.125 ;
        RECT 236.705 43.080 236.995 43.125 ;
        RECT 188.865 42.940 236.995 43.080 ;
        RECT 188.865 42.895 189.155 42.940 ;
        RECT 236.705 42.895 236.995 42.940 ;
        RECT 575.265 43.080 575.555 43.125 ;
        RECT 623.105 43.080 623.395 43.125 ;
        RECT 575.265 42.940 623.395 43.080 ;
        RECT 575.265 42.895 575.555 42.940 ;
        RECT 623.105 42.895 623.395 42.940 ;
      LAYER via ;
        RECT 46.740 44.580 47.000 44.840 ;
        RECT 1156.720 44.580 1156.980 44.840 ;
      LAYER met2 ;
        RECT 1156.780 44.870 1156.920 54.000 ;
        RECT 46.740 44.550 47.000 44.870 ;
        RECT 1156.720 44.550 1156.980 44.870 ;
        RECT 46.800 2.400 46.940 44.550 ;
        RECT 46.730 0.000 47.010 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 667.785 51.085 667.955 53.635 ;
        RECT 740.005 51.255 740.175 53.635 ;
        RECT 740.925 53.465 741.095 54.000 ;
        RECT 716.085 50.575 716.255 51.255 ;
        RECT 739.085 51.085 740.175 51.255 ;
        RECT 788.305 51.085 788.475 54.000 ;
        RECT 837.985 51.255 838.155 54.000 ;
        RECT 883.985 53.295 884.155 54.000 ;
        RECT 884.905 53.295 885.075 53.635 ;
        RECT 883.985 53.125 885.075 53.295 ;
        RECT 837.525 51.085 838.155 51.255 ;
        RECT 716.085 50.405 717.175 50.575 ;
        RECT 739.085 50.405 739.255 51.085 ;
        RECT 1174.705 50.745 1174.875 53.635 ;
        RECT 1175.625 53.465 1176.715 53.635 ;
        RECT 1176.545 51.085 1176.715 53.465 ;
      LAYER mcon ;
        RECT 667.785 53.465 667.955 53.635 ;
        RECT 740.005 53.465 740.175 53.635 ;
        RECT 716.085 51.085 716.255 51.255 ;
        RECT 884.905 53.465 885.075 53.635 ;
        RECT 1174.705 53.465 1174.875 53.635 ;
        RECT 717.005 50.405 717.175 50.575 ;
      LAYER met1 ;
        RECT 250.490 53.620 250.810 53.680 ;
        RECT 667.725 53.620 668.015 53.665 ;
        RECT 250.490 53.480 668.015 53.620 ;
        RECT 250.490 53.420 250.810 53.480 ;
        RECT 667.725 53.435 668.015 53.480 ;
        RECT 739.945 53.620 740.235 53.665 ;
        RECT 740.865 53.620 741.155 53.665 ;
        RECT 739.945 53.480 741.155 53.620 ;
        RECT 739.945 53.435 740.235 53.480 ;
        RECT 740.865 53.435 741.155 53.480 ;
        RECT 884.845 53.620 885.135 53.665 ;
        RECT 934.050 53.620 934.370 53.680 ;
        RECT 884.845 53.480 934.370 53.620 ;
        RECT 884.845 53.435 885.135 53.480 ;
        RECT 934.050 53.420 934.370 53.480 ;
        RECT 1174.645 53.620 1174.935 53.665 ;
        RECT 1175.565 53.620 1175.855 53.665 ;
        RECT 1174.645 53.480 1175.855 53.620 ;
        RECT 1174.645 53.435 1174.935 53.480 ;
        RECT 1175.565 53.435 1175.855 53.480 ;
        RECT 667.725 51.240 668.015 51.285 ;
        RECT 716.025 51.240 716.315 51.285 ;
        RECT 667.725 51.100 716.315 51.240 ;
        RECT 667.725 51.055 668.015 51.100 ;
        RECT 716.025 51.055 716.315 51.100 ;
        RECT 788.245 51.240 788.535 51.285 ;
        RECT 837.465 51.240 837.755 51.285 ;
        RECT 788.245 51.100 837.755 51.240 ;
        RECT 788.245 51.055 788.535 51.100 ;
        RECT 837.465 51.055 837.755 51.100 ;
        RECT 981.890 51.240 982.210 51.300 ;
        RECT 1176.485 51.240 1176.775 51.285 ;
        RECT 1198.090 51.240 1198.410 51.300 ;
        RECT 981.890 51.100 1127.940 51.240 ;
        RECT 981.890 51.040 982.210 51.100 ;
        RECT 1127.800 50.900 1127.940 51.100 ;
        RECT 1176.485 51.100 1198.410 51.240 ;
        RECT 1176.485 51.055 1176.775 51.100 ;
        RECT 1198.090 51.040 1198.410 51.100 ;
        RECT 1174.645 50.900 1174.935 50.945 ;
        RECT 1127.800 50.760 1174.935 50.900 ;
        RECT 1174.645 50.715 1174.935 50.760 ;
        RECT 716.945 50.560 717.235 50.605 ;
        RECT 739.025 50.560 739.315 50.605 ;
        RECT 716.945 50.420 739.315 50.560 ;
        RECT 716.945 50.375 717.235 50.420 ;
        RECT 739.025 50.375 739.315 50.420 ;
      LAYER via ;
        RECT 250.520 53.420 250.780 53.680 ;
        RECT 934.080 53.420 934.340 53.680 ;
        RECT 981.920 51.040 982.180 51.300 ;
        RECT 1198.120 51.040 1198.380 51.300 ;
      LAYER met2 ;
        RECT 250.520 53.390 250.780 53.710 ;
        RECT 934.080 53.565 934.340 53.710 ;
        RECT 250.580 16.900 250.720 53.390 ;
        RECT 934.070 53.195 934.350 53.565 ;
        RECT 981.910 53.195 982.190 53.565 ;
        RECT 981.980 51.330 982.120 53.195 ;
        RECT 1198.180 51.330 1198.320 54.000 ;
        RECT 981.920 51.010 982.180 51.330 ;
        RECT 1198.120 51.010 1198.380 51.330 ;
        RECT 249.200 16.760 250.720 16.900 ;
        RECT 249.200 2.400 249.340 16.760 ;
        RECT 249.130 0.000 249.410 2.400 ;
      LAYER via2 ;
        RECT 934.070 53.240 934.350 53.520 ;
        RECT 981.910 53.240 982.190 53.520 ;
      LAYER met3 ;
        RECT 934.045 53.530 934.375 53.545 ;
        RECT 981.885 53.530 982.215 53.545 ;
        RECT 934.045 53.230 982.215 53.530 ;
        RECT 934.045 53.215 934.375 53.230 ;
        RECT 981.885 53.215 982.215 53.230 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 644.325 50.915 644.495 53.975 ;
        RECT 669.625 51.935 669.795 52.615 ;
        RECT 691.705 52.445 692.335 52.615 ;
        RECT 668.245 51.765 669.795 51.935 ;
        RECT 668.245 50.915 668.415 51.765 ;
        RECT 644.325 50.745 644.955 50.915 ;
        RECT 666.865 50.745 668.415 50.915 ;
        RECT 692.165 50.745 692.335 52.445 ;
        RECT 692.625 50.745 692.795 54.000 ;
        RECT 740.465 53.805 740.635 54.000 ;
        RECT 741.385 53.805 741.555 54.000 ;
        RECT 788.765 50.745 788.935 54.000 ;
        RECT 885.365 53.805 885.535 54.000 ;
        RECT 934.585 53.805 934.755 54.000 ;
        RECT 981.045 50.745 981.215 54.000 ;
        RECT 1177.005 50.745 1177.175 53.975 ;
      LAYER mcon ;
        RECT 644.325 53.805 644.495 53.975 ;
        RECT 669.625 52.445 669.795 52.615 ;
        RECT 644.785 50.745 644.955 50.915 ;
        RECT 1177.005 53.805 1177.175 53.975 ;
      LAYER met1 ;
        RECT 266.590 53.960 266.910 54.000 ;
        RECT 644.265 53.960 644.555 54.000 ;
        RECT 266.590 53.820 644.555 53.960 ;
        RECT 266.590 53.760 266.910 53.820 ;
        RECT 644.265 53.775 644.555 53.820 ;
        RECT 740.405 53.960 740.695 54.000 ;
        RECT 741.325 53.960 741.615 54.000 ;
        RECT 740.405 53.820 741.615 53.960 ;
        RECT 740.405 53.775 740.695 53.820 ;
        RECT 741.325 53.775 741.615 53.820 ;
        RECT 885.305 53.960 885.595 54.000 ;
        RECT 934.525 53.960 934.815 54.000 ;
        RECT 885.305 53.820 934.815 53.960 ;
        RECT 885.305 53.775 885.595 53.820 ;
        RECT 934.525 53.775 934.815 53.820 ;
        RECT 1175.090 53.960 1175.410 54.000 ;
        RECT 1176.945 53.960 1177.235 54.000 ;
        RECT 1175.090 53.820 1177.235 53.960 ;
        RECT 1175.090 53.760 1175.410 53.820 ;
        RECT 1176.945 53.775 1177.235 53.820 ;
        RECT 669.565 52.600 669.855 52.645 ;
        RECT 691.645 52.600 691.935 52.645 ;
        RECT 669.565 52.460 691.935 52.600 ;
        RECT 669.565 52.415 669.855 52.460 ;
        RECT 691.645 52.415 691.935 52.460 ;
        RECT 644.725 50.900 645.015 50.945 ;
        RECT 666.805 50.900 667.095 50.945 ;
        RECT 644.725 50.760 667.095 50.900 ;
        RECT 644.725 50.715 645.015 50.760 ;
        RECT 666.805 50.715 667.095 50.760 ;
        RECT 692.105 50.900 692.395 50.945 ;
        RECT 692.565 50.900 692.855 50.945 ;
        RECT 692.105 50.760 692.855 50.900 ;
        RECT 692.105 50.715 692.395 50.760 ;
        RECT 692.565 50.715 692.855 50.760 ;
        RECT 788.705 50.900 788.995 50.945 ;
        RECT 837.910 50.900 838.230 50.960 ;
        RECT 788.705 50.760 838.230 50.900 ;
        RECT 788.705 50.715 788.995 50.760 ;
        RECT 837.910 50.700 838.230 50.760 ;
        RECT 980.985 50.900 981.275 50.945 ;
        RECT 1127.250 50.900 1127.570 50.960 ;
        RECT 980.985 50.760 1127.570 50.900 ;
        RECT 980.985 50.715 981.275 50.760 ;
        RECT 1127.250 50.700 1127.570 50.760 ;
        RECT 1176.945 50.900 1177.235 50.945 ;
        RECT 1204.530 50.900 1204.850 50.960 ;
        RECT 1176.945 50.760 1204.850 50.900 ;
        RECT 1176.945 50.715 1177.235 50.760 ;
        RECT 1204.530 50.700 1204.850 50.760 ;
      LAYER via ;
        RECT 266.620 53.760 266.880 54.000 ;
        RECT 1175.120 53.760 1175.380 54.000 ;
        RECT 837.940 50.700 838.200 50.960 ;
        RECT 1127.280 50.700 1127.540 50.960 ;
        RECT 1204.560 50.700 1204.820 50.960 ;
      LAYER met2 ;
        RECT 266.620 53.730 266.880 54.000 ;
        RECT 266.680 2.400 266.820 53.730 ;
        RECT 838.000 50.990 838.140 54.000 ;
        RECT 1175.120 53.730 1175.380 54.000 ;
        RECT 1175.180 53.565 1175.320 53.730 ;
        RECT 1127.270 53.195 1127.550 53.565 ;
        RECT 1175.110 53.195 1175.390 53.565 ;
        RECT 1127.340 50.990 1127.480 53.195 ;
        RECT 1204.620 50.990 1204.760 54.000 ;
        RECT 837.940 50.670 838.200 50.990 ;
        RECT 1127.280 50.670 1127.540 50.990 ;
        RECT 1204.560 50.670 1204.820 50.990 ;
        RECT 266.610 0.000 266.890 2.400 ;
      LAYER via2 ;
        RECT 1127.270 53.240 1127.550 53.520 ;
        RECT 1175.110 53.240 1175.390 53.520 ;
      LAYER met3 ;
        RECT 1127.245 53.530 1127.575 53.545 ;
        RECT 1175.085 53.530 1175.415 53.545 ;
        RECT 1127.245 53.230 1175.415 53.530 ;
        RECT 1127.245 53.215 1127.575 53.230 ;
        RECT 1175.085 53.215 1175.415 53.230 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 691.245 50.575 691.415 54.000 ;
        RECT 691.245 50.405 691.875 50.575 ;
        RECT 1127.785 50.405 1127.955 54.000 ;
      LAYER mcon ;
        RECT 691.705 50.405 691.875 50.575 ;
      LAYER met1 ;
        RECT 716.470 51.240 716.790 51.300 ;
        RECT 716.470 51.100 788.000 51.240 ;
        RECT 716.470 51.040 716.790 51.100 ;
        RECT 787.860 50.900 788.000 51.100 ;
        RECT 838.460 51.100 980.740 51.240 ;
        RECT 787.860 50.760 788.460 50.900 ;
        RECT 691.645 50.560 691.935 50.605 ;
        RECT 716.470 50.560 716.790 50.620 ;
        RECT 691.645 50.420 716.790 50.560 ;
        RECT 788.320 50.560 788.460 50.760 ;
        RECT 838.460 50.560 838.600 51.100 ;
        RECT 788.320 50.420 838.600 50.560 ;
        RECT 980.600 50.560 980.740 51.100 ;
        RECT 1127.725 50.560 1128.015 50.605 ;
        RECT 980.600 50.420 1128.015 50.560 ;
        RECT 691.645 50.375 691.935 50.420 ;
        RECT 716.470 50.360 716.790 50.420 ;
        RECT 1127.725 50.375 1128.015 50.420 ;
      LAYER via ;
        RECT 716.500 51.040 716.760 51.300 ;
        RECT 716.500 50.360 716.760 50.620 ;
      LAYER met2 ;
        RECT 284.620 2.400 284.760 54.000 ;
        RECT 716.500 51.010 716.760 51.330 ;
        RECT 716.560 50.650 716.700 51.010 ;
        RECT 716.500 50.330 716.760 50.650 ;
        RECT 284.550 0.000 284.830 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1161.825 51.085 1162.455 51.255 ;
        RECT 690.785 48.195 690.955 50.915 ;
        RECT 690.785 48.025 691.875 48.195 ;
        RECT 740.465 47.685 740.635 50.915 ;
      LAYER mcon ;
        RECT 1162.285 51.085 1162.455 51.255 ;
        RECT 690.785 50.745 690.955 50.915 ;
        RECT 740.465 50.745 740.635 50.915 ;
        RECT 691.705 48.025 691.875 48.195 ;
      LAYER met1 ;
        RECT 302.470 51.240 302.790 51.300 ;
        RECT 1128.170 51.240 1128.490 51.300 ;
        RECT 1161.765 51.240 1162.055 51.285 ;
        RECT 302.470 51.100 667.480 51.240 ;
        RECT 302.470 51.040 302.790 51.100 ;
        RECT 667.340 50.900 667.480 51.100 ;
        RECT 1128.170 51.100 1162.055 51.240 ;
        RECT 1128.170 51.040 1128.490 51.100 ;
        RECT 1161.765 51.055 1162.055 51.100 ;
        RECT 1162.210 51.240 1162.530 51.300 ;
        RECT 1162.210 51.100 1162.725 51.240 ;
        RECT 1162.210 51.040 1162.530 51.100 ;
        RECT 690.725 50.900 691.015 50.945 ;
        RECT 667.340 50.760 691.015 50.900 ;
        RECT 690.725 50.715 691.015 50.760 ;
        RECT 740.405 50.900 740.695 50.945 ;
        RECT 787.310 50.900 787.630 50.960 ;
        RECT 740.405 50.760 787.630 50.900 ;
        RECT 740.405 50.715 740.695 50.760 ;
        RECT 787.310 50.700 787.630 50.760 ;
        RECT 839.290 50.900 839.610 50.960 ;
        RECT 979.590 50.900 979.910 50.960 ;
        RECT 839.290 50.760 979.910 50.900 ;
        RECT 839.290 50.700 839.610 50.760 ;
        RECT 979.590 50.700 979.910 50.760 ;
        RECT 1209.590 50.560 1209.910 50.620 ;
        RECT 1211.890 50.560 1212.210 50.620 ;
        RECT 1209.590 50.420 1212.210 50.560 ;
        RECT 1209.590 50.360 1209.910 50.420 ;
        RECT 1211.890 50.360 1212.210 50.420 ;
        RECT 691.645 48.180 691.935 48.225 ;
        RECT 691.645 48.040 693.240 48.180 ;
        RECT 691.645 47.995 691.935 48.040 ;
        RECT 693.100 47.840 693.240 48.040 ;
        RECT 740.405 47.840 740.695 47.885 ;
        RECT 693.100 47.700 740.695 47.840 ;
        RECT 740.405 47.655 740.695 47.700 ;
      LAYER via ;
        RECT 302.500 51.040 302.760 51.300 ;
        RECT 1128.200 51.040 1128.460 51.300 ;
        RECT 1162.240 51.040 1162.500 51.300 ;
        RECT 787.340 50.700 787.600 50.960 ;
        RECT 839.320 50.700 839.580 50.960 ;
        RECT 979.620 50.700 979.880 50.960 ;
        RECT 1209.620 50.360 1209.880 50.620 ;
        RECT 1211.920 50.360 1212.180 50.620 ;
      LAYER met2 ;
        RECT 789.170 51.835 789.450 52.205 ;
        RECT 839.310 51.835 839.590 52.205 ;
        RECT 982.370 51.835 982.650 52.205 ;
        RECT 1031.590 51.835 1031.870 52.205 ;
        RECT 1080.810 51.835 1081.090 52.205 ;
        RECT 1128.190 51.835 1128.470 52.205 ;
        RECT 302.500 51.010 302.760 51.330 ;
        RECT 302.560 2.400 302.700 51.010 ;
        RECT 787.340 50.845 787.600 50.990 ;
        RECT 789.240 50.845 789.380 51.835 ;
        RECT 839.380 50.990 839.520 51.835 ;
        RECT 787.330 50.475 787.610 50.845 ;
        RECT 789.170 50.475 789.450 50.845 ;
        RECT 839.320 50.670 839.580 50.990 ;
        RECT 979.620 50.845 979.880 50.990 ;
        RECT 982.440 50.845 982.580 51.835 ;
        RECT 1031.660 50.845 1031.800 51.835 ;
        RECT 1080.880 50.845 1081.020 51.835 ;
        RECT 1128.260 51.330 1128.400 51.835 ;
        RECT 1128.200 51.010 1128.460 51.330 ;
        RECT 1162.240 51.010 1162.500 51.330 ;
        RECT 979.610 50.475 979.890 50.845 ;
        RECT 982.370 50.475 982.650 50.845 ;
        RECT 1031.590 50.475 1031.870 50.845 ;
        RECT 1080.810 50.475 1081.090 50.845 ;
        RECT 1162.300 50.165 1162.440 51.010 ;
        RECT 1211.980 50.650 1212.120 54.000 ;
        RECT 1209.620 50.330 1209.880 50.650 ;
        RECT 1211.920 50.330 1212.180 50.650 ;
        RECT 1209.680 50.165 1209.820 50.330 ;
        RECT 1162.230 49.795 1162.510 50.165 ;
        RECT 1209.610 49.795 1209.890 50.165 ;
        RECT 302.490 0.000 302.770 2.400 ;
      LAYER via2 ;
        RECT 789.170 51.880 789.450 52.160 ;
        RECT 839.310 51.880 839.590 52.160 ;
        RECT 982.370 51.880 982.650 52.160 ;
        RECT 1031.590 51.880 1031.870 52.160 ;
        RECT 1080.810 51.880 1081.090 52.160 ;
        RECT 1128.190 51.880 1128.470 52.160 ;
        RECT 787.330 50.520 787.610 50.800 ;
        RECT 789.170 50.520 789.450 50.800 ;
        RECT 979.610 50.520 979.890 50.800 ;
        RECT 982.370 50.520 982.650 50.800 ;
        RECT 1031.590 50.520 1031.870 50.800 ;
        RECT 1080.810 50.520 1081.090 50.800 ;
        RECT 1162.230 49.840 1162.510 50.120 ;
        RECT 1209.610 49.840 1209.890 50.120 ;
      LAYER met3 ;
        RECT 789.145 52.170 789.475 52.185 ;
        RECT 839.285 52.170 839.615 52.185 ;
        RECT 789.145 51.870 839.615 52.170 ;
        RECT 789.145 51.855 789.475 51.870 ;
        RECT 839.285 51.855 839.615 51.870 ;
        RECT 982.345 52.170 982.675 52.185 ;
        RECT 1031.565 52.170 1031.895 52.185 ;
        RECT 982.345 51.870 1031.895 52.170 ;
        RECT 982.345 51.855 982.675 51.870 ;
        RECT 1031.565 51.855 1031.895 51.870 ;
        RECT 1080.785 52.170 1081.115 52.185 ;
        RECT 1128.165 52.170 1128.495 52.185 ;
        RECT 1080.785 51.870 1128.495 52.170 ;
        RECT 1080.785 51.855 1081.115 51.870 ;
        RECT 1128.165 51.855 1128.495 51.870 ;
        RECT 787.305 50.810 787.635 50.825 ;
        RECT 789.145 50.810 789.475 50.825 ;
        RECT 787.305 50.510 789.475 50.810 ;
        RECT 787.305 50.495 787.635 50.510 ;
        RECT 789.145 50.495 789.475 50.510 ;
        RECT 979.585 50.810 979.915 50.825 ;
        RECT 982.345 50.810 982.675 50.825 ;
        RECT 979.585 50.510 982.675 50.810 ;
        RECT 979.585 50.495 979.915 50.510 ;
        RECT 982.345 50.495 982.675 50.510 ;
        RECT 1031.565 50.810 1031.895 50.825 ;
        RECT 1080.785 50.810 1081.115 50.825 ;
        RECT 1031.565 50.510 1081.115 50.810 ;
        RECT 1031.565 50.495 1031.895 50.510 ;
        RECT 1080.785 50.495 1081.115 50.510 ;
        RECT 1162.205 50.130 1162.535 50.145 ;
        RECT 1209.585 50.130 1209.915 50.145 ;
        RECT 1162.205 49.830 1209.915 50.130 ;
        RECT 1162.205 49.815 1162.535 49.830 ;
        RECT 1209.585 49.815 1209.915 49.830 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1191.725 53.125 1191.895 54.000 ;
        RECT 692.625 48.025 693.715 48.195 ;
        RECT 739.545 48.025 739.715 50.575 ;
        RECT 692.625 47.685 692.795 48.025 ;
      LAYER mcon ;
        RECT 739.545 50.405 739.715 50.575 ;
        RECT 693.545 48.025 693.715 48.195 ;
      LAYER met1 ;
        RECT 1191.665 53.280 1191.955 53.325 ;
        RECT 1218.790 53.280 1219.110 53.340 ;
        RECT 1191.665 53.140 1219.110 53.280 ;
        RECT 1191.665 53.095 1191.955 53.140 ;
        RECT 1218.790 53.080 1219.110 53.140 ;
        RECT 326.390 50.900 326.710 50.960 ;
        RECT 644.250 50.900 644.570 50.960 ;
        RECT 326.390 50.760 644.570 50.900 ;
        RECT 326.390 50.700 326.710 50.760 ;
        RECT 644.250 50.700 644.570 50.760 ;
        RECT 739.485 50.560 739.775 50.605 ;
        RECT 787.770 50.560 788.090 50.620 ;
        RECT 739.485 50.420 788.090 50.560 ;
        RECT 739.485 50.375 739.775 50.420 ;
        RECT 787.770 50.360 788.090 50.420 ;
        RECT 838.830 50.560 839.150 50.620 ;
        RECT 980.050 50.560 980.370 50.620 ;
        RECT 838.830 50.420 980.370 50.560 ;
        RECT 838.830 50.360 839.150 50.420 ;
        RECT 980.050 50.360 980.370 50.420 ;
        RECT 693.485 48.180 693.775 48.225 ;
        RECT 739.485 48.180 739.775 48.225 ;
        RECT 693.485 48.040 739.775 48.180 ;
        RECT 693.485 47.995 693.775 48.040 ;
        RECT 739.485 47.995 739.775 48.040 ;
        RECT 644.250 47.840 644.570 47.900 ;
        RECT 692.565 47.840 692.855 47.885 ;
        RECT 644.250 47.700 692.855 47.840 ;
        RECT 644.250 47.640 644.570 47.700 ;
        RECT 692.565 47.655 692.855 47.700 ;
        RECT 320.410 16.900 320.730 16.960 ;
        RECT 325.930 16.900 326.250 16.960 ;
        RECT 320.410 16.760 326.250 16.900 ;
        RECT 320.410 16.700 320.730 16.760 ;
        RECT 325.930 16.700 326.250 16.760 ;
      LAYER via ;
        RECT 1218.820 53.080 1219.080 53.340 ;
        RECT 326.420 50.700 326.680 50.960 ;
        RECT 644.280 50.700 644.540 50.960 ;
        RECT 787.800 50.360 788.060 50.620 ;
        RECT 838.860 50.360 839.120 50.620 ;
        RECT 980.080 50.360 980.340 50.620 ;
        RECT 644.280 47.640 644.540 47.900 ;
        RECT 320.440 16.700 320.700 16.960 ;
        RECT 325.960 16.700 326.220 16.960 ;
      LAYER met2 ;
        RECT 326.420 50.670 326.680 50.990 ;
        RECT 644.280 50.670 644.540 50.990 ;
        RECT 326.480 17.410 326.620 50.670 ;
        RECT 644.340 47.930 644.480 50.670 ;
        RECT 787.800 50.330 788.060 50.650 ;
        RECT 838.850 50.475 839.130 50.845 ;
        RECT 838.860 50.330 839.120 50.475 ;
        RECT 980.080 50.330 980.340 50.650 ;
        RECT 787.860 50.165 788.000 50.330 ;
        RECT 980.140 50.165 980.280 50.330 ;
        RECT 787.790 49.795 788.070 50.165 ;
        RECT 980.070 49.795 980.350 50.165 ;
        RECT 1079.960 49.485 1080.100 54.000 ;
        RECT 1218.880 53.370 1219.020 54.000 ;
        RECT 1218.820 53.050 1219.080 53.370 ;
        RECT 1079.890 49.115 1080.170 49.485 ;
        RECT 644.280 47.610 644.540 47.930 ;
        RECT 326.020 17.270 326.620 17.410 ;
        RECT 326.020 16.990 326.160 17.270 ;
        RECT 320.440 16.670 320.700 16.990 ;
        RECT 325.960 16.670 326.220 16.990 ;
        RECT 320.500 2.400 320.640 16.670 ;
        RECT 320.430 0.000 320.710 2.400 ;
      LAYER via2 ;
        RECT 838.850 50.520 839.130 50.800 ;
        RECT 787.790 49.840 788.070 50.120 ;
        RECT 980.070 49.840 980.350 50.120 ;
        RECT 1079.890 49.160 1080.170 49.440 ;
      LAYER met3 ;
        RECT 838.825 50.810 839.155 50.825 ;
        RECT 791.230 50.510 839.155 50.810 ;
        RECT 787.765 50.130 788.095 50.145 ;
        RECT 791.230 50.130 791.530 50.510 ;
        RECT 838.825 50.495 839.155 50.510 ;
        RECT 983.510 50.510 1030.730 50.810 ;
        RECT 787.765 49.830 791.530 50.130 ;
        RECT 980.045 50.130 980.375 50.145 ;
        RECT 983.510 50.130 983.810 50.510 ;
        RECT 980.045 49.830 983.810 50.130 ;
        RECT 787.765 49.815 788.095 49.830 ;
        RECT 980.045 49.815 980.375 49.830 ;
        RECT 1030.430 49.450 1030.730 50.510 ;
        RECT 1079.865 49.450 1080.195 49.465 ;
        RECT 1030.430 49.150 1080.195 49.450 ;
        RECT 1079.865 49.135 1080.195 49.150 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 740.005 48.025 740.175 50.915 ;
        RECT 741.385 44.285 741.555 48.195 ;
        RECT 789.225 44.285 789.395 54.000 ;
        RECT 982.885 44.965 983.055 54.000 ;
      LAYER mcon ;
        RECT 740.005 50.745 740.175 50.915 ;
        RECT 741.385 48.025 741.555 48.195 ;
      LAYER met1 ;
        RECT 1192.570 53.960 1192.890 54.000 ;
        RECT 1220.630 53.960 1220.950 54.000 ;
        RECT 1192.570 53.820 1220.950 53.960 ;
        RECT 1192.570 53.760 1192.890 53.820 ;
        RECT 1220.630 53.760 1220.950 53.820 ;
        RECT 693.010 50.900 693.330 50.960 ;
        RECT 739.945 50.900 740.235 50.945 ;
        RECT 693.010 50.760 740.235 50.900 ;
        RECT 693.010 50.700 693.330 50.760 ;
        RECT 739.945 50.715 740.235 50.760 ;
        RECT 340.190 50.560 340.510 50.620 ;
        RECT 691.170 50.560 691.490 50.620 ;
        RECT 340.190 50.420 691.490 50.560 ;
        RECT 340.190 50.360 340.510 50.420 ;
        RECT 691.170 50.360 691.490 50.420 ;
        RECT 1128.170 50.560 1128.490 50.620 ;
        RECT 1175.090 50.560 1175.410 50.620 ;
        RECT 1128.170 50.420 1175.410 50.560 ;
        RECT 1128.170 50.360 1128.490 50.420 ;
        RECT 1175.090 50.360 1175.410 50.420 ;
        RECT 739.945 48.180 740.235 48.225 ;
        RECT 741.325 48.180 741.615 48.225 ;
        RECT 739.945 48.040 741.615 48.180 ;
        RECT 739.945 47.995 740.235 48.040 ;
        RECT 741.325 47.995 741.615 48.040 ;
        RECT 958.890 45.120 959.210 45.180 ;
        RECT 982.825 45.120 983.115 45.165 ;
        RECT 958.890 44.980 983.115 45.120 ;
        RECT 958.890 44.920 959.210 44.980 ;
        RECT 982.825 44.935 983.115 44.980 ;
        RECT 741.325 44.440 741.615 44.485 ;
        RECT 789.165 44.440 789.455 44.485 ;
        RECT 741.325 44.300 789.455 44.440 ;
        RECT 741.325 44.255 741.615 44.300 ;
        RECT 789.165 44.255 789.455 44.300 ;
      LAYER via ;
        RECT 1192.600 53.760 1192.860 54.000 ;
        RECT 1220.660 53.760 1220.920 54.000 ;
        RECT 693.040 50.700 693.300 50.960 ;
        RECT 340.220 50.360 340.480 50.620 ;
        RECT 691.200 50.360 691.460 50.620 ;
        RECT 1128.200 50.360 1128.460 50.620 ;
        RECT 1175.120 50.360 1175.380 50.620 ;
        RECT 958.920 44.920 959.180 45.180 ;
      LAYER met2 ;
        RECT 693.040 50.845 693.300 50.990 ;
        RECT 340.220 50.330 340.480 50.650 ;
        RECT 691.190 50.475 691.470 50.845 ;
        RECT 693.030 50.475 693.310 50.845 ;
        RECT 691.200 50.330 691.460 50.475 ;
        RECT 340.280 3.130 340.420 50.330 ;
        RECT 837.540 50.165 837.680 54.000 ;
        RECT 958.910 50.475 959.190 50.845 ;
        RECT 837.470 49.795 837.750 50.165 ;
        RECT 958.980 45.210 959.120 50.475 ;
        RECT 1079.040 50.165 1079.180 54.000 ;
        RECT 1192.600 53.730 1192.860 54.000 ;
        RECT 1220.660 53.730 1220.920 54.000 ;
        RECT 1192.660 50.845 1192.800 53.730 ;
        RECT 1128.200 50.330 1128.460 50.650 ;
        RECT 1175.110 50.475 1175.390 50.845 ;
        RECT 1192.590 50.475 1192.870 50.845 ;
        RECT 1175.120 50.330 1175.380 50.475 ;
        RECT 1128.260 50.165 1128.400 50.330 ;
        RECT 1078.970 49.795 1079.250 50.165 ;
        RECT 1128.190 49.795 1128.470 50.165 ;
        RECT 958.920 44.890 959.180 45.210 ;
        RECT 338.440 2.990 340.420 3.130 ;
        RECT 338.440 2.400 338.580 2.990 ;
        RECT 338.370 0.000 338.650 2.400 ;
      LAYER via2 ;
        RECT 691.190 50.520 691.470 50.800 ;
        RECT 693.030 50.520 693.310 50.800 ;
        RECT 958.910 50.520 959.190 50.800 ;
        RECT 837.470 49.840 837.750 50.120 ;
        RECT 1175.110 50.520 1175.390 50.800 ;
        RECT 1192.590 50.520 1192.870 50.800 ;
        RECT 1078.970 49.840 1079.250 50.120 ;
        RECT 1128.190 49.840 1128.470 50.120 ;
      LAYER met3 ;
        RECT 691.165 50.810 691.495 50.825 ;
        RECT 693.005 50.810 693.335 50.825 ;
        RECT 691.165 50.510 693.335 50.810 ;
        RECT 691.165 50.495 691.495 50.510 ;
        RECT 693.005 50.495 693.335 50.510 ;
        RECT 885.950 50.810 886.330 50.820 ;
        RECT 958.885 50.810 959.215 50.825 ;
        RECT 885.950 50.510 959.215 50.810 ;
        RECT 885.950 50.500 886.330 50.510 ;
        RECT 958.885 50.495 959.215 50.510 ;
        RECT 1175.085 50.810 1175.415 50.825 ;
        RECT 1192.565 50.810 1192.895 50.825 ;
        RECT 1175.085 50.510 1192.895 50.810 ;
        RECT 1175.085 50.495 1175.415 50.510 ;
        RECT 1192.565 50.495 1192.895 50.510 ;
        RECT 837.445 50.130 837.775 50.145 ;
        RECT 885.030 50.130 885.410 50.140 ;
        RECT 837.445 49.830 885.410 50.130 ;
        RECT 837.445 49.815 837.775 49.830 ;
        RECT 885.030 49.820 885.410 49.830 ;
        RECT 1078.945 50.130 1079.275 50.145 ;
        RECT 1128.165 50.130 1128.495 50.145 ;
        RECT 1078.945 49.830 1128.495 50.130 ;
        RECT 1078.945 49.815 1079.275 49.830 ;
        RECT 1128.165 49.815 1128.495 49.830 ;
      LAYER via3 ;
        RECT 885.980 50.500 886.300 50.820 ;
        RECT 885.060 49.820 885.380 50.140 ;
      LAYER met4 ;
        RECT 885.975 50.495 886.305 50.825 ;
        RECT 885.055 49.815 885.385 50.145 ;
        RECT 885.070 49.450 885.370 49.815 ;
        RECT 885.990 49.450 886.290 50.495 ;
        RECT 885.070 49.150 886.290 49.450 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 355.830 15.880 356.150 15.940 ;
        RECT 360.890 15.880 361.210 15.940 ;
        RECT 355.830 15.740 361.210 15.880 ;
        RECT 355.830 15.680 356.150 15.740 ;
        RECT 360.890 15.680 361.210 15.740 ;
      LAYER via ;
        RECT 355.860 15.680 356.120 15.940 ;
        RECT 360.920 15.680 361.180 15.940 ;
      LAYER met2 ;
        RECT 360.980 15.970 361.120 54.000 ;
        RECT 355.860 15.650 356.120 15.970 ;
        RECT 360.920 15.650 361.180 15.970 ;
        RECT 355.920 2.400 356.060 15.650 ;
        RECT 355.850 0.000 356.130 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 373.770 2.960 374.090 3.020 ;
        RECT 374.690 2.960 375.010 3.020 ;
        RECT 373.770 2.820 375.010 2.960 ;
        RECT 373.770 2.760 374.090 2.820 ;
        RECT 374.690 2.760 375.010 2.820 ;
      LAYER via ;
        RECT 373.800 2.760 374.060 3.020 ;
        RECT 374.720 2.760 374.980 3.020 ;
      LAYER met2 ;
        RECT 374.780 3.050 374.920 54.000 ;
        RECT 373.800 2.730 374.060 3.050 ;
        RECT 374.720 2.730 374.980 3.050 ;
        RECT 373.860 2.400 374.000 2.730 ;
        RECT 373.790 0.000 374.070 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 391.710 15.540 392.030 15.600 ;
        RECT 395.390 15.540 395.710 15.600 ;
        RECT 391.710 15.400 395.710 15.540 ;
        RECT 391.710 15.340 392.030 15.400 ;
        RECT 395.390 15.340 395.710 15.400 ;
      LAYER via ;
        RECT 391.740 15.340 392.000 15.600 ;
        RECT 395.420 15.340 395.680 15.600 ;
      LAYER met2 ;
        RECT 395.480 15.630 395.620 54.000 ;
        RECT 391.740 15.310 392.000 15.630 ;
        RECT 395.420 15.310 395.680 15.630 ;
        RECT 391.800 2.400 391.940 15.310 ;
        RECT 391.730 0.000 392.010 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 409.650 17.580 409.970 17.640 ;
        RECT 415.170 17.580 415.490 17.640 ;
        RECT 409.650 17.440 415.490 17.580 ;
        RECT 409.650 17.380 409.970 17.440 ;
        RECT 415.170 17.380 415.490 17.440 ;
      LAYER via ;
        RECT 409.680 17.380 409.940 17.640 ;
        RECT 415.200 17.380 415.460 17.640 ;
      LAYER met2 ;
        RECT 415.720 18.090 415.860 54.000 ;
        RECT 415.260 17.950 415.860 18.090 ;
        RECT 415.260 17.670 415.400 17.950 ;
        RECT 409.680 17.350 409.940 17.670 ;
        RECT 415.200 17.350 415.460 17.670 ;
        RECT 409.740 2.400 409.880 17.350 ;
        RECT 409.670 0.000 409.950 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.180 3.130 71.320 54.000 ;
        RECT 70.720 2.990 71.320 3.130 ;
        RECT 70.720 2.400 70.860 2.990 ;
        RECT 70.650 0.000 70.930 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 427.130 15.200 427.450 15.260 ;
        RECT 429.890 15.200 430.210 15.260 ;
        RECT 427.130 15.060 430.210 15.200 ;
        RECT 427.130 15.000 427.450 15.060 ;
        RECT 429.890 15.000 430.210 15.060 ;
      LAYER via ;
        RECT 427.160 15.000 427.420 15.260 ;
        RECT 429.920 15.000 430.180 15.260 ;
      LAYER met2 ;
        RECT 429.980 15.290 430.120 54.000 ;
        RECT 427.160 14.970 427.420 15.290 ;
        RECT 429.920 14.970 430.180 15.290 ;
        RECT 427.220 2.400 427.360 14.970 ;
        RECT 427.150 0.000 427.430 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 445.070 15.200 445.390 15.260 ;
        RECT 450.590 15.200 450.910 15.260 ;
        RECT 445.070 15.060 450.910 15.200 ;
        RECT 445.070 15.000 445.390 15.060 ;
        RECT 450.590 15.000 450.910 15.060 ;
      LAYER via ;
        RECT 445.100 15.000 445.360 15.260 ;
        RECT 450.620 15.000 450.880 15.260 ;
      LAYER met2 ;
        RECT 450.680 15.290 450.820 54.000 ;
        RECT 445.100 14.970 445.360 15.290 ;
        RECT 450.620 14.970 450.880 15.290 ;
        RECT 445.160 2.400 445.300 14.970 ;
        RECT 445.090 0.000 445.370 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 463.100 2.400 463.240 54.000 ;
        RECT 463.030 0.000 463.310 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 480.950 17.580 481.270 17.640 ;
        RECT 485.090 17.580 485.410 17.640 ;
        RECT 480.950 17.440 485.410 17.580 ;
        RECT 480.950 17.380 481.270 17.440 ;
        RECT 485.090 17.380 485.410 17.440 ;
      LAYER via ;
        RECT 480.980 17.380 481.240 17.640 ;
        RECT 485.120 17.380 485.380 17.640 ;
      LAYER met2 ;
        RECT 485.180 17.670 485.320 54.000 ;
        RECT 480.980 17.350 481.240 17.670 ;
        RECT 485.120 17.350 485.380 17.670 ;
        RECT 481.040 2.400 481.180 17.350 ;
        RECT 480.970 0.000 481.250 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 497.510 15.200 497.830 15.260 ;
        RECT 498.890 15.200 499.210 15.260 ;
        RECT 497.510 15.060 499.210 15.200 ;
        RECT 497.510 15.000 497.830 15.060 ;
        RECT 498.890 15.000 499.210 15.060 ;
      LAYER via ;
        RECT 497.540 15.000 497.800 15.260 ;
        RECT 498.920 15.000 499.180 15.260 ;
      LAYER met2 ;
        RECT 497.600 15.290 497.740 54.000 ;
        RECT 497.540 14.970 497.800 15.290 ;
        RECT 498.920 14.970 499.180 15.290 ;
        RECT 498.980 2.400 499.120 14.970 ;
        RECT 498.910 0.000 499.190 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 516.370 14.520 516.690 14.580 ;
        RECT 519.590 14.520 519.910 14.580 ;
        RECT 516.370 14.380 519.910 14.520 ;
        RECT 516.370 14.320 516.690 14.380 ;
        RECT 519.590 14.320 519.910 14.380 ;
      LAYER via ;
        RECT 516.400 14.320 516.660 14.580 ;
        RECT 519.620 14.320 519.880 14.580 ;
      LAYER met2 ;
        RECT 519.680 14.610 519.820 54.000 ;
        RECT 516.400 14.290 516.660 14.610 ;
        RECT 519.620 14.290 519.880 14.610 ;
        RECT 516.460 2.400 516.600 14.290 ;
        RECT 516.390 0.000 516.670 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 534.310 14.860 534.630 14.920 ;
        RECT 539.830 14.860 540.150 14.920 ;
        RECT 534.310 14.720 540.150 14.860 ;
        RECT 534.310 14.660 534.630 14.720 ;
        RECT 539.830 14.660 540.150 14.720 ;
      LAYER via ;
        RECT 534.340 14.660 534.600 14.920 ;
        RECT 539.860 14.660 540.120 14.920 ;
      LAYER met2 ;
        RECT 539.920 14.950 540.060 54.000 ;
        RECT 534.340 14.630 534.600 14.950 ;
        RECT 539.860 14.630 540.120 14.950 ;
        RECT 534.400 2.400 534.540 14.630 ;
        RECT 534.330 0.000 534.610 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 554.180 17.410 554.320 54.000 ;
        RECT 552.340 17.270 554.320 17.410 ;
        RECT 552.340 2.400 552.480 17.270 ;
        RECT 552.270 0.000 552.550 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 570.190 17.580 570.510 17.640 ;
        RECT 574.790 17.580 575.110 17.640 ;
        RECT 570.190 17.440 575.110 17.580 ;
        RECT 570.190 17.380 570.510 17.440 ;
        RECT 574.790 17.380 575.110 17.440 ;
      LAYER via ;
        RECT 570.220 17.380 570.480 17.640 ;
        RECT 574.820 17.380 575.080 17.640 ;
      LAYER met2 ;
        RECT 574.880 17.670 575.020 54.000 ;
        RECT 570.220 17.350 570.480 17.670 ;
        RECT 574.820 17.350 575.080 17.670 ;
        RECT 570.280 2.400 570.420 17.350 ;
        RECT 570.210 0.000 570.490 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 588.680 17.410 588.820 54.000 ;
        RECT 588.220 17.270 588.820 17.410 ;
        RECT 588.220 2.400 588.360 17.270 ;
        RECT 588.150 0.000 588.430 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 94.090 17.580 94.410 17.640 ;
        RECT 98.690 17.580 99.010 17.640 ;
        RECT 94.090 17.440 99.010 17.580 ;
        RECT 94.090 17.380 94.410 17.440 ;
        RECT 98.690 17.380 99.010 17.440 ;
      LAYER via ;
        RECT 94.120 17.380 94.380 17.640 ;
        RECT 98.720 17.380 98.980 17.640 ;
      LAYER met2 ;
        RECT 98.780 17.670 98.920 54.000 ;
        RECT 94.120 17.350 94.380 17.670 ;
        RECT 98.720 17.350 98.980 17.670 ;
        RECT 94.180 2.400 94.320 17.350 ;
        RECT 94.110 0.000 94.390 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 605.610 17.580 605.930 17.640 ;
        RECT 609.290 17.580 609.610 17.640 ;
        RECT 605.610 17.440 609.610 17.580 ;
        RECT 605.610 17.380 605.930 17.440 ;
        RECT 609.290 17.380 609.610 17.440 ;
      LAYER via ;
        RECT 605.640 17.380 605.900 17.640 ;
        RECT 609.320 17.380 609.580 17.640 ;
      LAYER met2 ;
        RECT 609.380 17.670 609.520 54.000 ;
        RECT 605.640 17.350 605.900 17.670 ;
        RECT 609.320 17.350 609.580 17.670 ;
        RECT 605.700 2.400 605.840 17.350 ;
        RECT 605.630 0.000 605.910 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 623.550 17.580 623.870 17.640 ;
        RECT 629.070 17.580 629.390 17.640 ;
        RECT 623.550 17.440 629.390 17.580 ;
        RECT 623.550 17.380 623.870 17.440 ;
        RECT 629.070 17.380 629.390 17.440 ;
      LAYER via ;
        RECT 623.580 17.380 623.840 17.640 ;
        RECT 629.100 17.380 629.360 17.640 ;
      LAYER met2 ;
        RECT 629.620 18.090 629.760 54.000 ;
        RECT 629.160 17.950 629.760 18.090 ;
        RECT 629.160 17.670 629.300 17.950 ;
        RECT 623.580 17.350 623.840 17.670 ;
        RECT 629.100 17.350 629.360 17.670 ;
        RECT 623.640 2.400 623.780 17.350 ;
        RECT 623.570 0.000 623.850 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 118.010 2.960 118.330 3.020 ;
        RECT 119.390 2.960 119.710 3.020 ;
        RECT 118.010 2.820 119.710 2.960 ;
        RECT 118.010 2.760 118.330 2.820 ;
        RECT 119.390 2.760 119.710 2.820 ;
      LAYER via ;
        RECT 118.040 2.760 118.300 3.020 ;
        RECT 119.420 2.760 119.680 3.020 ;
      LAYER met2 ;
        RECT 119.480 3.050 119.620 54.000 ;
        RECT 118.040 2.730 118.300 3.050 ;
        RECT 119.420 2.730 119.680 3.050 ;
        RECT 118.100 2.400 118.240 2.730 ;
        RECT 118.030 0.000 118.310 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 141.930 15.880 142.250 15.940 ;
        RECT 146.990 15.880 147.310 15.940 ;
        RECT 141.930 15.740 147.310 15.880 ;
        RECT 141.930 15.680 142.250 15.740 ;
        RECT 146.990 15.680 147.310 15.740 ;
      LAYER via ;
        RECT 141.960 15.680 142.220 15.940 ;
        RECT 147.020 15.680 147.280 15.940 ;
      LAYER met2 ;
        RECT 147.080 15.970 147.220 54.000 ;
        RECT 141.960 15.650 142.220 15.970 ;
        RECT 147.020 15.650 147.280 15.970 ;
        RECT 142.020 2.400 142.160 15.650 ;
        RECT 141.950 0.000 142.230 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1184.840 20.245 1184.980 54.000 ;
        RECT 159.890 19.875 160.170 20.245 ;
        RECT 1184.770 19.875 1185.050 20.245 ;
        RECT 159.960 2.400 160.100 19.875 ;
        RECT 159.890 0.000 160.170 2.400 ;
      LAYER via2 ;
        RECT 159.890 19.920 160.170 20.200 ;
        RECT 1184.770 19.920 1185.050 20.200 ;
      LAYER met3 ;
        RECT 159.865 20.210 160.195 20.225 ;
        RECT 1184.745 20.210 1185.075 20.225 ;
        RECT 159.865 19.910 1185.075 20.210 ;
        RECT 159.865 19.895 160.195 19.910 ;
        RECT 1184.745 19.895 1185.075 19.910 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 739.545 21.165 740.635 21.335 ;
        RECT 739.545 20.825 739.715 21.165 ;
        RECT 182.025 15.725 182.195 17.595 ;
        RECT 229.865 15.725 230.035 17.595 ;
        RECT 281.385 15.725 281.555 17.595 ;
        RECT 326.465 15.725 326.635 17.595 ;
        RECT 375.225 14.705 375.395 17.595 ;
        RECT 423.065 14.705 423.235 17.595 ;
        RECT 468.605 14.365 468.775 17.595 ;
        RECT 519.665 14.875 519.835 17.595 ;
        RECT 740.465 17.425 740.635 21.165 ;
        RECT 519.205 14.705 519.835 14.875 ;
      LAYER mcon ;
        RECT 182.025 17.425 182.195 17.595 ;
        RECT 229.865 17.425 230.035 17.595 ;
        RECT 281.385 17.425 281.555 17.595 ;
        RECT 326.465 17.425 326.635 17.595 ;
        RECT 375.225 17.425 375.395 17.595 ;
        RECT 423.065 17.425 423.235 17.595 ;
        RECT 468.605 17.425 468.775 17.595 ;
        RECT 519.665 17.425 519.835 17.595 ;
      LAYER met1 ;
        RECT 644.250 21.320 644.570 21.380 ;
        RECT 644.250 21.180 672.080 21.320 ;
        RECT 644.250 21.120 644.570 21.180 ;
        RECT 671.940 20.980 672.080 21.180 ;
        RECT 739.485 20.980 739.775 21.025 ;
        RECT 671.940 20.840 739.775 20.980 ;
        RECT 739.485 20.795 739.775 20.840 ;
        RECT 177.350 17.580 177.670 17.640 ;
        RECT 181.965 17.580 182.255 17.625 ;
        RECT 177.350 17.440 182.255 17.580 ;
        RECT 177.350 17.380 177.670 17.440 ;
        RECT 181.965 17.395 182.255 17.440 ;
        RECT 229.805 17.580 230.095 17.625 ;
        RECT 281.325 17.580 281.615 17.625 ;
        RECT 229.805 17.440 281.615 17.580 ;
        RECT 229.805 17.395 230.095 17.440 ;
        RECT 281.325 17.395 281.615 17.440 ;
        RECT 326.405 17.580 326.695 17.625 ;
        RECT 375.165 17.580 375.455 17.625 ;
        RECT 326.405 17.440 375.455 17.580 ;
        RECT 326.405 17.395 326.695 17.440 ;
        RECT 375.165 17.395 375.455 17.440 ;
        RECT 423.005 17.580 423.295 17.625 ;
        RECT 468.545 17.580 468.835 17.625 ;
        RECT 423.005 17.440 468.835 17.580 ;
        RECT 423.005 17.395 423.295 17.440 ;
        RECT 468.545 17.395 468.835 17.440 ;
        RECT 519.605 17.580 519.895 17.625 ;
        RECT 740.405 17.580 740.695 17.625 ;
        RECT 788.230 17.580 788.550 17.640 ;
        RECT 519.605 17.440 569.960 17.580 ;
        RECT 519.605 17.395 519.895 17.440 ;
        RECT 569.820 17.240 569.960 17.440 ;
        RECT 740.405 17.440 788.550 17.580 ;
        RECT 740.405 17.395 740.695 17.440 ;
        RECT 788.230 17.380 788.550 17.440 ;
        RECT 1031.110 17.580 1031.430 17.640 ;
        RECT 1183.370 17.580 1183.690 17.640 ;
        RECT 1031.110 17.440 1183.690 17.580 ;
        RECT 1031.110 17.380 1031.430 17.440 ;
        RECT 1183.370 17.380 1183.690 17.440 ;
        RECT 644.250 17.240 644.570 17.300 ;
        RECT 569.820 17.100 644.570 17.240 ;
        RECT 644.250 17.040 644.570 17.100 ;
        RECT 790.530 17.240 790.850 17.300 ;
        RECT 932.670 17.240 932.990 17.300 ;
        RECT 790.530 17.100 932.990 17.240 ;
        RECT 790.530 17.040 790.850 17.100 ;
        RECT 932.670 17.040 932.990 17.100 ;
        RECT 181.965 15.880 182.255 15.925 ;
        RECT 229.805 15.880 230.095 15.925 ;
        RECT 181.965 15.740 230.095 15.880 ;
        RECT 181.965 15.695 182.255 15.740 ;
        RECT 229.805 15.695 230.095 15.740 ;
        RECT 281.325 15.880 281.615 15.925 ;
        RECT 326.405 15.880 326.695 15.925 ;
        RECT 281.325 15.740 326.695 15.880 ;
        RECT 281.325 15.695 281.615 15.740 ;
        RECT 326.405 15.695 326.695 15.740 ;
        RECT 935.890 15.880 936.210 15.940 ;
        RECT 980.970 15.880 981.290 15.940 ;
        RECT 935.890 15.740 981.290 15.880 ;
        RECT 935.890 15.680 936.210 15.740 ;
        RECT 980.970 15.680 981.290 15.740 ;
        RECT 983.730 15.880 984.050 15.940 ;
        RECT 1029.270 15.880 1029.590 15.940 ;
        RECT 983.730 15.740 1029.590 15.880 ;
        RECT 983.730 15.680 984.050 15.740 ;
        RECT 1029.270 15.680 1029.590 15.740 ;
        RECT 375.165 14.860 375.455 14.905 ;
        RECT 423.005 14.860 423.295 14.905 ;
        RECT 519.145 14.860 519.435 14.905 ;
        RECT 375.165 14.720 423.295 14.860 ;
        RECT 375.165 14.675 375.455 14.720 ;
        RECT 423.005 14.675 423.295 14.720 ;
        RECT 513.700 14.720 519.435 14.860 ;
        RECT 468.545 14.520 468.835 14.565 ;
        RECT 513.700 14.520 513.840 14.720 ;
        RECT 519.145 14.675 519.435 14.720 ;
        RECT 468.545 14.380 513.840 14.520 ;
        RECT 468.545 14.335 468.835 14.380 ;
      LAYER via ;
        RECT 644.280 21.120 644.540 21.380 ;
        RECT 177.380 17.380 177.640 17.640 ;
        RECT 788.260 17.380 788.520 17.640 ;
        RECT 1031.140 17.380 1031.400 17.640 ;
        RECT 1183.400 17.380 1183.660 17.640 ;
        RECT 644.280 17.040 644.540 17.300 ;
        RECT 790.560 17.040 790.820 17.300 ;
        RECT 932.700 17.040 932.960 17.300 ;
        RECT 935.920 15.680 936.180 15.940 ;
        RECT 981.000 15.680 981.260 15.940 ;
        RECT 983.760 15.680 984.020 15.940 ;
        RECT 1029.300 15.680 1029.560 15.940 ;
      LAYER met2 ;
        RECT 644.280 21.090 644.540 21.410 ;
        RECT 177.380 17.350 177.640 17.670 ;
        RECT 177.440 2.400 177.580 17.350 ;
        RECT 644.340 17.330 644.480 21.090 ;
        RECT 1183.460 17.670 1183.600 54.000 ;
        RECT 788.260 17.350 788.520 17.670 ;
        RECT 1031.140 17.350 1031.400 17.670 ;
        RECT 1183.400 17.350 1183.660 17.670 ;
        RECT 644.280 17.010 644.540 17.330 ;
        RECT 788.320 16.165 788.460 17.350 ;
        RECT 790.560 17.010 790.820 17.330 ;
        RECT 932.700 17.010 932.960 17.330 ;
        RECT 790.620 16.165 790.760 17.010 ;
        RECT 932.760 16.165 932.900 17.010 ;
        RECT 1031.200 16.165 1031.340 17.350 ;
        RECT 788.250 15.795 788.530 16.165 ;
        RECT 790.550 15.795 790.830 16.165 ;
        RECT 932.690 15.795 932.970 16.165 ;
        RECT 935.910 15.795 936.190 16.165 ;
        RECT 980.990 15.795 981.270 16.165 ;
        RECT 983.750 15.795 984.030 16.165 ;
        RECT 1029.290 15.795 1029.570 16.165 ;
        RECT 1031.130 15.795 1031.410 16.165 ;
        RECT 935.920 15.650 936.180 15.795 ;
        RECT 981.000 15.650 981.260 15.795 ;
        RECT 983.760 15.650 984.020 15.795 ;
        RECT 1029.300 15.650 1029.560 15.795 ;
        RECT 177.370 0.000 177.650 2.400 ;
      LAYER via2 ;
        RECT 788.250 15.840 788.530 16.120 ;
        RECT 790.550 15.840 790.830 16.120 ;
        RECT 932.690 15.840 932.970 16.120 ;
        RECT 935.910 15.840 936.190 16.120 ;
        RECT 980.990 15.840 981.270 16.120 ;
        RECT 983.750 15.840 984.030 16.120 ;
        RECT 1029.290 15.840 1029.570 16.120 ;
        RECT 1031.130 15.840 1031.410 16.120 ;
      LAYER met3 ;
        RECT 788.225 16.130 788.555 16.145 ;
        RECT 790.525 16.130 790.855 16.145 ;
        RECT 788.225 15.830 790.855 16.130 ;
        RECT 788.225 15.815 788.555 15.830 ;
        RECT 790.525 15.815 790.855 15.830 ;
        RECT 932.665 16.130 932.995 16.145 ;
        RECT 935.885 16.130 936.215 16.145 ;
        RECT 932.665 15.830 936.215 16.130 ;
        RECT 932.665 15.815 932.995 15.830 ;
        RECT 935.885 15.815 936.215 15.830 ;
        RECT 980.965 16.130 981.295 16.145 ;
        RECT 983.725 16.130 984.055 16.145 ;
        RECT 980.965 15.830 984.055 16.130 ;
        RECT 980.965 15.815 981.295 15.830 ;
        RECT 983.725 15.815 984.055 15.830 ;
        RECT 1029.265 16.130 1029.595 16.145 ;
        RECT 1031.105 16.130 1031.435 16.145 ;
        RECT 1029.265 15.830 1031.435 16.130 ;
        RECT 1029.265 15.815 1029.595 15.830 ;
        RECT 1031.105 15.815 1031.435 15.830 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 906.065 17.765 907.615 17.935 ;
      LAYER mcon ;
        RECT 907.445 17.765 907.615 17.935 ;
      LAYER met1 ;
        RECT 194.830 18.260 195.150 18.320 ;
        RECT 1174.170 18.260 1174.490 18.320 ;
        RECT 194.830 18.120 223.580 18.260 ;
        RECT 194.830 18.060 195.150 18.120 ;
        RECT 223.440 17.920 223.580 18.120 ;
        RECT 1127.800 18.120 1174.490 18.260 ;
        RECT 906.005 17.920 906.295 17.965 ;
        RECT 223.440 17.780 906.295 17.920 ;
        RECT 906.005 17.735 906.295 17.780 ;
        RECT 907.385 17.920 907.675 17.965 ;
        RECT 1127.800 17.920 1127.940 18.120 ;
        RECT 1174.170 18.060 1174.490 18.120 ;
        RECT 907.385 17.780 1127.940 17.920 ;
        RECT 1176.930 17.920 1177.250 17.980 ;
        RECT 1192.110 17.920 1192.430 17.980 ;
        RECT 1176.930 17.780 1192.430 17.920 ;
        RECT 907.385 17.735 907.675 17.780 ;
        RECT 1176.930 17.720 1177.250 17.780 ;
        RECT 1192.110 17.720 1192.430 17.780 ;
      LAYER via ;
        RECT 194.860 18.060 195.120 18.320 ;
        RECT 1174.200 18.060 1174.460 18.320 ;
        RECT 1176.960 17.720 1177.220 17.980 ;
        RECT 1192.140 17.720 1192.400 17.980 ;
      LAYER met2 ;
        RECT 1191.740 53.960 1191.880 54.000 ;
        RECT 1191.740 53.820 1192.340 53.960 ;
        RECT 194.860 18.030 195.120 18.350 ;
        RECT 1174.200 18.030 1174.460 18.350 ;
        RECT 194.920 9.250 195.060 18.030 ;
        RECT 1174.260 16.845 1174.400 18.030 ;
        RECT 1192.200 18.010 1192.340 53.820 ;
        RECT 1176.960 17.690 1177.220 18.010 ;
        RECT 1192.140 17.690 1192.400 18.010 ;
        RECT 1177.020 16.845 1177.160 17.690 ;
        RECT 1174.190 16.475 1174.470 16.845 ;
        RECT 1176.950 16.475 1177.230 16.845 ;
        RECT 194.920 9.110 195.520 9.250 ;
        RECT 195.380 2.400 195.520 9.110 ;
        RECT 195.310 0.000 195.590 2.400 ;
      LAYER via2 ;
        RECT 1174.190 16.520 1174.470 16.800 ;
        RECT 1176.950 16.520 1177.230 16.800 ;
      LAYER met3 ;
        RECT 1174.165 16.810 1174.495 16.825 ;
        RECT 1176.925 16.810 1177.255 16.825 ;
        RECT 1174.165 16.510 1177.255 16.810 ;
        RECT 1174.165 16.495 1174.495 16.510 ;
        RECT 1176.925 16.495 1177.255 16.510 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1151.705 18.445 1151.875 19.975 ;
        RECT 1164.585 19.805 1164.755 39.355 ;
      LAYER mcon ;
        RECT 1164.585 39.185 1164.755 39.355 ;
        RECT 1151.705 19.805 1151.875 19.975 ;
      LAYER met1 ;
        RECT 1164.525 39.340 1164.815 39.385 ;
        RECT 1189.350 39.340 1189.670 39.400 ;
        RECT 1164.525 39.200 1189.670 39.340 ;
        RECT 1164.525 39.155 1164.815 39.200 ;
        RECT 1189.350 39.140 1189.670 39.200 ;
        RECT 1151.645 19.960 1151.935 20.005 ;
        RECT 1164.525 19.960 1164.815 20.005 ;
        RECT 1151.645 19.820 1164.815 19.960 ;
        RECT 1151.645 19.775 1151.935 19.820 ;
        RECT 1164.525 19.775 1164.815 19.820 ;
        RECT 213.230 18.600 213.550 18.660 ;
        RECT 1151.645 18.600 1151.935 18.645 ;
        RECT 213.230 18.460 1151.935 18.600 ;
        RECT 213.230 18.400 213.550 18.460 ;
        RECT 1151.645 18.415 1151.935 18.460 ;
      LAYER via ;
        RECT 1189.380 39.140 1189.640 39.400 ;
        RECT 213.260 18.400 213.520 18.660 ;
      LAYER met2 ;
        RECT 1189.440 39.430 1189.580 54.000 ;
        RECT 1189.380 39.110 1189.640 39.430 ;
        RECT 213.260 18.370 213.520 18.690 ;
        RECT 213.320 2.400 213.460 18.370 ;
        RECT 213.250 0.000 213.530 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1174.705 19.465 1175.335 19.635 ;
        RECT 1175.165 17.765 1175.335 19.465 ;
        RECT 1176.545 17.765 1176.715 18.615 ;
      LAYER mcon ;
        RECT 1176.545 18.445 1176.715 18.615 ;
      LAYER met1 ;
        RECT 231.170 19.620 231.490 19.680 ;
        RECT 1174.645 19.620 1174.935 19.665 ;
        RECT 231.170 19.480 1174.935 19.620 ;
        RECT 231.170 19.420 231.490 19.480 ;
        RECT 1174.645 19.435 1174.935 19.480 ;
        RECT 1176.485 18.600 1176.775 18.645 ;
        RECT 1198.550 18.600 1198.870 18.660 ;
        RECT 1176.485 18.460 1198.870 18.600 ;
        RECT 1176.485 18.415 1176.775 18.460 ;
        RECT 1198.550 18.400 1198.870 18.460 ;
        RECT 1175.105 17.920 1175.395 17.965 ;
        RECT 1176.485 17.920 1176.775 17.965 ;
        RECT 1175.105 17.780 1176.775 17.920 ;
        RECT 1175.105 17.735 1175.395 17.780 ;
        RECT 1176.485 17.735 1176.775 17.780 ;
      LAYER via ;
        RECT 231.200 19.420 231.460 19.680 ;
        RECT 1198.580 18.400 1198.840 18.660 ;
      LAYER met2 ;
        RECT 231.200 19.390 231.460 19.710 ;
        RECT 231.260 2.400 231.400 19.390 ;
        RECT 1198.640 18.690 1198.780 54.000 ;
        RECT 1198.580 18.370 1198.840 18.690 ;
        RECT 231.190 0.000 231.470 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 52.690 17.580 53.010 17.640 ;
        RECT 57.290 17.580 57.610 17.640 ;
        RECT 52.690 17.440 57.610 17.580 ;
        RECT 52.690 17.380 53.010 17.440 ;
        RECT 57.290 17.380 57.610 17.440 ;
      LAYER via ;
        RECT 52.720 17.380 52.980 17.640 ;
        RECT 57.320 17.380 57.580 17.640 ;
      LAYER met2 ;
        RECT 57.380 17.670 57.520 54.000 ;
        RECT 52.720 17.350 52.980 17.670 ;
        RECT 57.320 17.350 57.580 17.670 ;
        RECT 52.780 2.400 52.920 17.350 ;
        RECT 52.710 0.000 52.990 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 255.090 20.300 255.410 20.360 ;
        RECT 1140.590 20.300 1140.910 20.360 ;
        RECT 255.090 20.160 1140.910 20.300 ;
        RECT 255.090 20.100 255.410 20.160 ;
        RECT 1140.590 20.100 1140.910 20.160 ;
        RECT 1152.090 18.600 1152.410 18.660 ;
        RECT 1176.010 18.600 1176.330 18.660 ;
        RECT 1152.090 18.460 1176.330 18.600 ;
        RECT 1152.090 18.400 1152.410 18.460 ;
        RECT 1176.010 18.400 1176.330 18.460 ;
        RECT 1183.830 17.580 1184.150 17.640 ;
        RECT 1205.450 17.580 1205.770 17.640 ;
        RECT 1183.830 17.440 1205.770 17.580 ;
        RECT 1183.830 17.380 1184.150 17.440 ;
        RECT 1205.450 17.380 1205.770 17.440 ;
      LAYER via ;
        RECT 255.120 20.100 255.380 20.360 ;
        RECT 1140.620 20.100 1140.880 20.360 ;
        RECT 1152.120 18.400 1152.380 18.660 ;
        RECT 1176.040 18.400 1176.300 18.660 ;
        RECT 1183.860 17.380 1184.120 17.640 ;
        RECT 1205.480 17.380 1205.740 17.640 ;
      LAYER met2 ;
        RECT 255.120 20.070 255.380 20.390 ;
        RECT 1140.620 20.070 1140.880 20.390 ;
        RECT 255.180 2.400 255.320 20.070 ;
        RECT 1140.680 18.205 1140.820 20.070 ;
        RECT 1152.120 18.370 1152.380 18.690 ;
        RECT 1176.040 18.370 1176.300 18.690 ;
        RECT 1152.180 18.205 1152.320 18.370 ;
        RECT 1176.100 18.205 1176.240 18.370 ;
        RECT 1140.610 17.835 1140.890 18.205 ;
        RECT 1152.110 17.835 1152.390 18.205 ;
        RECT 1176.030 17.835 1176.310 18.205 ;
        RECT 1183.850 17.835 1184.130 18.205 ;
        RECT 1183.920 17.670 1184.060 17.835 ;
        RECT 1205.540 17.670 1205.680 54.000 ;
        RECT 1183.860 17.350 1184.120 17.670 ;
        RECT 1205.480 17.350 1205.740 17.670 ;
        RECT 255.110 0.000 255.390 2.400 ;
      LAYER via2 ;
        RECT 1140.610 17.880 1140.890 18.160 ;
        RECT 1152.110 17.880 1152.390 18.160 ;
        RECT 1176.030 17.880 1176.310 18.160 ;
        RECT 1183.850 17.880 1184.130 18.160 ;
      LAYER met3 ;
        RECT 1140.585 18.170 1140.915 18.185 ;
        RECT 1152.085 18.170 1152.415 18.185 ;
        RECT 1140.585 17.870 1152.415 18.170 ;
        RECT 1140.585 17.855 1140.915 17.870 ;
        RECT 1152.085 17.855 1152.415 17.870 ;
        RECT 1176.005 18.170 1176.335 18.185 ;
        RECT 1183.825 18.170 1184.155 18.185 ;
        RECT 1176.005 17.870 1184.155 18.170 ;
        RECT 1176.005 17.855 1176.335 17.870 ;
        RECT 1183.825 17.855 1184.155 17.870 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 272.570 14.860 272.890 14.920 ;
        RECT 278.090 14.860 278.410 14.920 ;
        RECT 272.570 14.720 278.410 14.860 ;
        RECT 272.570 14.660 272.890 14.720 ;
        RECT 278.090 14.660 278.410 14.720 ;
      LAYER via ;
        RECT 272.600 14.660 272.860 14.920 ;
        RECT 278.120 14.660 278.380 14.920 ;
      LAYER met2 ;
        RECT 278.180 14.950 278.320 54.000 ;
        RECT 272.600 14.630 272.860 14.950 ;
        RECT 278.120 14.630 278.380 14.950 ;
        RECT 272.660 2.400 272.800 14.630 ;
        RECT 272.590 0.000 272.870 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 290.510 20.640 290.830 20.700 ;
        RECT 1175.550 20.640 1175.870 20.700 ;
        RECT 290.510 20.500 1175.870 20.640 ;
        RECT 290.510 20.440 290.830 20.500 ;
        RECT 1175.550 20.440 1175.870 20.500 ;
        RECT 1190.270 20.640 1190.590 20.700 ;
        RECT 1213.730 20.640 1214.050 20.700 ;
        RECT 1190.270 20.500 1214.050 20.640 ;
        RECT 1190.270 20.440 1190.590 20.500 ;
        RECT 1213.730 20.440 1214.050 20.500 ;
      LAYER via ;
        RECT 290.540 20.440 290.800 20.700 ;
        RECT 1175.580 20.440 1175.840 20.700 ;
        RECT 1190.300 20.440 1190.560 20.700 ;
        RECT 1213.760 20.440 1214.020 20.700 ;
      LAYER met2 ;
        RECT 290.540 20.410 290.800 20.730 ;
        RECT 1175.570 20.555 1175.850 20.925 ;
        RECT 1190.290 20.555 1190.570 20.925 ;
        RECT 1213.820 20.730 1213.960 54.000 ;
        RECT 1175.580 20.410 1175.840 20.555 ;
        RECT 1190.300 20.410 1190.560 20.555 ;
        RECT 1213.760 20.410 1214.020 20.730 ;
        RECT 290.600 2.400 290.740 20.410 ;
        RECT 290.530 0.000 290.810 2.400 ;
      LAYER via2 ;
        RECT 1175.570 20.600 1175.850 20.880 ;
        RECT 1190.290 20.600 1190.570 20.880 ;
      LAYER met3 ;
        RECT 1175.545 20.890 1175.875 20.905 ;
        RECT 1190.265 20.890 1190.595 20.905 ;
        RECT 1175.545 20.590 1190.595 20.890 ;
        RECT 1175.545 20.575 1175.875 20.590 ;
        RECT 1190.265 20.575 1190.595 20.590 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 308.450 16.900 308.770 16.960 ;
        RECT 312.590 16.900 312.910 16.960 ;
        RECT 308.450 16.760 312.910 16.900 ;
        RECT 308.450 16.700 308.770 16.760 ;
        RECT 312.590 16.700 312.910 16.760 ;
      LAYER via ;
        RECT 308.480 16.700 308.740 16.960 ;
        RECT 312.620 16.700 312.880 16.960 ;
      LAYER met2 ;
        RECT 312.680 16.990 312.820 54.000 ;
        RECT 308.480 16.670 308.740 16.990 ;
        RECT 312.620 16.670 312.880 16.990 ;
        RECT 308.540 2.400 308.680 16.670 ;
        RECT 308.470 0.000 308.750 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 326.390 16.900 326.710 16.960 ;
        RECT 1175.550 16.900 1175.870 16.960 ;
        RECT 326.390 16.760 1175.870 16.900 ;
        RECT 326.390 16.700 326.710 16.760 ;
        RECT 1175.550 16.700 1175.870 16.760 ;
        RECT 1185.670 16.900 1185.990 16.960 ;
        RECT 1219.250 16.900 1219.570 16.960 ;
        RECT 1185.670 16.760 1219.570 16.900 ;
        RECT 1185.670 16.700 1185.990 16.760 ;
        RECT 1219.250 16.700 1219.570 16.760 ;
      LAYER via ;
        RECT 326.420 16.700 326.680 16.960 ;
        RECT 1175.580 16.700 1175.840 16.960 ;
        RECT 1185.700 16.700 1185.960 16.960 ;
        RECT 1219.280 16.700 1219.540 16.960 ;
      LAYER met2 ;
        RECT 1175.570 17.155 1175.850 17.525 ;
        RECT 1185.690 17.155 1185.970 17.525 ;
        RECT 1175.640 16.990 1175.780 17.155 ;
        RECT 1185.760 16.990 1185.900 17.155 ;
        RECT 1219.340 16.990 1219.480 54.000 ;
        RECT 326.420 16.670 326.680 16.990 ;
        RECT 1175.580 16.670 1175.840 16.990 ;
        RECT 1185.700 16.670 1185.960 16.990 ;
        RECT 1219.280 16.670 1219.540 16.990 ;
        RECT 326.480 2.400 326.620 16.670 ;
        RECT 326.410 0.000 326.690 2.400 ;
      LAYER via2 ;
        RECT 1175.570 17.200 1175.850 17.480 ;
        RECT 1185.690 17.200 1185.970 17.480 ;
      LAYER met3 ;
        RECT 1175.545 17.490 1175.875 17.505 ;
        RECT 1185.665 17.490 1185.995 17.505 ;
        RECT 1175.545 17.190 1185.995 17.490 ;
        RECT 1175.545 17.175 1175.875 17.190 ;
        RECT 1185.665 17.175 1185.995 17.190 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 343.870 15.880 344.190 15.940 ;
        RECT 347.090 15.880 347.410 15.940 ;
        RECT 343.870 15.740 347.410 15.880 ;
        RECT 343.870 15.680 344.190 15.740 ;
        RECT 347.090 15.680 347.410 15.740 ;
      LAYER via ;
        RECT 343.900 15.680 344.160 15.940 ;
        RECT 347.120 15.680 347.380 15.940 ;
      LAYER met2 ;
        RECT 347.180 15.970 347.320 54.000 ;
        RECT 343.900 15.650 344.160 15.970 ;
        RECT 347.120 15.650 347.380 15.970 ;
        RECT 343.960 2.400 344.100 15.650 ;
        RECT 343.890 0.000 344.170 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 361.810 15.880 362.130 15.940 ;
        RECT 1225.690 15.880 1226.010 15.940 ;
        RECT 361.810 15.740 935.200 15.880 ;
        RECT 361.810 15.680 362.130 15.740 ;
        RECT 935.060 15.540 935.200 15.740 ;
        RECT 981.520 15.740 983.040 15.880 ;
        RECT 981.520 15.540 981.660 15.740 ;
        RECT 935.060 15.400 981.660 15.540 ;
        RECT 982.900 15.540 983.040 15.740 ;
        RECT 1029.820 15.740 1226.010 15.880 ;
        RECT 1029.820 15.540 1029.960 15.740 ;
        RECT 1225.690 15.680 1226.010 15.740 ;
        RECT 982.900 15.400 1029.960 15.540 ;
      LAYER via ;
        RECT 361.840 15.680 362.100 15.940 ;
        RECT 1225.720 15.680 1225.980 15.940 ;
      LAYER met2 ;
        RECT 1225.780 15.970 1225.920 54.000 ;
        RECT 361.840 15.650 362.100 15.970 ;
        RECT 1225.720 15.650 1225.980 15.970 ;
        RECT 361.900 2.400 362.040 15.650 ;
        RECT 361.830 0.000 362.110 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 381.680 16.730 381.820 54.000 ;
        RECT 379.840 16.590 381.820 16.730 ;
        RECT 379.840 2.400 379.980 16.590 ;
        RECT 379.770 0.000 380.050 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 934.585 15.385 935.215 15.555 ;
        RECT 935.045 15.045 935.215 15.385 ;
        RECT 1029.805 15.385 1030.435 15.555 ;
        RECT 981.045 15.045 983.055 15.215 ;
        RECT 1029.805 15.045 1029.975 15.385 ;
      LAYER mcon ;
        RECT 1030.265 15.385 1030.435 15.555 ;
        RECT 982.885 15.045 983.055 15.215 ;
      LAYER met1 ;
        RECT 934.525 15.540 934.815 15.585 ;
        RECT 426.760 15.400 934.815 15.540 ;
        RECT 397.690 15.200 398.010 15.260 ;
        RECT 426.760 15.200 426.900 15.400 ;
        RECT 934.525 15.355 934.815 15.400 ;
        RECT 1030.205 15.540 1030.495 15.585 ;
        RECT 1233.050 15.540 1233.370 15.600 ;
        RECT 1030.205 15.400 1233.370 15.540 ;
        RECT 1030.205 15.355 1030.495 15.400 ;
        RECT 1233.050 15.340 1233.370 15.400 ;
        RECT 397.690 15.060 426.900 15.200 ;
        RECT 934.985 15.200 935.275 15.245 ;
        RECT 980.985 15.200 981.275 15.245 ;
        RECT 934.985 15.060 981.275 15.200 ;
        RECT 397.690 15.000 398.010 15.060 ;
        RECT 934.985 15.015 935.275 15.060 ;
        RECT 980.985 15.015 981.275 15.060 ;
        RECT 982.825 15.200 983.115 15.245 ;
        RECT 1029.745 15.200 1030.035 15.245 ;
        RECT 982.825 15.060 1030.035 15.200 ;
        RECT 982.825 15.015 983.115 15.060 ;
        RECT 1029.745 15.015 1030.035 15.060 ;
      LAYER via ;
        RECT 397.720 15.000 397.980 15.260 ;
        RECT 1233.080 15.340 1233.340 15.600 ;
      LAYER met2 ;
        RECT 1233.140 15.630 1233.280 54.000 ;
        RECT 1233.080 15.310 1233.340 15.630 ;
        RECT 397.720 14.970 397.980 15.290 ;
        RECT 397.780 2.400 397.920 14.970 ;
        RECT 397.710 0.000 397.990 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 416.180 17.410 416.320 54.000 ;
        RECT 415.720 17.270 416.320 17.410 ;
        RECT 415.720 2.400 415.860 17.270 ;
        RECT 415.650 0.000 415.930 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 291.060 17.950 292.120 18.090 ;
        RECT 291.060 17.525 291.200 17.950 ;
        RECT 291.980 17.525 292.120 17.950 ;
        RECT 76.630 17.155 76.910 17.525 ;
        RECT 290.990 17.155 291.270 17.525 ;
        RECT 291.910 17.155 292.190 17.525 ;
        RECT 76.700 2.400 76.840 17.155 ;
        RECT 1163.680 16.845 1163.820 54.000 ;
        RECT 1163.610 16.475 1163.890 16.845 ;
        RECT 76.630 0.000 76.910 2.400 ;
      LAYER via2 ;
        RECT 76.630 17.200 76.910 17.480 ;
        RECT 290.990 17.200 291.270 17.480 ;
        RECT 291.910 17.200 292.190 17.480 ;
        RECT 1163.610 16.520 1163.890 16.800 ;
      LAYER met3 ;
        RECT 76.605 17.490 76.935 17.505 ;
        RECT 290.965 17.490 291.295 17.505 ;
        RECT 76.605 17.190 291.295 17.490 ;
        RECT 76.605 17.175 76.935 17.190 ;
        RECT 290.965 17.175 291.295 17.190 ;
        RECT 291.885 17.490 292.215 17.505 ;
        RECT 291.885 17.190 1139.290 17.490 ;
        RECT 291.885 17.175 292.215 17.190 ;
        RECT 1138.990 16.810 1139.290 17.190 ;
        RECT 1163.585 16.810 1163.915 16.825 ;
        RECT 1138.990 16.510 1163.915 16.810 ;
        RECT 1163.585 16.495 1163.915 16.510 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 433.110 15.200 433.430 15.260 ;
        RECT 436.790 15.200 437.110 15.260 ;
        RECT 433.110 15.060 437.110 15.200 ;
        RECT 433.110 15.000 433.430 15.060 ;
        RECT 436.790 15.000 437.110 15.060 ;
      LAYER via ;
        RECT 433.140 15.000 433.400 15.260 ;
        RECT 436.820 15.000 437.080 15.260 ;
      LAYER met2 ;
        RECT 436.880 15.290 437.020 54.000 ;
        RECT 433.140 14.970 433.400 15.290 ;
        RECT 436.820 14.970 437.080 15.290 ;
        RECT 433.200 2.400 433.340 14.970 ;
        RECT 433.130 0.000 433.410 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 934.050 15.200 934.370 15.260 ;
        RECT 513.240 15.060 934.370 15.200 ;
        RECT 451.050 14.860 451.370 14.920 ;
        RECT 513.240 14.860 513.380 15.060 ;
        RECT 934.050 15.000 934.370 15.060 ;
        RECT 1038.470 15.200 1038.790 15.260 ;
        RECT 1239.490 15.200 1239.810 15.260 ;
        RECT 1038.470 15.060 1239.810 15.200 ;
        RECT 1038.470 15.000 1038.790 15.060 ;
        RECT 1239.490 15.000 1239.810 15.060 ;
        RECT 451.050 14.720 513.380 14.860 ;
        RECT 935.430 14.860 935.750 14.920 ;
        RECT 979.590 14.860 979.910 14.920 ;
        RECT 935.430 14.720 979.910 14.860 ;
        RECT 451.050 14.660 451.370 14.720 ;
        RECT 935.430 14.660 935.750 14.720 ;
        RECT 979.590 14.660 979.910 14.720 ;
      LAYER via ;
        RECT 451.080 14.660 451.340 14.920 ;
        RECT 934.080 15.000 934.340 15.260 ;
        RECT 1038.500 15.000 1038.760 15.260 ;
        RECT 1239.520 15.000 1239.780 15.260 ;
        RECT 935.460 14.660 935.720 14.920 ;
        RECT 979.620 14.660 979.880 14.920 ;
      LAYER met2 ;
        RECT 934.140 15.290 935.660 15.370 ;
        RECT 1239.580 15.290 1239.720 54.000 ;
        RECT 934.080 15.230 935.660 15.290 ;
        RECT 934.080 14.970 934.340 15.230 ;
        RECT 935.520 14.950 935.660 15.230 ;
        RECT 1038.500 14.970 1038.760 15.290 ;
        RECT 1239.520 14.970 1239.780 15.290 ;
        RECT 451.080 14.630 451.340 14.950 ;
        RECT 935.460 14.630 935.720 14.950 ;
        RECT 979.620 14.805 979.880 14.950 ;
        RECT 1038.560 14.805 1038.700 14.970 ;
        RECT 451.140 2.400 451.280 14.630 ;
        RECT 979.610 14.435 979.890 14.805 ;
        RECT 1038.490 14.435 1038.770 14.805 ;
        RECT 451.070 0.000 451.350 2.400 ;
      LAYER via2 ;
        RECT 979.610 14.480 979.890 14.760 ;
        RECT 1038.490 14.480 1038.770 14.760 ;
      LAYER met3 ;
        RECT 979.585 14.770 979.915 14.785 ;
        RECT 1038.465 14.770 1038.795 14.785 ;
        RECT 979.585 14.470 1038.795 14.770 ;
        RECT 979.585 14.455 979.915 14.470 ;
        RECT 1038.465 14.455 1038.795 14.470 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 468.990 17.580 469.310 17.640 ;
        RECT 471.290 17.580 471.610 17.640 ;
        RECT 468.990 17.440 471.610 17.580 ;
        RECT 468.990 17.380 469.310 17.440 ;
        RECT 471.290 17.380 471.610 17.440 ;
      LAYER via ;
        RECT 469.020 17.380 469.280 17.640 ;
        RECT 471.320 17.380 471.580 17.640 ;
      LAYER met2 ;
        RECT 471.380 17.670 471.520 54.000 ;
        RECT 469.020 17.350 469.280 17.670 ;
        RECT 471.320 17.350 471.580 17.670 ;
        RECT 469.080 2.400 469.220 17.350 ;
        RECT 469.010 0.000 469.290 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 981.045 13.005 981.215 14.535 ;
        RECT 992.545 13.005 992.715 14.875 ;
        RECT 1029.345 14.705 1030.895 14.875 ;
      LAYER mcon ;
        RECT 992.545 14.705 992.715 14.875 ;
        RECT 1030.725 14.705 1030.895 14.875 ;
        RECT 981.045 14.365 981.215 14.535 ;
      LAYER met1 ;
        RECT 992.485 14.860 992.775 14.905 ;
        RECT 1029.285 14.860 1029.575 14.905 ;
        RECT 543.600 14.720 935.200 14.860 ;
        RECT 486.930 14.180 487.250 14.240 ;
        RECT 543.600 14.180 543.740 14.720 ;
        RECT 935.060 14.520 935.200 14.720 ;
        RECT 992.485 14.720 1029.575 14.860 ;
        RECT 992.485 14.675 992.775 14.720 ;
        RECT 1029.285 14.675 1029.575 14.720 ;
        RECT 1030.665 14.860 1030.955 14.905 ;
        RECT 1253.290 14.860 1253.610 14.920 ;
        RECT 1030.665 14.720 1253.610 14.860 ;
        RECT 1030.665 14.675 1030.955 14.720 ;
        RECT 1253.290 14.660 1253.610 14.720 ;
        RECT 980.985 14.520 981.275 14.565 ;
        RECT 935.060 14.380 981.275 14.520 ;
        RECT 980.985 14.335 981.275 14.380 ;
        RECT 486.930 14.040 543.740 14.180 ;
        RECT 486.930 13.980 487.250 14.040 ;
        RECT 980.985 13.160 981.275 13.205 ;
        RECT 992.485 13.160 992.775 13.205 ;
        RECT 980.985 13.020 992.775 13.160 ;
        RECT 980.985 12.975 981.275 13.020 ;
        RECT 992.485 12.975 992.775 13.020 ;
      LAYER via ;
        RECT 486.960 13.980 487.220 14.240 ;
        RECT 1253.320 14.660 1253.580 14.920 ;
      LAYER met2 ;
        RECT 1253.380 14.950 1253.520 54.000 ;
        RECT 1253.320 14.630 1253.580 14.950 ;
        RECT 486.960 13.950 487.220 14.270 ;
        RECT 487.020 2.400 487.160 13.950 ;
        RECT 486.950 0.000 487.230 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 505.880 16.730 506.020 54.000 ;
        RECT 504.960 16.590 506.020 16.730 ;
        RECT 504.960 2.400 505.100 16.590 ;
        RECT 504.890 0.000 505.170 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 543.125 14.195 543.295 14.535 ;
        RECT 934.125 14.195 934.295 14.535 ;
        RECT 981.505 14.365 982.595 14.535 ;
        RECT 543.125 14.025 544.215 14.195 ;
        RECT 563.825 14.025 567.215 14.195 ;
        RECT 934.125 14.025 935.215 14.195 ;
        RECT 981.505 14.025 981.675 14.365 ;
      LAYER mcon ;
        RECT 543.125 14.365 543.295 14.535 ;
        RECT 934.125 14.365 934.295 14.535 ;
        RECT 982.425 14.365 982.595 14.535 ;
        RECT 544.045 14.025 544.215 14.195 ;
        RECT 567.045 14.025 567.215 14.195 ;
        RECT 935.045 14.025 935.215 14.195 ;
      LAYER met1 ;
        RECT 522.350 14.520 522.670 14.580 ;
        RECT 543.065 14.520 543.355 14.565 ;
        RECT 934.065 14.520 934.355 14.565 ;
        RECT 522.350 14.380 543.355 14.520 ;
        RECT 522.350 14.320 522.670 14.380 ;
        RECT 543.065 14.335 543.355 14.380 ;
        RECT 567.980 14.380 934.355 14.520 ;
        RECT 543.985 14.180 544.275 14.225 ;
        RECT 563.765 14.180 564.055 14.225 ;
        RECT 543.985 14.040 564.055 14.180 ;
        RECT 543.985 13.995 544.275 14.040 ;
        RECT 563.765 13.995 564.055 14.040 ;
        RECT 566.985 14.180 567.275 14.225 ;
        RECT 567.980 14.180 568.120 14.380 ;
        RECT 934.065 14.335 934.355 14.380 ;
        RECT 982.365 14.520 982.655 14.565 ;
        RECT 1260.650 14.520 1260.970 14.580 ;
        RECT 982.365 14.380 1260.970 14.520 ;
        RECT 982.365 14.335 982.655 14.380 ;
        RECT 1260.650 14.320 1260.970 14.380 ;
        RECT 566.985 14.040 568.120 14.180 ;
        RECT 934.985 14.180 935.275 14.225 ;
        RECT 981.445 14.180 981.735 14.225 ;
        RECT 934.985 14.040 981.735 14.180 ;
        RECT 566.985 13.995 567.275 14.040 ;
        RECT 934.985 13.995 935.275 14.040 ;
        RECT 981.445 13.995 981.735 14.040 ;
      LAYER via ;
        RECT 522.380 14.320 522.640 14.580 ;
        RECT 1260.680 14.320 1260.940 14.580 ;
      LAYER met2 ;
        RECT 1260.740 14.610 1260.880 54.000 ;
        RECT 522.380 14.290 522.640 14.610 ;
        RECT 1260.680 14.290 1260.940 14.610 ;
        RECT 522.440 2.400 522.580 14.290 ;
        RECT 522.370 0.000 522.650 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 540.380 2.400 540.520 54.000 ;
        RECT 540.310 0.000 540.590 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 935.505 14.535 935.675 17.255 ;
        RECT 567.505 13.005 567.675 14.535 ;
        RECT 934.585 14.365 935.675 14.535 ;
        RECT 568.425 13.005 568.595 14.195 ;
      LAYER mcon ;
        RECT 935.505 17.085 935.675 17.255 ;
        RECT 567.505 14.365 567.675 14.535 ;
        RECT 568.425 14.025 568.595 14.195 ;
      LAYER met1 ;
        RECT 935.445 17.240 935.735 17.285 ;
        RECT 981.430 17.240 981.750 17.300 ;
        RECT 935.445 17.100 981.750 17.240 ;
        RECT 935.445 17.055 935.735 17.100 ;
        RECT 981.430 17.040 981.750 17.100 ;
        RECT 558.230 14.520 558.550 14.580 ;
        RECT 567.445 14.520 567.735 14.565 ;
        RECT 558.230 14.380 567.735 14.520 ;
        RECT 558.230 14.320 558.550 14.380 ;
        RECT 567.445 14.335 567.735 14.380 ;
        RECT 934.525 14.335 934.815 14.565 ;
        RECT 568.365 14.180 568.655 14.225 ;
        RECT 934.600 14.180 934.740 14.335 ;
        RECT 568.365 14.040 934.740 14.180 ;
        RECT 981.890 14.180 982.210 14.240 ;
        RECT 1267.090 14.180 1267.410 14.240 ;
        RECT 981.890 14.040 1267.410 14.180 ;
        RECT 568.365 13.995 568.655 14.040 ;
        RECT 981.890 13.980 982.210 14.040 ;
        RECT 1267.090 13.980 1267.410 14.040 ;
        RECT 567.445 13.160 567.735 13.205 ;
        RECT 568.365 13.160 568.655 13.205 ;
        RECT 567.445 13.020 568.655 13.160 ;
        RECT 567.445 12.975 567.735 13.020 ;
        RECT 568.365 12.975 568.655 13.020 ;
      LAYER via ;
        RECT 981.460 17.040 981.720 17.300 ;
        RECT 558.260 14.320 558.520 14.580 ;
        RECT 981.920 13.980 982.180 14.240 ;
        RECT 1267.120 13.980 1267.380 14.240 ;
      LAYER met2 ;
        RECT 981.460 17.010 981.720 17.330 ;
        RECT 558.260 14.290 558.520 14.610 ;
        RECT 558.320 2.400 558.460 14.290 ;
        RECT 981.520 14.180 981.660 17.010 ;
        RECT 1267.180 14.270 1267.320 54.000 ;
        RECT 981.920 14.180 982.180 14.270 ;
        RECT 981.520 14.040 982.180 14.180 ;
        RECT 981.920 13.950 982.180 14.040 ;
        RECT 1267.120 13.950 1267.380 14.270 ;
        RECT 558.250 0.000 558.530 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 576.170 17.580 576.490 17.640 ;
        RECT 581.690 17.580 582.010 17.640 ;
        RECT 576.170 17.440 582.010 17.580 ;
        RECT 576.170 17.380 576.490 17.440 ;
        RECT 581.690 17.380 582.010 17.440 ;
      LAYER via ;
        RECT 576.200 17.380 576.460 17.640 ;
        RECT 581.720 17.380 581.980 17.640 ;
      LAYER met2 ;
        RECT 581.780 17.670 581.920 54.000 ;
        RECT 576.200 17.350 576.460 17.670 ;
        RECT 581.720 17.350 581.980 17.670 ;
        RECT 576.260 2.400 576.400 17.350 ;
        RECT 576.190 0.000 576.470 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 885.825 21.165 887.375 21.335 ;
        RECT 664.565 14.025 666.575 14.195 ;
        RECT 664.565 12.665 664.735 14.025 ;
        RECT 666.405 12.665 666.575 14.025 ;
        RECT 712.865 12.665 713.035 17.255 ;
        RECT 761.625 12.665 761.795 17.255 ;
        RECT 809.465 12.665 809.635 17.595 ;
        RECT 885.825 17.425 885.995 21.165 ;
        RECT 954.825 12.665 954.995 21.335 ;
        RECT 1002.665 14.025 1003.295 14.195 ;
        RECT 1002.665 12.665 1002.835 14.025 ;
        RECT 1003.125 12.665 1003.295 14.025 ;
        RECT 1050.965 12.665 1051.135 17.255 ;
        RECT 1126.865 17.085 1127.495 17.255 ;
      LAYER mcon ;
        RECT 887.205 21.165 887.375 21.335 ;
        RECT 954.825 21.165 954.995 21.335 ;
        RECT 809.465 17.425 809.635 17.595 ;
        RECT 712.865 17.085 713.035 17.255 ;
        RECT 761.625 17.085 761.795 17.255 ;
        RECT 1050.965 17.085 1051.135 17.255 ;
        RECT 1127.325 17.085 1127.495 17.255 ;
      LAYER met1 ;
        RECT 887.145 21.320 887.435 21.365 ;
        RECT 954.765 21.320 955.055 21.365 ;
        RECT 887.145 21.180 955.055 21.320 ;
        RECT 887.145 21.135 887.435 21.180 ;
        RECT 954.765 21.135 955.055 21.180 ;
        RECT 809.405 17.580 809.695 17.625 ;
        RECT 885.765 17.580 886.055 17.625 ;
        RECT 809.405 17.440 886.055 17.580 ;
        RECT 809.405 17.395 809.695 17.440 ;
        RECT 885.765 17.395 886.055 17.440 ;
        RECT 712.805 17.240 713.095 17.285 ;
        RECT 761.565 17.240 761.855 17.285 ;
        RECT 712.805 17.100 761.855 17.240 ;
        RECT 712.805 17.055 713.095 17.100 ;
        RECT 761.565 17.055 761.855 17.100 ;
        RECT 1050.905 17.240 1051.195 17.285 ;
        RECT 1126.805 17.240 1127.095 17.285 ;
        RECT 1050.905 17.100 1127.095 17.240 ;
        RECT 1050.905 17.055 1051.195 17.100 ;
        RECT 1126.805 17.055 1127.095 17.100 ;
        RECT 1127.265 17.240 1127.555 17.285 ;
        RECT 1273.530 17.240 1273.850 17.300 ;
        RECT 1127.265 17.100 1273.850 17.240 ;
        RECT 1127.265 17.055 1127.555 17.100 ;
        RECT 1273.530 17.040 1273.850 17.100 ;
        RECT 593.650 12.820 593.970 12.880 ;
        RECT 664.505 12.820 664.795 12.865 ;
        RECT 593.650 12.680 664.795 12.820 ;
        RECT 593.650 12.620 593.970 12.680 ;
        RECT 664.505 12.635 664.795 12.680 ;
        RECT 666.345 12.820 666.635 12.865 ;
        RECT 712.805 12.820 713.095 12.865 ;
        RECT 666.345 12.680 713.095 12.820 ;
        RECT 666.345 12.635 666.635 12.680 ;
        RECT 712.805 12.635 713.095 12.680 ;
        RECT 761.565 12.820 761.855 12.865 ;
        RECT 809.405 12.820 809.695 12.865 ;
        RECT 761.565 12.680 809.695 12.820 ;
        RECT 761.565 12.635 761.855 12.680 ;
        RECT 809.405 12.635 809.695 12.680 ;
        RECT 954.765 12.820 955.055 12.865 ;
        RECT 1002.605 12.820 1002.895 12.865 ;
        RECT 954.765 12.680 1002.895 12.820 ;
        RECT 954.765 12.635 955.055 12.680 ;
        RECT 1002.605 12.635 1002.895 12.680 ;
        RECT 1003.065 12.820 1003.355 12.865 ;
        RECT 1050.905 12.820 1051.195 12.865 ;
        RECT 1003.065 12.680 1051.195 12.820 ;
        RECT 1003.065 12.635 1003.355 12.680 ;
        RECT 1050.905 12.635 1051.195 12.680 ;
      LAYER via ;
        RECT 1273.560 17.040 1273.820 17.300 ;
        RECT 593.680 12.620 593.940 12.880 ;
      LAYER met2 ;
        RECT 1272.700 46.650 1272.840 54.000 ;
        RECT 1272.700 46.510 1273.760 46.650 ;
        RECT 1273.620 17.330 1273.760 46.510 ;
        RECT 1273.560 17.010 1273.820 17.330 ;
        RECT 593.680 12.590 593.940 12.910 ;
        RECT 593.740 2.400 593.880 12.590 ;
        RECT 593.670 0.000 593.950 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 100.070 17.580 100.390 17.640 ;
        RECT 105.590 17.580 105.910 17.640 ;
        RECT 100.070 17.440 105.910 17.580 ;
        RECT 100.070 17.380 100.390 17.440 ;
        RECT 105.590 17.380 105.910 17.440 ;
      LAYER via ;
        RECT 100.100 17.380 100.360 17.640 ;
        RECT 105.620 17.380 105.880 17.640 ;
      LAYER met2 ;
        RECT 105.680 17.670 105.820 54.000 ;
        RECT 100.100 17.350 100.360 17.670 ;
        RECT 105.620 17.350 105.880 17.670 ;
        RECT 100.160 2.400 100.300 17.350 ;
        RECT 100.090 0.000 100.370 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 616.725 13.005 616.895 20.995 ;
        RECT 644.785 17.425 644.955 20.995 ;
        RECT 692.165 17.595 692.335 19.975 ;
        RECT 1099.265 17.935 1099.435 19.975 ;
        RECT 1099.265 17.765 1099.895 17.935 ;
        RECT 691.705 17.425 692.335 17.595 ;
        RECT 1099.725 12.665 1099.895 17.765 ;
        RECT 1148.485 12.665 1148.655 20.315 ;
        RECT 1247.845 17.425 1248.015 18.615 ;
      LAYER mcon ;
        RECT 616.725 20.825 616.895 20.995 ;
        RECT 644.785 20.825 644.955 20.995 ;
        RECT 1148.485 20.145 1148.655 20.315 ;
        RECT 692.165 19.805 692.335 19.975 ;
        RECT 1099.265 19.805 1099.435 19.975 ;
        RECT 1247.845 18.445 1248.015 18.615 ;
      LAYER met1 ;
        RECT 616.665 20.980 616.955 21.025 ;
        RECT 644.725 20.980 645.015 21.025 ;
        RECT 616.665 20.840 645.015 20.980 ;
        RECT 616.665 20.795 616.955 20.840 ;
        RECT 644.725 20.795 645.015 20.840 ;
        RECT 1148.425 20.300 1148.715 20.345 ;
        RECT 1150.710 20.300 1151.030 20.360 ;
        RECT 1148.425 20.160 1151.030 20.300 ;
        RECT 1148.425 20.115 1148.715 20.160 ;
        RECT 1150.710 20.100 1151.030 20.160 ;
        RECT 692.105 19.960 692.395 20.005 ;
        RECT 1078.950 19.960 1079.270 20.020 ;
        RECT 692.105 19.820 1079.270 19.960 ;
        RECT 692.105 19.775 692.395 19.820 ;
        RECT 1078.950 19.760 1079.270 19.820 ;
        RECT 1098.730 19.960 1099.050 20.020 ;
        RECT 1099.205 19.960 1099.495 20.005 ;
        RECT 1098.730 19.820 1099.495 19.960 ;
        RECT 1098.730 19.760 1099.050 19.820 ;
        RECT 1099.205 19.775 1099.495 19.820 ;
        RECT 1247.785 18.600 1248.075 18.645 ;
        RECT 1273.990 18.600 1274.310 18.660 ;
        RECT 1247.785 18.460 1274.310 18.600 ;
        RECT 1247.785 18.415 1248.075 18.460 ;
        RECT 1273.990 18.400 1274.310 18.460 ;
        RECT 1174.630 18.260 1174.950 18.320 ;
        RECT 1174.630 18.120 1206.140 18.260 ;
        RECT 1174.630 18.060 1174.950 18.120 ;
        RECT 644.725 17.580 645.015 17.625 ;
        RECT 691.645 17.580 691.935 17.625 ;
        RECT 644.725 17.440 691.935 17.580 ;
        RECT 1206.000 17.580 1206.140 18.120 ;
        RECT 1247.785 17.580 1248.075 17.625 ;
        RECT 1206.000 17.440 1248.075 17.580 ;
        RECT 644.725 17.395 645.015 17.440 ;
        RECT 691.645 17.395 691.935 17.440 ;
        RECT 1247.785 17.395 1248.075 17.440 ;
        RECT 611.590 13.160 611.910 13.220 ;
        RECT 616.665 13.160 616.955 13.205 ;
        RECT 611.590 13.020 616.955 13.160 ;
        RECT 611.590 12.960 611.910 13.020 ;
        RECT 616.665 12.975 616.955 13.020 ;
        RECT 1099.665 12.820 1099.955 12.865 ;
        RECT 1148.425 12.820 1148.715 12.865 ;
        RECT 1099.665 12.680 1148.715 12.820 ;
        RECT 1099.665 12.635 1099.955 12.680 ;
        RECT 1148.425 12.635 1148.715 12.680 ;
      LAYER via ;
        RECT 1150.740 20.100 1151.000 20.360 ;
        RECT 1078.980 19.760 1079.240 20.020 ;
        RECT 1098.760 19.760 1099.020 20.020 ;
        RECT 1274.020 18.400 1274.280 18.660 ;
        RECT 1174.660 18.060 1174.920 18.320 ;
        RECT 611.620 12.960 611.880 13.220 ;
      LAYER met2 ;
        RECT 1078.970 20.555 1079.250 20.925 ;
        RECT 1098.750 20.555 1099.030 20.925 ;
        RECT 1150.730 20.555 1151.010 20.925 ;
        RECT 1174.650 20.555 1174.930 20.925 ;
        RECT 1079.040 20.050 1079.180 20.555 ;
        RECT 1098.820 20.050 1098.960 20.555 ;
        RECT 1150.800 20.390 1150.940 20.555 ;
        RECT 1150.740 20.070 1151.000 20.390 ;
        RECT 1078.980 19.730 1079.240 20.050 ;
        RECT 1098.760 19.730 1099.020 20.050 ;
        RECT 1174.720 18.350 1174.860 20.555 ;
        RECT 1274.080 18.690 1274.220 54.000 ;
        RECT 1274.020 18.370 1274.280 18.690 ;
        RECT 1174.660 18.030 1174.920 18.350 ;
        RECT 611.620 12.930 611.880 13.250 ;
        RECT 611.680 2.400 611.820 12.930 ;
        RECT 611.610 0.000 611.890 2.400 ;
      LAYER via2 ;
        RECT 1078.970 20.600 1079.250 20.880 ;
        RECT 1098.750 20.600 1099.030 20.880 ;
        RECT 1150.730 20.600 1151.010 20.880 ;
        RECT 1174.650 20.600 1174.930 20.880 ;
      LAYER met3 ;
        RECT 1078.945 20.890 1079.275 20.905 ;
        RECT 1098.725 20.890 1099.055 20.905 ;
        RECT 1078.945 20.590 1099.055 20.890 ;
        RECT 1078.945 20.575 1079.275 20.590 ;
        RECT 1098.725 20.575 1099.055 20.590 ;
        RECT 1150.705 20.890 1151.035 20.905 ;
        RECT 1174.625 20.890 1174.955 20.905 ;
        RECT 1150.705 20.590 1174.955 20.890 ;
        RECT 1150.705 20.575 1151.035 20.590 ;
        RECT 1174.625 20.575 1174.955 20.590 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 630.080 17.410 630.220 54.000 ;
        RECT 629.620 17.270 630.220 17.410 ;
        RECT 629.620 2.400 629.760 17.270 ;
        RECT 629.550 0.000 629.830 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1177.940 18.885 1178.080 54.000 ;
        RECT 124.010 18.515 124.290 18.885 ;
        RECT 1177.870 18.515 1178.150 18.885 ;
        RECT 124.080 2.400 124.220 18.515 ;
        RECT 124.010 0.000 124.290 2.400 ;
      LAYER via2 ;
        RECT 124.010 18.560 124.290 18.840 ;
        RECT 1177.870 18.560 1178.150 18.840 ;
      LAYER met3 ;
        RECT 123.985 18.850 124.315 18.865 ;
        RECT 1177.845 18.850 1178.175 18.865 ;
        RECT 123.985 18.550 1178.175 18.850 ;
        RECT 123.985 18.535 124.315 18.550 ;
        RECT 1177.845 18.535 1178.175 18.550 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 147.910 17.920 148.230 17.980 ;
        RECT 153.890 17.920 154.210 17.980 ;
        RECT 147.910 17.780 154.210 17.920 ;
        RECT 147.910 17.720 148.230 17.780 ;
        RECT 153.890 17.720 154.210 17.780 ;
      LAYER via ;
        RECT 147.940 17.720 148.200 17.980 ;
        RECT 153.920 17.720 154.180 17.980 ;
      LAYER met2 ;
        RECT 153.980 18.010 154.120 54.000 ;
        RECT 147.940 17.690 148.200 18.010 ;
        RECT 153.920 17.690 154.180 18.010 ;
        RECT 148.000 2.400 148.140 17.690 ;
        RECT 147.930 0.000 148.210 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 837.525 21.165 838.615 21.335 ;
        RECT 200.885 15.385 201.055 16.915 ;
        RECT 229.405 15.385 229.575 17.255 ;
        RECT 281.845 15.385 282.015 17.255 ;
        RECT 326.005 15.385 326.175 17.595 ;
        RECT 641.105 17.425 644.495 17.595 ;
        RECT 644.325 17.255 644.495 17.425 ;
        RECT 375.685 14.365 375.855 17.255 ;
        RECT 422.605 14.365 422.775 17.255 ;
        RECT 644.325 17.085 645.415 17.255 ;
        RECT 664.105 13.005 664.275 17.255 ;
        RECT 666.865 13.005 667.035 17.255 ;
        RECT 711.945 13.005 712.115 17.255 ;
        RECT 713.785 13.005 713.955 18.275 ;
        RECT 742.305 18.105 747.995 18.275 ;
        RECT 760.705 13.005 760.875 18.275 ;
        RECT 762.545 13.005 762.715 17.255 ;
        RECT 808.085 13.005 808.255 17.595 ;
        RECT 810.385 13.005 810.555 18.275 ;
        RECT 813.605 18.105 816.995 18.275 ;
        RECT 831.545 18.105 837.235 18.275 ;
        RECT 837.525 18.105 837.695 21.165 ;
        RECT 838.445 20.825 838.615 21.165 ;
        RECT 857.305 13.005 857.475 20.995 ;
        RECT 858.685 13.005 858.855 20.995 ;
        RECT 884.445 17.935 884.615 20.995 ;
        RECT 885.365 17.935 885.535 18.275 ;
        RECT 884.445 17.765 885.535 17.935 ;
        RECT 905.605 13.005 905.775 18.275 ;
        RECT 906.985 13.005 907.155 17.595 ;
        RECT 953.905 13.005 954.075 20.995 ;
        RECT 955.285 13.005 955.455 20.995 ;
        RECT 1001.285 13.005 1001.455 20.995 ;
        RECT 1003.585 13.005 1003.755 20.995 ;
        RECT 1087.305 19.805 1087.475 21.335 ;
        RECT 1092.825 19.805 1092.995 21.335 ;
        RECT 1098.345 19.805 1098.975 19.975 ;
        RECT 1049.585 13.005 1049.755 17.255 ;
        RECT 1051.885 13.005 1052.055 18.275 ;
        RECT 1098.805 13.005 1098.975 19.805 ;
      LAYER mcon ;
        RECT 1087.305 21.165 1087.475 21.335 ;
        RECT 857.305 20.825 857.475 20.995 ;
        RECT 713.785 18.105 713.955 18.275 ;
        RECT 747.825 18.105 747.995 18.275 ;
        RECT 760.705 18.105 760.875 18.275 ;
        RECT 326.005 17.425 326.175 17.595 ;
        RECT 229.405 17.085 229.575 17.255 ;
        RECT 200.885 16.745 201.055 16.915 ;
        RECT 281.845 17.085 282.015 17.255 ;
        RECT 375.685 17.085 375.855 17.255 ;
        RECT 422.605 17.085 422.775 17.255 ;
        RECT 645.245 17.085 645.415 17.255 ;
        RECT 664.105 17.085 664.275 17.255 ;
        RECT 666.865 17.085 667.035 17.255 ;
        RECT 711.945 17.085 712.115 17.255 ;
        RECT 810.385 18.105 810.555 18.275 ;
        RECT 816.825 18.105 816.995 18.275 ;
        RECT 837.065 18.105 837.235 18.275 ;
        RECT 808.085 17.425 808.255 17.595 ;
        RECT 762.545 17.085 762.715 17.255 ;
        RECT 858.685 20.825 858.855 20.995 ;
        RECT 884.445 20.825 884.615 20.995 ;
        RECT 953.905 20.825 954.075 20.995 ;
        RECT 885.365 18.105 885.535 18.275 ;
        RECT 905.605 18.105 905.775 18.275 ;
        RECT 906.985 17.425 907.155 17.595 ;
        RECT 955.285 20.825 955.455 20.995 ;
        RECT 1001.285 20.825 1001.455 20.995 ;
        RECT 1003.585 20.825 1003.755 20.995 ;
        RECT 1092.825 21.165 1092.995 21.335 ;
        RECT 1051.885 18.105 1052.055 18.275 ;
        RECT 1049.585 17.085 1049.755 17.255 ;
      LAYER met1 ;
        RECT 1087.245 21.320 1087.535 21.365 ;
        RECT 1092.765 21.320 1093.055 21.365 ;
        RECT 1087.245 21.180 1093.055 21.320 ;
        RECT 1087.245 21.135 1087.535 21.180 ;
        RECT 1092.765 21.135 1093.055 21.180 ;
        RECT 838.385 20.980 838.675 21.025 ;
        RECT 857.245 20.980 857.535 21.025 ;
        RECT 838.385 20.840 857.535 20.980 ;
        RECT 838.385 20.795 838.675 20.840 ;
        RECT 857.245 20.795 857.535 20.840 ;
        RECT 858.625 20.980 858.915 21.025 ;
        RECT 884.385 20.980 884.675 21.025 ;
        RECT 858.625 20.840 884.675 20.980 ;
        RECT 858.625 20.795 858.915 20.840 ;
        RECT 884.385 20.795 884.675 20.840 ;
        RECT 934.050 20.980 934.370 21.040 ;
        RECT 953.845 20.980 954.135 21.025 ;
        RECT 934.050 20.840 954.135 20.980 ;
        RECT 934.050 20.780 934.370 20.840 ;
        RECT 953.845 20.795 954.135 20.840 ;
        RECT 955.225 20.980 955.515 21.025 ;
        RECT 981.890 20.980 982.210 21.040 ;
        RECT 955.225 20.840 982.210 20.980 ;
        RECT 955.225 20.795 955.515 20.840 ;
        RECT 981.890 20.780 982.210 20.840 ;
        RECT 982.350 20.980 982.670 21.040 ;
        RECT 1001.225 20.980 1001.515 21.025 ;
        RECT 982.350 20.840 1001.515 20.980 ;
        RECT 982.350 20.780 982.670 20.840 ;
        RECT 1001.225 20.795 1001.515 20.840 ;
        RECT 1003.525 20.980 1003.815 21.025 ;
        RECT 1030.190 20.980 1030.510 21.040 ;
        RECT 1003.525 20.840 1030.510 20.980 ;
        RECT 1003.525 20.795 1003.815 20.840 ;
        RECT 1030.190 20.780 1030.510 20.840 ;
        RECT 1079.410 19.960 1079.730 20.020 ;
        RECT 1087.245 19.960 1087.535 20.005 ;
        RECT 1079.410 19.820 1087.535 19.960 ;
        RECT 1079.410 19.760 1079.730 19.820 ;
        RECT 1087.245 19.775 1087.535 19.820 ;
        RECT 1092.765 19.960 1093.055 20.005 ;
        RECT 1098.285 19.960 1098.575 20.005 ;
        RECT 1092.765 19.820 1098.575 19.960 ;
        RECT 1092.765 19.775 1093.055 19.820 ;
        RECT 1098.285 19.775 1098.575 19.820 ;
        RECT 713.725 18.260 714.015 18.305 ;
        RECT 742.245 18.260 742.535 18.305 ;
        RECT 713.725 18.120 742.535 18.260 ;
        RECT 713.725 18.075 714.015 18.120 ;
        RECT 742.245 18.075 742.535 18.120 ;
        RECT 747.765 18.260 748.055 18.305 ;
        RECT 760.645 18.260 760.935 18.305 ;
        RECT 747.765 18.120 760.935 18.260 ;
        RECT 747.765 18.075 748.055 18.120 ;
        RECT 760.645 18.075 760.935 18.120 ;
        RECT 810.325 18.260 810.615 18.305 ;
        RECT 813.545 18.260 813.835 18.305 ;
        RECT 810.325 18.120 813.835 18.260 ;
        RECT 810.325 18.075 810.615 18.120 ;
        RECT 813.545 18.075 813.835 18.120 ;
        RECT 816.765 18.260 817.055 18.305 ;
        RECT 831.485 18.260 831.775 18.305 ;
        RECT 816.765 18.120 831.775 18.260 ;
        RECT 816.765 18.075 817.055 18.120 ;
        RECT 831.485 18.075 831.775 18.120 ;
        RECT 837.005 18.260 837.295 18.305 ;
        RECT 837.465 18.260 837.755 18.305 ;
        RECT 837.005 18.120 837.755 18.260 ;
        RECT 837.005 18.075 837.295 18.120 ;
        RECT 837.465 18.075 837.755 18.120 ;
        RECT 885.305 18.260 885.595 18.305 ;
        RECT 905.545 18.260 905.835 18.305 ;
        RECT 885.305 18.120 905.835 18.260 ;
        RECT 885.305 18.075 885.595 18.120 ;
        RECT 905.545 18.075 905.835 18.120 ;
        RECT 1051.825 18.260 1052.115 18.305 ;
        RECT 1078.950 18.260 1079.270 18.320 ;
        RECT 1051.825 18.120 1079.270 18.260 ;
        RECT 1051.825 18.075 1052.115 18.120 ;
        RECT 1078.950 18.060 1079.270 18.120 ;
        RECT 1100.110 18.260 1100.430 18.320 ;
        RECT 1122.650 18.260 1122.970 18.320 ;
        RECT 1100.110 18.120 1122.970 18.260 ;
        RECT 1100.110 18.060 1100.430 18.120 ;
        RECT 1122.650 18.060 1122.970 18.120 ;
        RECT 1128.170 17.920 1128.490 17.980 ;
        RECT 1173.710 17.920 1174.030 17.980 ;
        RECT 1128.170 17.780 1174.030 17.920 ;
        RECT 1128.170 17.720 1128.490 17.780 ;
        RECT 1173.710 17.720 1174.030 17.780 ;
        RECT 325.945 17.395 326.235 17.625 ;
        RECT 630.450 17.580 630.770 17.640 ;
        RECT 641.045 17.580 641.335 17.625 ;
        RECT 808.025 17.580 808.315 17.625 ;
        RECT 630.450 17.440 641.335 17.580 ;
        RECT 229.345 17.240 229.635 17.285 ;
        RECT 281.785 17.240 282.075 17.285 ;
        RECT 229.345 17.100 282.075 17.240 ;
        RECT 326.020 17.240 326.160 17.395 ;
        RECT 630.450 17.380 630.770 17.440 ;
        RECT 641.045 17.395 641.335 17.440 ;
        RECT 789.700 17.440 808.315 17.580 ;
        RECT 375.625 17.240 375.915 17.285 ;
        RECT 326.020 17.100 375.915 17.240 ;
        RECT 229.345 17.055 229.635 17.100 ;
        RECT 281.785 17.055 282.075 17.100 ;
        RECT 375.625 17.055 375.915 17.100 ;
        RECT 422.545 17.240 422.835 17.285 ;
        RECT 498.430 17.240 498.750 17.300 ;
        RECT 422.545 17.100 498.750 17.240 ;
        RECT 422.545 17.055 422.835 17.100 ;
        RECT 498.430 17.040 498.750 17.100 ;
        RECT 519.130 17.240 519.450 17.300 ;
        RECT 569.270 17.240 569.590 17.300 ;
        RECT 519.130 17.100 569.590 17.240 ;
        RECT 519.130 17.040 519.450 17.100 ;
        RECT 569.270 17.040 569.590 17.100 ;
        RECT 645.185 17.240 645.475 17.285 ;
        RECT 664.045 17.240 664.335 17.285 ;
        RECT 645.185 17.100 664.335 17.240 ;
        RECT 645.185 17.055 645.475 17.100 ;
        RECT 664.045 17.055 664.335 17.100 ;
        RECT 666.805 17.240 667.095 17.285 ;
        RECT 711.885 17.240 712.175 17.285 ;
        RECT 666.805 17.100 712.175 17.240 ;
        RECT 666.805 17.055 667.095 17.100 ;
        RECT 711.885 17.055 712.175 17.100 ;
        RECT 762.485 17.240 762.775 17.285 ;
        RECT 789.700 17.240 789.840 17.440 ;
        RECT 808.025 17.395 808.315 17.440 ;
        RECT 906.925 17.580 907.215 17.625 ;
        RECT 906.925 17.440 933.360 17.580 ;
        RECT 906.925 17.395 907.215 17.440 ;
        RECT 762.485 17.100 789.840 17.240 ;
        RECT 933.220 17.240 933.360 17.440 ;
        RECT 934.050 17.240 934.370 17.300 ;
        RECT 933.220 17.100 934.370 17.240 ;
        RECT 762.485 17.055 762.775 17.100 ;
        RECT 934.050 17.040 934.370 17.100 ;
        RECT 981.890 17.240 982.210 17.300 ;
        RECT 982.350 17.240 982.670 17.300 ;
        RECT 981.890 17.100 982.670 17.240 ;
        RECT 981.890 17.040 982.210 17.100 ;
        RECT 982.350 17.040 982.670 17.100 ;
        RECT 1030.190 17.240 1030.510 17.300 ;
        RECT 1049.525 17.240 1049.815 17.285 ;
        RECT 1030.190 17.100 1049.815 17.240 ;
        RECT 1030.190 17.040 1030.510 17.100 ;
        RECT 1049.525 17.055 1049.815 17.100 ;
        RECT 165.850 16.900 166.170 16.960 ;
        RECT 200.825 16.900 201.115 16.945 ;
        RECT 165.850 16.760 201.115 16.900 ;
        RECT 165.850 16.700 166.170 16.760 ;
        RECT 200.825 16.715 201.115 16.760 ;
        RECT 1176.010 16.900 1176.330 16.960 ;
        RECT 1185.210 16.900 1185.530 16.960 ;
        RECT 1176.010 16.760 1185.530 16.900 ;
        RECT 1176.010 16.700 1176.330 16.760 ;
        RECT 1185.210 16.700 1185.530 16.760 ;
        RECT 200.825 15.540 201.115 15.585 ;
        RECT 229.345 15.540 229.635 15.585 ;
        RECT 200.825 15.400 229.635 15.540 ;
        RECT 200.825 15.355 201.115 15.400 ;
        RECT 229.345 15.355 229.635 15.400 ;
        RECT 281.785 15.540 282.075 15.585 ;
        RECT 325.945 15.540 326.235 15.585 ;
        RECT 281.785 15.400 326.235 15.540 ;
        RECT 281.785 15.355 282.075 15.400 ;
        RECT 325.945 15.355 326.235 15.400 ;
        RECT 375.625 14.520 375.915 14.565 ;
        RECT 422.545 14.520 422.835 14.565 ;
        RECT 375.625 14.380 422.835 14.520 ;
        RECT 375.625 14.335 375.915 14.380 ;
        RECT 422.545 14.335 422.835 14.380 ;
        RECT 664.045 13.160 664.335 13.205 ;
        RECT 666.805 13.160 667.095 13.205 ;
        RECT 664.045 13.020 667.095 13.160 ;
        RECT 664.045 12.975 664.335 13.020 ;
        RECT 666.805 12.975 667.095 13.020 ;
        RECT 711.885 13.160 712.175 13.205 ;
        RECT 713.725 13.160 714.015 13.205 ;
        RECT 711.885 13.020 714.015 13.160 ;
        RECT 711.885 12.975 712.175 13.020 ;
        RECT 713.725 12.975 714.015 13.020 ;
        RECT 760.645 13.160 760.935 13.205 ;
        RECT 762.485 13.160 762.775 13.205 ;
        RECT 760.645 13.020 762.775 13.160 ;
        RECT 760.645 12.975 760.935 13.020 ;
        RECT 762.485 12.975 762.775 13.020 ;
        RECT 808.025 13.160 808.315 13.205 ;
        RECT 810.325 13.160 810.615 13.205 ;
        RECT 808.025 13.020 810.615 13.160 ;
        RECT 808.025 12.975 808.315 13.020 ;
        RECT 810.325 12.975 810.615 13.020 ;
        RECT 857.245 13.160 857.535 13.205 ;
        RECT 858.625 13.160 858.915 13.205 ;
        RECT 857.245 13.020 858.915 13.160 ;
        RECT 857.245 12.975 857.535 13.020 ;
        RECT 858.625 12.975 858.915 13.020 ;
        RECT 905.545 13.160 905.835 13.205 ;
        RECT 906.925 13.160 907.215 13.205 ;
        RECT 905.545 13.020 907.215 13.160 ;
        RECT 905.545 12.975 905.835 13.020 ;
        RECT 906.925 12.975 907.215 13.020 ;
        RECT 953.845 13.160 954.135 13.205 ;
        RECT 955.225 13.160 955.515 13.205 ;
        RECT 953.845 13.020 955.515 13.160 ;
        RECT 953.845 12.975 954.135 13.020 ;
        RECT 955.225 12.975 955.515 13.020 ;
        RECT 1001.225 13.160 1001.515 13.205 ;
        RECT 1003.525 13.160 1003.815 13.205 ;
        RECT 1001.225 13.020 1003.815 13.160 ;
        RECT 1001.225 12.975 1001.515 13.020 ;
        RECT 1003.525 12.975 1003.815 13.020 ;
        RECT 1049.525 13.160 1049.815 13.205 ;
        RECT 1051.825 13.160 1052.115 13.205 ;
        RECT 1049.525 13.020 1052.115 13.160 ;
        RECT 1049.525 12.975 1049.815 13.020 ;
        RECT 1051.825 12.975 1052.115 13.020 ;
        RECT 1098.745 13.160 1099.035 13.205 ;
        RECT 1100.110 13.160 1100.430 13.220 ;
        RECT 1098.745 13.020 1100.430 13.160 ;
        RECT 1098.745 12.975 1099.035 13.020 ;
        RECT 1100.110 12.960 1100.430 13.020 ;
      LAYER via ;
        RECT 934.080 20.780 934.340 21.040 ;
        RECT 981.920 20.780 982.180 21.040 ;
        RECT 982.380 20.780 982.640 21.040 ;
        RECT 1030.220 20.780 1030.480 21.040 ;
        RECT 1079.440 19.760 1079.700 20.020 ;
        RECT 1078.980 18.060 1079.240 18.320 ;
        RECT 1100.140 18.060 1100.400 18.320 ;
        RECT 1122.680 18.060 1122.940 18.320 ;
        RECT 1128.200 17.720 1128.460 17.980 ;
        RECT 1173.740 17.720 1174.000 17.980 ;
        RECT 630.480 17.380 630.740 17.640 ;
        RECT 498.460 17.040 498.720 17.300 ;
        RECT 519.160 17.040 519.420 17.300 ;
        RECT 569.300 17.040 569.560 17.300 ;
        RECT 934.080 17.040 934.340 17.300 ;
        RECT 981.920 17.040 982.180 17.300 ;
        RECT 982.380 17.040 982.640 17.300 ;
        RECT 1030.220 17.040 1030.480 17.300 ;
        RECT 165.880 16.700 166.140 16.960 ;
        RECT 1176.040 16.700 1176.300 16.960 ;
        RECT 1185.240 16.700 1185.500 16.960 ;
        RECT 1100.140 12.960 1100.400 13.220 ;
      LAYER met2 ;
        RECT 934.080 20.750 934.340 21.070 ;
        RECT 981.920 20.750 982.180 21.070 ;
        RECT 982.380 20.750 982.640 21.070 ;
        RECT 1030.220 20.750 1030.480 21.070 ;
        RECT 630.480 17.350 630.740 17.670 ;
        RECT 498.460 17.010 498.720 17.330 ;
        RECT 519.160 17.010 519.420 17.330 ;
        RECT 569.300 17.010 569.560 17.330 ;
        RECT 165.880 16.670 166.140 16.990 ;
        RECT 165.940 2.400 166.080 16.670 ;
        RECT 498.520 16.165 498.660 17.010 ;
        RECT 519.220 16.165 519.360 17.010 ;
        RECT 569.360 16.165 569.500 17.010 ;
        RECT 630.540 16.165 630.680 17.350 ;
        RECT 934.140 17.330 934.280 20.750 ;
        RECT 981.980 17.330 982.120 20.750 ;
        RECT 982.440 17.330 982.580 20.750 ;
        RECT 1030.280 17.330 1030.420 20.750 ;
        RECT 1079.440 19.730 1079.700 20.050 ;
        RECT 1078.980 18.260 1079.240 18.350 ;
        RECT 1079.500 18.260 1079.640 19.730 ;
        RECT 1078.980 18.120 1079.640 18.260 ;
        RECT 1078.980 18.030 1079.240 18.120 ;
        RECT 1100.140 18.030 1100.400 18.350 ;
        RECT 1122.680 18.030 1122.940 18.350 ;
        RECT 934.080 17.010 934.340 17.330 ;
        RECT 981.920 17.010 982.180 17.330 ;
        RECT 982.380 17.010 982.640 17.330 ;
        RECT 1030.220 17.010 1030.480 17.330 ;
        RECT 498.450 15.795 498.730 16.165 ;
        RECT 519.150 15.795 519.430 16.165 ;
        RECT 569.290 15.795 569.570 16.165 ;
        RECT 630.470 15.795 630.750 16.165 ;
        RECT 1100.200 13.250 1100.340 18.030 ;
        RECT 1122.740 16.165 1122.880 18.030 ;
        RECT 1128.200 17.690 1128.460 18.010 ;
        RECT 1173.740 17.690 1174.000 18.010 ;
        RECT 1128.260 16.165 1128.400 17.690 ;
        RECT 1173.800 16.165 1173.940 17.690 ;
        RECT 1185.300 16.990 1185.440 54.000 ;
        RECT 1176.040 16.670 1176.300 16.990 ;
        RECT 1185.240 16.670 1185.500 16.990 ;
        RECT 1176.100 16.165 1176.240 16.670 ;
        RECT 1122.670 15.795 1122.950 16.165 ;
        RECT 1128.190 15.795 1128.470 16.165 ;
        RECT 1173.730 15.795 1174.010 16.165 ;
        RECT 1176.030 15.795 1176.310 16.165 ;
        RECT 1100.140 12.930 1100.400 13.250 ;
        RECT 165.870 0.000 166.150 2.400 ;
      LAYER via2 ;
        RECT 498.450 15.840 498.730 16.120 ;
        RECT 519.150 15.840 519.430 16.120 ;
        RECT 569.290 15.840 569.570 16.120 ;
        RECT 630.470 15.840 630.750 16.120 ;
        RECT 1122.670 15.840 1122.950 16.120 ;
        RECT 1128.190 15.840 1128.470 16.120 ;
        RECT 1173.730 15.840 1174.010 16.120 ;
        RECT 1176.030 15.840 1176.310 16.120 ;
      LAYER met3 ;
        RECT 498.425 16.130 498.755 16.145 ;
        RECT 519.125 16.130 519.455 16.145 ;
        RECT 498.425 15.830 519.455 16.130 ;
        RECT 498.425 15.815 498.755 15.830 ;
        RECT 519.125 15.815 519.455 15.830 ;
        RECT 569.265 16.130 569.595 16.145 ;
        RECT 630.445 16.130 630.775 16.145 ;
        RECT 569.265 15.830 630.775 16.130 ;
        RECT 569.265 15.815 569.595 15.830 ;
        RECT 630.445 15.815 630.775 15.830 ;
        RECT 1122.645 16.130 1122.975 16.145 ;
        RECT 1128.165 16.130 1128.495 16.145 ;
        RECT 1122.645 15.830 1128.495 16.130 ;
        RECT 1122.645 15.815 1122.975 15.830 ;
        RECT 1128.165 15.815 1128.495 15.830 ;
        RECT 1173.705 16.130 1174.035 16.145 ;
        RECT 1176.005 16.130 1176.335 16.145 ;
        RECT 1173.705 15.830 1176.335 16.130 ;
        RECT 1173.705 15.815 1174.035 15.830 ;
        RECT 1176.005 15.815 1176.335 15.830 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 183.330 17.920 183.650 17.980 ;
        RECT 188.390 17.920 188.710 17.980 ;
        RECT 183.330 17.780 188.710 17.920 ;
        RECT 183.330 17.720 183.650 17.780 ;
        RECT 188.390 17.720 188.710 17.780 ;
      LAYER via ;
        RECT 183.360 17.720 183.620 17.980 ;
        RECT 188.420 17.720 188.680 17.980 ;
      LAYER met2 ;
        RECT 188.480 18.010 188.620 54.000 ;
        RECT 183.360 17.690 183.620 18.010 ;
        RECT 188.420 17.690 188.680 18.010 ;
        RECT 183.420 2.400 183.560 17.690 ;
        RECT 183.350 0.000 183.630 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 223.885 16.745 224.055 18.275 ;
        RECT 694.465 17.425 694.635 18.275 ;
        RECT 740.005 17.425 740.175 20.995 ;
        RECT 761.165 18.105 761.335 20.995 ;
        RECT 795.665 18.105 795.835 20.995 ;
        RECT 837.985 18.105 838.155 20.995 ;
        RECT 884.905 18.105 885.075 20.995 ;
        RECT 886.285 17.425 886.455 20.995 ;
      LAYER mcon ;
        RECT 740.005 20.825 740.175 20.995 ;
        RECT 223.885 18.105 224.055 18.275 ;
        RECT 694.465 18.105 694.635 18.275 ;
        RECT 761.165 20.825 761.335 20.995 ;
        RECT 795.665 20.825 795.835 20.995 ;
        RECT 837.985 20.825 838.155 20.995 ;
        RECT 884.905 20.825 885.075 20.995 ;
        RECT 886.285 20.825 886.455 20.995 ;
      LAYER met1 ;
        RECT 739.945 20.980 740.235 21.025 ;
        RECT 761.105 20.980 761.395 21.025 ;
        RECT 739.945 20.840 761.395 20.980 ;
        RECT 739.945 20.795 740.235 20.840 ;
        RECT 761.105 20.795 761.395 20.840 ;
        RECT 795.605 20.980 795.895 21.025 ;
        RECT 837.925 20.980 838.215 21.025 ;
        RECT 795.605 20.840 838.215 20.980 ;
        RECT 795.605 20.795 795.895 20.840 ;
        RECT 837.925 20.795 838.215 20.840 ;
        RECT 884.845 20.980 885.135 21.025 ;
        RECT 886.225 20.980 886.515 21.025 ;
        RECT 884.845 20.840 886.515 20.980 ;
        RECT 884.845 20.795 885.135 20.840 ;
        RECT 886.225 20.795 886.515 20.840 ;
        RECT 1178.310 20.300 1178.630 20.360 ;
        RECT 1189.810 20.300 1190.130 20.360 ;
        RECT 1178.310 20.160 1190.130 20.300 ;
        RECT 1178.310 20.100 1178.630 20.160 ;
        RECT 1189.810 20.100 1190.130 20.160 ;
        RECT 223.825 18.260 224.115 18.305 ;
        RECT 694.405 18.260 694.695 18.305 ;
        RECT 223.825 18.120 694.695 18.260 ;
        RECT 223.825 18.075 224.115 18.120 ;
        RECT 694.405 18.075 694.695 18.120 ;
        RECT 761.105 18.260 761.395 18.305 ;
        RECT 795.605 18.260 795.895 18.305 ;
        RECT 761.105 18.120 795.895 18.260 ;
        RECT 761.105 18.075 761.395 18.120 ;
        RECT 795.605 18.075 795.895 18.120 ;
        RECT 837.925 18.260 838.215 18.305 ;
        RECT 884.845 18.260 885.135 18.305 ;
        RECT 1051.350 18.260 1051.670 18.320 ;
        RECT 837.925 18.120 885.135 18.260 ;
        RECT 837.925 18.075 838.215 18.120 ;
        RECT 884.845 18.075 885.135 18.120 ;
        RECT 906.540 18.120 1051.670 18.260 ;
        RECT 694.405 17.580 694.695 17.625 ;
        RECT 739.945 17.580 740.235 17.625 ;
        RECT 694.405 17.440 740.235 17.580 ;
        RECT 694.405 17.395 694.695 17.440 ;
        RECT 739.945 17.395 740.235 17.440 ;
        RECT 886.225 17.580 886.515 17.625 ;
        RECT 906.540 17.580 906.680 18.120 ;
        RECT 1051.350 18.060 1051.670 18.120 ;
        RECT 1125.870 18.260 1126.190 18.320 ;
        RECT 1127.250 18.260 1127.570 18.320 ;
        RECT 1125.870 18.120 1127.570 18.260 ;
        RECT 1125.870 18.060 1126.190 18.120 ;
        RECT 1127.250 18.060 1127.570 18.120 ;
        RECT 886.225 17.440 906.680 17.580 ;
        RECT 886.225 17.395 886.515 17.440 ;
        RECT 201.270 16.900 201.590 16.960 ;
        RECT 223.825 16.900 224.115 16.945 ;
        RECT 201.270 16.760 224.115 16.900 ;
        RECT 201.270 16.700 201.590 16.760 ;
        RECT 223.825 16.715 224.115 16.760 ;
      LAYER via ;
        RECT 1178.340 20.100 1178.600 20.360 ;
        RECT 1189.840 20.100 1190.100 20.360 ;
        RECT 1051.380 18.060 1051.640 18.320 ;
        RECT 1125.900 18.060 1126.160 18.320 ;
        RECT 1127.280 18.060 1127.540 18.320 ;
        RECT 201.300 16.700 201.560 16.960 ;
      LAYER met2 ;
        RECT 1127.270 21.235 1127.550 21.605 ;
        RECT 1178.330 21.235 1178.610 21.605 ;
        RECT 1127.340 18.350 1127.480 21.235 ;
        RECT 1178.400 20.390 1178.540 21.235 ;
        RECT 1189.900 20.390 1190.040 54.000 ;
        RECT 1178.340 20.070 1178.600 20.390 ;
        RECT 1189.840 20.070 1190.100 20.390 ;
        RECT 1051.380 18.030 1051.640 18.350 ;
        RECT 1125.900 18.030 1126.160 18.350 ;
        RECT 1127.280 18.030 1127.540 18.350 ;
        RECT 201.300 16.670 201.560 16.990 ;
        RECT 201.360 2.400 201.500 16.670 ;
        RECT 1051.440 15.485 1051.580 18.030 ;
        RECT 1125.960 15.485 1126.100 18.030 ;
        RECT 1051.370 15.115 1051.650 15.485 ;
        RECT 1125.890 15.115 1126.170 15.485 ;
        RECT 201.290 0.000 201.570 2.400 ;
      LAYER via2 ;
        RECT 1127.270 21.280 1127.550 21.560 ;
        RECT 1178.330 21.280 1178.610 21.560 ;
        RECT 1051.370 15.160 1051.650 15.440 ;
        RECT 1125.890 15.160 1126.170 15.440 ;
      LAYER met3 ;
        RECT 1127.245 21.570 1127.575 21.585 ;
        RECT 1178.305 21.570 1178.635 21.585 ;
        RECT 1127.245 21.270 1178.635 21.570 ;
        RECT 1127.245 21.255 1127.575 21.270 ;
        RECT 1178.305 21.255 1178.635 21.270 ;
        RECT 1051.345 15.450 1051.675 15.465 ;
        RECT 1125.865 15.450 1126.195 15.465 ;
        RECT 1051.345 15.150 1126.195 15.450 ;
        RECT 1051.345 15.135 1051.675 15.150 ;
        RECT 1125.865 15.135 1126.195 15.150 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 219.210 17.920 219.530 17.980 ;
        RECT 222.890 17.920 223.210 17.980 ;
        RECT 219.210 17.780 223.210 17.920 ;
        RECT 219.210 17.720 219.530 17.780 ;
        RECT 222.890 17.720 223.210 17.780 ;
      LAYER via ;
        RECT 219.240 17.720 219.500 17.980 ;
        RECT 222.920 17.720 223.180 17.980 ;
      LAYER met2 ;
        RECT 222.980 18.010 223.120 54.000 ;
        RECT 219.240 17.690 219.500 18.010 ;
        RECT 222.920 17.690 223.180 18.010 ;
        RECT 219.300 2.400 219.440 17.690 ;
        RECT 219.230 0.000 219.510 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 665.025 19.805 665.195 20.995 ;
        RECT 671.465 19.805 671.635 20.995 ;
        RECT 694.005 17.425 694.175 21.335 ;
        RECT 788.765 17.425 788.935 21.335 ;
        RECT 789.225 17.425 789.395 21.335 ;
        RECT 933.665 17.425 933.835 20.995 ;
        RECT 1030.725 17.425 1030.895 21.335 ;
        RECT 1079.485 18.105 1079.655 21.335 ;
        RECT 1099.725 18.105 1099.895 19.975 ;
      LAYER mcon ;
        RECT 694.005 21.165 694.175 21.335 ;
        RECT 665.025 20.825 665.195 20.995 ;
        RECT 671.465 20.825 671.635 20.995 ;
        RECT 788.765 21.165 788.935 21.335 ;
        RECT 789.225 21.165 789.395 21.335 ;
        RECT 1030.725 21.165 1030.895 21.335 ;
        RECT 933.665 20.825 933.835 20.995 ;
        RECT 1079.485 21.165 1079.655 21.335 ;
        RECT 1099.725 19.805 1099.895 19.975 ;
      LAYER met1 ;
        RECT 693.945 21.320 694.235 21.365 ;
        RECT 788.705 21.320 788.995 21.365 ;
        RECT 693.945 21.180 788.995 21.320 ;
        RECT 693.945 21.135 694.235 21.180 ;
        RECT 788.705 21.135 788.995 21.180 ;
        RECT 789.165 21.320 789.455 21.365 ;
        RECT 1030.665 21.320 1030.955 21.365 ;
        RECT 1079.425 21.320 1079.715 21.365 ;
        RECT 789.165 21.180 886.900 21.320 ;
        RECT 789.165 21.135 789.455 21.180 ;
        RECT 664.965 20.980 665.255 21.025 ;
        RECT 671.405 20.980 671.695 21.025 ;
        RECT 664.965 20.840 671.695 20.980 ;
        RECT 886.760 20.980 886.900 21.180 ;
        RECT 1030.665 21.180 1079.715 21.320 ;
        RECT 1030.665 21.135 1030.955 21.180 ;
        RECT 1079.425 21.135 1079.715 21.180 ;
        RECT 933.605 20.980 933.895 21.025 ;
        RECT 886.760 20.840 933.895 20.980 ;
        RECT 664.965 20.795 665.255 20.840 ;
        RECT 671.405 20.795 671.695 20.840 ;
        RECT 933.605 20.795 933.895 20.840 ;
        RECT 1151.260 20.160 1178.080 20.300 ;
        RECT 237.150 19.960 237.470 20.020 ;
        RECT 664.965 19.960 665.255 20.005 ;
        RECT 237.150 19.820 665.255 19.960 ;
        RECT 237.150 19.760 237.470 19.820 ;
        RECT 664.965 19.775 665.255 19.820 ;
        RECT 671.405 19.960 671.695 20.005 ;
        RECT 688.410 19.960 688.730 20.020 ;
        RECT 671.405 19.820 688.730 19.960 ;
        RECT 671.405 19.775 671.695 19.820 ;
        RECT 688.410 19.760 688.730 19.820 ;
        RECT 1099.665 19.960 1099.955 20.005 ;
        RECT 1151.260 19.960 1151.400 20.160 ;
        RECT 1099.665 19.820 1151.400 19.960 ;
        RECT 1177.940 19.960 1178.080 20.160 ;
        RECT 1196.710 19.960 1197.030 20.020 ;
        RECT 1177.940 19.820 1197.030 19.960 ;
        RECT 1099.665 19.775 1099.955 19.820 ;
        RECT 1196.710 19.760 1197.030 19.820 ;
        RECT 1079.425 18.260 1079.715 18.305 ;
        RECT 1099.665 18.260 1099.955 18.305 ;
        RECT 1079.425 18.120 1099.955 18.260 ;
        RECT 1079.425 18.075 1079.715 18.120 ;
        RECT 1099.665 18.075 1099.955 18.120 ;
        RECT 692.090 17.580 692.410 17.640 ;
        RECT 693.945 17.580 694.235 17.625 ;
        RECT 692.090 17.440 694.235 17.580 ;
        RECT 692.090 17.380 692.410 17.440 ;
        RECT 693.945 17.395 694.235 17.440 ;
        RECT 788.705 17.580 788.995 17.625 ;
        RECT 789.165 17.580 789.455 17.625 ;
        RECT 788.705 17.440 789.455 17.580 ;
        RECT 788.705 17.395 788.995 17.440 ;
        RECT 789.165 17.395 789.455 17.440 ;
        RECT 933.605 17.580 933.895 17.625 ;
        RECT 1030.665 17.580 1030.955 17.625 ;
        RECT 933.605 17.440 1030.955 17.580 ;
        RECT 933.605 17.395 933.895 17.440 ;
        RECT 1030.665 17.395 1030.955 17.440 ;
      LAYER via ;
        RECT 237.180 19.760 237.440 20.020 ;
        RECT 688.440 19.760 688.700 20.020 ;
        RECT 1196.740 19.760 1197.000 20.020 ;
        RECT 692.120 17.380 692.380 17.640 ;
      LAYER met2 ;
        RECT 688.500 20.670 689.560 20.810 ;
        RECT 688.500 20.050 688.640 20.670 ;
        RECT 237.180 19.730 237.440 20.050 ;
        RECT 688.440 19.730 688.700 20.050 ;
        RECT 237.240 2.400 237.380 19.730 ;
        RECT 689.420 17.580 689.560 20.670 ;
        RECT 1196.800 20.050 1196.940 54.000 ;
        RECT 1196.740 19.730 1197.000 20.050 ;
        RECT 692.120 17.580 692.380 17.670 ;
        RECT 689.420 17.440 692.380 17.580 ;
        RECT 692.120 17.350 692.380 17.440 ;
        RECT 237.170 0.000 237.450 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 58.670 17.580 58.990 17.640 ;
        RECT 64.190 17.580 64.510 17.640 ;
        RECT 58.670 17.440 64.510 17.580 ;
        RECT 58.670 17.380 58.990 17.440 ;
        RECT 64.190 17.380 64.510 17.440 ;
      LAYER via ;
        RECT 58.700 17.380 58.960 17.640 ;
        RECT 64.220 17.380 64.480 17.640 ;
      LAYER met2 ;
        RECT 64.280 17.670 64.420 54.000 ;
        RECT 58.700 17.350 58.960 17.670 ;
        RECT 64.220 17.350 64.480 17.670 ;
        RECT 58.760 2.400 58.900 17.350 ;
        RECT 58.690 0.000 58.970 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1165.060 45.290 1165.200 54.000 ;
        RECT 1164.600 45.150 1165.200 45.290 ;
        RECT 82.610 17.835 82.890 18.205 ;
        RECT 82.680 2.400 82.820 17.835 ;
        RECT 1164.600 17.525 1164.740 45.150 ;
        RECT 1164.530 17.155 1164.810 17.525 ;
        RECT 82.610 0.000 82.890 2.400 ;
      LAYER via2 ;
        RECT 82.610 17.880 82.890 18.160 ;
        RECT 1164.530 17.200 1164.810 17.480 ;
      LAYER met3 ;
        RECT 82.585 18.170 82.915 18.185 ;
        RECT 82.585 17.870 1140.210 18.170 ;
        RECT 82.585 17.855 82.915 17.870 ;
        RECT 1139.910 17.490 1140.210 17.870 ;
        RECT 1164.505 17.490 1164.835 17.505 ;
        RECT 1139.910 17.190 1164.835 17.490 ;
        RECT 1164.505 17.175 1164.835 17.190 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 106.050 15.540 106.370 15.600 ;
        RECT 112.490 15.540 112.810 15.600 ;
        RECT 106.050 15.400 112.810 15.540 ;
        RECT 106.050 15.340 106.370 15.400 ;
        RECT 112.490 15.340 112.810 15.400 ;
      LAYER via ;
        RECT 106.080 15.340 106.340 15.600 ;
        RECT 112.520 15.340 112.780 15.600 ;
      LAYER met2 ;
        RECT 112.580 15.630 112.720 54.000 ;
        RECT 106.080 15.310 106.340 15.630 ;
        RECT 112.520 15.310 112.780 15.630 ;
        RECT 106.140 2.400 106.280 15.310 ;
        RECT 106.070 0.000 106.350 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1176.100 53.960 1176.240 54.000 ;
        RECT 1176.100 53.820 1176.700 53.960 ;
        RECT 1176.560 21.490 1176.700 53.820 ;
        RECT 1176.100 21.350 1176.700 21.490 ;
        RECT 1176.100 19.565 1176.240 21.350 ;
        RECT 129.990 19.195 130.270 19.565 ;
        RECT 1176.030 19.195 1176.310 19.565 ;
        RECT 130.060 2.400 130.200 19.195 ;
        RECT 129.990 0.000 130.270 2.400 ;
      LAYER via2 ;
        RECT 129.990 19.240 130.270 19.520 ;
        RECT 1176.030 19.240 1176.310 19.520 ;
      LAYER met3 ;
        RECT 129.965 19.530 130.295 19.545 ;
        RECT 1176.005 19.530 1176.335 19.545 ;
        RECT 129.965 19.230 1176.335 19.530 ;
        RECT 129.965 19.215 130.295 19.230 ;
        RECT 1176.005 19.215 1176.335 19.230 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 28.770 2.960 29.090 3.020 ;
        RECT 29.690 2.960 30.010 3.020 ;
        RECT 28.770 2.820 30.010 2.960 ;
        RECT 28.770 2.760 29.090 2.820 ;
        RECT 29.690 2.760 30.010 2.820 ;
      LAYER via ;
        RECT 28.800 2.760 29.060 3.020 ;
        RECT 29.720 2.760 29.980 3.020 ;
      LAYER met2 ;
        RECT 29.710 1686.555 29.990 1686.925 ;
        RECT 29.780 3.050 29.920 1686.555 ;
        RECT 28.800 2.730 29.060 3.050 ;
        RECT 29.720 2.730 29.980 3.050 ;
        RECT 28.860 2.400 29.000 2.730 ;
        RECT 28.790 0.000 29.070 2.400 ;
      LAYER via2 ;
        RECT 29.710 1686.600 29.990 1686.880 ;
      LAYER met3 ;
        RECT 29.685 1686.890 30.015 1686.905 ;
        RECT 29.685 1686.590 54.000 1686.890 ;
        RECT 29.685 1686.575 30.015 1686.590 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1157.700 30.445 1157.840 54.000 ;
        RECT 1157.630 30.075 1157.910 30.445 ;
        RECT 34.770 16.475 35.050 16.845 ;
        RECT 290.990 16.475 291.270 16.845 ;
        RECT 291.910 16.475 292.190 16.845 ;
        RECT 740.870 16.475 741.150 16.845 ;
        RECT 1040.790 16.475 1041.070 16.845 ;
        RECT 34.840 2.400 34.980 16.475 ;
        RECT 291.060 16.050 291.200 16.475 ;
        RECT 291.980 16.050 292.120 16.475 ;
        RECT 291.060 15.910 292.120 16.050 ;
        RECT 740.410 15.370 740.690 15.485 ;
        RECT 740.940 15.370 741.080 16.475 ;
        RECT 740.410 15.230 741.080 15.370 ;
        RECT 740.410 15.115 740.690 15.230 ;
        RECT 1040.860 12.765 1041.000 16.475 ;
        RECT 1040.790 12.395 1041.070 12.765 ;
        RECT 34.770 0.000 35.050 2.400 ;
      LAYER via2 ;
        RECT 1157.630 30.120 1157.910 30.400 ;
        RECT 34.770 16.520 35.050 16.800 ;
        RECT 290.990 16.520 291.270 16.800 ;
        RECT 291.910 16.520 292.190 16.800 ;
        RECT 740.870 16.520 741.150 16.800 ;
        RECT 1040.790 16.520 1041.070 16.800 ;
        RECT 740.410 15.160 740.690 15.440 ;
        RECT 1040.790 12.440 1041.070 12.720 ;
      LAYER met3 ;
        RECT 1113.190 30.410 1113.570 30.420 ;
        RECT 1157.605 30.410 1157.935 30.425 ;
        RECT 1113.190 30.110 1157.935 30.410 ;
        RECT 1113.190 30.100 1113.570 30.110 ;
        RECT 1157.605 30.095 1157.935 30.110 ;
        RECT 34.745 16.810 35.075 16.825 ;
        RECT 290.965 16.810 291.295 16.825 ;
        RECT 34.745 16.510 291.295 16.810 ;
        RECT 34.745 16.495 35.075 16.510 ;
        RECT 290.965 16.495 291.295 16.510 ;
        RECT 291.885 16.810 292.215 16.825 ;
        RECT 726.790 16.810 727.170 16.820 ;
        RECT 291.885 16.510 727.170 16.810 ;
        RECT 291.885 16.495 292.215 16.510 ;
        RECT 726.790 16.500 727.170 16.510 ;
        RECT 740.845 16.810 741.175 16.825 ;
        RECT 1040.765 16.810 1041.095 16.825 ;
        RECT 740.845 16.510 1041.095 16.810 ;
        RECT 740.845 16.495 741.175 16.510 ;
        RECT 1040.765 16.495 1041.095 16.510 ;
        RECT 726.790 15.450 727.170 15.460 ;
        RECT 740.385 15.450 740.715 15.465 ;
        RECT 726.790 15.150 740.715 15.450 ;
        RECT 726.790 15.140 727.170 15.150 ;
        RECT 740.385 15.135 740.715 15.150 ;
        RECT 1113.190 14.090 1113.570 14.100 ;
        RECT 1064.470 13.790 1113.570 14.090 ;
        RECT 1040.765 12.730 1041.095 12.745 ;
        RECT 1064.470 12.730 1064.770 13.790 ;
        RECT 1113.190 13.780 1113.570 13.790 ;
        RECT 1040.765 12.430 1064.770 12.730 ;
        RECT 1040.765 12.415 1041.095 12.430 ;
      LAYER via3 ;
        RECT 1113.220 30.100 1113.540 30.420 ;
        RECT 726.820 16.500 727.140 16.820 ;
        RECT 726.820 15.140 727.140 15.460 ;
        RECT 1113.220 13.780 1113.540 14.100 ;
      LAYER met4 ;
        RECT 1113.215 30.095 1113.545 30.425 ;
        RECT 726.815 16.495 727.145 16.825 ;
        RECT 726.830 15.465 727.130 16.495 ;
        RECT 726.815 15.135 727.145 15.465 ;
        RECT 1113.230 14.105 1113.530 30.095 ;
        RECT 1113.215 13.775 1113.545 14.105 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 4.000 6.880 6.000 3512.800 ;
        RECT 2918.580 6.880 2920.580 3512.800 ;
      LAYER via4 ;
        RECT 4.410 3511.210 5.590 3512.390 ;
        RECT 4.410 3396.900 5.590 3398.080 ;
        RECT 4.410 3243.720 5.590 3244.900 ;
        RECT 4.410 3090.540 5.590 3091.720 ;
        RECT 4.410 2937.360 5.590 2938.540 ;
        RECT 4.410 2784.180 5.590 2785.360 ;
        RECT 4.410 2631.000 5.590 2632.180 ;
        RECT 4.410 2477.820 5.590 2479.000 ;
        RECT 4.410 2324.640 5.590 2325.820 ;
        RECT 4.410 2171.460 5.590 2172.640 ;
        RECT 4.410 2018.280 5.590 2019.460 ;
        RECT 4.410 1865.100 5.590 1866.280 ;
        RECT 4.410 1711.920 5.590 1713.100 ;
        RECT 4.410 1558.740 5.590 1559.920 ;
        RECT 4.410 1405.560 5.590 1406.740 ;
        RECT 4.410 1252.380 5.590 1253.560 ;
        RECT 4.410 1099.200 5.590 1100.380 ;
        RECT 4.410 946.020 5.590 947.200 ;
        RECT 4.410 792.840 5.590 794.020 ;
        RECT 4.410 639.660 5.590 640.840 ;
        RECT 4.410 486.480 5.590 487.660 ;
        RECT 4.410 333.300 5.590 334.480 ;
        RECT 4.410 180.120 5.590 181.300 ;
        RECT 4.410 26.940 5.590 28.120 ;
        RECT 4.410 7.290 5.590 8.470 ;
        RECT 2918.990 3511.210 2920.170 3512.390 ;
        RECT 2918.990 3396.900 2920.170 3398.080 ;
        RECT 2918.990 3243.720 2920.170 3244.900 ;
        RECT 2918.990 3090.540 2920.170 3091.720 ;
        RECT 2918.990 2937.360 2920.170 2938.540 ;
        RECT 2918.990 2784.180 2920.170 2785.360 ;
        RECT 2918.990 2631.000 2920.170 2632.180 ;
        RECT 2918.990 2477.820 2920.170 2479.000 ;
        RECT 2918.990 2324.640 2920.170 2325.820 ;
        RECT 2918.990 2171.460 2920.170 2172.640 ;
        RECT 2918.990 2018.280 2920.170 2019.460 ;
        RECT 2918.990 1865.100 2920.170 1866.280 ;
        RECT 2918.990 1711.920 2920.170 1713.100 ;
        RECT 2918.990 1558.740 2920.170 1559.920 ;
        RECT 2918.990 1405.560 2920.170 1406.740 ;
        RECT 2918.990 1252.380 2920.170 1253.560 ;
        RECT 2918.990 1099.200 2920.170 1100.380 ;
        RECT 2918.990 946.020 2920.170 947.200 ;
        RECT 2918.990 792.840 2920.170 794.020 ;
        RECT 2918.990 639.660 2920.170 640.840 ;
        RECT 2918.990 486.480 2920.170 487.660 ;
        RECT 2918.990 333.300 2920.170 334.480 ;
        RECT 2918.990 180.120 2920.170 181.300 ;
        RECT 2918.990 26.940 2920.170 28.120 ;
        RECT 2918.990 7.290 2920.170 8.470 ;
      LAYER met5 ;
        RECT 4.000 3510.800 2920.580 3512.800 ;
        RECT 0.000 3396.690 54.000 3398.290 ;
        RECT 2870.580 3396.690 2924.580 3398.290 ;
        RECT 0.000 3243.510 54.000 3245.110 ;
        RECT 2870.580 3243.510 2924.580 3245.110 ;
        RECT 0.000 3090.330 54.000 3091.930 ;
        RECT 2870.580 3090.330 2924.580 3091.930 ;
        RECT 0.000 2937.150 54.000 2938.750 ;
        RECT 2870.580 2937.150 2924.580 2938.750 ;
        RECT 0.000 2783.970 54.000 2785.570 ;
        RECT 2870.580 2783.970 2924.580 2785.570 ;
        RECT 0.000 2630.790 54.000 2632.390 ;
        RECT 2870.580 2630.790 2924.580 2632.390 ;
        RECT 0.000 2477.610 54.000 2479.210 ;
        RECT 2870.580 2477.610 2924.580 2479.210 ;
        RECT 0.000 2324.430 54.000 2326.030 ;
        RECT 2870.580 2324.430 2924.580 2326.030 ;
        RECT 0.000 2171.250 54.000 2172.850 ;
        RECT 2870.580 2171.250 2924.580 2172.850 ;
        RECT 0.000 2018.070 54.000 2019.670 ;
        RECT 2870.580 2018.070 2924.580 2019.670 ;
        RECT 0.000 1864.890 54.000 1866.490 ;
        RECT 2870.580 1864.890 2924.580 1866.490 ;
        RECT 0.000 1711.710 54.000 1713.310 ;
        RECT 2870.580 1711.710 2924.580 1713.310 ;
        RECT 0.000 1558.530 54.000 1560.130 ;
        RECT 2870.580 1558.530 2924.580 1560.130 ;
        RECT 0.000 1405.350 54.000 1406.950 ;
        RECT 2870.580 1405.350 2924.580 1406.950 ;
        RECT 0.000 1252.170 54.000 1253.770 ;
        RECT 2870.580 1252.170 2924.580 1253.770 ;
        RECT 0.000 1098.990 54.000 1100.590 ;
        RECT 2870.580 1098.990 2924.580 1100.590 ;
        RECT 0.000 945.810 54.000 947.410 ;
        RECT 2870.580 945.810 2924.580 947.410 ;
        RECT 0.000 792.630 54.000 794.230 ;
        RECT 2870.580 792.630 2924.580 794.230 ;
        RECT 0.000 639.450 54.000 641.050 ;
        RECT 2870.580 639.450 2924.580 641.050 ;
        RECT 0.000 486.270 54.000 487.870 ;
        RECT 2870.580 486.270 2924.580 487.870 ;
        RECT 0.000 333.090 54.000 334.690 ;
        RECT 2870.580 333.090 2924.580 334.690 ;
        RECT 0.000 179.910 54.000 181.510 ;
        RECT 2870.580 179.910 2924.580 181.510 ;
        RECT 0.000 26.730 2924.580 28.330 ;
        RECT 4.000 6.880 2920.580 8.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 0.000 2.880 2.000 3516.800 ;
        RECT 2922.580 2.880 2924.580 3516.800 ;
      LAYER via4 ;
        RECT 0.410 3515.210 1.590 3516.390 ;
        RECT 0.410 3473.490 1.590 3474.670 ;
        RECT 0.410 3320.310 1.590 3321.490 ;
        RECT 0.410 3167.130 1.590 3168.310 ;
        RECT 0.410 3013.950 1.590 3015.130 ;
        RECT 0.410 2860.770 1.590 2861.950 ;
        RECT 0.410 2707.590 1.590 2708.770 ;
        RECT 0.410 2554.410 1.590 2555.590 ;
        RECT 0.410 2401.230 1.590 2402.410 ;
        RECT 0.410 2248.050 1.590 2249.230 ;
        RECT 0.410 2094.870 1.590 2096.050 ;
        RECT 0.410 1941.690 1.590 1942.870 ;
        RECT 0.410 1788.510 1.590 1789.690 ;
        RECT 0.410 1635.330 1.590 1636.510 ;
        RECT 0.410 1482.150 1.590 1483.330 ;
        RECT 0.410 1328.970 1.590 1330.150 ;
        RECT 0.410 1175.790 1.590 1176.970 ;
        RECT 0.410 1022.610 1.590 1023.790 ;
        RECT 0.410 869.430 1.590 870.610 ;
        RECT 0.410 716.250 1.590 717.430 ;
        RECT 0.410 563.070 1.590 564.250 ;
        RECT 0.410 409.890 1.590 411.070 ;
        RECT 0.410 256.710 1.590 257.890 ;
        RECT 0.410 103.530 1.590 104.710 ;
        RECT 0.410 3.290 1.590 4.470 ;
        RECT 2922.990 3515.210 2924.170 3516.390 ;
        RECT 2922.990 3473.490 2924.170 3474.670 ;
        RECT 2922.990 3320.310 2924.170 3321.490 ;
        RECT 2922.990 3167.130 2924.170 3168.310 ;
        RECT 2922.990 3013.950 2924.170 3015.130 ;
        RECT 2922.990 2860.770 2924.170 2861.950 ;
        RECT 2922.990 2707.590 2924.170 2708.770 ;
        RECT 2922.990 2554.410 2924.170 2555.590 ;
        RECT 2922.990 2401.230 2924.170 2402.410 ;
        RECT 2922.990 2248.050 2924.170 2249.230 ;
        RECT 2922.990 2094.870 2924.170 2096.050 ;
        RECT 2922.990 1941.690 2924.170 1942.870 ;
        RECT 2922.990 1788.510 2924.170 1789.690 ;
        RECT 2922.990 1635.330 2924.170 1636.510 ;
        RECT 2922.990 1482.150 2924.170 1483.330 ;
        RECT 2922.990 1328.970 2924.170 1330.150 ;
        RECT 2922.990 1175.790 2924.170 1176.970 ;
        RECT 2922.990 1022.610 2924.170 1023.790 ;
        RECT 2922.990 869.430 2924.170 870.610 ;
        RECT 2922.990 716.250 2924.170 717.430 ;
        RECT 2922.990 563.070 2924.170 564.250 ;
        RECT 2922.990 409.890 2924.170 411.070 ;
        RECT 2922.990 256.710 2924.170 257.890 ;
        RECT 2922.990 103.530 2924.170 104.710 ;
        RECT 2922.990 3.290 2924.170 4.470 ;
      LAYER met5 ;
        RECT 0.000 3514.800 2924.580 3516.800 ;
        RECT 0.000 3473.280 2924.580 3474.880 ;
        RECT 0.000 3320.100 54.000 3321.700 ;
        RECT 2870.580 3320.100 2924.580 3321.700 ;
        RECT 0.000 3166.920 54.000 3168.520 ;
        RECT 2870.580 3166.920 2924.580 3168.520 ;
        RECT 0.000 3013.740 54.000 3015.340 ;
        RECT 2870.580 3013.740 2924.580 3015.340 ;
        RECT 0.000 2860.560 54.000 2862.160 ;
        RECT 2870.580 2860.560 2924.580 2862.160 ;
        RECT 0.000 2707.380 54.000 2708.980 ;
        RECT 2870.580 2707.380 2924.580 2708.980 ;
        RECT 0.000 2554.200 54.000 2555.800 ;
        RECT 2870.580 2554.200 2924.580 2555.800 ;
        RECT 0.000 2401.020 54.000 2402.620 ;
        RECT 2870.580 2401.020 2924.580 2402.620 ;
        RECT 0.000 2247.840 54.000 2249.440 ;
        RECT 2870.580 2247.840 2924.580 2249.440 ;
        RECT 0.000 2094.660 54.000 2096.260 ;
        RECT 2870.580 2094.660 2924.580 2096.260 ;
        RECT 0.000 1941.480 54.000 1943.080 ;
        RECT 2870.580 1941.480 2924.580 1943.080 ;
        RECT 0.000 1788.300 54.000 1789.900 ;
        RECT 2870.580 1788.300 2924.580 1789.900 ;
        RECT 0.000 1635.120 54.000 1636.720 ;
        RECT 2870.580 1635.120 2924.580 1636.720 ;
        RECT 0.000 1481.940 54.000 1483.540 ;
        RECT 2870.580 1481.940 2924.580 1483.540 ;
        RECT 0.000 1328.760 54.000 1330.360 ;
        RECT 2870.580 1328.760 2924.580 1330.360 ;
        RECT 0.000 1175.580 54.000 1177.180 ;
        RECT 2870.580 1175.580 2924.580 1177.180 ;
        RECT 0.000 1022.400 54.000 1024.000 ;
        RECT 2870.580 1022.400 2924.580 1024.000 ;
        RECT 0.000 869.220 54.000 870.820 ;
        RECT 2870.580 869.220 2924.580 870.820 ;
        RECT 0.000 716.040 54.000 717.640 ;
        RECT 2870.580 716.040 2924.580 717.640 ;
        RECT 0.000 562.860 54.000 564.460 ;
        RECT 2870.580 562.860 2924.580 564.460 ;
        RECT 0.000 409.680 54.000 411.280 ;
        RECT 2870.580 409.680 2924.580 411.280 ;
        RECT 0.000 256.500 54.000 258.100 ;
        RECT 2870.580 256.500 2924.580 258.100 ;
        RECT 0.000 103.320 54.000 104.920 ;
        RECT 2870.580 103.320 2924.580 104.920 ;
        RECT 0.000 2.880 2924.580 4.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 84.965 54.000 2868.135 3466.000 ;
      LAYER met1 ;
        RECT 8.000 3508.560 2916.580 3509.040 ;
        RECT 8.000 3505.840 2916.580 3506.320 ;
        RECT 8.000 3503.120 2916.580 3503.600 ;
        RECT 8.000 3500.400 2916.580 3500.880 ;
        RECT 8.000 3497.680 2916.580 3498.160 ;
        RECT 8.000 3494.960 2916.580 3495.440 ;
        RECT 8.000 3492.240 2916.580 3492.720 ;
        RECT 8.000 3489.520 2916.580 3490.000 ;
        RECT 8.000 3486.800 2916.580 3487.280 ;
        RECT 8.000 3484.080 2916.580 3484.560 ;
        RECT 8.000 3481.360 2916.580 3481.840 ;
        RECT 8.000 3478.640 2916.580 3479.120 ;
        RECT 8.000 3475.920 2916.580 3476.400 ;
        RECT 8.000 3473.200 2916.580 3473.680 ;
        RECT 8.000 3470.480 2916.580 3470.960 ;
        RECT 8.000 3467.760 2916.580 3468.240 ;
        RECT 54.000 3465.520 2870.580 3466.000 ;
        RECT 8.000 3465.040 2916.580 3465.520 ;
        RECT 54.000 3462.800 2870.580 3465.040 ;
        RECT 8.000 3462.320 2916.580 3462.800 ;
        RECT 54.000 3460.080 2870.580 3462.320 ;
        RECT 8.000 3459.600 2916.580 3460.080 ;
        RECT 54.000 3457.360 2870.580 3459.600 ;
        RECT 8.000 3456.880 2916.580 3457.360 ;
        RECT 54.000 3454.640 2870.580 3456.880 ;
        RECT 8.000 3454.160 2916.580 3454.640 ;
        RECT 54.000 3451.920 2870.580 3454.160 ;
        RECT 8.000 3451.440 2916.580 3451.920 ;
        RECT 54.000 3449.200 2870.580 3451.440 ;
        RECT 8.000 3448.720 2916.580 3449.200 ;
        RECT 54.000 3446.480 2870.580 3448.720 ;
        RECT 8.000 3446.000 2916.580 3446.480 ;
        RECT 54.000 3443.760 2870.580 3446.000 ;
        RECT 8.000 3443.280 2916.580 3443.760 ;
        RECT 54.000 3441.040 2870.580 3443.280 ;
        RECT 8.000 3440.560 2916.580 3441.040 ;
        RECT 54.000 3438.320 2870.580 3440.560 ;
        RECT 8.000 3437.840 2916.580 3438.320 ;
        RECT 54.000 3435.600 2870.580 3437.840 ;
        RECT 8.000 3435.120 2916.580 3435.600 ;
        RECT 54.000 3432.880 2870.580 3435.120 ;
        RECT 8.000 3432.400 2916.580 3432.880 ;
        RECT 54.000 3430.160 2870.580 3432.400 ;
        RECT 8.000 3429.680 2916.580 3430.160 ;
        RECT 54.000 3427.440 2870.580 3429.680 ;
        RECT 8.000 3426.960 2916.580 3427.440 ;
        RECT 54.000 3424.720 2870.580 3426.960 ;
        RECT 8.000 3424.240 2916.580 3424.720 ;
        RECT 54.000 3422.000 2870.580 3424.240 ;
        RECT 8.000 3421.520 2916.580 3422.000 ;
        RECT 54.000 3419.280 2870.580 3421.520 ;
        RECT 8.000 3418.800 2916.580 3419.280 ;
        RECT 54.000 3416.560 2870.580 3418.800 ;
        RECT 8.000 3416.080 2916.580 3416.560 ;
        RECT 54.000 3413.840 2870.580 3416.080 ;
        RECT 8.000 3413.360 2916.580 3413.840 ;
        RECT 54.000 3411.120 2870.580 3413.360 ;
        RECT 8.000 3410.640 2916.580 3411.120 ;
        RECT 54.000 3408.400 2870.580 3410.640 ;
        RECT 8.000 3407.920 2916.580 3408.400 ;
        RECT 54.000 3405.680 2870.580 3407.920 ;
        RECT 8.000 3405.200 2916.580 3405.680 ;
        RECT 54.000 3402.960 2870.580 3405.200 ;
        RECT 8.000 3402.480 2916.580 3402.960 ;
        RECT 54.000 3400.240 2870.580 3402.480 ;
        RECT 8.000 3399.760 2916.580 3400.240 ;
        RECT 54.000 3397.520 2870.580 3399.760 ;
        RECT 8.000 3397.040 2916.580 3397.520 ;
        RECT 54.000 3394.800 2870.580 3397.040 ;
        RECT 8.000 3394.320 2916.580 3394.800 ;
        RECT 54.000 3392.080 2870.580 3394.320 ;
        RECT 8.000 3391.600 2916.580 3392.080 ;
        RECT 54.000 3389.360 2870.580 3391.600 ;
        RECT 8.000 3388.880 2916.580 3389.360 ;
        RECT 54.000 3386.640 2870.580 3388.880 ;
        RECT 8.000 3386.160 2916.580 3386.640 ;
        RECT 54.000 3383.920 2870.580 3386.160 ;
        RECT 8.000 3383.440 2916.580 3383.920 ;
        RECT 54.000 3381.200 2870.580 3383.440 ;
        RECT 8.000 3380.720 2916.580 3381.200 ;
        RECT 54.000 3378.480 2870.580 3380.720 ;
        RECT 8.000 3378.000 2916.580 3378.480 ;
        RECT 54.000 3375.760 2870.580 3378.000 ;
        RECT 8.000 3375.280 2916.580 3375.760 ;
        RECT 54.000 3373.040 2870.580 3375.280 ;
        RECT 8.000 3372.560 2916.580 3373.040 ;
        RECT 54.000 3370.320 2870.580 3372.560 ;
        RECT 8.000 3369.840 2916.580 3370.320 ;
        RECT 54.000 3367.600 2870.580 3369.840 ;
        RECT 8.000 3367.120 2916.580 3367.600 ;
        RECT 54.000 3364.880 2870.580 3367.120 ;
        RECT 8.000 3364.400 2916.580 3364.880 ;
        RECT 54.000 3362.160 2870.580 3364.400 ;
        RECT 8.000 3361.680 2916.580 3362.160 ;
        RECT 54.000 3359.440 2870.580 3361.680 ;
        RECT 8.000 3358.960 2916.580 3359.440 ;
        RECT 54.000 3356.720 2870.580 3358.960 ;
        RECT 8.000 3356.240 2916.580 3356.720 ;
        RECT 54.000 3354.000 2870.580 3356.240 ;
        RECT 8.000 3353.520 2916.580 3354.000 ;
        RECT 54.000 3351.280 2870.580 3353.520 ;
        RECT 8.000 3350.800 2916.580 3351.280 ;
        RECT 54.000 3348.560 2870.580 3350.800 ;
        RECT 8.000 3348.080 2916.580 3348.560 ;
        RECT 54.000 3345.840 2870.580 3348.080 ;
        RECT 8.000 3345.360 2916.580 3345.840 ;
        RECT 54.000 3343.120 2870.580 3345.360 ;
        RECT 8.000 3342.640 2916.580 3343.120 ;
        RECT 54.000 3340.400 2870.580 3342.640 ;
        RECT 8.000 3339.920 2916.580 3340.400 ;
        RECT 54.000 3337.680 2870.580 3339.920 ;
        RECT 8.000 3337.200 2916.580 3337.680 ;
        RECT 54.000 3334.960 2870.580 3337.200 ;
        RECT 8.000 3334.480 2916.580 3334.960 ;
        RECT 54.000 3332.240 2870.580 3334.480 ;
        RECT 8.000 3331.760 2916.580 3332.240 ;
        RECT 54.000 3329.520 2870.580 3331.760 ;
        RECT 8.000 3329.040 2916.580 3329.520 ;
        RECT 54.000 3326.800 2870.580 3329.040 ;
        RECT 8.000 3326.320 2916.580 3326.800 ;
        RECT 54.000 3324.080 2870.580 3326.320 ;
        RECT 8.000 3323.600 2916.580 3324.080 ;
        RECT 54.000 3321.360 2870.580 3323.600 ;
        RECT 8.000 3320.880 2916.580 3321.360 ;
        RECT 54.000 3318.640 2870.580 3320.880 ;
        RECT 8.000 3318.160 2916.580 3318.640 ;
        RECT 54.000 3315.920 2870.580 3318.160 ;
        RECT 8.000 3315.440 2916.580 3315.920 ;
        RECT 54.000 3313.200 2870.580 3315.440 ;
        RECT 8.000 3312.720 2916.580 3313.200 ;
        RECT 54.000 3310.480 2870.580 3312.720 ;
        RECT 8.000 3310.000 2916.580 3310.480 ;
        RECT 54.000 3307.760 2870.580 3310.000 ;
        RECT 8.000 3307.280 2916.580 3307.760 ;
        RECT 54.000 3305.040 2870.580 3307.280 ;
        RECT 8.000 3304.560 2916.580 3305.040 ;
        RECT 54.000 3302.320 2870.580 3304.560 ;
        RECT 8.000 3301.840 2916.580 3302.320 ;
        RECT 54.000 3299.600 2870.580 3301.840 ;
        RECT 8.000 3299.120 2916.580 3299.600 ;
        RECT 54.000 3296.880 2870.580 3299.120 ;
        RECT 8.000 3296.400 2916.580 3296.880 ;
        RECT 54.000 3294.160 2870.580 3296.400 ;
        RECT 8.000 3293.680 2916.580 3294.160 ;
        RECT 54.000 3291.440 2870.580 3293.680 ;
        RECT 8.000 3290.960 2916.580 3291.440 ;
        RECT 54.000 3288.720 2870.580 3290.960 ;
        RECT 8.000 3288.240 2916.580 3288.720 ;
        RECT 54.000 3286.000 2870.580 3288.240 ;
        RECT 8.000 3285.520 2916.580 3286.000 ;
        RECT 54.000 3283.280 2870.580 3285.520 ;
        RECT 8.000 3282.800 2916.580 3283.280 ;
        RECT 54.000 3280.560 2870.580 3282.800 ;
        RECT 8.000 3280.080 2916.580 3280.560 ;
        RECT 54.000 3277.840 2870.580 3280.080 ;
        RECT 8.000 3277.360 2916.580 3277.840 ;
        RECT 54.000 3275.120 2870.580 3277.360 ;
        RECT 8.000 3274.640 2916.580 3275.120 ;
        RECT 54.000 3272.400 2870.580 3274.640 ;
        RECT 8.000 3271.920 2916.580 3272.400 ;
        RECT 54.000 3269.680 2870.580 3271.920 ;
        RECT 8.000 3269.200 2916.580 3269.680 ;
        RECT 54.000 3266.960 2870.580 3269.200 ;
        RECT 8.000 3266.480 2916.580 3266.960 ;
        RECT 54.000 3264.240 2870.580 3266.480 ;
        RECT 8.000 3263.760 2916.580 3264.240 ;
        RECT 54.000 3261.520 2870.580 3263.760 ;
        RECT 8.000 3261.040 2916.580 3261.520 ;
        RECT 54.000 3258.800 2870.580 3261.040 ;
        RECT 8.000 3258.320 2916.580 3258.800 ;
        RECT 54.000 3256.080 2870.580 3258.320 ;
        RECT 8.000 3255.600 2916.580 3256.080 ;
        RECT 54.000 3253.360 2870.580 3255.600 ;
        RECT 8.000 3252.880 2916.580 3253.360 ;
        RECT 54.000 3250.640 2870.580 3252.880 ;
        RECT 8.000 3250.160 2916.580 3250.640 ;
        RECT 54.000 3247.920 2870.580 3250.160 ;
        RECT 8.000 3247.440 2916.580 3247.920 ;
        RECT 54.000 3245.200 2870.580 3247.440 ;
        RECT 8.000 3244.720 2916.580 3245.200 ;
        RECT 54.000 3242.480 2870.580 3244.720 ;
        RECT 8.000 3242.000 2916.580 3242.480 ;
        RECT 54.000 3239.760 2870.580 3242.000 ;
        RECT 8.000 3239.280 2916.580 3239.760 ;
        RECT 54.000 3237.040 2870.580 3239.280 ;
        RECT 8.000 3236.560 2916.580 3237.040 ;
        RECT 54.000 3234.320 2870.580 3236.560 ;
        RECT 8.000 3233.840 2916.580 3234.320 ;
        RECT 54.000 3231.600 2870.580 3233.840 ;
        RECT 8.000 3231.120 2916.580 3231.600 ;
        RECT 54.000 3228.880 2870.580 3231.120 ;
        RECT 8.000 3228.400 2916.580 3228.880 ;
        RECT 54.000 3226.160 2870.580 3228.400 ;
        RECT 8.000 3225.680 2916.580 3226.160 ;
        RECT 54.000 3223.440 2870.580 3225.680 ;
        RECT 8.000 3222.960 2916.580 3223.440 ;
        RECT 54.000 3220.720 2870.580 3222.960 ;
        RECT 8.000 3220.240 2916.580 3220.720 ;
        RECT 54.000 3218.000 2870.580 3220.240 ;
        RECT 8.000 3217.520 2916.580 3218.000 ;
        RECT 54.000 3215.280 2870.580 3217.520 ;
        RECT 8.000 3214.800 2916.580 3215.280 ;
        RECT 54.000 3212.560 2870.580 3214.800 ;
        RECT 8.000 3212.080 2916.580 3212.560 ;
        RECT 54.000 3209.840 2870.580 3212.080 ;
        RECT 8.000 3209.360 2916.580 3209.840 ;
        RECT 54.000 3207.120 2870.580 3209.360 ;
        RECT 8.000 3206.640 2916.580 3207.120 ;
        RECT 54.000 3204.400 2870.580 3206.640 ;
        RECT 8.000 3203.920 2916.580 3204.400 ;
        RECT 54.000 3201.680 2870.580 3203.920 ;
        RECT 8.000 3201.200 2916.580 3201.680 ;
        RECT 54.000 3198.960 2870.580 3201.200 ;
        RECT 8.000 3198.480 2916.580 3198.960 ;
        RECT 54.000 3196.240 2870.580 3198.480 ;
        RECT 8.000 3195.760 2916.580 3196.240 ;
        RECT 54.000 3193.520 2870.580 3195.760 ;
        RECT 8.000 3193.040 2916.580 3193.520 ;
        RECT 54.000 3190.800 2870.580 3193.040 ;
        RECT 8.000 3190.320 2916.580 3190.800 ;
        RECT 54.000 3188.080 2870.580 3190.320 ;
        RECT 8.000 3187.600 2916.580 3188.080 ;
        RECT 54.000 3185.360 2870.580 3187.600 ;
        RECT 8.000 3184.880 2916.580 3185.360 ;
        RECT 54.000 3182.640 2870.580 3184.880 ;
        RECT 8.000 3182.160 2916.580 3182.640 ;
        RECT 54.000 3179.920 2870.580 3182.160 ;
        RECT 8.000 3179.440 2916.580 3179.920 ;
        RECT 54.000 3177.200 2870.580 3179.440 ;
        RECT 8.000 3176.720 2916.580 3177.200 ;
        RECT 54.000 3174.480 2870.580 3176.720 ;
        RECT 8.000 3174.000 2916.580 3174.480 ;
        RECT 54.000 3171.760 2870.580 3174.000 ;
        RECT 8.000 3171.280 2916.580 3171.760 ;
        RECT 54.000 3169.040 2870.580 3171.280 ;
        RECT 8.000 3168.560 2916.580 3169.040 ;
        RECT 54.000 3166.320 2870.580 3168.560 ;
        RECT 8.000 3165.840 2916.580 3166.320 ;
        RECT 54.000 3163.600 2870.580 3165.840 ;
        RECT 8.000 3163.120 2916.580 3163.600 ;
        RECT 54.000 3160.880 2870.580 3163.120 ;
        RECT 8.000 3160.400 2916.580 3160.880 ;
        RECT 54.000 3158.160 2870.580 3160.400 ;
        RECT 8.000 3157.680 2916.580 3158.160 ;
        RECT 54.000 3155.440 2870.580 3157.680 ;
        RECT 8.000 3154.960 2916.580 3155.440 ;
        RECT 54.000 3152.720 2870.580 3154.960 ;
        RECT 8.000 3152.240 2916.580 3152.720 ;
        RECT 54.000 3150.000 2870.580 3152.240 ;
        RECT 8.000 3149.520 2916.580 3150.000 ;
        RECT 54.000 3147.280 2870.580 3149.520 ;
        RECT 8.000 3146.800 2916.580 3147.280 ;
        RECT 54.000 3144.560 2870.580 3146.800 ;
        RECT 8.000 3144.080 2916.580 3144.560 ;
        RECT 54.000 3141.840 2870.580 3144.080 ;
        RECT 8.000 3141.360 2916.580 3141.840 ;
        RECT 54.000 3139.120 2870.580 3141.360 ;
        RECT 8.000 3138.640 2916.580 3139.120 ;
        RECT 54.000 3136.400 2870.580 3138.640 ;
        RECT 8.000 3135.920 2916.580 3136.400 ;
        RECT 54.000 3133.680 2870.580 3135.920 ;
        RECT 8.000 3133.200 2916.580 3133.680 ;
        RECT 54.000 3130.960 2870.580 3133.200 ;
        RECT 8.000 3130.480 2916.580 3130.960 ;
        RECT 54.000 3128.240 2870.580 3130.480 ;
        RECT 8.000 3127.760 2916.580 3128.240 ;
        RECT 54.000 3125.520 2870.580 3127.760 ;
        RECT 8.000 3125.040 2916.580 3125.520 ;
        RECT 54.000 3122.800 2870.580 3125.040 ;
        RECT 8.000 3122.320 2916.580 3122.800 ;
        RECT 54.000 3120.080 2870.580 3122.320 ;
        RECT 8.000 3119.600 2916.580 3120.080 ;
        RECT 54.000 3117.360 2870.580 3119.600 ;
        RECT 8.000 3116.880 2916.580 3117.360 ;
        RECT 54.000 3114.640 2870.580 3116.880 ;
        RECT 8.000 3114.160 2916.580 3114.640 ;
        RECT 54.000 3111.920 2870.580 3114.160 ;
        RECT 8.000 3111.440 2916.580 3111.920 ;
        RECT 54.000 3109.200 2870.580 3111.440 ;
        RECT 8.000 3108.720 2916.580 3109.200 ;
        RECT 54.000 3106.480 2870.580 3108.720 ;
        RECT 8.000 3106.000 2916.580 3106.480 ;
        RECT 54.000 3103.760 2870.580 3106.000 ;
        RECT 8.000 3103.280 2916.580 3103.760 ;
        RECT 54.000 3101.040 2870.580 3103.280 ;
        RECT 8.000 3100.560 2916.580 3101.040 ;
        RECT 54.000 3098.320 2870.580 3100.560 ;
        RECT 8.000 3097.840 2916.580 3098.320 ;
        RECT 54.000 3095.600 2870.580 3097.840 ;
        RECT 8.000 3095.120 2916.580 3095.600 ;
        RECT 54.000 3092.880 2870.580 3095.120 ;
        RECT 8.000 3092.400 2916.580 3092.880 ;
        RECT 54.000 3090.160 2870.580 3092.400 ;
        RECT 8.000 3089.680 2916.580 3090.160 ;
        RECT 54.000 3087.440 2870.580 3089.680 ;
        RECT 8.000 3086.960 2916.580 3087.440 ;
        RECT 54.000 3084.720 2870.580 3086.960 ;
        RECT 8.000 3084.240 2916.580 3084.720 ;
        RECT 54.000 3082.000 2870.580 3084.240 ;
        RECT 8.000 3081.520 2916.580 3082.000 ;
        RECT 54.000 3079.280 2870.580 3081.520 ;
        RECT 8.000 3078.800 2916.580 3079.280 ;
        RECT 54.000 3076.560 2870.580 3078.800 ;
        RECT 8.000 3076.080 2916.580 3076.560 ;
        RECT 54.000 3073.840 2870.580 3076.080 ;
        RECT 8.000 3073.360 2916.580 3073.840 ;
        RECT 54.000 3071.120 2870.580 3073.360 ;
        RECT 8.000 3070.640 2916.580 3071.120 ;
        RECT 54.000 3068.400 2870.580 3070.640 ;
        RECT 8.000 3067.920 2916.580 3068.400 ;
        RECT 54.000 3065.680 2870.580 3067.920 ;
        RECT 8.000 3065.200 2916.580 3065.680 ;
        RECT 54.000 3062.960 2870.580 3065.200 ;
        RECT 8.000 3062.480 2916.580 3062.960 ;
        RECT 54.000 3060.240 2870.580 3062.480 ;
        RECT 8.000 3059.760 2916.580 3060.240 ;
        RECT 54.000 3057.520 2870.580 3059.760 ;
        RECT 8.000 3057.040 2916.580 3057.520 ;
        RECT 54.000 3054.800 2870.580 3057.040 ;
        RECT 8.000 3054.320 2916.580 3054.800 ;
        RECT 54.000 3052.080 2870.580 3054.320 ;
        RECT 8.000 3051.600 2916.580 3052.080 ;
        RECT 54.000 3049.360 2870.580 3051.600 ;
        RECT 8.000 3048.880 2916.580 3049.360 ;
        RECT 54.000 3046.640 2870.580 3048.880 ;
        RECT 8.000 3046.160 2916.580 3046.640 ;
        RECT 54.000 3043.920 2870.580 3046.160 ;
        RECT 8.000 3043.440 2916.580 3043.920 ;
        RECT 54.000 3041.200 2870.580 3043.440 ;
        RECT 8.000 3040.720 2916.580 3041.200 ;
        RECT 54.000 3038.480 2870.580 3040.720 ;
        RECT 8.000 3038.000 2916.580 3038.480 ;
        RECT 54.000 3035.760 2870.580 3038.000 ;
        RECT 8.000 3035.280 2916.580 3035.760 ;
        RECT 54.000 3033.040 2870.580 3035.280 ;
        RECT 8.000 3032.560 2916.580 3033.040 ;
        RECT 54.000 3030.320 2870.580 3032.560 ;
        RECT 8.000 3029.840 2916.580 3030.320 ;
        RECT 54.000 3027.600 2870.580 3029.840 ;
        RECT 8.000 3027.120 2916.580 3027.600 ;
        RECT 54.000 3024.880 2870.580 3027.120 ;
        RECT 8.000 3024.400 2916.580 3024.880 ;
        RECT 54.000 3022.160 2870.580 3024.400 ;
        RECT 8.000 3021.680 2916.580 3022.160 ;
        RECT 54.000 3019.440 2870.580 3021.680 ;
        RECT 8.000 3018.960 2916.580 3019.440 ;
        RECT 54.000 3016.720 2870.580 3018.960 ;
        RECT 8.000 3016.240 2916.580 3016.720 ;
        RECT 54.000 3014.000 2870.580 3016.240 ;
        RECT 8.000 3013.520 2916.580 3014.000 ;
        RECT 54.000 3011.280 2870.580 3013.520 ;
        RECT 8.000 3010.800 2916.580 3011.280 ;
        RECT 54.000 3008.560 2870.580 3010.800 ;
        RECT 8.000 3008.080 2916.580 3008.560 ;
        RECT 54.000 3005.840 2870.580 3008.080 ;
        RECT 8.000 3005.360 2916.580 3005.840 ;
        RECT 54.000 3003.120 2870.580 3005.360 ;
        RECT 8.000 3002.640 2916.580 3003.120 ;
        RECT 54.000 3000.400 2870.580 3002.640 ;
        RECT 8.000 2999.920 2916.580 3000.400 ;
        RECT 54.000 2997.680 2870.580 2999.920 ;
        RECT 8.000 2997.200 2916.580 2997.680 ;
        RECT 54.000 2994.960 2870.580 2997.200 ;
        RECT 8.000 2994.480 2916.580 2994.960 ;
        RECT 54.000 2992.240 2870.580 2994.480 ;
        RECT 8.000 2991.760 2916.580 2992.240 ;
        RECT 54.000 2989.520 2870.580 2991.760 ;
        RECT 8.000 2989.040 2916.580 2989.520 ;
        RECT 54.000 2986.800 2870.580 2989.040 ;
        RECT 8.000 2986.320 2916.580 2986.800 ;
        RECT 54.000 2984.080 2870.580 2986.320 ;
        RECT 8.000 2983.600 2916.580 2984.080 ;
        RECT 54.000 2981.360 2870.580 2983.600 ;
        RECT 8.000 2980.880 2916.580 2981.360 ;
        RECT 54.000 2978.640 2870.580 2980.880 ;
        RECT 8.000 2978.160 2916.580 2978.640 ;
        RECT 54.000 2975.920 2870.580 2978.160 ;
        RECT 8.000 2975.440 2916.580 2975.920 ;
        RECT 54.000 2973.200 2870.580 2975.440 ;
        RECT 8.000 2972.720 2916.580 2973.200 ;
        RECT 54.000 2970.480 2870.580 2972.720 ;
        RECT 8.000 2970.000 2916.580 2970.480 ;
        RECT 54.000 2967.760 2870.580 2970.000 ;
        RECT 8.000 2967.280 2916.580 2967.760 ;
        RECT 54.000 2965.040 2870.580 2967.280 ;
        RECT 8.000 2964.560 2916.580 2965.040 ;
        RECT 54.000 2962.320 2870.580 2964.560 ;
        RECT 8.000 2961.840 2916.580 2962.320 ;
        RECT 54.000 2959.600 2870.580 2961.840 ;
        RECT 8.000 2959.120 2916.580 2959.600 ;
        RECT 54.000 2956.880 2870.580 2959.120 ;
        RECT 8.000 2956.400 2916.580 2956.880 ;
        RECT 54.000 2954.160 2870.580 2956.400 ;
        RECT 8.000 2953.680 2916.580 2954.160 ;
        RECT 54.000 2951.440 2870.580 2953.680 ;
        RECT 8.000 2950.960 2916.580 2951.440 ;
        RECT 54.000 2948.720 2870.580 2950.960 ;
        RECT 8.000 2948.240 2916.580 2948.720 ;
        RECT 54.000 2946.000 2870.580 2948.240 ;
        RECT 8.000 2945.520 2916.580 2946.000 ;
        RECT 54.000 2943.280 2870.580 2945.520 ;
        RECT 8.000 2942.800 2916.580 2943.280 ;
        RECT 54.000 2940.560 2870.580 2942.800 ;
        RECT 8.000 2940.080 2916.580 2940.560 ;
        RECT 54.000 2937.840 2870.580 2940.080 ;
        RECT 8.000 2937.360 2916.580 2937.840 ;
        RECT 54.000 2935.120 2870.580 2937.360 ;
        RECT 8.000 2934.640 2916.580 2935.120 ;
        RECT 54.000 2932.400 2870.580 2934.640 ;
        RECT 8.000 2931.920 2916.580 2932.400 ;
        RECT 54.000 2929.680 2870.580 2931.920 ;
        RECT 8.000 2929.200 2916.580 2929.680 ;
        RECT 54.000 2926.960 2870.580 2929.200 ;
        RECT 8.000 2926.480 2916.580 2926.960 ;
        RECT 54.000 2924.240 2870.580 2926.480 ;
        RECT 8.000 2923.760 2916.580 2924.240 ;
        RECT 54.000 2921.520 2870.580 2923.760 ;
        RECT 8.000 2921.040 2916.580 2921.520 ;
        RECT 54.000 2918.800 2870.580 2921.040 ;
        RECT 8.000 2918.320 2916.580 2918.800 ;
        RECT 54.000 2916.080 2870.580 2918.320 ;
        RECT 8.000 2915.600 2916.580 2916.080 ;
        RECT 54.000 2913.360 2870.580 2915.600 ;
        RECT 8.000 2912.880 2916.580 2913.360 ;
        RECT 54.000 2910.640 2870.580 2912.880 ;
        RECT 8.000 2910.160 2916.580 2910.640 ;
        RECT 54.000 2907.920 2870.580 2910.160 ;
        RECT 8.000 2907.440 2916.580 2907.920 ;
        RECT 54.000 2905.200 2870.580 2907.440 ;
        RECT 8.000 2904.720 2916.580 2905.200 ;
        RECT 54.000 2902.480 2870.580 2904.720 ;
        RECT 8.000 2902.000 2916.580 2902.480 ;
        RECT 54.000 2899.760 2870.580 2902.000 ;
        RECT 8.000 2899.280 2916.580 2899.760 ;
        RECT 54.000 2897.040 2870.580 2899.280 ;
        RECT 8.000 2896.560 2916.580 2897.040 ;
        RECT 54.000 2894.320 2870.580 2896.560 ;
        RECT 8.000 2893.840 2916.580 2894.320 ;
        RECT 54.000 2891.600 2870.580 2893.840 ;
        RECT 8.000 2891.120 2916.580 2891.600 ;
        RECT 54.000 2888.880 2870.580 2891.120 ;
        RECT 8.000 2888.400 2916.580 2888.880 ;
        RECT 54.000 2886.160 2870.580 2888.400 ;
        RECT 8.000 2885.680 2916.580 2886.160 ;
        RECT 54.000 2883.440 2870.580 2885.680 ;
        RECT 8.000 2882.960 2916.580 2883.440 ;
        RECT 54.000 2880.720 2870.580 2882.960 ;
        RECT 8.000 2880.240 2916.580 2880.720 ;
        RECT 54.000 2878.000 2870.580 2880.240 ;
        RECT 8.000 2877.520 2916.580 2878.000 ;
        RECT 54.000 2875.280 2870.580 2877.520 ;
        RECT 8.000 2874.800 2916.580 2875.280 ;
        RECT 54.000 2872.560 2870.580 2874.800 ;
        RECT 8.000 2872.080 2916.580 2872.560 ;
        RECT 54.000 2869.840 2870.580 2872.080 ;
        RECT 8.000 2869.360 2916.580 2869.840 ;
        RECT 54.000 2867.120 2870.580 2869.360 ;
        RECT 8.000 2866.640 2916.580 2867.120 ;
        RECT 54.000 2864.400 2870.580 2866.640 ;
        RECT 8.000 2863.920 2916.580 2864.400 ;
        RECT 54.000 2861.680 2870.580 2863.920 ;
        RECT 8.000 2861.200 2916.580 2861.680 ;
        RECT 54.000 2858.960 2870.580 2861.200 ;
        RECT 8.000 2858.480 2916.580 2858.960 ;
        RECT 54.000 2856.240 2870.580 2858.480 ;
        RECT 8.000 2855.760 2916.580 2856.240 ;
        RECT 54.000 2853.520 2870.580 2855.760 ;
        RECT 8.000 2853.040 2916.580 2853.520 ;
        RECT 54.000 2850.800 2870.580 2853.040 ;
        RECT 8.000 2850.320 2916.580 2850.800 ;
        RECT 54.000 2848.080 2870.580 2850.320 ;
        RECT 8.000 2847.600 2916.580 2848.080 ;
        RECT 54.000 2845.360 2870.580 2847.600 ;
        RECT 8.000 2844.880 2916.580 2845.360 ;
        RECT 54.000 2842.640 2870.580 2844.880 ;
        RECT 8.000 2842.160 2916.580 2842.640 ;
        RECT 54.000 2839.920 2870.580 2842.160 ;
        RECT 8.000 2839.440 2916.580 2839.920 ;
        RECT 54.000 2837.200 2870.580 2839.440 ;
        RECT 8.000 2836.720 2916.580 2837.200 ;
        RECT 54.000 2834.480 2870.580 2836.720 ;
        RECT 8.000 2834.000 2916.580 2834.480 ;
        RECT 54.000 2831.760 2870.580 2834.000 ;
        RECT 8.000 2831.280 2916.580 2831.760 ;
        RECT 54.000 2829.040 2870.580 2831.280 ;
        RECT 8.000 2828.560 2916.580 2829.040 ;
        RECT 54.000 2826.320 2870.580 2828.560 ;
        RECT 8.000 2825.840 2916.580 2826.320 ;
        RECT 54.000 2823.600 2870.580 2825.840 ;
        RECT 8.000 2823.120 2916.580 2823.600 ;
        RECT 54.000 2820.880 2870.580 2823.120 ;
        RECT 8.000 2820.400 2916.580 2820.880 ;
        RECT 54.000 2818.160 2870.580 2820.400 ;
        RECT 8.000 2817.680 2916.580 2818.160 ;
        RECT 54.000 2815.440 2870.580 2817.680 ;
        RECT 8.000 2814.960 2916.580 2815.440 ;
        RECT 54.000 2812.720 2870.580 2814.960 ;
        RECT 8.000 2812.240 2916.580 2812.720 ;
        RECT 54.000 2810.000 2870.580 2812.240 ;
        RECT 8.000 2809.520 2916.580 2810.000 ;
        RECT 54.000 2807.280 2870.580 2809.520 ;
        RECT 8.000 2806.800 2916.580 2807.280 ;
        RECT 54.000 2804.560 2870.580 2806.800 ;
        RECT 8.000 2804.080 2916.580 2804.560 ;
        RECT 54.000 2801.840 2870.580 2804.080 ;
        RECT 8.000 2801.360 2916.580 2801.840 ;
        RECT 54.000 2799.120 2870.580 2801.360 ;
        RECT 8.000 2798.640 2916.580 2799.120 ;
        RECT 54.000 2796.400 2870.580 2798.640 ;
        RECT 8.000 2795.920 2916.580 2796.400 ;
        RECT 54.000 2793.680 2870.580 2795.920 ;
        RECT 8.000 2793.200 2916.580 2793.680 ;
        RECT 54.000 2790.960 2870.580 2793.200 ;
        RECT 8.000 2790.480 2916.580 2790.960 ;
        RECT 54.000 2788.240 2870.580 2790.480 ;
        RECT 8.000 2787.760 2916.580 2788.240 ;
        RECT 54.000 2785.520 2870.580 2787.760 ;
        RECT 8.000 2785.040 2916.580 2785.520 ;
        RECT 54.000 2782.800 2870.580 2785.040 ;
        RECT 8.000 2782.320 2916.580 2782.800 ;
        RECT 54.000 2780.080 2870.580 2782.320 ;
        RECT 8.000 2779.600 2916.580 2780.080 ;
        RECT 54.000 2777.360 2870.580 2779.600 ;
        RECT 8.000 2776.880 2916.580 2777.360 ;
        RECT 54.000 2774.640 2870.580 2776.880 ;
        RECT 8.000 2774.160 2916.580 2774.640 ;
        RECT 54.000 2771.920 2870.580 2774.160 ;
        RECT 8.000 2771.440 2916.580 2771.920 ;
        RECT 54.000 2769.200 2870.580 2771.440 ;
        RECT 8.000 2768.720 2916.580 2769.200 ;
        RECT 54.000 2766.480 2870.580 2768.720 ;
        RECT 8.000 2766.000 2916.580 2766.480 ;
        RECT 54.000 2763.760 2870.580 2766.000 ;
        RECT 8.000 2763.280 2916.580 2763.760 ;
        RECT 54.000 2761.040 2870.580 2763.280 ;
        RECT 8.000 2760.560 2916.580 2761.040 ;
        RECT 54.000 2758.320 2870.580 2760.560 ;
        RECT 8.000 2757.840 2916.580 2758.320 ;
        RECT 54.000 2755.600 2870.580 2757.840 ;
        RECT 8.000 2755.120 2916.580 2755.600 ;
        RECT 54.000 2752.880 2870.580 2755.120 ;
        RECT 8.000 2752.400 2916.580 2752.880 ;
        RECT 54.000 2750.160 2870.580 2752.400 ;
        RECT 8.000 2749.680 2916.580 2750.160 ;
        RECT 54.000 2747.440 2870.580 2749.680 ;
        RECT 8.000 2746.960 2916.580 2747.440 ;
        RECT 54.000 2744.720 2870.580 2746.960 ;
        RECT 8.000 2744.240 2916.580 2744.720 ;
        RECT 54.000 2742.000 2870.580 2744.240 ;
        RECT 8.000 2741.520 2916.580 2742.000 ;
        RECT 54.000 2739.280 2870.580 2741.520 ;
        RECT 8.000 2738.800 2916.580 2739.280 ;
        RECT 54.000 2736.560 2870.580 2738.800 ;
        RECT 8.000 2736.080 2916.580 2736.560 ;
        RECT 54.000 2733.840 2870.580 2736.080 ;
        RECT 8.000 2733.360 2916.580 2733.840 ;
        RECT 54.000 2731.120 2870.580 2733.360 ;
        RECT 8.000 2730.640 2916.580 2731.120 ;
        RECT 54.000 2728.400 2870.580 2730.640 ;
        RECT 8.000 2727.920 2916.580 2728.400 ;
        RECT 54.000 2725.680 2870.580 2727.920 ;
        RECT 8.000 2725.200 2916.580 2725.680 ;
        RECT 54.000 2722.960 2870.580 2725.200 ;
        RECT 8.000 2722.480 2916.580 2722.960 ;
        RECT 54.000 2720.240 2870.580 2722.480 ;
        RECT 8.000 2719.760 2916.580 2720.240 ;
        RECT 54.000 2717.520 2870.580 2719.760 ;
        RECT 8.000 2717.040 2916.580 2717.520 ;
        RECT 54.000 2714.800 2870.580 2717.040 ;
        RECT 8.000 2714.320 2916.580 2714.800 ;
        RECT 54.000 2712.080 2870.580 2714.320 ;
        RECT 8.000 2711.600 2916.580 2712.080 ;
        RECT 54.000 2709.360 2870.580 2711.600 ;
        RECT 8.000 2708.880 2916.580 2709.360 ;
        RECT 54.000 2706.640 2870.580 2708.880 ;
        RECT 8.000 2706.160 2916.580 2706.640 ;
        RECT 54.000 2703.920 2870.580 2706.160 ;
        RECT 8.000 2703.440 2916.580 2703.920 ;
        RECT 54.000 2701.200 2870.580 2703.440 ;
        RECT 8.000 2700.720 2916.580 2701.200 ;
        RECT 54.000 2698.480 2870.580 2700.720 ;
        RECT 8.000 2698.000 2916.580 2698.480 ;
        RECT 54.000 2695.760 2870.580 2698.000 ;
        RECT 8.000 2695.280 2916.580 2695.760 ;
        RECT 54.000 2693.040 2870.580 2695.280 ;
        RECT 8.000 2692.560 2916.580 2693.040 ;
        RECT 54.000 2690.320 2870.580 2692.560 ;
        RECT 8.000 2689.840 2916.580 2690.320 ;
        RECT 54.000 2687.600 2870.580 2689.840 ;
        RECT 8.000 2687.120 2916.580 2687.600 ;
        RECT 54.000 2684.880 2870.580 2687.120 ;
        RECT 8.000 2684.400 2916.580 2684.880 ;
        RECT 54.000 2682.160 2870.580 2684.400 ;
        RECT 8.000 2681.680 2916.580 2682.160 ;
        RECT 54.000 2679.440 2870.580 2681.680 ;
        RECT 8.000 2678.960 2916.580 2679.440 ;
        RECT 54.000 2676.720 2870.580 2678.960 ;
        RECT 8.000 2676.240 2916.580 2676.720 ;
        RECT 54.000 2674.000 2870.580 2676.240 ;
        RECT 8.000 2673.520 2916.580 2674.000 ;
        RECT 54.000 2671.280 2870.580 2673.520 ;
        RECT 8.000 2670.800 2916.580 2671.280 ;
        RECT 54.000 2668.560 2870.580 2670.800 ;
        RECT 8.000 2668.080 2916.580 2668.560 ;
        RECT 54.000 2665.840 2870.580 2668.080 ;
        RECT 8.000 2665.360 2916.580 2665.840 ;
        RECT 54.000 2663.120 2870.580 2665.360 ;
        RECT 8.000 2662.640 2916.580 2663.120 ;
        RECT 54.000 2660.400 2870.580 2662.640 ;
        RECT 8.000 2659.920 2916.580 2660.400 ;
        RECT 54.000 2657.680 2870.580 2659.920 ;
        RECT 8.000 2657.200 2916.580 2657.680 ;
        RECT 54.000 2654.960 2870.580 2657.200 ;
        RECT 8.000 2654.480 2916.580 2654.960 ;
        RECT 54.000 2652.240 2870.580 2654.480 ;
        RECT 8.000 2651.760 2916.580 2652.240 ;
        RECT 54.000 2649.520 2870.580 2651.760 ;
        RECT 8.000 2649.040 2916.580 2649.520 ;
        RECT 54.000 2646.800 2870.580 2649.040 ;
        RECT 8.000 2646.320 2916.580 2646.800 ;
        RECT 54.000 2644.080 2870.580 2646.320 ;
        RECT 8.000 2643.600 2916.580 2644.080 ;
        RECT 54.000 2641.360 2870.580 2643.600 ;
        RECT 8.000 2640.880 2916.580 2641.360 ;
        RECT 54.000 2638.640 2870.580 2640.880 ;
        RECT 8.000 2638.160 2916.580 2638.640 ;
        RECT 54.000 2635.920 2870.580 2638.160 ;
        RECT 8.000 2635.440 2916.580 2635.920 ;
        RECT 54.000 2633.200 2870.580 2635.440 ;
        RECT 8.000 2632.720 2916.580 2633.200 ;
        RECT 54.000 2630.480 2870.580 2632.720 ;
        RECT 8.000 2630.000 2916.580 2630.480 ;
        RECT 54.000 2627.760 2870.580 2630.000 ;
        RECT 8.000 2627.280 2916.580 2627.760 ;
        RECT 54.000 2625.040 2870.580 2627.280 ;
        RECT 8.000 2624.560 2916.580 2625.040 ;
        RECT 54.000 2622.320 2870.580 2624.560 ;
        RECT 8.000 2621.840 2916.580 2622.320 ;
        RECT 54.000 2619.600 2870.580 2621.840 ;
        RECT 8.000 2619.120 2916.580 2619.600 ;
        RECT 54.000 2616.880 2870.580 2619.120 ;
        RECT 8.000 2616.400 2916.580 2616.880 ;
        RECT 54.000 2614.160 2870.580 2616.400 ;
        RECT 8.000 2613.680 2916.580 2614.160 ;
        RECT 54.000 2611.440 2870.580 2613.680 ;
        RECT 8.000 2610.960 2916.580 2611.440 ;
        RECT 54.000 2608.720 2870.580 2610.960 ;
        RECT 8.000 2608.240 2916.580 2608.720 ;
        RECT 54.000 2606.000 2870.580 2608.240 ;
        RECT 8.000 2605.520 2916.580 2606.000 ;
        RECT 54.000 2603.280 2870.580 2605.520 ;
        RECT 8.000 2602.800 2916.580 2603.280 ;
        RECT 54.000 2600.560 2870.580 2602.800 ;
        RECT 8.000 2600.080 2916.580 2600.560 ;
        RECT 54.000 2597.840 2870.580 2600.080 ;
        RECT 8.000 2597.360 2916.580 2597.840 ;
        RECT 54.000 2595.120 2870.580 2597.360 ;
        RECT 8.000 2594.640 2916.580 2595.120 ;
        RECT 54.000 2592.400 2870.580 2594.640 ;
        RECT 8.000 2591.920 2916.580 2592.400 ;
        RECT 54.000 2589.680 2870.580 2591.920 ;
        RECT 8.000 2589.200 2916.580 2589.680 ;
        RECT 54.000 2586.960 2870.580 2589.200 ;
        RECT 8.000 2586.480 2916.580 2586.960 ;
        RECT 54.000 2584.240 2870.580 2586.480 ;
        RECT 8.000 2583.760 2916.580 2584.240 ;
        RECT 54.000 2581.520 2870.580 2583.760 ;
        RECT 8.000 2581.040 2916.580 2581.520 ;
        RECT 54.000 2578.800 2870.580 2581.040 ;
        RECT 8.000 2578.320 2916.580 2578.800 ;
        RECT 54.000 2576.080 2870.580 2578.320 ;
        RECT 8.000 2575.600 2916.580 2576.080 ;
        RECT 54.000 2573.360 2870.580 2575.600 ;
        RECT 8.000 2572.880 2916.580 2573.360 ;
        RECT 54.000 2570.640 2870.580 2572.880 ;
        RECT 8.000 2570.160 2916.580 2570.640 ;
        RECT 54.000 2567.920 2870.580 2570.160 ;
        RECT 8.000 2567.440 2916.580 2567.920 ;
        RECT 54.000 2565.200 2870.580 2567.440 ;
        RECT 8.000 2564.720 2916.580 2565.200 ;
        RECT 54.000 2562.480 2870.580 2564.720 ;
        RECT 8.000 2562.000 2916.580 2562.480 ;
        RECT 54.000 2559.760 2870.580 2562.000 ;
        RECT 8.000 2559.280 2916.580 2559.760 ;
        RECT 54.000 2557.040 2870.580 2559.280 ;
        RECT 8.000 2556.560 2916.580 2557.040 ;
        RECT 54.000 2554.320 2870.580 2556.560 ;
        RECT 8.000 2553.840 2916.580 2554.320 ;
        RECT 54.000 2551.600 2870.580 2553.840 ;
        RECT 8.000 2551.120 2916.580 2551.600 ;
        RECT 54.000 2548.880 2870.580 2551.120 ;
        RECT 8.000 2548.400 2916.580 2548.880 ;
        RECT 54.000 2546.160 2870.580 2548.400 ;
        RECT 8.000 2545.680 2916.580 2546.160 ;
        RECT 54.000 2543.440 2870.580 2545.680 ;
        RECT 8.000 2542.960 2916.580 2543.440 ;
        RECT 54.000 2540.720 2870.580 2542.960 ;
        RECT 8.000 2540.240 2916.580 2540.720 ;
        RECT 54.000 2538.000 2870.580 2540.240 ;
        RECT 8.000 2537.520 2916.580 2538.000 ;
        RECT 54.000 2535.280 2870.580 2537.520 ;
        RECT 8.000 2534.800 2916.580 2535.280 ;
        RECT 54.000 2532.560 2870.580 2534.800 ;
        RECT 8.000 2532.080 2916.580 2532.560 ;
        RECT 54.000 2529.840 2870.580 2532.080 ;
        RECT 8.000 2529.360 2916.580 2529.840 ;
        RECT 54.000 2527.120 2870.580 2529.360 ;
        RECT 8.000 2526.640 2916.580 2527.120 ;
        RECT 54.000 2524.400 2870.580 2526.640 ;
        RECT 8.000 2523.920 2916.580 2524.400 ;
        RECT 54.000 2521.680 2870.580 2523.920 ;
        RECT 8.000 2521.200 2916.580 2521.680 ;
        RECT 54.000 2518.960 2870.580 2521.200 ;
        RECT 8.000 2518.480 2916.580 2518.960 ;
        RECT 54.000 2516.240 2870.580 2518.480 ;
        RECT 8.000 2515.760 2916.580 2516.240 ;
        RECT 54.000 2513.520 2870.580 2515.760 ;
        RECT 8.000 2513.040 2916.580 2513.520 ;
        RECT 54.000 2510.800 2870.580 2513.040 ;
        RECT 8.000 2510.320 2916.580 2510.800 ;
        RECT 54.000 2508.080 2870.580 2510.320 ;
        RECT 8.000 2507.600 2916.580 2508.080 ;
        RECT 54.000 2505.360 2870.580 2507.600 ;
        RECT 8.000 2504.880 2916.580 2505.360 ;
        RECT 54.000 2502.640 2870.580 2504.880 ;
        RECT 8.000 2502.160 2916.580 2502.640 ;
        RECT 54.000 2499.920 2870.580 2502.160 ;
        RECT 8.000 2499.440 2916.580 2499.920 ;
        RECT 54.000 2497.200 2870.580 2499.440 ;
        RECT 8.000 2496.720 2916.580 2497.200 ;
        RECT 54.000 2494.480 2870.580 2496.720 ;
        RECT 8.000 2494.000 2916.580 2494.480 ;
        RECT 54.000 2491.760 2870.580 2494.000 ;
        RECT 8.000 2491.280 2916.580 2491.760 ;
        RECT 54.000 2489.040 2870.580 2491.280 ;
        RECT 8.000 2488.560 2916.580 2489.040 ;
        RECT 54.000 2486.320 2870.580 2488.560 ;
        RECT 8.000 2485.840 2916.580 2486.320 ;
        RECT 54.000 2483.600 2870.580 2485.840 ;
        RECT 8.000 2483.120 2916.580 2483.600 ;
        RECT 54.000 2480.880 2870.580 2483.120 ;
        RECT 8.000 2480.400 2916.580 2480.880 ;
        RECT 54.000 2478.160 2870.580 2480.400 ;
        RECT 8.000 2477.680 2916.580 2478.160 ;
        RECT 54.000 2475.440 2870.580 2477.680 ;
        RECT 8.000 2474.960 2916.580 2475.440 ;
        RECT 54.000 2472.720 2870.580 2474.960 ;
        RECT 8.000 2472.240 2916.580 2472.720 ;
        RECT 54.000 2470.000 2870.580 2472.240 ;
        RECT 8.000 2469.520 2916.580 2470.000 ;
        RECT 54.000 2467.280 2870.580 2469.520 ;
        RECT 8.000 2466.800 2916.580 2467.280 ;
        RECT 54.000 2464.560 2870.580 2466.800 ;
        RECT 8.000 2464.080 2916.580 2464.560 ;
        RECT 54.000 2461.840 2870.580 2464.080 ;
        RECT 8.000 2461.360 2916.580 2461.840 ;
        RECT 54.000 2459.120 2870.580 2461.360 ;
        RECT 8.000 2458.640 2916.580 2459.120 ;
        RECT 54.000 2456.400 2870.580 2458.640 ;
        RECT 8.000 2455.920 2916.580 2456.400 ;
        RECT 54.000 2453.680 2870.580 2455.920 ;
        RECT 8.000 2453.200 2916.580 2453.680 ;
        RECT 54.000 2450.960 2870.580 2453.200 ;
        RECT 8.000 2450.480 2916.580 2450.960 ;
        RECT 54.000 2448.240 2870.580 2450.480 ;
        RECT 8.000 2447.760 2916.580 2448.240 ;
        RECT 54.000 2445.520 2870.580 2447.760 ;
        RECT 8.000 2445.040 2916.580 2445.520 ;
        RECT 54.000 2442.800 2870.580 2445.040 ;
        RECT 8.000 2442.320 2916.580 2442.800 ;
        RECT 54.000 2440.080 2870.580 2442.320 ;
        RECT 8.000 2439.600 2916.580 2440.080 ;
        RECT 54.000 2437.360 2870.580 2439.600 ;
        RECT 8.000 2436.880 2916.580 2437.360 ;
        RECT 54.000 2434.640 2870.580 2436.880 ;
        RECT 8.000 2434.160 2916.580 2434.640 ;
        RECT 54.000 2431.920 2870.580 2434.160 ;
        RECT 8.000 2431.440 2916.580 2431.920 ;
        RECT 54.000 2429.200 2870.580 2431.440 ;
        RECT 8.000 2428.720 2916.580 2429.200 ;
        RECT 54.000 2426.480 2870.580 2428.720 ;
        RECT 8.000 2426.000 2916.580 2426.480 ;
        RECT 54.000 2423.760 2870.580 2426.000 ;
        RECT 8.000 2423.280 2916.580 2423.760 ;
        RECT 54.000 2421.040 2870.580 2423.280 ;
        RECT 8.000 2420.560 2916.580 2421.040 ;
        RECT 54.000 2418.320 2870.580 2420.560 ;
        RECT 8.000 2417.840 2916.580 2418.320 ;
        RECT 54.000 2415.600 2870.580 2417.840 ;
        RECT 8.000 2415.120 2916.580 2415.600 ;
        RECT 54.000 2412.880 2870.580 2415.120 ;
        RECT 8.000 2412.400 2916.580 2412.880 ;
        RECT 54.000 2410.160 2870.580 2412.400 ;
        RECT 8.000 2409.680 2916.580 2410.160 ;
        RECT 54.000 2407.440 2870.580 2409.680 ;
        RECT 8.000 2406.960 2916.580 2407.440 ;
        RECT 54.000 2404.720 2870.580 2406.960 ;
        RECT 8.000 2404.240 2916.580 2404.720 ;
        RECT 54.000 2402.000 2870.580 2404.240 ;
        RECT 8.000 2401.520 2916.580 2402.000 ;
        RECT 54.000 2399.280 2870.580 2401.520 ;
        RECT 8.000 2398.800 2916.580 2399.280 ;
        RECT 54.000 2396.560 2870.580 2398.800 ;
        RECT 8.000 2396.080 2916.580 2396.560 ;
        RECT 54.000 2393.840 2870.580 2396.080 ;
        RECT 8.000 2393.360 2916.580 2393.840 ;
        RECT 54.000 2391.120 2870.580 2393.360 ;
        RECT 8.000 2390.640 2916.580 2391.120 ;
        RECT 54.000 2388.400 2870.580 2390.640 ;
        RECT 8.000 2387.920 2916.580 2388.400 ;
        RECT 54.000 2385.680 2870.580 2387.920 ;
        RECT 8.000 2385.200 2916.580 2385.680 ;
        RECT 54.000 2382.960 2870.580 2385.200 ;
        RECT 8.000 2382.480 2916.580 2382.960 ;
        RECT 54.000 2380.240 2870.580 2382.480 ;
        RECT 8.000 2379.760 2916.580 2380.240 ;
        RECT 54.000 2377.520 2870.580 2379.760 ;
        RECT 8.000 2377.040 2916.580 2377.520 ;
        RECT 54.000 2374.800 2870.580 2377.040 ;
        RECT 8.000 2374.320 2916.580 2374.800 ;
        RECT 54.000 2372.080 2870.580 2374.320 ;
        RECT 8.000 2371.600 2916.580 2372.080 ;
        RECT 54.000 2369.360 2870.580 2371.600 ;
        RECT 8.000 2368.880 2916.580 2369.360 ;
        RECT 54.000 2366.640 2870.580 2368.880 ;
        RECT 8.000 2366.160 2916.580 2366.640 ;
        RECT 54.000 2363.920 2870.580 2366.160 ;
        RECT 8.000 2363.440 2916.580 2363.920 ;
        RECT 54.000 2361.200 2870.580 2363.440 ;
        RECT 8.000 2360.720 2916.580 2361.200 ;
        RECT 54.000 2358.480 2870.580 2360.720 ;
        RECT 8.000 2358.000 2916.580 2358.480 ;
        RECT 54.000 2355.760 2870.580 2358.000 ;
        RECT 8.000 2355.280 2916.580 2355.760 ;
        RECT 54.000 2353.040 2870.580 2355.280 ;
        RECT 8.000 2352.560 2916.580 2353.040 ;
        RECT 54.000 2350.320 2870.580 2352.560 ;
        RECT 8.000 2349.840 2916.580 2350.320 ;
        RECT 54.000 2347.600 2870.580 2349.840 ;
        RECT 8.000 2347.120 2916.580 2347.600 ;
        RECT 54.000 2344.880 2870.580 2347.120 ;
        RECT 8.000 2344.400 2916.580 2344.880 ;
        RECT 54.000 2342.160 2870.580 2344.400 ;
        RECT 8.000 2341.680 2916.580 2342.160 ;
        RECT 54.000 2339.440 2870.580 2341.680 ;
        RECT 8.000 2338.960 2916.580 2339.440 ;
        RECT 54.000 2336.720 2870.580 2338.960 ;
        RECT 8.000 2336.240 2916.580 2336.720 ;
        RECT 54.000 2334.000 2870.580 2336.240 ;
        RECT 8.000 2333.520 2916.580 2334.000 ;
        RECT 54.000 2331.280 2870.580 2333.520 ;
        RECT 8.000 2330.800 2916.580 2331.280 ;
        RECT 54.000 2328.560 2870.580 2330.800 ;
        RECT 8.000 2328.080 2916.580 2328.560 ;
        RECT 54.000 2325.840 2870.580 2328.080 ;
        RECT 8.000 2325.360 2916.580 2325.840 ;
        RECT 54.000 2323.120 2870.580 2325.360 ;
        RECT 8.000 2322.640 2916.580 2323.120 ;
        RECT 54.000 2320.400 2870.580 2322.640 ;
        RECT 8.000 2319.920 2916.580 2320.400 ;
        RECT 54.000 2317.680 2870.580 2319.920 ;
        RECT 8.000 2317.200 2916.580 2317.680 ;
        RECT 54.000 2314.960 2870.580 2317.200 ;
        RECT 8.000 2314.480 2916.580 2314.960 ;
        RECT 54.000 2312.240 2870.580 2314.480 ;
        RECT 8.000 2311.760 2916.580 2312.240 ;
        RECT 54.000 2309.520 2870.580 2311.760 ;
        RECT 8.000 2309.040 2916.580 2309.520 ;
        RECT 54.000 2306.800 2870.580 2309.040 ;
        RECT 8.000 2306.320 2916.580 2306.800 ;
        RECT 54.000 2304.080 2870.580 2306.320 ;
        RECT 8.000 2303.600 2916.580 2304.080 ;
        RECT 54.000 2301.360 2870.580 2303.600 ;
        RECT 8.000 2300.880 2916.580 2301.360 ;
        RECT 54.000 2298.640 2870.580 2300.880 ;
        RECT 8.000 2298.160 2916.580 2298.640 ;
        RECT 54.000 2295.920 2870.580 2298.160 ;
        RECT 8.000 2295.440 2916.580 2295.920 ;
        RECT 54.000 2293.200 2870.580 2295.440 ;
        RECT 8.000 2292.720 2916.580 2293.200 ;
        RECT 54.000 2290.480 2870.580 2292.720 ;
        RECT 8.000 2290.000 2916.580 2290.480 ;
        RECT 54.000 2287.760 2870.580 2290.000 ;
        RECT 8.000 2287.280 2916.580 2287.760 ;
        RECT 54.000 2285.040 2870.580 2287.280 ;
        RECT 8.000 2284.560 2916.580 2285.040 ;
        RECT 54.000 2282.320 2870.580 2284.560 ;
        RECT 8.000 2281.840 2916.580 2282.320 ;
        RECT 54.000 2279.600 2870.580 2281.840 ;
        RECT 8.000 2279.120 2916.580 2279.600 ;
        RECT 54.000 2276.880 2870.580 2279.120 ;
        RECT 8.000 2276.400 2916.580 2276.880 ;
        RECT 54.000 2274.160 2870.580 2276.400 ;
        RECT 8.000 2273.680 2916.580 2274.160 ;
        RECT 54.000 2271.440 2870.580 2273.680 ;
        RECT 8.000 2270.960 2916.580 2271.440 ;
        RECT 54.000 2268.720 2870.580 2270.960 ;
        RECT 8.000 2268.240 2916.580 2268.720 ;
        RECT 54.000 2266.000 2870.580 2268.240 ;
        RECT 8.000 2265.520 2916.580 2266.000 ;
        RECT 54.000 2263.280 2870.580 2265.520 ;
        RECT 8.000 2262.800 2916.580 2263.280 ;
        RECT 54.000 2260.560 2870.580 2262.800 ;
        RECT 8.000 2260.080 2916.580 2260.560 ;
        RECT 54.000 2257.840 2870.580 2260.080 ;
        RECT 8.000 2257.360 2916.580 2257.840 ;
        RECT 54.000 2255.120 2870.580 2257.360 ;
        RECT 8.000 2254.640 2916.580 2255.120 ;
        RECT 54.000 2252.400 2870.580 2254.640 ;
        RECT 8.000 2251.920 2916.580 2252.400 ;
        RECT 54.000 2249.680 2870.580 2251.920 ;
        RECT 8.000 2249.200 2916.580 2249.680 ;
        RECT 54.000 2246.960 2870.580 2249.200 ;
        RECT 8.000 2246.480 2916.580 2246.960 ;
        RECT 54.000 2244.240 2870.580 2246.480 ;
        RECT 8.000 2243.760 2916.580 2244.240 ;
        RECT 54.000 2241.520 2870.580 2243.760 ;
        RECT 8.000 2241.040 2916.580 2241.520 ;
        RECT 54.000 2238.800 2870.580 2241.040 ;
        RECT 8.000 2238.320 2916.580 2238.800 ;
        RECT 54.000 2236.080 2870.580 2238.320 ;
        RECT 8.000 2235.600 2916.580 2236.080 ;
        RECT 54.000 2233.360 2870.580 2235.600 ;
        RECT 8.000 2232.880 2916.580 2233.360 ;
        RECT 54.000 2230.640 2870.580 2232.880 ;
        RECT 8.000 2230.160 2916.580 2230.640 ;
        RECT 54.000 2227.920 2870.580 2230.160 ;
        RECT 8.000 2227.440 2916.580 2227.920 ;
        RECT 54.000 2225.200 2870.580 2227.440 ;
        RECT 8.000 2224.720 2916.580 2225.200 ;
        RECT 54.000 2222.480 2870.580 2224.720 ;
        RECT 8.000 2222.000 2916.580 2222.480 ;
        RECT 54.000 2219.760 2870.580 2222.000 ;
        RECT 8.000 2219.280 2916.580 2219.760 ;
        RECT 54.000 2217.040 2870.580 2219.280 ;
        RECT 8.000 2216.560 2916.580 2217.040 ;
        RECT 54.000 2214.320 2870.580 2216.560 ;
        RECT 8.000 2213.840 2916.580 2214.320 ;
        RECT 54.000 2211.600 2870.580 2213.840 ;
        RECT 8.000 2211.120 2916.580 2211.600 ;
        RECT 54.000 2208.880 2870.580 2211.120 ;
        RECT 8.000 2208.400 2916.580 2208.880 ;
        RECT 54.000 2206.160 2870.580 2208.400 ;
        RECT 8.000 2205.680 2916.580 2206.160 ;
        RECT 54.000 2203.440 2870.580 2205.680 ;
        RECT 8.000 2202.960 2916.580 2203.440 ;
        RECT 54.000 2200.720 2870.580 2202.960 ;
        RECT 8.000 2200.240 2916.580 2200.720 ;
        RECT 54.000 2198.000 2870.580 2200.240 ;
        RECT 8.000 2197.520 2916.580 2198.000 ;
        RECT 54.000 2195.280 2870.580 2197.520 ;
        RECT 8.000 2194.800 2916.580 2195.280 ;
        RECT 54.000 2192.560 2870.580 2194.800 ;
        RECT 8.000 2192.080 2916.580 2192.560 ;
        RECT 54.000 2189.840 2870.580 2192.080 ;
        RECT 8.000 2189.360 2916.580 2189.840 ;
        RECT 54.000 2187.120 2870.580 2189.360 ;
        RECT 8.000 2186.640 2916.580 2187.120 ;
        RECT 54.000 2184.400 2870.580 2186.640 ;
        RECT 8.000 2183.920 2916.580 2184.400 ;
        RECT 54.000 2181.680 2870.580 2183.920 ;
        RECT 8.000 2181.200 2916.580 2181.680 ;
        RECT 54.000 2178.960 2870.580 2181.200 ;
        RECT 8.000 2178.480 2916.580 2178.960 ;
        RECT 54.000 2176.240 2870.580 2178.480 ;
        RECT 8.000 2175.760 2916.580 2176.240 ;
        RECT 54.000 2173.520 2870.580 2175.760 ;
        RECT 8.000 2173.040 2916.580 2173.520 ;
        RECT 54.000 2170.800 2870.580 2173.040 ;
        RECT 8.000 2170.320 2916.580 2170.800 ;
        RECT 54.000 2168.080 2870.580 2170.320 ;
        RECT 8.000 2167.600 2916.580 2168.080 ;
        RECT 54.000 2165.360 2870.580 2167.600 ;
        RECT 8.000 2164.880 2916.580 2165.360 ;
        RECT 54.000 2162.640 2870.580 2164.880 ;
        RECT 8.000 2162.160 2916.580 2162.640 ;
        RECT 54.000 2159.920 2870.580 2162.160 ;
        RECT 8.000 2159.440 2916.580 2159.920 ;
        RECT 54.000 2157.200 2870.580 2159.440 ;
        RECT 8.000 2156.720 2916.580 2157.200 ;
        RECT 54.000 2154.480 2870.580 2156.720 ;
        RECT 8.000 2154.000 2916.580 2154.480 ;
        RECT 54.000 2151.760 2870.580 2154.000 ;
        RECT 8.000 2151.280 2916.580 2151.760 ;
        RECT 54.000 2149.040 2870.580 2151.280 ;
        RECT 8.000 2148.560 2916.580 2149.040 ;
        RECT 54.000 2146.320 2870.580 2148.560 ;
        RECT 8.000 2145.840 2916.580 2146.320 ;
        RECT 54.000 2143.600 2870.580 2145.840 ;
        RECT 8.000 2143.120 2916.580 2143.600 ;
        RECT 54.000 2140.880 2870.580 2143.120 ;
        RECT 8.000 2140.400 2916.580 2140.880 ;
        RECT 54.000 2138.160 2870.580 2140.400 ;
        RECT 8.000 2137.680 2916.580 2138.160 ;
        RECT 54.000 2135.440 2870.580 2137.680 ;
        RECT 8.000 2134.960 2916.580 2135.440 ;
        RECT 54.000 2132.720 2870.580 2134.960 ;
        RECT 8.000 2132.240 2916.580 2132.720 ;
        RECT 54.000 2130.000 2870.580 2132.240 ;
        RECT 8.000 2129.520 2916.580 2130.000 ;
        RECT 54.000 2127.280 2870.580 2129.520 ;
        RECT 8.000 2126.800 2916.580 2127.280 ;
        RECT 54.000 2124.560 2870.580 2126.800 ;
        RECT 8.000 2124.080 2916.580 2124.560 ;
        RECT 54.000 2121.840 2870.580 2124.080 ;
        RECT 8.000 2121.360 2916.580 2121.840 ;
        RECT 54.000 2119.120 2870.580 2121.360 ;
        RECT 8.000 2118.640 2916.580 2119.120 ;
        RECT 54.000 2116.400 2870.580 2118.640 ;
        RECT 8.000 2115.920 2916.580 2116.400 ;
        RECT 54.000 2113.680 2870.580 2115.920 ;
        RECT 8.000 2113.200 2916.580 2113.680 ;
        RECT 54.000 2110.960 2870.580 2113.200 ;
        RECT 8.000 2110.480 2916.580 2110.960 ;
        RECT 54.000 2108.240 2870.580 2110.480 ;
        RECT 8.000 2107.760 2916.580 2108.240 ;
        RECT 54.000 2105.520 2870.580 2107.760 ;
        RECT 8.000 2105.040 2916.580 2105.520 ;
        RECT 54.000 2102.800 2870.580 2105.040 ;
        RECT 8.000 2102.320 2916.580 2102.800 ;
        RECT 54.000 2100.080 2870.580 2102.320 ;
        RECT 8.000 2099.600 2916.580 2100.080 ;
        RECT 54.000 2097.360 2870.580 2099.600 ;
        RECT 8.000 2096.880 2916.580 2097.360 ;
        RECT 54.000 2094.640 2870.580 2096.880 ;
        RECT 8.000 2094.160 2916.580 2094.640 ;
        RECT 54.000 2091.920 2870.580 2094.160 ;
        RECT 8.000 2091.440 2916.580 2091.920 ;
        RECT 54.000 2089.200 2870.580 2091.440 ;
        RECT 8.000 2088.720 2916.580 2089.200 ;
        RECT 54.000 2086.480 2870.580 2088.720 ;
        RECT 8.000 2086.000 2916.580 2086.480 ;
        RECT 54.000 2083.760 2870.580 2086.000 ;
        RECT 8.000 2083.280 2916.580 2083.760 ;
        RECT 54.000 2081.040 2870.580 2083.280 ;
        RECT 8.000 2080.560 2916.580 2081.040 ;
        RECT 54.000 2078.320 2870.580 2080.560 ;
        RECT 8.000 2077.840 2916.580 2078.320 ;
        RECT 54.000 2075.600 2870.580 2077.840 ;
        RECT 8.000 2075.120 2916.580 2075.600 ;
        RECT 54.000 2072.880 2870.580 2075.120 ;
        RECT 8.000 2072.400 2916.580 2072.880 ;
        RECT 54.000 2070.160 2870.580 2072.400 ;
        RECT 8.000 2069.680 2916.580 2070.160 ;
        RECT 54.000 2067.440 2870.580 2069.680 ;
        RECT 8.000 2066.960 2916.580 2067.440 ;
        RECT 54.000 2064.720 2870.580 2066.960 ;
        RECT 8.000 2064.240 2916.580 2064.720 ;
        RECT 54.000 2062.000 2870.580 2064.240 ;
        RECT 8.000 2061.520 2916.580 2062.000 ;
        RECT 54.000 2059.280 2870.580 2061.520 ;
        RECT 8.000 2058.800 2916.580 2059.280 ;
        RECT 54.000 2056.560 2870.580 2058.800 ;
        RECT 8.000 2056.080 2916.580 2056.560 ;
        RECT 54.000 2053.840 2870.580 2056.080 ;
        RECT 8.000 2053.360 2916.580 2053.840 ;
        RECT 54.000 2051.120 2870.580 2053.360 ;
        RECT 8.000 2050.640 2916.580 2051.120 ;
        RECT 54.000 2048.400 2870.580 2050.640 ;
        RECT 8.000 2047.920 2916.580 2048.400 ;
        RECT 54.000 2045.680 2870.580 2047.920 ;
        RECT 8.000 2045.200 2916.580 2045.680 ;
        RECT 54.000 2042.960 2870.580 2045.200 ;
        RECT 8.000 2042.480 2916.580 2042.960 ;
        RECT 54.000 2040.240 2870.580 2042.480 ;
        RECT 8.000 2039.760 2916.580 2040.240 ;
        RECT 54.000 2037.520 2870.580 2039.760 ;
        RECT 8.000 2037.040 2916.580 2037.520 ;
        RECT 54.000 2034.800 2870.580 2037.040 ;
        RECT 8.000 2034.320 2916.580 2034.800 ;
        RECT 54.000 2032.080 2870.580 2034.320 ;
        RECT 8.000 2031.600 2916.580 2032.080 ;
        RECT 54.000 2029.360 2870.580 2031.600 ;
        RECT 8.000 2028.880 2916.580 2029.360 ;
        RECT 54.000 2026.640 2870.580 2028.880 ;
        RECT 8.000 2026.160 2916.580 2026.640 ;
        RECT 54.000 2023.920 2870.580 2026.160 ;
        RECT 8.000 2023.440 2916.580 2023.920 ;
        RECT 54.000 2021.200 2870.580 2023.440 ;
        RECT 8.000 2020.720 2916.580 2021.200 ;
        RECT 54.000 2018.480 2870.580 2020.720 ;
        RECT 8.000 2018.000 2916.580 2018.480 ;
        RECT 54.000 2015.760 2870.580 2018.000 ;
        RECT 8.000 2015.280 2916.580 2015.760 ;
        RECT 54.000 2013.040 2870.580 2015.280 ;
        RECT 8.000 2012.560 2916.580 2013.040 ;
        RECT 54.000 2010.320 2870.580 2012.560 ;
        RECT 8.000 2009.840 2916.580 2010.320 ;
        RECT 54.000 2007.600 2870.580 2009.840 ;
        RECT 8.000 2007.120 2916.580 2007.600 ;
        RECT 54.000 2004.880 2870.580 2007.120 ;
        RECT 8.000 2004.400 2916.580 2004.880 ;
        RECT 54.000 2002.160 2870.580 2004.400 ;
        RECT 8.000 2001.680 2916.580 2002.160 ;
        RECT 54.000 1999.440 2870.580 2001.680 ;
        RECT 8.000 1998.960 2916.580 1999.440 ;
        RECT 54.000 1996.720 2870.580 1998.960 ;
        RECT 8.000 1996.240 2916.580 1996.720 ;
        RECT 54.000 1994.000 2870.580 1996.240 ;
        RECT 8.000 1993.520 2916.580 1994.000 ;
        RECT 54.000 1991.280 2870.580 1993.520 ;
        RECT 8.000 1990.800 2916.580 1991.280 ;
        RECT 54.000 1988.560 2870.580 1990.800 ;
        RECT 8.000 1988.080 2916.580 1988.560 ;
        RECT 54.000 1985.840 2870.580 1988.080 ;
        RECT 8.000 1985.360 2916.580 1985.840 ;
        RECT 54.000 1983.120 2870.580 1985.360 ;
        RECT 8.000 1982.640 2916.580 1983.120 ;
        RECT 54.000 1980.400 2870.580 1982.640 ;
        RECT 8.000 1979.920 2916.580 1980.400 ;
        RECT 54.000 1977.680 2870.580 1979.920 ;
        RECT 8.000 1977.200 2916.580 1977.680 ;
        RECT 54.000 1974.960 2870.580 1977.200 ;
        RECT 8.000 1974.480 2916.580 1974.960 ;
        RECT 54.000 1972.240 2870.580 1974.480 ;
        RECT 8.000 1971.760 2916.580 1972.240 ;
        RECT 54.000 1969.520 2870.580 1971.760 ;
        RECT 8.000 1969.040 2916.580 1969.520 ;
        RECT 54.000 1966.800 2870.580 1969.040 ;
        RECT 8.000 1966.320 2916.580 1966.800 ;
        RECT 54.000 1964.080 2870.580 1966.320 ;
        RECT 8.000 1963.600 2916.580 1964.080 ;
        RECT 54.000 1961.360 2870.580 1963.600 ;
        RECT 8.000 1960.880 2916.580 1961.360 ;
        RECT 54.000 1958.640 2870.580 1960.880 ;
        RECT 8.000 1958.160 2916.580 1958.640 ;
        RECT 54.000 1955.920 2870.580 1958.160 ;
        RECT 8.000 1955.440 2916.580 1955.920 ;
        RECT 54.000 1953.200 2870.580 1955.440 ;
        RECT 8.000 1952.720 2916.580 1953.200 ;
        RECT 54.000 1950.480 2870.580 1952.720 ;
        RECT 8.000 1950.000 2916.580 1950.480 ;
        RECT 54.000 1947.760 2870.580 1950.000 ;
        RECT 8.000 1947.280 2916.580 1947.760 ;
        RECT 54.000 1945.040 2870.580 1947.280 ;
        RECT 8.000 1944.560 2916.580 1945.040 ;
        RECT 54.000 1942.320 2870.580 1944.560 ;
        RECT 8.000 1941.840 2916.580 1942.320 ;
        RECT 54.000 1939.600 2870.580 1941.840 ;
        RECT 8.000 1939.120 2916.580 1939.600 ;
        RECT 54.000 1936.880 2870.580 1939.120 ;
        RECT 8.000 1936.400 2916.580 1936.880 ;
        RECT 54.000 1934.160 2870.580 1936.400 ;
        RECT 8.000 1933.680 2916.580 1934.160 ;
        RECT 54.000 1931.440 2870.580 1933.680 ;
        RECT 8.000 1930.960 2916.580 1931.440 ;
        RECT 54.000 1928.720 2870.580 1930.960 ;
        RECT 8.000 1928.240 2916.580 1928.720 ;
        RECT 54.000 1926.000 2870.580 1928.240 ;
        RECT 8.000 1925.520 2916.580 1926.000 ;
        RECT 54.000 1923.280 2870.580 1925.520 ;
        RECT 8.000 1922.800 2916.580 1923.280 ;
        RECT 54.000 1920.560 2870.580 1922.800 ;
        RECT 8.000 1920.080 2916.580 1920.560 ;
        RECT 54.000 1917.840 2870.580 1920.080 ;
        RECT 8.000 1917.360 2916.580 1917.840 ;
        RECT 54.000 1915.120 2870.580 1917.360 ;
        RECT 8.000 1914.640 2916.580 1915.120 ;
        RECT 54.000 1912.400 2870.580 1914.640 ;
        RECT 8.000 1911.920 2916.580 1912.400 ;
        RECT 54.000 1909.680 2870.580 1911.920 ;
        RECT 8.000 1909.200 2916.580 1909.680 ;
        RECT 54.000 1906.960 2870.580 1909.200 ;
        RECT 8.000 1906.480 2916.580 1906.960 ;
        RECT 54.000 1904.240 2870.580 1906.480 ;
        RECT 8.000 1903.760 2916.580 1904.240 ;
        RECT 54.000 1901.520 2870.580 1903.760 ;
        RECT 8.000 1901.040 2916.580 1901.520 ;
        RECT 54.000 1898.800 2870.580 1901.040 ;
        RECT 8.000 1898.320 2916.580 1898.800 ;
        RECT 54.000 1896.080 2870.580 1898.320 ;
        RECT 8.000 1895.600 2916.580 1896.080 ;
        RECT 54.000 1893.360 2870.580 1895.600 ;
        RECT 8.000 1892.880 2916.580 1893.360 ;
        RECT 54.000 1890.640 2870.580 1892.880 ;
        RECT 8.000 1890.160 2916.580 1890.640 ;
        RECT 54.000 1887.920 2870.580 1890.160 ;
        RECT 8.000 1887.440 2916.580 1887.920 ;
        RECT 54.000 1885.200 2870.580 1887.440 ;
        RECT 8.000 1884.720 2916.580 1885.200 ;
        RECT 54.000 1882.480 2870.580 1884.720 ;
        RECT 8.000 1882.000 2916.580 1882.480 ;
        RECT 54.000 1879.760 2870.580 1882.000 ;
        RECT 8.000 1879.280 2916.580 1879.760 ;
        RECT 54.000 1877.040 2870.580 1879.280 ;
        RECT 8.000 1876.560 2916.580 1877.040 ;
        RECT 54.000 1874.320 2870.580 1876.560 ;
        RECT 8.000 1873.840 2916.580 1874.320 ;
        RECT 54.000 1871.600 2870.580 1873.840 ;
        RECT 8.000 1871.120 2916.580 1871.600 ;
        RECT 54.000 1868.880 2870.580 1871.120 ;
        RECT 8.000 1868.400 2916.580 1868.880 ;
        RECT 54.000 1866.160 2870.580 1868.400 ;
        RECT 8.000 1865.680 2916.580 1866.160 ;
        RECT 54.000 1863.440 2870.580 1865.680 ;
        RECT 8.000 1862.960 2916.580 1863.440 ;
        RECT 54.000 1860.720 2870.580 1862.960 ;
        RECT 8.000 1860.240 2916.580 1860.720 ;
        RECT 54.000 1858.000 2870.580 1860.240 ;
        RECT 8.000 1857.520 2916.580 1858.000 ;
        RECT 54.000 1855.280 2870.580 1857.520 ;
        RECT 8.000 1854.800 2916.580 1855.280 ;
        RECT 54.000 1852.560 2870.580 1854.800 ;
        RECT 8.000 1852.080 2916.580 1852.560 ;
        RECT 54.000 1849.840 2870.580 1852.080 ;
        RECT 8.000 1849.360 2916.580 1849.840 ;
        RECT 54.000 1847.120 2870.580 1849.360 ;
        RECT 8.000 1846.640 2916.580 1847.120 ;
        RECT 54.000 1844.400 2870.580 1846.640 ;
        RECT 8.000 1843.920 2916.580 1844.400 ;
        RECT 54.000 1841.680 2870.580 1843.920 ;
        RECT 8.000 1841.200 2916.580 1841.680 ;
        RECT 54.000 1838.960 2870.580 1841.200 ;
        RECT 8.000 1838.480 2916.580 1838.960 ;
        RECT 54.000 1836.240 2870.580 1838.480 ;
        RECT 8.000 1835.760 2916.580 1836.240 ;
        RECT 54.000 1833.520 2870.580 1835.760 ;
        RECT 8.000 1833.040 2916.580 1833.520 ;
        RECT 54.000 1830.800 2870.580 1833.040 ;
        RECT 8.000 1830.320 2916.580 1830.800 ;
        RECT 54.000 1828.080 2870.580 1830.320 ;
        RECT 8.000 1827.600 2916.580 1828.080 ;
        RECT 54.000 1825.360 2870.580 1827.600 ;
        RECT 8.000 1824.880 2916.580 1825.360 ;
        RECT 54.000 1822.640 2870.580 1824.880 ;
        RECT 8.000 1822.160 2916.580 1822.640 ;
        RECT 54.000 1819.920 2870.580 1822.160 ;
        RECT 8.000 1819.440 2916.580 1819.920 ;
        RECT 54.000 1817.200 2870.580 1819.440 ;
        RECT 8.000 1816.720 2916.580 1817.200 ;
        RECT 54.000 1814.480 2870.580 1816.720 ;
        RECT 8.000 1814.000 2916.580 1814.480 ;
        RECT 54.000 1811.760 2870.580 1814.000 ;
        RECT 8.000 1811.280 2916.580 1811.760 ;
        RECT 54.000 1809.040 2870.580 1811.280 ;
        RECT 8.000 1808.560 2916.580 1809.040 ;
        RECT 54.000 1806.320 2870.580 1808.560 ;
        RECT 8.000 1805.840 2916.580 1806.320 ;
        RECT 54.000 1803.600 2870.580 1805.840 ;
        RECT 8.000 1803.120 2916.580 1803.600 ;
        RECT 54.000 1800.880 2870.580 1803.120 ;
        RECT 8.000 1800.400 2916.580 1800.880 ;
        RECT 54.000 1798.160 2870.580 1800.400 ;
        RECT 8.000 1797.680 2916.580 1798.160 ;
        RECT 54.000 1795.440 2870.580 1797.680 ;
        RECT 8.000 1794.960 2916.580 1795.440 ;
        RECT 54.000 1792.720 2870.580 1794.960 ;
        RECT 8.000 1792.240 2916.580 1792.720 ;
        RECT 54.000 1790.000 2870.580 1792.240 ;
        RECT 8.000 1789.520 2916.580 1790.000 ;
        RECT 54.000 1787.280 2870.580 1789.520 ;
        RECT 8.000 1786.800 2916.580 1787.280 ;
        RECT 54.000 1784.560 2870.580 1786.800 ;
        RECT 8.000 1784.080 2916.580 1784.560 ;
        RECT 54.000 1781.840 2870.580 1784.080 ;
        RECT 8.000 1781.360 2916.580 1781.840 ;
        RECT 54.000 1779.120 2870.580 1781.360 ;
        RECT 8.000 1778.640 2916.580 1779.120 ;
        RECT 54.000 1776.400 2870.580 1778.640 ;
        RECT 8.000 1775.920 2916.580 1776.400 ;
        RECT 54.000 1773.680 2870.580 1775.920 ;
        RECT 8.000 1773.200 2916.580 1773.680 ;
        RECT 54.000 1770.960 2870.580 1773.200 ;
        RECT 8.000 1770.480 2916.580 1770.960 ;
        RECT 54.000 1768.240 2870.580 1770.480 ;
        RECT 8.000 1767.760 2916.580 1768.240 ;
        RECT 54.000 1765.520 2870.580 1767.760 ;
        RECT 8.000 1765.040 2916.580 1765.520 ;
        RECT 54.000 1762.800 2870.580 1765.040 ;
        RECT 8.000 1762.320 2916.580 1762.800 ;
        RECT 54.000 1760.080 2870.580 1762.320 ;
        RECT 8.000 1759.600 2916.580 1760.080 ;
        RECT 54.000 1757.360 2870.580 1759.600 ;
        RECT 8.000 1756.880 2916.580 1757.360 ;
        RECT 54.000 1754.640 2870.580 1756.880 ;
        RECT 8.000 1754.160 2916.580 1754.640 ;
        RECT 54.000 1751.920 2870.580 1754.160 ;
        RECT 8.000 1751.440 2916.580 1751.920 ;
        RECT 54.000 1749.200 2870.580 1751.440 ;
        RECT 8.000 1748.720 2916.580 1749.200 ;
        RECT 54.000 1746.480 2870.580 1748.720 ;
        RECT 8.000 1746.000 2916.580 1746.480 ;
        RECT 54.000 1743.760 2870.580 1746.000 ;
        RECT 8.000 1743.280 2916.580 1743.760 ;
        RECT 54.000 1741.040 2870.580 1743.280 ;
        RECT 8.000 1740.560 2916.580 1741.040 ;
        RECT 54.000 1738.320 2870.580 1740.560 ;
        RECT 8.000 1737.840 2916.580 1738.320 ;
        RECT 54.000 1735.600 2870.580 1737.840 ;
        RECT 8.000 1735.120 2916.580 1735.600 ;
        RECT 54.000 1732.880 2870.580 1735.120 ;
        RECT 8.000 1732.400 2916.580 1732.880 ;
        RECT 54.000 1730.160 2870.580 1732.400 ;
        RECT 8.000 1729.680 2916.580 1730.160 ;
        RECT 54.000 1727.440 2870.580 1729.680 ;
        RECT 8.000 1726.960 2916.580 1727.440 ;
        RECT 54.000 1724.720 2870.580 1726.960 ;
        RECT 8.000 1724.240 2916.580 1724.720 ;
        RECT 54.000 1722.000 2870.580 1724.240 ;
        RECT 8.000 1721.520 2916.580 1722.000 ;
        RECT 54.000 1719.280 2870.580 1721.520 ;
        RECT 8.000 1718.800 2916.580 1719.280 ;
        RECT 54.000 1716.560 2870.580 1718.800 ;
        RECT 8.000 1716.080 2916.580 1716.560 ;
        RECT 54.000 1713.840 2870.580 1716.080 ;
        RECT 8.000 1713.360 2916.580 1713.840 ;
        RECT 54.000 1711.120 2870.580 1713.360 ;
        RECT 8.000 1710.640 2916.580 1711.120 ;
        RECT 54.000 1708.400 2870.580 1710.640 ;
        RECT 8.000 1707.920 2916.580 1708.400 ;
        RECT 54.000 1705.680 2870.580 1707.920 ;
        RECT 8.000 1705.200 2916.580 1705.680 ;
        RECT 54.000 1702.960 2870.580 1705.200 ;
        RECT 8.000 1702.480 2916.580 1702.960 ;
        RECT 54.000 1700.240 2870.580 1702.480 ;
        RECT 8.000 1699.760 2916.580 1700.240 ;
        RECT 54.000 1697.520 2870.580 1699.760 ;
        RECT 8.000 1697.040 2916.580 1697.520 ;
        RECT 54.000 1694.800 2870.580 1697.040 ;
        RECT 8.000 1694.320 2916.580 1694.800 ;
        RECT 54.000 1692.080 2870.580 1694.320 ;
        RECT 8.000 1691.600 2916.580 1692.080 ;
        RECT 54.000 1689.360 2870.580 1691.600 ;
        RECT 8.000 1688.880 2916.580 1689.360 ;
        RECT 54.000 1686.640 2870.580 1688.880 ;
        RECT 8.000 1686.160 2916.580 1686.640 ;
        RECT 54.000 1683.920 2870.580 1686.160 ;
        RECT 8.000 1683.440 2916.580 1683.920 ;
        RECT 54.000 1681.200 2870.580 1683.440 ;
        RECT 8.000 1680.720 2916.580 1681.200 ;
        RECT 54.000 1678.480 2870.580 1680.720 ;
        RECT 8.000 1678.000 2916.580 1678.480 ;
        RECT 54.000 1675.760 2870.580 1678.000 ;
        RECT 8.000 1675.280 2916.580 1675.760 ;
        RECT 54.000 1673.040 2870.580 1675.280 ;
        RECT 8.000 1672.560 2916.580 1673.040 ;
        RECT 54.000 1670.320 2870.580 1672.560 ;
        RECT 8.000 1669.840 2916.580 1670.320 ;
        RECT 54.000 1667.600 2870.580 1669.840 ;
        RECT 8.000 1667.120 2916.580 1667.600 ;
        RECT 54.000 1664.880 2870.580 1667.120 ;
        RECT 8.000 1664.400 2916.580 1664.880 ;
        RECT 54.000 1662.160 2870.580 1664.400 ;
        RECT 8.000 1661.680 2916.580 1662.160 ;
        RECT 54.000 1659.440 2870.580 1661.680 ;
        RECT 8.000 1658.960 2916.580 1659.440 ;
        RECT 54.000 1656.720 2870.580 1658.960 ;
        RECT 8.000 1656.240 2916.580 1656.720 ;
        RECT 54.000 1654.000 2870.580 1656.240 ;
        RECT 8.000 1653.520 2916.580 1654.000 ;
        RECT 54.000 1651.280 2870.580 1653.520 ;
        RECT 8.000 1650.800 2916.580 1651.280 ;
        RECT 54.000 1648.560 2870.580 1650.800 ;
        RECT 8.000 1648.080 2916.580 1648.560 ;
        RECT 54.000 1645.840 2870.580 1648.080 ;
        RECT 8.000 1645.360 2916.580 1645.840 ;
        RECT 54.000 1643.120 2870.580 1645.360 ;
        RECT 8.000 1642.640 2916.580 1643.120 ;
        RECT 54.000 1640.400 2870.580 1642.640 ;
        RECT 8.000 1639.920 2916.580 1640.400 ;
        RECT 54.000 1637.680 2870.580 1639.920 ;
        RECT 8.000 1637.200 2916.580 1637.680 ;
        RECT 54.000 1634.960 2870.580 1637.200 ;
        RECT 8.000 1634.480 2916.580 1634.960 ;
        RECT 54.000 1632.240 2870.580 1634.480 ;
        RECT 8.000 1631.760 2916.580 1632.240 ;
        RECT 54.000 1629.520 2870.580 1631.760 ;
        RECT 8.000 1629.040 2916.580 1629.520 ;
        RECT 54.000 1626.800 2870.580 1629.040 ;
        RECT 8.000 1626.320 2916.580 1626.800 ;
        RECT 54.000 1624.080 2870.580 1626.320 ;
        RECT 8.000 1623.600 2916.580 1624.080 ;
        RECT 54.000 1621.360 2870.580 1623.600 ;
        RECT 8.000 1620.880 2916.580 1621.360 ;
        RECT 54.000 1618.640 2870.580 1620.880 ;
        RECT 8.000 1618.160 2916.580 1618.640 ;
        RECT 54.000 1615.920 2870.580 1618.160 ;
        RECT 8.000 1615.440 2916.580 1615.920 ;
        RECT 54.000 1613.200 2870.580 1615.440 ;
        RECT 8.000 1612.720 2916.580 1613.200 ;
        RECT 54.000 1610.480 2870.580 1612.720 ;
        RECT 8.000 1610.000 2916.580 1610.480 ;
        RECT 54.000 1607.760 2870.580 1610.000 ;
        RECT 8.000 1607.280 2916.580 1607.760 ;
        RECT 54.000 1605.040 2870.580 1607.280 ;
        RECT 8.000 1604.560 2916.580 1605.040 ;
        RECT 54.000 1602.320 2870.580 1604.560 ;
        RECT 8.000 1601.840 2916.580 1602.320 ;
        RECT 54.000 1599.600 2870.580 1601.840 ;
        RECT 8.000 1599.120 2916.580 1599.600 ;
        RECT 54.000 1596.880 2870.580 1599.120 ;
        RECT 8.000 1596.400 2916.580 1596.880 ;
        RECT 54.000 1594.160 2870.580 1596.400 ;
        RECT 8.000 1593.680 2916.580 1594.160 ;
        RECT 54.000 1591.440 2870.580 1593.680 ;
        RECT 8.000 1590.960 2916.580 1591.440 ;
        RECT 54.000 1588.720 2870.580 1590.960 ;
        RECT 8.000 1588.240 2916.580 1588.720 ;
        RECT 54.000 1586.000 2870.580 1588.240 ;
        RECT 8.000 1585.520 2916.580 1586.000 ;
        RECT 54.000 1583.280 2870.580 1585.520 ;
        RECT 8.000 1582.800 2916.580 1583.280 ;
        RECT 54.000 1580.560 2870.580 1582.800 ;
        RECT 8.000 1580.080 2916.580 1580.560 ;
        RECT 54.000 1577.840 2870.580 1580.080 ;
        RECT 8.000 1577.360 2916.580 1577.840 ;
        RECT 54.000 1575.120 2870.580 1577.360 ;
        RECT 8.000 1574.640 2916.580 1575.120 ;
        RECT 54.000 1572.400 2870.580 1574.640 ;
        RECT 8.000 1571.920 2916.580 1572.400 ;
        RECT 54.000 1569.680 2870.580 1571.920 ;
        RECT 8.000 1569.200 2916.580 1569.680 ;
        RECT 54.000 1566.960 2870.580 1569.200 ;
        RECT 8.000 1566.480 2916.580 1566.960 ;
        RECT 54.000 1564.240 2870.580 1566.480 ;
        RECT 8.000 1563.760 2916.580 1564.240 ;
        RECT 54.000 1561.520 2870.580 1563.760 ;
        RECT 8.000 1561.040 2916.580 1561.520 ;
        RECT 54.000 1558.800 2870.580 1561.040 ;
        RECT 8.000 1558.320 2916.580 1558.800 ;
        RECT 54.000 1556.080 2870.580 1558.320 ;
        RECT 8.000 1555.600 2916.580 1556.080 ;
        RECT 54.000 1553.360 2870.580 1555.600 ;
        RECT 8.000 1552.880 2916.580 1553.360 ;
        RECT 54.000 1550.640 2870.580 1552.880 ;
        RECT 8.000 1550.160 2916.580 1550.640 ;
        RECT 54.000 1547.920 2870.580 1550.160 ;
        RECT 8.000 1547.440 2916.580 1547.920 ;
        RECT 54.000 1545.200 2870.580 1547.440 ;
        RECT 8.000 1544.720 2916.580 1545.200 ;
        RECT 54.000 1542.480 2870.580 1544.720 ;
        RECT 8.000 1542.000 2916.580 1542.480 ;
        RECT 54.000 1539.760 2870.580 1542.000 ;
        RECT 8.000 1539.280 2916.580 1539.760 ;
        RECT 54.000 1537.040 2870.580 1539.280 ;
        RECT 8.000 1536.560 2916.580 1537.040 ;
        RECT 54.000 1534.320 2870.580 1536.560 ;
        RECT 8.000 1533.840 2916.580 1534.320 ;
        RECT 54.000 1531.600 2870.580 1533.840 ;
        RECT 8.000 1531.120 2916.580 1531.600 ;
        RECT 54.000 1528.880 2870.580 1531.120 ;
        RECT 8.000 1528.400 2916.580 1528.880 ;
        RECT 54.000 1526.160 2870.580 1528.400 ;
        RECT 8.000 1525.680 2916.580 1526.160 ;
        RECT 54.000 1523.440 2870.580 1525.680 ;
        RECT 8.000 1522.960 2916.580 1523.440 ;
        RECT 54.000 1520.720 2870.580 1522.960 ;
        RECT 8.000 1520.240 2916.580 1520.720 ;
        RECT 54.000 1518.000 2870.580 1520.240 ;
        RECT 8.000 1517.520 2916.580 1518.000 ;
        RECT 54.000 1515.280 2870.580 1517.520 ;
        RECT 8.000 1514.800 2916.580 1515.280 ;
        RECT 54.000 1512.560 2870.580 1514.800 ;
        RECT 8.000 1512.080 2916.580 1512.560 ;
        RECT 54.000 1509.840 2870.580 1512.080 ;
        RECT 8.000 1509.360 2916.580 1509.840 ;
        RECT 54.000 1507.120 2870.580 1509.360 ;
        RECT 8.000 1506.640 2916.580 1507.120 ;
        RECT 54.000 1504.400 2870.580 1506.640 ;
        RECT 8.000 1503.920 2916.580 1504.400 ;
        RECT 54.000 1501.680 2870.580 1503.920 ;
        RECT 8.000 1501.200 2916.580 1501.680 ;
        RECT 54.000 1498.960 2870.580 1501.200 ;
        RECT 8.000 1498.480 2916.580 1498.960 ;
        RECT 54.000 1496.240 2870.580 1498.480 ;
        RECT 8.000 1495.760 2916.580 1496.240 ;
        RECT 54.000 1493.520 2870.580 1495.760 ;
        RECT 8.000 1493.040 2916.580 1493.520 ;
        RECT 54.000 1490.800 2870.580 1493.040 ;
        RECT 8.000 1490.320 2916.580 1490.800 ;
        RECT 54.000 1488.080 2870.580 1490.320 ;
        RECT 8.000 1487.600 2916.580 1488.080 ;
        RECT 54.000 1485.360 2870.580 1487.600 ;
        RECT 8.000 1484.880 2916.580 1485.360 ;
        RECT 54.000 1482.640 2870.580 1484.880 ;
        RECT 8.000 1482.160 2916.580 1482.640 ;
        RECT 54.000 1479.920 2870.580 1482.160 ;
        RECT 8.000 1479.440 2916.580 1479.920 ;
        RECT 54.000 1477.200 2870.580 1479.440 ;
        RECT 8.000 1476.720 2916.580 1477.200 ;
        RECT 54.000 1474.480 2870.580 1476.720 ;
        RECT 8.000 1474.000 2916.580 1474.480 ;
        RECT 54.000 1471.760 2870.580 1474.000 ;
        RECT 8.000 1471.280 2916.580 1471.760 ;
        RECT 54.000 1469.040 2870.580 1471.280 ;
        RECT 8.000 1468.560 2916.580 1469.040 ;
        RECT 54.000 1466.320 2870.580 1468.560 ;
        RECT 8.000 1465.840 2916.580 1466.320 ;
        RECT 54.000 1463.600 2870.580 1465.840 ;
        RECT 8.000 1463.120 2916.580 1463.600 ;
        RECT 54.000 1460.880 2870.580 1463.120 ;
        RECT 8.000 1460.400 2916.580 1460.880 ;
        RECT 54.000 1458.160 2870.580 1460.400 ;
        RECT 8.000 1457.680 2916.580 1458.160 ;
        RECT 54.000 1455.440 2870.580 1457.680 ;
        RECT 8.000 1454.960 2916.580 1455.440 ;
        RECT 54.000 1452.720 2870.580 1454.960 ;
        RECT 8.000 1452.240 2916.580 1452.720 ;
        RECT 54.000 1450.000 2870.580 1452.240 ;
        RECT 8.000 1449.520 2916.580 1450.000 ;
        RECT 54.000 1447.280 2870.580 1449.520 ;
        RECT 8.000 1446.800 2916.580 1447.280 ;
        RECT 54.000 1444.560 2870.580 1446.800 ;
        RECT 8.000 1444.080 2916.580 1444.560 ;
        RECT 54.000 1441.840 2870.580 1444.080 ;
        RECT 8.000 1441.360 2916.580 1441.840 ;
        RECT 54.000 1439.120 2870.580 1441.360 ;
        RECT 8.000 1438.640 2916.580 1439.120 ;
        RECT 54.000 1436.400 2870.580 1438.640 ;
        RECT 8.000 1435.920 2916.580 1436.400 ;
        RECT 54.000 1433.680 2870.580 1435.920 ;
        RECT 8.000 1433.200 2916.580 1433.680 ;
        RECT 54.000 1430.960 2870.580 1433.200 ;
        RECT 8.000 1430.480 2916.580 1430.960 ;
        RECT 54.000 1428.240 2870.580 1430.480 ;
        RECT 8.000 1427.760 2916.580 1428.240 ;
        RECT 54.000 1425.520 2870.580 1427.760 ;
        RECT 8.000 1425.040 2916.580 1425.520 ;
        RECT 54.000 1422.800 2870.580 1425.040 ;
        RECT 8.000 1422.320 2916.580 1422.800 ;
        RECT 54.000 1420.080 2870.580 1422.320 ;
        RECT 8.000 1419.600 2916.580 1420.080 ;
        RECT 54.000 1417.360 2870.580 1419.600 ;
        RECT 8.000 1416.880 2916.580 1417.360 ;
        RECT 54.000 1414.640 2870.580 1416.880 ;
        RECT 8.000 1414.160 2916.580 1414.640 ;
        RECT 54.000 1411.920 2870.580 1414.160 ;
        RECT 8.000 1411.440 2916.580 1411.920 ;
        RECT 54.000 1409.200 2870.580 1411.440 ;
        RECT 8.000 1408.720 2916.580 1409.200 ;
        RECT 54.000 1406.480 2870.580 1408.720 ;
        RECT 8.000 1406.000 2916.580 1406.480 ;
        RECT 54.000 1403.760 2870.580 1406.000 ;
        RECT 8.000 1403.280 2916.580 1403.760 ;
        RECT 54.000 1401.040 2870.580 1403.280 ;
        RECT 8.000 1400.560 2916.580 1401.040 ;
        RECT 54.000 1398.320 2870.580 1400.560 ;
        RECT 8.000 1397.840 2916.580 1398.320 ;
        RECT 54.000 1395.600 2870.580 1397.840 ;
        RECT 8.000 1395.120 2916.580 1395.600 ;
        RECT 54.000 1392.880 2870.580 1395.120 ;
        RECT 8.000 1392.400 2916.580 1392.880 ;
        RECT 54.000 1390.160 2870.580 1392.400 ;
        RECT 8.000 1389.680 2916.580 1390.160 ;
        RECT 54.000 1387.440 2870.580 1389.680 ;
        RECT 8.000 1386.960 2916.580 1387.440 ;
        RECT 54.000 1384.720 2870.580 1386.960 ;
        RECT 8.000 1384.240 2916.580 1384.720 ;
        RECT 54.000 1382.000 2870.580 1384.240 ;
        RECT 8.000 1381.520 2916.580 1382.000 ;
        RECT 54.000 1379.280 2870.580 1381.520 ;
        RECT 8.000 1378.800 2916.580 1379.280 ;
        RECT 54.000 1376.560 2870.580 1378.800 ;
        RECT 8.000 1376.080 2916.580 1376.560 ;
        RECT 54.000 1373.840 2870.580 1376.080 ;
        RECT 8.000 1373.360 2916.580 1373.840 ;
        RECT 54.000 1371.120 2870.580 1373.360 ;
        RECT 8.000 1370.640 2916.580 1371.120 ;
        RECT 54.000 1368.400 2870.580 1370.640 ;
        RECT 8.000 1367.920 2916.580 1368.400 ;
        RECT 54.000 1365.680 2870.580 1367.920 ;
        RECT 8.000 1365.200 2916.580 1365.680 ;
        RECT 54.000 1362.960 2870.580 1365.200 ;
        RECT 8.000 1362.480 2916.580 1362.960 ;
        RECT 54.000 1360.240 2870.580 1362.480 ;
        RECT 8.000 1359.760 2916.580 1360.240 ;
        RECT 54.000 1357.520 2870.580 1359.760 ;
        RECT 8.000 1357.040 2916.580 1357.520 ;
        RECT 54.000 1354.800 2870.580 1357.040 ;
        RECT 8.000 1354.320 2916.580 1354.800 ;
        RECT 54.000 1352.080 2870.580 1354.320 ;
        RECT 8.000 1351.600 2916.580 1352.080 ;
        RECT 54.000 1349.360 2870.580 1351.600 ;
        RECT 8.000 1348.880 2916.580 1349.360 ;
        RECT 54.000 1346.640 2870.580 1348.880 ;
        RECT 8.000 1346.160 2916.580 1346.640 ;
        RECT 54.000 1343.920 2870.580 1346.160 ;
        RECT 8.000 1343.440 2916.580 1343.920 ;
        RECT 54.000 1341.200 2870.580 1343.440 ;
        RECT 8.000 1340.720 2916.580 1341.200 ;
        RECT 54.000 1338.480 2870.580 1340.720 ;
        RECT 8.000 1338.000 2916.580 1338.480 ;
        RECT 54.000 1335.760 2870.580 1338.000 ;
        RECT 8.000 1335.280 2916.580 1335.760 ;
        RECT 54.000 1333.040 2870.580 1335.280 ;
        RECT 8.000 1332.560 2916.580 1333.040 ;
        RECT 54.000 1330.320 2870.580 1332.560 ;
        RECT 8.000 1329.840 2916.580 1330.320 ;
        RECT 54.000 1327.600 2870.580 1329.840 ;
        RECT 8.000 1327.120 2916.580 1327.600 ;
        RECT 54.000 1324.880 2870.580 1327.120 ;
        RECT 8.000 1324.400 2916.580 1324.880 ;
        RECT 54.000 1322.160 2870.580 1324.400 ;
        RECT 8.000 1321.680 2916.580 1322.160 ;
        RECT 54.000 1319.440 2870.580 1321.680 ;
        RECT 8.000 1318.960 2916.580 1319.440 ;
        RECT 54.000 1316.720 2870.580 1318.960 ;
        RECT 8.000 1316.240 2916.580 1316.720 ;
        RECT 54.000 1314.000 2870.580 1316.240 ;
        RECT 8.000 1313.520 2916.580 1314.000 ;
        RECT 54.000 1311.280 2870.580 1313.520 ;
        RECT 8.000 1310.800 2916.580 1311.280 ;
        RECT 54.000 1308.560 2870.580 1310.800 ;
        RECT 8.000 1308.080 2916.580 1308.560 ;
        RECT 54.000 1305.840 2870.580 1308.080 ;
        RECT 8.000 1305.360 2916.580 1305.840 ;
        RECT 54.000 1303.120 2870.580 1305.360 ;
        RECT 8.000 1302.640 2916.580 1303.120 ;
        RECT 54.000 1300.400 2870.580 1302.640 ;
        RECT 8.000 1299.920 2916.580 1300.400 ;
        RECT 54.000 1297.680 2870.580 1299.920 ;
        RECT 8.000 1297.200 2916.580 1297.680 ;
        RECT 54.000 1294.960 2870.580 1297.200 ;
        RECT 8.000 1294.480 2916.580 1294.960 ;
        RECT 54.000 1292.240 2870.580 1294.480 ;
        RECT 8.000 1291.760 2916.580 1292.240 ;
        RECT 54.000 1289.520 2870.580 1291.760 ;
        RECT 8.000 1289.040 2916.580 1289.520 ;
        RECT 54.000 1286.800 2870.580 1289.040 ;
        RECT 8.000 1286.320 2916.580 1286.800 ;
        RECT 54.000 1284.080 2870.580 1286.320 ;
        RECT 8.000 1283.600 2916.580 1284.080 ;
        RECT 54.000 1281.360 2870.580 1283.600 ;
        RECT 8.000 1280.880 2916.580 1281.360 ;
        RECT 54.000 1278.640 2870.580 1280.880 ;
        RECT 8.000 1278.160 2916.580 1278.640 ;
        RECT 54.000 1275.920 2870.580 1278.160 ;
        RECT 8.000 1275.440 2916.580 1275.920 ;
        RECT 54.000 1273.200 2870.580 1275.440 ;
        RECT 8.000 1272.720 2916.580 1273.200 ;
        RECT 54.000 1270.480 2870.580 1272.720 ;
        RECT 8.000 1270.000 2916.580 1270.480 ;
        RECT 54.000 1267.760 2870.580 1270.000 ;
        RECT 8.000 1267.280 2916.580 1267.760 ;
        RECT 54.000 1265.040 2870.580 1267.280 ;
        RECT 8.000 1264.560 2916.580 1265.040 ;
        RECT 54.000 1262.320 2870.580 1264.560 ;
        RECT 8.000 1261.840 2916.580 1262.320 ;
        RECT 54.000 1259.600 2870.580 1261.840 ;
        RECT 8.000 1259.120 2916.580 1259.600 ;
        RECT 54.000 1256.880 2870.580 1259.120 ;
        RECT 8.000 1256.400 2916.580 1256.880 ;
        RECT 54.000 1254.160 2870.580 1256.400 ;
        RECT 8.000 1253.680 2916.580 1254.160 ;
        RECT 54.000 1251.440 2870.580 1253.680 ;
        RECT 8.000 1250.960 2916.580 1251.440 ;
        RECT 54.000 1248.720 2870.580 1250.960 ;
        RECT 8.000 1248.240 2916.580 1248.720 ;
        RECT 54.000 1246.000 2870.580 1248.240 ;
        RECT 8.000 1245.520 2916.580 1246.000 ;
        RECT 54.000 1243.280 2870.580 1245.520 ;
        RECT 8.000 1242.800 2916.580 1243.280 ;
        RECT 54.000 1240.560 2870.580 1242.800 ;
        RECT 8.000 1240.080 2916.580 1240.560 ;
        RECT 54.000 1237.840 2870.580 1240.080 ;
        RECT 8.000 1237.360 2916.580 1237.840 ;
        RECT 54.000 1235.120 2870.580 1237.360 ;
        RECT 8.000 1234.640 2916.580 1235.120 ;
        RECT 54.000 1232.400 2870.580 1234.640 ;
        RECT 8.000 1231.920 2916.580 1232.400 ;
        RECT 54.000 1229.680 2870.580 1231.920 ;
        RECT 8.000 1229.200 2916.580 1229.680 ;
        RECT 54.000 1226.960 2870.580 1229.200 ;
        RECT 8.000 1226.480 2916.580 1226.960 ;
        RECT 54.000 1224.240 2870.580 1226.480 ;
        RECT 8.000 1223.760 2916.580 1224.240 ;
        RECT 54.000 1221.520 2870.580 1223.760 ;
        RECT 8.000 1221.040 2916.580 1221.520 ;
        RECT 54.000 1218.800 2870.580 1221.040 ;
        RECT 8.000 1218.320 2916.580 1218.800 ;
        RECT 54.000 1216.080 2870.580 1218.320 ;
        RECT 8.000 1215.600 2916.580 1216.080 ;
        RECT 54.000 1213.360 2870.580 1215.600 ;
        RECT 8.000 1212.880 2916.580 1213.360 ;
        RECT 54.000 1210.640 2870.580 1212.880 ;
        RECT 8.000 1210.160 2916.580 1210.640 ;
        RECT 54.000 1207.920 2870.580 1210.160 ;
        RECT 8.000 1207.440 2916.580 1207.920 ;
        RECT 54.000 1205.200 2870.580 1207.440 ;
        RECT 8.000 1204.720 2916.580 1205.200 ;
        RECT 54.000 1202.480 2870.580 1204.720 ;
        RECT 8.000 1202.000 2916.580 1202.480 ;
        RECT 54.000 1199.760 2870.580 1202.000 ;
        RECT 8.000 1199.280 2916.580 1199.760 ;
        RECT 54.000 1197.040 2870.580 1199.280 ;
        RECT 8.000 1196.560 2916.580 1197.040 ;
        RECT 54.000 1194.320 2870.580 1196.560 ;
        RECT 8.000 1193.840 2916.580 1194.320 ;
        RECT 54.000 1191.600 2870.580 1193.840 ;
        RECT 8.000 1191.120 2916.580 1191.600 ;
        RECT 54.000 1188.880 2870.580 1191.120 ;
        RECT 8.000 1188.400 2916.580 1188.880 ;
        RECT 54.000 1186.160 2870.580 1188.400 ;
        RECT 8.000 1185.680 2916.580 1186.160 ;
        RECT 54.000 1183.440 2870.580 1185.680 ;
        RECT 8.000 1182.960 2916.580 1183.440 ;
        RECT 54.000 1180.720 2870.580 1182.960 ;
        RECT 8.000 1180.240 2916.580 1180.720 ;
        RECT 54.000 1178.000 2870.580 1180.240 ;
        RECT 8.000 1177.520 2916.580 1178.000 ;
        RECT 54.000 1175.280 2870.580 1177.520 ;
        RECT 8.000 1174.800 2916.580 1175.280 ;
        RECT 54.000 1172.560 2870.580 1174.800 ;
        RECT 8.000 1172.080 2916.580 1172.560 ;
        RECT 54.000 1169.840 2870.580 1172.080 ;
        RECT 8.000 1169.360 2916.580 1169.840 ;
        RECT 54.000 1167.120 2870.580 1169.360 ;
        RECT 8.000 1166.640 2916.580 1167.120 ;
        RECT 54.000 1164.400 2870.580 1166.640 ;
        RECT 8.000 1163.920 2916.580 1164.400 ;
        RECT 54.000 1161.680 2870.580 1163.920 ;
        RECT 8.000 1161.200 2916.580 1161.680 ;
        RECT 54.000 1158.960 2870.580 1161.200 ;
        RECT 8.000 1158.480 2916.580 1158.960 ;
        RECT 54.000 1156.240 2870.580 1158.480 ;
        RECT 8.000 1155.760 2916.580 1156.240 ;
        RECT 54.000 1153.520 2870.580 1155.760 ;
        RECT 8.000 1153.040 2916.580 1153.520 ;
        RECT 54.000 1150.800 2870.580 1153.040 ;
        RECT 8.000 1150.320 2916.580 1150.800 ;
        RECT 54.000 1148.080 2870.580 1150.320 ;
        RECT 8.000 1147.600 2916.580 1148.080 ;
        RECT 54.000 1145.360 2870.580 1147.600 ;
        RECT 8.000 1144.880 2916.580 1145.360 ;
        RECT 54.000 1142.640 2870.580 1144.880 ;
        RECT 8.000 1142.160 2916.580 1142.640 ;
        RECT 54.000 1139.920 2870.580 1142.160 ;
        RECT 8.000 1139.440 2916.580 1139.920 ;
        RECT 54.000 1137.200 2870.580 1139.440 ;
        RECT 8.000 1136.720 2916.580 1137.200 ;
        RECT 54.000 1134.480 2870.580 1136.720 ;
        RECT 8.000 1134.000 2916.580 1134.480 ;
        RECT 54.000 1131.760 2870.580 1134.000 ;
        RECT 8.000 1131.280 2916.580 1131.760 ;
        RECT 54.000 1129.040 2870.580 1131.280 ;
        RECT 8.000 1128.560 2916.580 1129.040 ;
        RECT 54.000 1126.320 2870.580 1128.560 ;
        RECT 8.000 1125.840 2916.580 1126.320 ;
        RECT 54.000 1123.600 2870.580 1125.840 ;
        RECT 8.000 1123.120 2916.580 1123.600 ;
        RECT 54.000 1120.880 2870.580 1123.120 ;
        RECT 8.000 1120.400 2916.580 1120.880 ;
        RECT 54.000 1118.160 2870.580 1120.400 ;
        RECT 8.000 1117.680 2916.580 1118.160 ;
        RECT 54.000 1115.440 2870.580 1117.680 ;
        RECT 8.000 1114.960 2916.580 1115.440 ;
        RECT 54.000 1112.720 2870.580 1114.960 ;
        RECT 8.000 1112.240 2916.580 1112.720 ;
        RECT 54.000 1110.000 2870.580 1112.240 ;
        RECT 8.000 1109.520 2916.580 1110.000 ;
        RECT 54.000 1107.280 2870.580 1109.520 ;
        RECT 8.000 1106.800 2916.580 1107.280 ;
        RECT 54.000 1104.560 2870.580 1106.800 ;
        RECT 8.000 1104.080 2916.580 1104.560 ;
        RECT 54.000 1101.840 2870.580 1104.080 ;
        RECT 8.000 1101.360 2916.580 1101.840 ;
        RECT 54.000 1099.120 2870.580 1101.360 ;
        RECT 8.000 1098.640 2916.580 1099.120 ;
        RECT 54.000 1096.400 2870.580 1098.640 ;
        RECT 8.000 1095.920 2916.580 1096.400 ;
        RECT 54.000 1093.680 2870.580 1095.920 ;
        RECT 8.000 1093.200 2916.580 1093.680 ;
        RECT 54.000 1090.960 2870.580 1093.200 ;
        RECT 8.000 1090.480 2916.580 1090.960 ;
        RECT 54.000 1088.240 2870.580 1090.480 ;
        RECT 8.000 1087.760 2916.580 1088.240 ;
        RECT 54.000 1085.520 2870.580 1087.760 ;
        RECT 8.000 1085.040 2916.580 1085.520 ;
        RECT 54.000 1082.800 2870.580 1085.040 ;
        RECT 8.000 1082.320 2916.580 1082.800 ;
        RECT 54.000 1080.080 2870.580 1082.320 ;
        RECT 8.000 1079.600 2916.580 1080.080 ;
        RECT 54.000 1077.360 2870.580 1079.600 ;
        RECT 8.000 1076.880 2916.580 1077.360 ;
        RECT 54.000 1074.640 2870.580 1076.880 ;
        RECT 8.000 1074.160 2916.580 1074.640 ;
        RECT 54.000 1071.920 2870.580 1074.160 ;
        RECT 8.000 1071.440 2916.580 1071.920 ;
        RECT 54.000 1069.200 2870.580 1071.440 ;
        RECT 8.000 1068.720 2916.580 1069.200 ;
        RECT 54.000 1066.480 2870.580 1068.720 ;
        RECT 8.000 1066.000 2916.580 1066.480 ;
        RECT 54.000 1063.760 2870.580 1066.000 ;
        RECT 8.000 1063.280 2916.580 1063.760 ;
        RECT 54.000 1061.040 2870.580 1063.280 ;
        RECT 8.000 1060.560 2916.580 1061.040 ;
        RECT 54.000 1058.320 2870.580 1060.560 ;
        RECT 8.000 1057.840 2916.580 1058.320 ;
        RECT 54.000 1055.600 2870.580 1057.840 ;
        RECT 8.000 1055.120 2916.580 1055.600 ;
        RECT 54.000 1052.880 2870.580 1055.120 ;
        RECT 8.000 1052.400 2916.580 1052.880 ;
        RECT 54.000 1050.160 2870.580 1052.400 ;
        RECT 8.000 1049.680 2916.580 1050.160 ;
        RECT 54.000 1047.440 2870.580 1049.680 ;
        RECT 8.000 1046.960 2916.580 1047.440 ;
        RECT 54.000 1044.720 2870.580 1046.960 ;
        RECT 8.000 1044.240 2916.580 1044.720 ;
        RECT 54.000 1042.000 2870.580 1044.240 ;
        RECT 8.000 1041.520 2916.580 1042.000 ;
        RECT 54.000 1039.280 2870.580 1041.520 ;
        RECT 8.000 1038.800 2916.580 1039.280 ;
        RECT 54.000 1036.560 2870.580 1038.800 ;
        RECT 8.000 1036.080 2916.580 1036.560 ;
        RECT 54.000 1033.840 2870.580 1036.080 ;
        RECT 8.000 1033.360 2916.580 1033.840 ;
        RECT 54.000 1031.120 2870.580 1033.360 ;
        RECT 8.000 1030.640 2916.580 1031.120 ;
        RECT 54.000 1028.400 2870.580 1030.640 ;
        RECT 8.000 1027.920 2916.580 1028.400 ;
        RECT 54.000 1025.680 2870.580 1027.920 ;
        RECT 8.000 1025.200 2916.580 1025.680 ;
        RECT 54.000 1022.960 2870.580 1025.200 ;
        RECT 8.000 1022.480 2916.580 1022.960 ;
        RECT 54.000 1020.240 2870.580 1022.480 ;
        RECT 8.000 1019.760 2916.580 1020.240 ;
        RECT 54.000 1017.520 2870.580 1019.760 ;
        RECT 8.000 1017.040 2916.580 1017.520 ;
        RECT 54.000 1014.800 2870.580 1017.040 ;
        RECT 8.000 1014.320 2916.580 1014.800 ;
        RECT 54.000 1012.080 2870.580 1014.320 ;
        RECT 8.000 1011.600 2916.580 1012.080 ;
        RECT 54.000 1009.360 2870.580 1011.600 ;
        RECT 8.000 1008.880 2916.580 1009.360 ;
        RECT 54.000 1006.640 2870.580 1008.880 ;
        RECT 8.000 1006.160 2916.580 1006.640 ;
        RECT 54.000 1003.920 2870.580 1006.160 ;
        RECT 8.000 1003.440 2916.580 1003.920 ;
        RECT 54.000 1001.200 2870.580 1003.440 ;
        RECT 8.000 1000.720 2916.580 1001.200 ;
        RECT 54.000 998.480 2870.580 1000.720 ;
        RECT 8.000 998.000 2916.580 998.480 ;
        RECT 54.000 995.760 2870.580 998.000 ;
        RECT 8.000 995.280 2916.580 995.760 ;
        RECT 54.000 993.040 2870.580 995.280 ;
        RECT 8.000 992.560 2916.580 993.040 ;
        RECT 54.000 990.320 2870.580 992.560 ;
        RECT 8.000 989.840 2916.580 990.320 ;
        RECT 54.000 987.600 2870.580 989.840 ;
        RECT 8.000 987.120 2916.580 987.600 ;
        RECT 54.000 984.880 2870.580 987.120 ;
        RECT 8.000 984.400 2916.580 984.880 ;
        RECT 54.000 982.160 2870.580 984.400 ;
        RECT 8.000 981.680 2916.580 982.160 ;
        RECT 54.000 979.440 2870.580 981.680 ;
        RECT 8.000 978.960 2916.580 979.440 ;
        RECT 54.000 976.720 2870.580 978.960 ;
        RECT 8.000 976.240 2916.580 976.720 ;
        RECT 54.000 974.000 2870.580 976.240 ;
        RECT 8.000 973.520 2916.580 974.000 ;
        RECT 54.000 971.280 2870.580 973.520 ;
        RECT 8.000 970.800 2916.580 971.280 ;
        RECT 54.000 968.560 2870.580 970.800 ;
        RECT 8.000 968.080 2916.580 968.560 ;
        RECT 54.000 965.840 2870.580 968.080 ;
        RECT 8.000 965.360 2916.580 965.840 ;
        RECT 54.000 963.120 2870.580 965.360 ;
        RECT 8.000 962.640 2916.580 963.120 ;
        RECT 54.000 960.400 2870.580 962.640 ;
        RECT 8.000 959.920 2916.580 960.400 ;
        RECT 54.000 957.680 2870.580 959.920 ;
        RECT 8.000 957.200 2916.580 957.680 ;
        RECT 54.000 954.960 2870.580 957.200 ;
        RECT 8.000 954.480 2916.580 954.960 ;
        RECT 54.000 952.240 2870.580 954.480 ;
        RECT 8.000 951.760 2916.580 952.240 ;
        RECT 54.000 949.520 2870.580 951.760 ;
        RECT 8.000 949.040 2916.580 949.520 ;
        RECT 54.000 946.800 2870.580 949.040 ;
        RECT 8.000 946.320 2916.580 946.800 ;
        RECT 54.000 944.080 2870.580 946.320 ;
        RECT 8.000 943.600 2916.580 944.080 ;
        RECT 54.000 941.360 2870.580 943.600 ;
        RECT 8.000 940.880 2916.580 941.360 ;
        RECT 54.000 938.640 2870.580 940.880 ;
        RECT 8.000 938.160 2916.580 938.640 ;
        RECT 54.000 935.920 2870.580 938.160 ;
        RECT 8.000 935.440 2916.580 935.920 ;
        RECT 54.000 933.200 2870.580 935.440 ;
        RECT 8.000 932.720 2916.580 933.200 ;
        RECT 54.000 930.480 2870.580 932.720 ;
        RECT 8.000 930.000 2916.580 930.480 ;
        RECT 54.000 927.760 2870.580 930.000 ;
        RECT 8.000 927.280 2916.580 927.760 ;
        RECT 54.000 925.040 2870.580 927.280 ;
        RECT 8.000 924.560 2916.580 925.040 ;
        RECT 54.000 922.320 2870.580 924.560 ;
        RECT 8.000 921.840 2916.580 922.320 ;
        RECT 54.000 919.600 2870.580 921.840 ;
        RECT 8.000 919.120 2916.580 919.600 ;
        RECT 54.000 916.880 2870.580 919.120 ;
        RECT 8.000 916.400 2916.580 916.880 ;
        RECT 54.000 914.160 2870.580 916.400 ;
        RECT 8.000 913.680 2916.580 914.160 ;
        RECT 54.000 911.440 2870.580 913.680 ;
        RECT 8.000 910.960 2916.580 911.440 ;
        RECT 54.000 908.720 2870.580 910.960 ;
        RECT 8.000 908.240 2916.580 908.720 ;
        RECT 54.000 906.000 2870.580 908.240 ;
        RECT 8.000 905.520 2916.580 906.000 ;
        RECT 54.000 903.280 2870.580 905.520 ;
        RECT 8.000 902.800 2916.580 903.280 ;
        RECT 54.000 900.560 2870.580 902.800 ;
        RECT 8.000 900.080 2916.580 900.560 ;
        RECT 54.000 897.840 2870.580 900.080 ;
        RECT 8.000 897.360 2916.580 897.840 ;
        RECT 54.000 895.120 2870.580 897.360 ;
        RECT 8.000 894.640 2916.580 895.120 ;
        RECT 54.000 892.400 2870.580 894.640 ;
        RECT 8.000 891.920 2916.580 892.400 ;
        RECT 54.000 889.680 2870.580 891.920 ;
        RECT 8.000 889.200 2916.580 889.680 ;
        RECT 54.000 886.960 2870.580 889.200 ;
        RECT 8.000 886.480 2916.580 886.960 ;
        RECT 54.000 884.240 2870.580 886.480 ;
        RECT 8.000 883.760 2916.580 884.240 ;
        RECT 54.000 881.520 2870.580 883.760 ;
        RECT 8.000 881.040 2916.580 881.520 ;
        RECT 54.000 878.800 2870.580 881.040 ;
        RECT 8.000 878.320 2916.580 878.800 ;
        RECT 54.000 876.080 2870.580 878.320 ;
        RECT 8.000 875.600 2916.580 876.080 ;
        RECT 54.000 873.360 2870.580 875.600 ;
        RECT 8.000 872.880 2916.580 873.360 ;
        RECT 54.000 870.640 2870.580 872.880 ;
        RECT 8.000 870.160 2916.580 870.640 ;
        RECT 54.000 867.920 2870.580 870.160 ;
        RECT 8.000 867.440 2916.580 867.920 ;
        RECT 54.000 865.200 2870.580 867.440 ;
        RECT 8.000 864.720 2916.580 865.200 ;
        RECT 54.000 862.480 2870.580 864.720 ;
        RECT 8.000 862.000 2916.580 862.480 ;
        RECT 54.000 859.760 2870.580 862.000 ;
        RECT 8.000 859.280 2916.580 859.760 ;
        RECT 54.000 857.040 2870.580 859.280 ;
        RECT 8.000 856.560 2916.580 857.040 ;
        RECT 54.000 854.320 2870.580 856.560 ;
        RECT 8.000 853.840 2916.580 854.320 ;
        RECT 54.000 851.600 2870.580 853.840 ;
        RECT 8.000 851.120 2916.580 851.600 ;
        RECT 54.000 848.880 2870.580 851.120 ;
        RECT 8.000 848.400 2916.580 848.880 ;
        RECT 54.000 846.160 2870.580 848.400 ;
        RECT 8.000 845.680 2916.580 846.160 ;
        RECT 54.000 843.440 2870.580 845.680 ;
        RECT 8.000 842.960 2916.580 843.440 ;
        RECT 54.000 840.720 2870.580 842.960 ;
        RECT 8.000 840.240 2916.580 840.720 ;
        RECT 54.000 838.000 2870.580 840.240 ;
        RECT 8.000 837.520 2916.580 838.000 ;
        RECT 54.000 835.280 2870.580 837.520 ;
        RECT 8.000 834.800 2916.580 835.280 ;
        RECT 54.000 832.560 2870.580 834.800 ;
        RECT 8.000 832.080 2916.580 832.560 ;
        RECT 54.000 829.840 2870.580 832.080 ;
        RECT 8.000 829.360 2916.580 829.840 ;
        RECT 54.000 827.120 2870.580 829.360 ;
        RECT 8.000 826.640 2916.580 827.120 ;
        RECT 54.000 824.400 2870.580 826.640 ;
        RECT 8.000 823.920 2916.580 824.400 ;
        RECT 54.000 821.680 2870.580 823.920 ;
        RECT 8.000 821.200 2916.580 821.680 ;
        RECT 54.000 818.960 2870.580 821.200 ;
        RECT 8.000 818.480 2916.580 818.960 ;
        RECT 54.000 816.240 2870.580 818.480 ;
        RECT 8.000 815.760 2916.580 816.240 ;
        RECT 54.000 813.520 2870.580 815.760 ;
        RECT 8.000 813.040 2916.580 813.520 ;
        RECT 54.000 810.800 2870.580 813.040 ;
        RECT 8.000 810.320 2916.580 810.800 ;
        RECT 54.000 808.080 2870.580 810.320 ;
        RECT 8.000 807.600 2916.580 808.080 ;
        RECT 54.000 805.360 2870.580 807.600 ;
        RECT 8.000 804.880 2916.580 805.360 ;
        RECT 54.000 802.640 2870.580 804.880 ;
        RECT 8.000 802.160 2916.580 802.640 ;
        RECT 54.000 799.920 2870.580 802.160 ;
        RECT 8.000 799.440 2916.580 799.920 ;
        RECT 54.000 797.200 2870.580 799.440 ;
        RECT 8.000 796.720 2916.580 797.200 ;
        RECT 54.000 794.480 2870.580 796.720 ;
        RECT 8.000 794.000 2916.580 794.480 ;
        RECT 54.000 791.760 2870.580 794.000 ;
        RECT 8.000 791.280 2916.580 791.760 ;
        RECT 54.000 789.040 2870.580 791.280 ;
        RECT 8.000 788.560 2916.580 789.040 ;
        RECT 54.000 786.320 2870.580 788.560 ;
        RECT 8.000 785.840 2916.580 786.320 ;
        RECT 54.000 783.600 2870.580 785.840 ;
        RECT 8.000 783.120 2916.580 783.600 ;
        RECT 54.000 780.880 2870.580 783.120 ;
        RECT 8.000 780.400 2916.580 780.880 ;
        RECT 54.000 778.160 2870.580 780.400 ;
        RECT 8.000 777.680 2916.580 778.160 ;
        RECT 54.000 775.440 2870.580 777.680 ;
        RECT 8.000 774.960 2916.580 775.440 ;
        RECT 54.000 772.720 2870.580 774.960 ;
        RECT 8.000 772.240 2916.580 772.720 ;
        RECT 54.000 770.000 2870.580 772.240 ;
        RECT 8.000 769.520 2916.580 770.000 ;
        RECT 54.000 767.280 2870.580 769.520 ;
        RECT 8.000 766.800 2916.580 767.280 ;
        RECT 54.000 764.560 2870.580 766.800 ;
        RECT 8.000 764.080 2916.580 764.560 ;
        RECT 54.000 761.840 2870.580 764.080 ;
        RECT 8.000 761.360 2916.580 761.840 ;
        RECT 54.000 759.120 2870.580 761.360 ;
        RECT 8.000 758.640 2916.580 759.120 ;
        RECT 54.000 756.400 2870.580 758.640 ;
        RECT 8.000 755.920 2916.580 756.400 ;
        RECT 54.000 753.680 2870.580 755.920 ;
        RECT 8.000 753.200 2916.580 753.680 ;
        RECT 54.000 750.960 2870.580 753.200 ;
        RECT 8.000 750.480 2916.580 750.960 ;
        RECT 54.000 748.240 2870.580 750.480 ;
        RECT 8.000 747.760 2916.580 748.240 ;
        RECT 54.000 745.520 2870.580 747.760 ;
        RECT 8.000 745.040 2916.580 745.520 ;
        RECT 54.000 742.800 2870.580 745.040 ;
        RECT 8.000 742.320 2916.580 742.800 ;
        RECT 54.000 740.080 2870.580 742.320 ;
        RECT 8.000 739.600 2916.580 740.080 ;
        RECT 54.000 737.360 2870.580 739.600 ;
        RECT 8.000 736.880 2916.580 737.360 ;
        RECT 54.000 734.640 2870.580 736.880 ;
        RECT 8.000 734.160 2916.580 734.640 ;
        RECT 54.000 731.920 2870.580 734.160 ;
        RECT 8.000 731.440 2916.580 731.920 ;
        RECT 54.000 729.200 2870.580 731.440 ;
        RECT 8.000 728.720 2916.580 729.200 ;
        RECT 54.000 726.480 2870.580 728.720 ;
        RECT 8.000 726.000 2916.580 726.480 ;
        RECT 54.000 723.760 2870.580 726.000 ;
        RECT 8.000 723.280 2916.580 723.760 ;
        RECT 54.000 721.040 2870.580 723.280 ;
        RECT 8.000 720.560 2916.580 721.040 ;
        RECT 54.000 718.320 2870.580 720.560 ;
        RECT 8.000 717.840 2916.580 718.320 ;
        RECT 54.000 715.600 2870.580 717.840 ;
        RECT 8.000 715.120 2916.580 715.600 ;
        RECT 54.000 712.880 2870.580 715.120 ;
        RECT 8.000 712.400 2916.580 712.880 ;
        RECT 54.000 710.160 2870.580 712.400 ;
        RECT 8.000 709.680 2916.580 710.160 ;
        RECT 54.000 707.440 2870.580 709.680 ;
        RECT 8.000 706.960 2916.580 707.440 ;
        RECT 54.000 704.720 2870.580 706.960 ;
        RECT 8.000 704.240 2916.580 704.720 ;
        RECT 54.000 702.000 2870.580 704.240 ;
        RECT 8.000 701.520 2916.580 702.000 ;
        RECT 54.000 699.280 2870.580 701.520 ;
        RECT 8.000 698.800 2916.580 699.280 ;
        RECT 54.000 696.560 2870.580 698.800 ;
        RECT 8.000 696.080 2916.580 696.560 ;
        RECT 54.000 693.840 2870.580 696.080 ;
        RECT 8.000 693.360 2916.580 693.840 ;
        RECT 54.000 691.120 2870.580 693.360 ;
        RECT 8.000 690.640 2916.580 691.120 ;
        RECT 54.000 688.400 2870.580 690.640 ;
        RECT 8.000 687.920 2916.580 688.400 ;
        RECT 54.000 685.680 2870.580 687.920 ;
        RECT 8.000 685.200 2916.580 685.680 ;
        RECT 54.000 682.960 2870.580 685.200 ;
        RECT 8.000 682.480 2916.580 682.960 ;
        RECT 54.000 680.240 2870.580 682.480 ;
        RECT 8.000 679.760 2916.580 680.240 ;
        RECT 54.000 677.520 2870.580 679.760 ;
        RECT 8.000 677.040 2916.580 677.520 ;
        RECT 54.000 674.800 2870.580 677.040 ;
        RECT 8.000 674.320 2916.580 674.800 ;
        RECT 54.000 672.080 2870.580 674.320 ;
        RECT 8.000 671.600 2916.580 672.080 ;
        RECT 54.000 669.360 2870.580 671.600 ;
        RECT 8.000 668.880 2916.580 669.360 ;
        RECT 54.000 666.640 2870.580 668.880 ;
        RECT 8.000 666.160 2916.580 666.640 ;
        RECT 54.000 663.920 2870.580 666.160 ;
        RECT 8.000 663.440 2916.580 663.920 ;
        RECT 54.000 661.200 2870.580 663.440 ;
        RECT 8.000 660.720 2916.580 661.200 ;
        RECT 54.000 658.480 2870.580 660.720 ;
        RECT 8.000 658.000 2916.580 658.480 ;
        RECT 54.000 655.760 2870.580 658.000 ;
        RECT 8.000 655.280 2916.580 655.760 ;
        RECT 54.000 653.040 2870.580 655.280 ;
        RECT 8.000 652.560 2916.580 653.040 ;
        RECT 54.000 650.320 2870.580 652.560 ;
        RECT 8.000 649.840 2916.580 650.320 ;
        RECT 54.000 647.600 2870.580 649.840 ;
        RECT 8.000 647.120 2916.580 647.600 ;
        RECT 54.000 644.880 2870.580 647.120 ;
        RECT 8.000 644.400 2916.580 644.880 ;
        RECT 54.000 642.160 2870.580 644.400 ;
        RECT 8.000 641.680 2916.580 642.160 ;
        RECT 54.000 639.440 2870.580 641.680 ;
        RECT 8.000 638.960 2916.580 639.440 ;
        RECT 54.000 636.720 2870.580 638.960 ;
        RECT 8.000 636.240 2916.580 636.720 ;
        RECT 54.000 634.000 2870.580 636.240 ;
        RECT 8.000 633.520 2916.580 634.000 ;
        RECT 54.000 631.280 2870.580 633.520 ;
        RECT 8.000 630.800 2916.580 631.280 ;
        RECT 54.000 628.560 2870.580 630.800 ;
        RECT 8.000 628.080 2916.580 628.560 ;
        RECT 54.000 625.840 2870.580 628.080 ;
        RECT 8.000 625.360 2916.580 625.840 ;
        RECT 54.000 623.120 2870.580 625.360 ;
        RECT 8.000 622.640 2916.580 623.120 ;
        RECT 54.000 620.400 2870.580 622.640 ;
        RECT 8.000 619.920 2916.580 620.400 ;
        RECT 54.000 617.680 2870.580 619.920 ;
        RECT 8.000 617.200 2916.580 617.680 ;
        RECT 54.000 614.960 2870.580 617.200 ;
        RECT 8.000 614.480 2916.580 614.960 ;
        RECT 54.000 612.240 2870.580 614.480 ;
        RECT 8.000 611.760 2916.580 612.240 ;
        RECT 54.000 609.520 2870.580 611.760 ;
        RECT 8.000 609.040 2916.580 609.520 ;
        RECT 54.000 606.800 2870.580 609.040 ;
        RECT 8.000 606.320 2916.580 606.800 ;
        RECT 54.000 604.080 2870.580 606.320 ;
        RECT 8.000 603.600 2916.580 604.080 ;
        RECT 54.000 601.360 2870.580 603.600 ;
        RECT 8.000 600.880 2916.580 601.360 ;
        RECT 54.000 598.640 2870.580 600.880 ;
        RECT 8.000 598.160 2916.580 598.640 ;
        RECT 54.000 595.920 2870.580 598.160 ;
        RECT 8.000 595.440 2916.580 595.920 ;
        RECT 54.000 593.200 2870.580 595.440 ;
        RECT 8.000 592.720 2916.580 593.200 ;
        RECT 54.000 590.480 2870.580 592.720 ;
        RECT 8.000 590.000 2916.580 590.480 ;
        RECT 54.000 587.760 2870.580 590.000 ;
        RECT 8.000 587.280 2916.580 587.760 ;
        RECT 54.000 585.040 2870.580 587.280 ;
        RECT 8.000 584.560 2916.580 585.040 ;
        RECT 54.000 582.320 2870.580 584.560 ;
        RECT 8.000 581.840 2916.580 582.320 ;
        RECT 54.000 579.600 2870.580 581.840 ;
        RECT 8.000 579.120 2916.580 579.600 ;
        RECT 54.000 576.880 2870.580 579.120 ;
        RECT 8.000 576.400 2916.580 576.880 ;
        RECT 54.000 574.160 2870.580 576.400 ;
        RECT 8.000 573.680 2916.580 574.160 ;
        RECT 54.000 571.440 2870.580 573.680 ;
        RECT 8.000 570.960 2916.580 571.440 ;
        RECT 54.000 568.720 2870.580 570.960 ;
        RECT 8.000 568.240 2916.580 568.720 ;
        RECT 54.000 566.000 2870.580 568.240 ;
        RECT 8.000 565.520 2916.580 566.000 ;
        RECT 54.000 563.280 2870.580 565.520 ;
        RECT 8.000 562.800 2916.580 563.280 ;
        RECT 54.000 560.560 2870.580 562.800 ;
        RECT 8.000 560.080 2916.580 560.560 ;
        RECT 54.000 557.840 2870.580 560.080 ;
        RECT 8.000 557.360 2916.580 557.840 ;
        RECT 54.000 555.120 2870.580 557.360 ;
        RECT 8.000 554.640 2916.580 555.120 ;
        RECT 54.000 552.400 2870.580 554.640 ;
        RECT 8.000 551.920 2916.580 552.400 ;
        RECT 54.000 549.680 2870.580 551.920 ;
        RECT 8.000 549.200 2916.580 549.680 ;
        RECT 54.000 546.960 2870.580 549.200 ;
        RECT 8.000 546.480 2916.580 546.960 ;
        RECT 54.000 544.240 2870.580 546.480 ;
        RECT 8.000 543.760 2916.580 544.240 ;
        RECT 54.000 541.520 2870.580 543.760 ;
        RECT 8.000 541.040 2916.580 541.520 ;
        RECT 54.000 538.800 2870.580 541.040 ;
        RECT 8.000 538.320 2916.580 538.800 ;
        RECT 54.000 536.080 2870.580 538.320 ;
        RECT 8.000 535.600 2916.580 536.080 ;
        RECT 54.000 533.360 2870.580 535.600 ;
        RECT 8.000 532.880 2916.580 533.360 ;
        RECT 54.000 530.640 2870.580 532.880 ;
        RECT 8.000 530.160 2916.580 530.640 ;
        RECT 54.000 527.920 2870.580 530.160 ;
        RECT 8.000 527.440 2916.580 527.920 ;
        RECT 54.000 525.200 2870.580 527.440 ;
        RECT 8.000 524.720 2916.580 525.200 ;
        RECT 54.000 522.480 2870.580 524.720 ;
        RECT 8.000 522.000 2916.580 522.480 ;
        RECT 54.000 519.760 2870.580 522.000 ;
        RECT 8.000 519.280 2916.580 519.760 ;
        RECT 54.000 517.040 2870.580 519.280 ;
        RECT 8.000 516.560 2916.580 517.040 ;
        RECT 54.000 514.320 2870.580 516.560 ;
        RECT 8.000 513.840 2916.580 514.320 ;
        RECT 54.000 511.600 2870.580 513.840 ;
        RECT 8.000 511.120 2916.580 511.600 ;
        RECT 54.000 508.880 2870.580 511.120 ;
        RECT 8.000 508.400 2916.580 508.880 ;
        RECT 54.000 506.160 2870.580 508.400 ;
        RECT 8.000 505.680 2916.580 506.160 ;
        RECT 54.000 503.440 2870.580 505.680 ;
        RECT 8.000 502.960 2916.580 503.440 ;
        RECT 54.000 500.720 2870.580 502.960 ;
        RECT 8.000 500.240 2916.580 500.720 ;
        RECT 54.000 498.000 2870.580 500.240 ;
        RECT 8.000 497.520 2916.580 498.000 ;
        RECT 54.000 495.280 2870.580 497.520 ;
        RECT 8.000 494.800 2916.580 495.280 ;
        RECT 54.000 492.560 2870.580 494.800 ;
        RECT 8.000 492.080 2916.580 492.560 ;
        RECT 54.000 489.840 2870.580 492.080 ;
        RECT 8.000 489.360 2916.580 489.840 ;
        RECT 54.000 487.120 2870.580 489.360 ;
        RECT 8.000 486.640 2916.580 487.120 ;
        RECT 54.000 484.400 2870.580 486.640 ;
        RECT 8.000 483.920 2916.580 484.400 ;
        RECT 54.000 481.680 2870.580 483.920 ;
        RECT 8.000 481.200 2916.580 481.680 ;
        RECT 54.000 478.960 2870.580 481.200 ;
        RECT 8.000 478.480 2916.580 478.960 ;
        RECT 54.000 476.240 2870.580 478.480 ;
        RECT 8.000 475.760 2916.580 476.240 ;
        RECT 54.000 473.520 2870.580 475.760 ;
        RECT 8.000 473.040 2916.580 473.520 ;
        RECT 54.000 470.800 2870.580 473.040 ;
        RECT 8.000 470.320 2916.580 470.800 ;
        RECT 54.000 468.080 2870.580 470.320 ;
        RECT 8.000 467.600 2916.580 468.080 ;
        RECT 54.000 465.360 2870.580 467.600 ;
        RECT 8.000 464.880 2916.580 465.360 ;
        RECT 54.000 462.640 2870.580 464.880 ;
        RECT 8.000 462.160 2916.580 462.640 ;
        RECT 54.000 459.920 2870.580 462.160 ;
        RECT 8.000 459.440 2916.580 459.920 ;
        RECT 54.000 457.200 2870.580 459.440 ;
        RECT 8.000 456.720 2916.580 457.200 ;
        RECT 54.000 454.480 2870.580 456.720 ;
        RECT 8.000 454.000 2916.580 454.480 ;
        RECT 54.000 451.760 2870.580 454.000 ;
        RECT 8.000 451.280 2916.580 451.760 ;
        RECT 54.000 449.040 2870.580 451.280 ;
        RECT 8.000 448.560 2916.580 449.040 ;
        RECT 54.000 446.320 2870.580 448.560 ;
        RECT 8.000 445.840 2916.580 446.320 ;
        RECT 54.000 443.600 2870.580 445.840 ;
        RECT 8.000 443.120 2916.580 443.600 ;
        RECT 54.000 440.880 2870.580 443.120 ;
        RECT 8.000 440.400 2916.580 440.880 ;
        RECT 54.000 438.160 2870.580 440.400 ;
        RECT 8.000 437.680 2916.580 438.160 ;
        RECT 54.000 435.440 2870.580 437.680 ;
        RECT 8.000 434.960 2916.580 435.440 ;
        RECT 54.000 432.720 2870.580 434.960 ;
        RECT 8.000 432.240 2916.580 432.720 ;
        RECT 54.000 430.000 2870.580 432.240 ;
        RECT 8.000 429.520 2916.580 430.000 ;
        RECT 54.000 427.280 2870.580 429.520 ;
        RECT 8.000 426.800 2916.580 427.280 ;
        RECT 54.000 424.560 2870.580 426.800 ;
        RECT 8.000 424.080 2916.580 424.560 ;
        RECT 54.000 421.840 2870.580 424.080 ;
        RECT 8.000 421.360 2916.580 421.840 ;
        RECT 54.000 419.120 2870.580 421.360 ;
        RECT 8.000 418.640 2916.580 419.120 ;
        RECT 54.000 416.400 2870.580 418.640 ;
        RECT 8.000 415.920 2916.580 416.400 ;
        RECT 54.000 413.680 2870.580 415.920 ;
        RECT 8.000 413.200 2916.580 413.680 ;
        RECT 54.000 410.960 2870.580 413.200 ;
        RECT 8.000 410.480 2916.580 410.960 ;
        RECT 54.000 408.240 2870.580 410.480 ;
        RECT 8.000 407.760 2916.580 408.240 ;
        RECT 54.000 405.520 2870.580 407.760 ;
        RECT 8.000 405.040 2916.580 405.520 ;
        RECT 54.000 402.800 2870.580 405.040 ;
        RECT 8.000 402.320 2916.580 402.800 ;
        RECT 54.000 400.080 2870.580 402.320 ;
        RECT 8.000 399.600 2916.580 400.080 ;
        RECT 54.000 397.360 2870.580 399.600 ;
        RECT 8.000 396.880 2916.580 397.360 ;
        RECT 54.000 394.640 2870.580 396.880 ;
        RECT 8.000 394.160 2916.580 394.640 ;
        RECT 54.000 391.920 2870.580 394.160 ;
        RECT 8.000 391.440 2916.580 391.920 ;
        RECT 54.000 389.200 2870.580 391.440 ;
        RECT 8.000 388.720 2916.580 389.200 ;
        RECT 54.000 386.480 2870.580 388.720 ;
        RECT 8.000 386.000 2916.580 386.480 ;
        RECT 54.000 383.760 2870.580 386.000 ;
        RECT 8.000 383.280 2916.580 383.760 ;
        RECT 54.000 381.040 2870.580 383.280 ;
        RECT 8.000 380.560 2916.580 381.040 ;
        RECT 54.000 378.320 2870.580 380.560 ;
        RECT 8.000 377.840 2916.580 378.320 ;
        RECT 54.000 375.600 2870.580 377.840 ;
        RECT 8.000 375.120 2916.580 375.600 ;
        RECT 54.000 372.880 2870.580 375.120 ;
        RECT 8.000 372.400 2916.580 372.880 ;
        RECT 54.000 370.160 2870.580 372.400 ;
        RECT 8.000 369.680 2916.580 370.160 ;
        RECT 54.000 367.440 2870.580 369.680 ;
        RECT 8.000 366.960 2916.580 367.440 ;
        RECT 54.000 364.720 2870.580 366.960 ;
        RECT 8.000 364.240 2916.580 364.720 ;
        RECT 54.000 362.000 2870.580 364.240 ;
        RECT 8.000 361.520 2916.580 362.000 ;
        RECT 54.000 359.280 2870.580 361.520 ;
        RECT 8.000 358.800 2916.580 359.280 ;
        RECT 54.000 356.560 2870.580 358.800 ;
        RECT 8.000 356.080 2916.580 356.560 ;
        RECT 54.000 353.840 2870.580 356.080 ;
        RECT 8.000 353.360 2916.580 353.840 ;
        RECT 54.000 351.120 2870.580 353.360 ;
        RECT 8.000 350.640 2916.580 351.120 ;
        RECT 54.000 348.400 2870.580 350.640 ;
        RECT 8.000 347.920 2916.580 348.400 ;
        RECT 54.000 345.680 2870.580 347.920 ;
        RECT 8.000 345.200 2916.580 345.680 ;
        RECT 54.000 342.960 2870.580 345.200 ;
        RECT 8.000 342.480 2916.580 342.960 ;
        RECT 54.000 340.240 2870.580 342.480 ;
        RECT 8.000 339.760 2916.580 340.240 ;
        RECT 54.000 337.520 2870.580 339.760 ;
        RECT 8.000 337.040 2916.580 337.520 ;
        RECT 54.000 334.800 2870.580 337.040 ;
        RECT 8.000 334.320 2916.580 334.800 ;
        RECT 54.000 332.080 2870.580 334.320 ;
        RECT 8.000 331.600 2916.580 332.080 ;
        RECT 54.000 329.360 2870.580 331.600 ;
        RECT 8.000 328.880 2916.580 329.360 ;
        RECT 54.000 326.640 2870.580 328.880 ;
        RECT 8.000 326.160 2916.580 326.640 ;
        RECT 54.000 323.920 2870.580 326.160 ;
        RECT 8.000 323.440 2916.580 323.920 ;
        RECT 54.000 321.200 2870.580 323.440 ;
        RECT 8.000 320.720 2916.580 321.200 ;
        RECT 54.000 318.480 2870.580 320.720 ;
        RECT 8.000 318.000 2916.580 318.480 ;
        RECT 54.000 315.760 2870.580 318.000 ;
        RECT 8.000 315.280 2916.580 315.760 ;
        RECT 54.000 313.040 2870.580 315.280 ;
        RECT 8.000 312.560 2916.580 313.040 ;
        RECT 54.000 310.320 2870.580 312.560 ;
        RECT 8.000 309.840 2916.580 310.320 ;
        RECT 54.000 307.600 2870.580 309.840 ;
        RECT 8.000 307.120 2916.580 307.600 ;
        RECT 54.000 304.880 2870.580 307.120 ;
        RECT 8.000 304.400 2916.580 304.880 ;
        RECT 54.000 302.160 2870.580 304.400 ;
        RECT 8.000 301.680 2916.580 302.160 ;
        RECT 54.000 299.440 2870.580 301.680 ;
        RECT 8.000 298.960 2916.580 299.440 ;
        RECT 54.000 296.720 2870.580 298.960 ;
        RECT 8.000 296.240 2916.580 296.720 ;
        RECT 54.000 294.000 2870.580 296.240 ;
        RECT 8.000 293.520 2916.580 294.000 ;
        RECT 54.000 291.280 2870.580 293.520 ;
        RECT 8.000 290.800 2916.580 291.280 ;
        RECT 54.000 288.560 2870.580 290.800 ;
        RECT 8.000 288.080 2916.580 288.560 ;
        RECT 54.000 285.840 2870.580 288.080 ;
        RECT 8.000 285.360 2916.580 285.840 ;
        RECT 54.000 283.120 2870.580 285.360 ;
        RECT 8.000 282.640 2916.580 283.120 ;
        RECT 54.000 280.400 2870.580 282.640 ;
        RECT 8.000 279.920 2916.580 280.400 ;
        RECT 54.000 277.680 2870.580 279.920 ;
        RECT 8.000 277.200 2916.580 277.680 ;
        RECT 54.000 274.960 2870.580 277.200 ;
        RECT 8.000 274.480 2916.580 274.960 ;
        RECT 54.000 272.240 2870.580 274.480 ;
        RECT 8.000 271.760 2916.580 272.240 ;
        RECT 54.000 269.520 2870.580 271.760 ;
        RECT 8.000 269.040 2916.580 269.520 ;
        RECT 54.000 266.800 2870.580 269.040 ;
        RECT 8.000 266.320 2916.580 266.800 ;
        RECT 54.000 264.080 2870.580 266.320 ;
        RECT 8.000 263.600 2916.580 264.080 ;
        RECT 54.000 261.360 2870.580 263.600 ;
        RECT 8.000 260.880 2916.580 261.360 ;
        RECT 54.000 258.640 2870.580 260.880 ;
        RECT 8.000 258.160 2916.580 258.640 ;
        RECT 54.000 255.920 2870.580 258.160 ;
        RECT 8.000 255.440 2916.580 255.920 ;
        RECT 54.000 253.200 2870.580 255.440 ;
        RECT 8.000 252.720 2916.580 253.200 ;
        RECT 54.000 250.480 2870.580 252.720 ;
        RECT 8.000 250.000 2916.580 250.480 ;
        RECT 54.000 247.760 2870.580 250.000 ;
        RECT 8.000 247.280 2916.580 247.760 ;
        RECT 54.000 245.040 2870.580 247.280 ;
        RECT 8.000 244.560 2916.580 245.040 ;
        RECT 54.000 242.320 2870.580 244.560 ;
        RECT 8.000 241.840 2916.580 242.320 ;
        RECT 54.000 239.600 2870.580 241.840 ;
        RECT 8.000 239.120 2916.580 239.600 ;
        RECT 54.000 236.880 2870.580 239.120 ;
        RECT 8.000 236.400 2916.580 236.880 ;
        RECT 54.000 234.160 2870.580 236.400 ;
        RECT 8.000 233.680 2916.580 234.160 ;
        RECT 54.000 231.440 2870.580 233.680 ;
        RECT 8.000 230.960 2916.580 231.440 ;
        RECT 54.000 228.720 2870.580 230.960 ;
        RECT 8.000 228.240 2916.580 228.720 ;
        RECT 54.000 226.000 2870.580 228.240 ;
        RECT 8.000 225.520 2916.580 226.000 ;
        RECT 54.000 223.280 2870.580 225.520 ;
        RECT 8.000 222.800 2916.580 223.280 ;
        RECT 54.000 220.560 2870.580 222.800 ;
        RECT 8.000 220.080 2916.580 220.560 ;
        RECT 54.000 217.840 2870.580 220.080 ;
        RECT 8.000 217.360 2916.580 217.840 ;
        RECT 54.000 215.120 2870.580 217.360 ;
        RECT 8.000 214.640 2916.580 215.120 ;
        RECT 54.000 212.400 2870.580 214.640 ;
        RECT 8.000 211.920 2916.580 212.400 ;
        RECT 54.000 209.680 2870.580 211.920 ;
        RECT 8.000 209.200 2916.580 209.680 ;
        RECT 54.000 206.960 2870.580 209.200 ;
        RECT 8.000 206.480 2916.580 206.960 ;
        RECT 54.000 204.240 2870.580 206.480 ;
        RECT 8.000 203.760 2916.580 204.240 ;
        RECT 54.000 201.520 2870.580 203.760 ;
        RECT 8.000 201.040 2916.580 201.520 ;
        RECT 54.000 198.800 2870.580 201.040 ;
        RECT 8.000 198.320 2916.580 198.800 ;
        RECT 54.000 196.080 2870.580 198.320 ;
        RECT 8.000 195.600 2916.580 196.080 ;
        RECT 54.000 193.360 2870.580 195.600 ;
        RECT 8.000 192.880 2916.580 193.360 ;
        RECT 54.000 190.640 2870.580 192.880 ;
        RECT 8.000 190.160 2916.580 190.640 ;
        RECT 54.000 187.920 2870.580 190.160 ;
        RECT 8.000 187.440 2916.580 187.920 ;
        RECT 54.000 185.200 2870.580 187.440 ;
        RECT 8.000 184.720 2916.580 185.200 ;
        RECT 54.000 182.480 2870.580 184.720 ;
        RECT 8.000 182.000 2916.580 182.480 ;
        RECT 54.000 179.760 2870.580 182.000 ;
        RECT 8.000 179.280 2916.580 179.760 ;
        RECT 54.000 177.040 2870.580 179.280 ;
        RECT 8.000 176.560 2916.580 177.040 ;
        RECT 54.000 174.320 2870.580 176.560 ;
        RECT 8.000 173.840 2916.580 174.320 ;
        RECT 54.000 171.600 2870.580 173.840 ;
        RECT 8.000 171.120 2916.580 171.600 ;
        RECT 54.000 168.880 2870.580 171.120 ;
        RECT 8.000 168.400 2916.580 168.880 ;
        RECT 54.000 166.160 2870.580 168.400 ;
        RECT 8.000 165.680 2916.580 166.160 ;
        RECT 54.000 163.440 2870.580 165.680 ;
        RECT 8.000 162.960 2916.580 163.440 ;
        RECT 54.000 160.720 2870.580 162.960 ;
        RECT 8.000 160.240 2916.580 160.720 ;
        RECT 54.000 158.000 2870.580 160.240 ;
        RECT 8.000 157.520 2916.580 158.000 ;
        RECT 54.000 155.280 2870.580 157.520 ;
        RECT 8.000 154.800 2916.580 155.280 ;
        RECT 54.000 152.560 2870.580 154.800 ;
        RECT 8.000 152.080 2916.580 152.560 ;
        RECT 54.000 149.840 2870.580 152.080 ;
        RECT 8.000 149.360 2916.580 149.840 ;
        RECT 54.000 147.120 2870.580 149.360 ;
        RECT 8.000 146.640 2916.580 147.120 ;
        RECT 54.000 144.400 2870.580 146.640 ;
        RECT 8.000 143.920 2916.580 144.400 ;
        RECT 54.000 141.680 2870.580 143.920 ;
        RECT 8.000 141.200 2916.580 141.680 ;
        RECT 54.000 138.960 2870.580 141.200 ;
        RECT 8.000 138.480 2916.580 138.960 ;
        RECT 54.000 136.240 2870.580 138.480 ;
        RECT 8.000 135.760 2916.580 136.240 ;
        RECT 54.000 133.520 2870.580 135.760 ;
        RECT 8.000 133.040 2916.580 133.520 ;
        RECT 54.000 130.800 2870.580 133.040 ;
        RECT 8.000 130.320 2916.580 130.800 ;
        RECT 54.000 128.080 2870.580 130.320 ;
        RECT 8.000 127.600 2916.580 128.080 ;
        RECT 54.000 125.360 2870.580 127.600 ;
        RECT 8.000 124.880 2916.580 125.360 ;
        RECT 54.000 122.640 2870.580 124.880 ;
        RECT 8.000 122.160 2916.580 122.640 ;
        RECT 54.000 119.920 2870.580 122.160 ;
        RECT 8.000 119.440 2916.580 119.920 ;
        RECT 54.000 117.200 2870.580 119.440 ;
        RECT 8.000 116.720 2916.580 117.200 ;
        RECT 54.000 114.480 2870.580 116.720 ;
        RECT 8.000 114.000 2916.580 114.480 ;
        RECT 54.000 111.760 2870.580 114.000 ;
        RECT 8.000 111.280 2916.580 111.760 ;
        RECT 54.000 109.040 2870.580 111.280 ;
        RECT 8.000 108.560 2916.580 109.040 ;
        RECT 54.000 106.320 2870.580 108.560 ;
        RECT 8.000 105.840 2916.580 106.320 ;
        RECT 54.000 103.600 2870.580 105.840 ;
        RECT 8.000 103.120 2916.580 103.600 ;
        RECT 54.000 100.880 2870.580 103.120 ;
        RECT 8.000 100.400 2916.580 100.880 ;
        RECT 54.000 98.160 2870.580 100.400 ;
        RECT 8.000 97.680 2916.580 98.160 ;
        RECT 54.000 95.440 2870.580 97.680 ;
        RECT 8.000 94.960 2916.580 95.440 ;
        RECT 54.000 92.720 2870.580 94.960 ;
        RECT 8.000 92.240 2916.580 92.720 ;
        RECT 54.000 90.000 2870.580 92.240 ;
        RECT 8.000 89.520 2916.580 90.000 ;
        RECT 54.000 87.280 2870.580 89.520 ;
        RECT 8.000 86.800 2916.580 87.280 ;
        RECT 54.000 84.560 2870.580 86.800 ;
        RECT 8.000 84.080 2916.580 84.560 ;
        RECT 54.000 81.840 2870.580 84.080 ;
        RECT 8.000 81.360 2916.580 81.840 ;
        RECT 54.000 79.120 2870.580 81.360 ;
        RECT 8.000 78.640 2916.580 79.120 ;
        RECT 54.000 76.400 2870.580 78.640 ;
        RECT 8.000 75.920 2916.580 76.400 ;
        RECT 54.000 73.680 2870.580 75.920 ;
        RECT 8.000 73.200 2916.580 73.680 ;
        RECT 54.000 70.960 2870.580 73.200 ;
        RECT 8.000 70.480 2916.580 70.960 ;
        RECT 54.000 68.240 2870.580 70.480 ;
        RECT 8.000 67.760 2916.580 68.240 ;
        RECT 54.000 65.520 2870.580 67.760 ;
        RECT 8.000 65.040 2916.580 65.520 ;
        RECT 54.000 62.800 2870.580 65.040 ;
        RECT 8.000 62.320 2916.580 62.800 ;
        RECT 54.000 60.080 2870.580 62.320 ;
        RECT 8.000 59.600 2916.580 60.080 ;
        RECT 54.000 57.360 2870.580 59.600 ;
        RECT 8.000 56.880 2916.580 57.360 ;
        RECT 54.000 54.640 2870.580 56.880 ;
        RECT 8.000 54.160 2916.580 54.640 ;
        RECT 54.000 54.000 2870.580 54.160 ;
        RECT 8.000 51.440 2916.580 51.920 ;
        RECT 8.000 48.720 2916.580 49.200 ;
        RECT 8.000 46.000 2916.580 46.480 ;
        RECT 8.000 43.280 2916.580 43.760 ;
        RECT 8.000 40.560 2916.580 41.040 ;
        RECT 8.000 37.840 2916.580 38.320 ;
        RECT 8.000 35.120 2916.580 35.600 ;
        RECT 8.000 32.400 2916.580 32.880 ;
        RECT 8.000 29.680 2916.580 30.160 ;
        RECT 8.000 26.960 2916.580 27.440 ;
        RECT 8.000 24.240 2916.580 24.720 ;
        RECT 8.000 21.520 2916.580 22.000 ;
        RECT 8.000 18.800 2916.580 19.280 ;
        RECT 8.000 16.080 2916.580 16.560 ;
        RECT 8.000 13.360 2916.580 13.840 ;
        RECT 8.000 10.640 2916.580 11.120 ;
      LAYER met2 ;
        RECT 57.320 54.000 2869.110 3466.000 ;
      LAYER met3 ;
        RECT 54.000 82.455 2870.580 3091.105 ;
      LAYER met4 ;
        RECT 457.255 54.000 2804.505 3091.105 ;
      LAYER met5 ;
        RECT 54.000 103.320 2870.580 3398.290 ;
  END
END user_project_wrapper
END LIBRARY

