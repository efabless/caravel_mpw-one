magic
tech sky130A
magscale 1 2
timestamp 1623348570
<< checkpaint >>
rect -1285 -1260 1388 1302
use sky130_fd_pr__dfm1sd__example_55959141808258  sky130_fd_pr__dfm1sd__example_55959141808258_0
timestamp 1623348570
transform 1 0 100 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 128 13 128 13 0 FreeSans 300 0 0 0 D
flabel comment s -25 42 -25 42 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 314296
string GDS_START 313524
<< end >>
