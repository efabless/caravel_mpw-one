magic
tech sky130A
magscale 1 2
timestamp 1606790299
<< obsli1 >>
rect 11000 10983 30136 30057
<< obsm1 >>
rect 10462 10952 30136 30088
<< metal2 >>
rect 10650 31576 10706 32376
rect 12490 31576 12546 32376
rect 14514 31576 14570 32376
rect 16354 31576 16410 32376
rect 18194 31576 18250 32376
rect 20218 31576 20274 32376
rect 22058 31576 22114 32376
rect 23898 31576 23954 32376
rect 25922 31576 25978 32376
rect 27762 31576 27818 32376
rect 29602 31576 29658 32376
rect 10466 8824 10522 9624
rect 12306 8824 12362 9624
rect 14146 8824 14202 9624
rect 15986 8824 16042 9624
rect 18010 8824 18066 9624
rect 19850 8824 19906 9624
rect 21690 8824 21746 9624
rect 23714 8824 23770 9624
rect 25554 8824 25610 9624
rect 27394 8824 27450 9624
rect 29418 8824 29474 9624
<< obsm2 >>
rect 10468 31520 10594 31576
rect 10762 31520 12434 31576
rect 12602 31520 14458 31576
rect 14626 31520 16298 31576
rect 16466 31520 18138 31576
rect 18306 31520 20162 31576
rect 20330 31520 22002 31576
rect 22170 31520 23842 31576
rect 24010 31520 25866 31576
rect 26034 31520 27706 31576
rect 27874 31520 29546 31576
rect 29714 31520 30024 31576
rect 10468 9680 30024 31520
rect 10578 9624 12250 9680
rect 12418 9624 14090 9680
rect 14258 9624 15930 9680
rect 16098 9624 17954 9680
rect 18122 9624 19794 9680
rect 19962 9624 21634 9680
rect 21802 9624 23658 9680
rect 23826 9624 25498 9680
rect 25666 9624 27338 9680
rect 27506 9624 29362 9680
rect 29530 9624 30024 9680
<< metal3 >>
rect 30504 30048 31304 30168
rect 9896 29232 10696 29352
rect 30504 27328 31304 27448
rect 9896 26240 10696 26360
rect 30504 24608 31304 24728
rect 9896 23520 10696 23640
rect 30504 21616 31304 21736
rect 9896 20800 10696 20920
rect 30504 18896 31304 19016
rect 9896 17808 10696 17928
rect 30504 16176 31304 16296
rect 9896 15088 10696 15208
rect 30504 13184 31304 13304
rect 9896 12368 10696 12488
rect 30504 10464 31304 10584
<< obsm3 >>
rect 0 30248 41136 41040
rect 0 29968 30424 30248
rect 31384 29968 41136 30248
rect 0 29432 41136 29968
rect 0 29152 9816 29432
rect 10776 29152 41136 29432
rect 0 27528 41136 29152
rect 0 27248 30424 27528
rect 31384 27248 41136 27528
rect 0 26440 41136 27248
rect 0 26160 9816 26440
rect 10776 26160 41136 26440
rect 0 24808 41136 26160
rect 0 24528 30424 24808
rect 31384 24528 41136 24808
rect 0 23720 41136 24528
rect 0 23440 9816 23720
rect 10776 23440 41136 23720
rect 0 21816 41136 23440
rect 0 21536 30424 21816
rect 31384 21536 41136 21816
rect 0 21000 41136 21536
rect 0 20720 9816 21000
rect 10776 20720 41136 21000
rect 0 19096 41136 20720
rect 0 18816 30424 19096
rect 31384 18816 41136 19096
rect 0 18008 41136 18816
rect 0 17728 9816 18008
rect 10776 17728 41136 18008
rect 0 16376 41136 17728
rect 0 16096 30424 16376
rect 31384 16096 41136 16376
rect 0 15288 41136 16096
rect 0 15008 9816 15288
rect 10776 15008 41136 15288
rect 0 13384 41136 15008
rect 0 13104 30424 13384
rect 31384 13104 41136 13384
rect 0 12568 41136 13104
rect 0 12288 9816 12568
rect 10776 12288 41136 12568
rect 0 10664 41136 12288
rect 0 10384 30424 10664
rect 31384 10384 41136 10664
rect 0 0 41136 10384
<< metal4 >>
rect 0 0 4000 41040
rect 5000 5000 9000 36040
<< obsm4 >>
rect 14104 0 41136 41040
<< labels >>
rlabel metal2 s 27762 31576 27818 32376 6 clockp[0]
port 1 nsew
rlabel metal2 s 21690 8824 21746 9624 6 clockp[1]
port 2 nsew
rlabel metal2 s 12306 8824 12362 9624 6 dco
port 3 nsew
rlabel metal2 s 10466 8824 10522 9624 6 div[0]
port 4 nsew
rlabel metal3 s 9896 17808 10696 17928 6 div[1]
port 5 nsew
rlabel metal2 s 27394 8824 27450 9624 6 div[2]
port 6 nsew
rlabel metal3 s 30504 10464 31304 10584 6 div[3]
port 7 nsew
rlabel metal3 s 9896 12368 10696 12488 6 div[4]
port 8 nsew
rlabel metal2 s 20218 31576 20274 32376 6 enable
port 9 nsew
rlabel metal2 s 14514 31576 14570 32376 6 ext_trim[0]
port 10 nsew
rlabel metal2 s 23898 31576 23954 32376 6 ext_trim[10]
port 11 nsew
rlabel metal3 s 9896 23520 10696 23640 6 ext_trim[11]
port 12 nsew
rlabel metal3 s 30504 13184 31304 13304 6 ext_trim[12]
port 13 nsew
rlabel metal2 s 29418 8824 29474 9624 6 ext_trim[13]
port 14 nsew
rlabel metal3 s 9896 20800 10696 20920 6 ext_trim[14]
port 15 nsew
rlabel metal2 s 14146 8824 14202 9624 6 ext_trim[15]
port 16 nsew
rlabel metal3 s 30504 27328 31304 27448 6 ext_trim[16]
port 17 nsew
rlabel metal3 s 9896 26240 10696 26360 6 ext_trim[17]
port 18 nsew
rlabel metal2 s 29602 31576 29658 32376 6 ext_trim[18]
port 19 nsew
rlabel metal2 s 18194 31576 18250 32376 6 ext_trim[19]
port 20 nsew
rlabel metal3 s 30504 24608 31304 24728 6 ext_trim[1]
port 21 nsew
rlabel metal2 s 25554 8824 25610 9624 6 ext_trim[20]
port 22 nsew
rlabel metal3 s 9896 29232 10696 29352 6 ext_trim[21]
port 23 nsew
rlabel metal3 s 30504 21616 31304 21736 6 ext_trim[22]
port 24 nsew
rlabel metal3 s 9896 15088 10696 15208 6 ext_trim[23]
port 25 nsew
rlabel metal2 s 19850 8824 19906 9624 6 ext_trim[24]
port 26 nsew
rlabel metal3 s 30504 16176 31304 16296 6 ext_trim[25]
port 27 nsew
rlabel metal3 s 30504 18896 31304 19016 6 ext_trim[2]
port 28 nsew
rlabel metal2 s 12490 31576 12546 32376 6 ext_trim[3]
port 29 nsew
rlabel metal2 s 25922 31576 25978 32376 6 ext_trim[4]
port 30 nsew
rlabel metal2 s 23714 8824 23770 9624 6 ext_trim[5]
port 31 nsew
rlabel metal2 s 22058 31576 22114 32376 6 ext_trim[6]
port 32 nsew
rlabel metal2 s 10650 31576 10706 32376 6 ext_trim[7]
port 33 nsew
rlabel metal2 s 16354 31576 16410 32376 6 ext_trim[8]
port 34 nsew
rlabel metal3 s 30504 30048 31304 30168 6 ext_trim[9]
port 35 nsew
rlabel metal2 s 18010 8824 18066 9624 6 osc
port 36 nsew
rlabel metal2 s 15986 8824 16042 9624 6 resetb
port 37 nsew
rlabel metal4 s 5000 5000 9000 36040 6 VPWR
port 38 nsew power default
rlabel metal4 s 0 0 4000 41040 6 VGND
port 39 nsew ground default
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 41136 41040
string LEFview TRUE
string GDS_FILE digital_pll.gds
string GDS_END 2654930
string GDS_START 265824
<< end >>

