magic
tech sky130A
magscale 12 1
timestamp 1598776550
<< metal5 >>
rect 0 0 15 105
<< properties >>
string FIXED_BBOX 0 -30 30 105
<< end >>
