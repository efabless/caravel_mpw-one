* NGSPICE file created from gpio_control_block.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_8 abstract view
.subckt sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

.subckt gpio_control_block mgmt_gpio_in mgmt_gpio_oeb mgmt_gpio_out one pad_gpio_ana_en
+ pad_gpio_ana_pol pad_gpio_ana_sel pad_gpio_dm[0] pad_gpio_dm[1] pad_gpio_dm[2] pad_gpio_holdover
+ pad_gpio_ib_mode_sel pad_gpio_in pad_gpio_inenb pad_gpio_out pad_gpio_outenb pad_gpio_slow_sel
+ pad_gpio_vtrip_sel resetn serial_clock serial_data_in serial_data_out user_gpio_in
+ user_gpio_oeb user_gpio_out zero vccd vssd1 vccd1
X_062_ _065_/A vssd1 vssd1 vccd vccd _062_/X sky130_fd_sc_hd__buf_2
XFILLER_13_3 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_6
X_045_ _047_/A vssd1 vssd1 vccd vccd _045_/X sky130_fd_sc_hd__buf_2
XFILLER_15_32 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
X_044_ _047_/A vssd1 vssd1 vccd vccd _044_/X sky130_fd_sc_hd__buf_2
X_061_ _065_/A vssd1 vssd1 vccd vccd _061_/X sky130_fd_sc_hd__buf_2
XFILLER_0_15 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_8
X_060_ _084_/A vssd1 vssd1 vccd vccd _065_/A sky130_fd_sc_hd__buf_2
X_043_ _084_/A vssd1 vssd1 vccd vccd _047_/A sky130_fd_sc_hd__buf_2
XFILLER_12_57 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_042_ _066_/A vssd1 vssd1 vccd vccd _084_/A sky130_fd_sc_hd__buf_2
X_111_ _083_/A _111_/D _084_/X vssd1 vssd1 vccd vccd serial_data_out sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_59 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
X_041_ _083_/A resetn vssd1 vssd1 vccd vccd _066_/A sky130_fd_sc_hd__or2_4
X_110_ _110_/CLK _110_/D _047_/A vssd1 vssd1 vccd vccd _111_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_1_3 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_29 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
XPHY_0 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_099_ _083_/A serial_data_in _056_/X vssd1 vssd1 vccd vccd _100_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_1_62 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_9 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_40 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
Xconst_source vssd1 vssd1 vccd vccd one zero sky130_fd_sc_hd__conb_1
XFILLER_4_62 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
X_098_ _083_/X _107_/D _057_/X vssd1 vssd1 vccd vccd pad_gpio_ana_pol sky130_fd_sc_hd__dfrtp_4
XPHY_2 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__tapvpwrvgnd_1_0 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_097_ _083_/X _106_/D _058_/X vssd1 vssd1 vccd vccd pad_gpio_ana_sel sky130_fd_sc_hd__dfrtp_4
XFILLER_10_62 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
XPHY_3 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_30 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_62 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_7 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_096_ _083_/X _105_/D _059_/X vssd1 vssd1 vccd vccd pad_gpio_ana_en sky130_fd_sc_hd__dfrtp_4
XPHY_4 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_079_ pad_gpio_dm[0] _079_/B vssd1 vssd1 vccd vccd _079_/Y sky130_fd_sc_hd__nand2_4
X_095_ _083_/X serial_data_out _061_/X vssd1 vssd1 vccd vccd pad_gpio_dm[2] sky130_fd_sc_hd__dfstp_4
X_078_ mgmt_gpio_out _079_/B vssd1 vssd1 vccd vccd _078_/X sky130_fd_sc_hd__or2_4
XFILLER_16_63 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_094_ _083_/X _111_/D _062_/X vssd1 vssd1 vccd vccd pad_gpio_dm[1] sky130_fd_sc_hd__dfstp_4
XPHY_6 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_077_ mgmt_gpio_oeb _077_/B pad_gpio_dm[1] vssd1 vssd1 vccd vccd _079_/B sky130_fd_sc_hd__and3_4
X_093_ _083_/X _110_/D _063_/X vssd1 vssd1 vccd vccd pad_gpio_dm[0] sky130_fd_sc_hd__dfrtp_4
X_076_ pad_gpio_dm[2] vssd1 vssd1 vccd vccd _077_/B sky130_fd_sc_hd__inv_2
XFILLER_16_32 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_4
X_059_ _059_/A vssd1 vssd1 vccd vccd _059_/X sky130_fd_sc_hd__buf_2
XPHY_7 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
Xgpio_in_buf _081_/Y gpio_in_buf/TE vssd1 vssd1 vccd vccd user_gpio_in sky130_fd_sc_hd__einvp_8
X_092_ _083_/X _101_/D _064_/X vssd1 vssd1 vccd vccd _092_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_1_36 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
X_075_ _092_/Q mgmt_gpio_oeb _086_/Q user_gpio_oeb _074_/Y vssd1 vssd1 vccd vccd pad_gpio_outenb
+ sky130_fd_sc_hd__a32o_4
X_058_ _059_/A vssd1 vssd1 vccd vccd _058_/X sky130_fd_sc_hd__buf_2
XPHY_8 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_074_ _086_/Q vssd1 vssd1 vccd vccd _074_/Y sky130_fd_sc_hd__inv_2
X_091_ _083_/X _104_/D _065_/X vssd1 vssd1 vccd vccd pad_gpio_ib_mode_sel sky130_fd_sc_hd__dfrtp_4
X_057_ _059_/A vssd1 vssd1 vccd vccd _057_/X sky130_fd_sc_hd__buf_2
XPHY_9 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_36 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_109_ _110_/CLK _109_/D _044_/X vssd1 vssd1 vccd vccd _110_/D sky130_fd_sc_hd__dfrtp_4
X_090_ _083_/X _103_/D _067_/X vssd1 vssd1 vccd vccd pad_gpio_inenb sky130_fd_sc_hd__dfrtp_4
XFILLER_6_3 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
X_056_ _059_/A vssd1 vssd1 vccd vccd _056_/X sky130_fd_sc_hd__buf_2
X_073_ _073_/A pad_gpio_inenb vssd1 vssd1 vccd vccd _073_/X sky130_fd_sc_hd__or2_4
X_108_ _110_/CLK _108_/D _045_/X vssd1 vssd1 vccd vccd _109_/D sky130_fd_sc_hd__dfrtp_4
X_072_ _092_/Q vssd1 vssd1 vccd vccd _073_/A sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0_serial_clock clkbuf_0_serial_clock/X vssd1 vssd1 vccd vccd _083_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_16_36 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_055_ _059_/A vssd1 vssd1 vccd vccd _055_/X sky130_fd_sc_hd__buf_2
XFILLER_16_6 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_12
X_107_ _110_/CLK _107_/D _046_/X vssd1 vssd1 vccd vccd _108_/D sky130_fd_sc_hd__dfrtp_4
X_071_ _071_/A vssd1 vssd1 vccd vccd _071_/X sky130_fd_sc_hd__buf_2
XFILLER_2_50 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
X_054_ _084_/A vssd1 vssd1 vccd vccd _059_/A sky130_fd_sc_hd__buf_2
X_106_ _110_/CLK _106_/D _047_/X vssd1 vssd1 vccd vccd _107_/D sky130_fd_sc_hd__dfrtp_4
X_070_ _071_/A vssd1 vssd1 vccd vccd _070_/X sky130_fd_sc_hd__buf_2
XFILLER_4_3 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_62 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
X_053_ _053_/A vssd1 vssd1 vccd vccd _053_/X sky130_fd_sc_hd__buf_2
X_105_ _110_/CLK _105_/D _049_/X vssd1 vssd1 vccd vccd _106_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_8_50 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_41 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_052_ _053_/A vssd1 vssd1 vccd vccd _052_/X sky130_fd_sc_hd__buf_2
X_104_ _110_/CLK _104_/D _050_/X vssd1 vssd1 vccd vccd _105_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_12_3 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_62 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_30 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_051_ _053_/A vssd1 vssd1 vccd vccd _051_/X sky130_fd_sc_hd__buf_2
XFILLER_16_18 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
X_103_ _110_/CLK _103_/D _051_/X vssd1 vssd1 vccd vccd _104_/D sky130_fd_sc_hd__dfrtp_4
XPHY_50 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_62 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_30 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_102_ _110_/CLK _102_/D _052_/X vssd1 vssd1 vccd vccd _103_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_2_3 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_12
X_050_ _053_/A vssd1 vssd1 vccd vccd _050_/X sky130_fd_sc_hd__buf_2
Xgpio_logic_high vssd1 vssd1 vccd1 vccd1 gpio_in_buf/TE gpio_logic_high/LO sky130_fd_sc_hd__conb_1
XFILLER_5_32 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
XPHY_51 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_101_ _083_/A _101_/D _053_/X vssd1 vssd1 vccd vccd _102_/D sky130_fd_sc_hd__dfrtp_4
XPHY_52 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_100_ _083_/A _100_/D _055_/X vssd1 vssd1 vccd vccd _101_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_11_32 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
XPHY_31 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_12
XPHY_32 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_089_ _083_/X _109_/D _068_/X vssd1 vssd1 vccd vccd pad_gpio_vtrip_sel sky130_fd_sc_hd__dfrtp_4
Xclkbuf_1_0_0_serial_clock clkbuf_0_serial_clock/X vssd1 vssd1 vccd vccd _110_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XPHY_33 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_15 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
Xclkbuf_0_serial_clock serial_clock vssd1 vssd1 vccd vccd clkbuf_0_serial_clock/X
+ sky130_fd_sc_hd__clkbuf_16
X_088_ _083_/X _108_/D _069_/X vssd1 vssd1 vccd vccd pad_gpio_slow_sel sky130_fd_sc_hd__dfrtp_4
XFILLER_5_37 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_57 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
XPHY_12 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_087_ _083_/X _102_/D _070_/X vssd1 vssd1 vccd vccd pad_gpio_holdover sky130_fd_sc_hd__dfrtp_4
XPHY_24 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_3 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
XPHY_35 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_086_ _083_/X _100_/D _071_/X vssd1 vssd1 vccd vccd _086_/Q sky130_fd_sc_hd__dfstp_4
X_069_ _071_/A vssd1 vssd1 vccd vccd _069_/X sky130_fd_sc_hd__buf_2
XPHY_25 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_085_ pad_gpio_in _073_/X vssd1 vssd1 vccd vccd mgmt_gpio_in sky130_fd_sc_hd__ebufn_2
X_068_ _071_/A vssd1 vssd1 vccd vccd _068_/X sky130_fd_sc_hd__buf_2
XPHY_48 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_26 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_067_ _071_/A vssd1 vssd1 vccd vccd _067_/X sky130_fd_sc_hd__buf_2
XFILLER_0_63 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_084_ _084_/A vssd1 vssd1 vccd vccd _084_/X sky130_fd_sc_hd__buf_2
XPHY_27 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_0 mgmt_gpio_out vssd1 vssd1 vccd vccd sky130_fd_sc_hd__diode_2
XPHY_38 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_62 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
XPHY_16 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_083_ _083_/A _083_/B vssd1 vssd1 vccd vccd _083_/X sky130_fd_sc_hd__and2_4
XFILLER_3_30 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_066_ _066_/A vssd1 vssd1 vccd vccd _071_/A sky130_fd_sc_hd__buf_2
XFILLER_9_62 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
X_049_ _053_/A vssd1 vssd1 vccd vccd _049_/X sky130_fd_sc_hd__buf_2
XANTENNA_1 serial_data_in vssd1 vssd1 vccd vccd sky130_fd_sc_hd__diode_2
XPHY_28 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_082_ resetn vssd1 vssd1 vccd vccd _083_/B sky130_fd_sc_hd__inv_2
XFILLER_12_62 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_32 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_6
X_065_ _065_/A vssd1 vssd1 vccd vccd _065_/X sky130_fd_sc_hd__buf_2
XFILLER_15_3 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_048_ _084_/A vssd1 vssd1 vccd vccd _053_/A sky130_fd_sc_hd__buf_2
XPHY_29 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_081_ pad_gpio_in vssd1 vssd1 vccd vccd _081_/Y sky130_fd_sc_hd__inv_2
X_064_ _065_/A vssd1 vssd1 vccd vccd _064_/X sky130_fd_sc_hd__buf_2
XPHY_19 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_047_ _047_/A vssd1 vssd1 vccd vccd _047_/X sky130_fd_sc_hd__buf_2
X_080_ _086_/Q _078_/X _079_/Y _074_/Y user_gpio_out vssd1 vssd1 vccd vccd pad_gpio_out
+ sky130_fd_sc_hd__a32o_4
X_063_ _065_/A vssd1 vssd1 vccd vccd _063_/X sky130_fd_sc_hd__buf_2
XFILLER_0_23 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
X_046_ _047_/A vssd1 vssd1 vccd vccd _046_/X sky130_fd_sc_hd__buf_2
.ends

