magic
tech sky130A
magscale 12 1
timestamp 1598768910
<< metal5 >>
rect 0 90 45 105
rect 15 0 30 90
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
