magic
tech sky130A
magscale 1 2
timestamp 1606789160
<< checkpaint >>
rect -1260 -1260 35194 19604
<< locali >>
rect 11325 9257 11383 9291
rect 11291 8883 11325 9053
rect 11291 7183 11325 7421
<< viali >>
rect 7151 15581 7185 15615
rect 7519 15241 7553 15275
rect 7703 15037 7737 15071
rect 6323 14629 6357 14663
rect 7427 14629 7461 14663
rect 6507 14493 6541 14527
rect 7611 14493 7645 14527
rect 6231 14153 6265 14187
rect 7335 14153 7369 14187
rect 7703 14085 7737 14119
rect 4759 13677 4793 13711
rect 4667 13541 4701 13575
rect 5679 13541 5713 13575
rect 7703 13541 7737 13575
rect 5955 13473 5989 13507
rect 4759 13201 4793 13235
rect 4207 13065 4241 13099
rect 4575 13065 4609 13099
rect 5771 12997 5805 13031
rect 6047 12997 6081 13031
rect 7795 12997 7829 13031
rect 4023 12861 4057 12895
rect 5955 12521 5989 12555
rect 7703 12521 7737 12555
rect 3195 12453 3229 12487
rect 4483 12453 4517 12487
rect 5679 12453 5713 12487
rect 4299 12385 4333 12419
rect 3379 12317 3413 12351
rect 4575 12317 4609 12351
rect 3103 12045 3137 12079
rect 5771 11977 5805 12011
rect 2827 11909 2861 11943
rect 4851 11909 4885 11943
rect 6047 11909 6081 11943
rect 7795 11909 7829 11943
rect 7979 11773 8013 11807
rect 4483 11433 4517 11467
rect 5955 11433 5989 11467
rect 1815 11365 1849 11399
rect 3011 11365 3045 11399
rect 4391 11365 4425 11399
rect 4759 11365 4793 11399
rect 5679 11365 5713 11399
rect 7703 11297 7737 11331
rect 1999 11229 2033 11263
rect 3195 11229 3229 11263
rect 1907 11025 1941 11059
rect 4851 10957 4885 10991
rect 6047 10957 6081 10991
rect 619 10889 653 10923
rect 1723 10889 1757 10923
rect 2827 10821 2861 10855
rect 5771 10821 5805 10855
rect 7795 10821 7829 10855
rect 803 10753 837 10787
rect 3090 10685 3124 10719
rect 1539 10345 1573 10379
rect 3287 10345 3321 10379
rect 7335 10345 7369 10379
rect 435 10277 469 10311
rect 1631 10277 1665 10311
rect 3747 10277 3781 10311
rect 3931 10277 3965 10311
rect 4207 10277 4241 10311
rect 4483 10277 4517 10311
rect 4759 10277 4793 10311
rect 5587 10277 5621 10311
rect 5955 10277 5989 10311
rect 2091 10209 2125 10243
rect 619 10141 653 10175
rect 1907 9937 1941 9971
rect 619 9801 653 9835
rect 1723 9801 1757 9835
rect 2827 9801 2861 9835
rect 5771 9801 5805 9835
rect 3103 9733 3137 9767
rect 4851 9733 4885 9767
rect 6047 9733 6081 9767
rect 7795 9733 7829 9767
rect 803 9665 837 9699
rect 5035 9325 5069 9359
rect 11291 9257 11325 9291
rect 11383 9257 11417 9291
rect 699 9189 733 9223
rect 1815 9189 1849 9223
rect 3747 9189 3781 9223
rect 5587 9189 5621 9223
rect 5955 9189 5989 9223
rect 895 9053 929 9087
rect 1999 9053 2033 9087
rect 7703 9053 7737 9087
rect 11291 9053 11325 9087
rect 1907 8849 1941 8883
rect 11291 8849 11325 8883
rect 6047 8781 6081 8815
rect 619 8713 653 8747
rect 1723 8713 1757 8747
rect 5771 8713 5805 8747
rect 2827 8645 2861 8679
rect 3103 8645 3137 8679
rect 4851 8645 4885 8679
rect 7795 8645 7829 8679
rect 803 8509 837 8543
rect 1999 8305 2033 8339
rect 895 8237 929 8271
rect 3287 8169 3321 8203
rect 4667 8169 4701 8203
rect 5587 8169 5621 8203
rect 5955 8169 5989 8203
rect 699 8101 733 8135
rect 1815 8101 1849 8135
rect 3011 8101 3045 8135
rect 3747 8101 3781 8135
rect 4023 8101 4057 8135
rect 4115 8101 4149 8135
rect 4575 8101 4609 8135
rect 7703 8033 7737 8067
rect 3103 7965 3137 7999
rect 803 7761 837 7795
rect 3103 7693 3137 7727
rect 6047 7693 6081 7727
rect 619 7625 653 7659
rect 1723 7625 1757 7659
rect 2827 7625 2861 7659
rect 5771 7625 5805 7659
rect 4851 7557 4885 7591
rect 7795 7557 7829 7591
rect 1907 7421 1941 7455
rect 11291 7421 11325 7455
rect 2735 7217 2769 7251
rect 4575 7217 4609 7251
rect 1999 7149 2033 7183
rect 11291 7149 11325 7183
rect 3655 7081 3689 7115
rect 711 7013 745 7047
rect 1815 7013 1849 7047
rect 2551 7013 2585 7047
rect 3563 7013 3597 7047
rect 3931 7013 3965 7047
rect 4115 7013 4149 7047
rect 4391 7013 4425 7047
rect 5679 7013 5713 7047
rect 4299 6945 4333 6979
rect 5955 6945 5989 6979
rect 7703 6945 7737 6979
rect 895 6877 929 6911
rect 1723 6537 1757 6571
rect 2827 6537 2861 6571
rect 5771 6537 5805 6571
rect 3103 6469 3137 6503
rect 4851 6469 4885 6503
rect 6047 6469 6081 6503
rect 7795 6469 7829 6503
rect 1907 6333 1941 6367
rect 1999 6129 2033 6163
rect 3379 6129 3413 6163
rect 4575 6129 4609 6163
rect 5955 5993 5989 6027
rect 1907 5925 1941 5959
rect 3195 5925 3229 5959
rect 4299 5925 4333 5959
rect 4483 5925 4517 5959
rect 5679 5925 5713 5959
rect 7703 5857 7737 5891
rect 4851 5517 4885 5551
rect 2827 5449 2861 5483
rect 5771 5449 5805 5483
rect 3103 5381 3137 5415
rect 6047 5381 6081 5415
rect 7795 5381 7829 5415
rect 3655 5041 3689 5075
rect 5679 4905 5713 4939
rect 5955 4905 5989 4939
rect 3471 4837 3505 4871
rect 4575 4837 4609 4871
rect 7703 4769 7737 4803
rect 4759 4701 4793 4735
rect 3747 4497 3781 4531
rect 3931 4361 3965 4395
rect 4575 4361 4609 4395
rect 5771 4293 5805 4327
rect 7795 4293 7829 4327
rect 4759 4225 4793 4259
rect 6034 4157 6068 4191
rect 5942 3953 5976 3987
rect 5679 3817 5713 3851
rect 7703 3817 7737 3851
rect 6323 3409 6357 3443
rect 6139 3273 6173 3307
rect 7335 3273 7369 3307
rect 7243 3205 7277 3239
rect 7519 3069 7553 3103
rect 7611 2865 7645 2899
rect 7427 2661 7461 2695
rect 7519 2185 7553 2219
rect 7703 2049 7737 2083
<< metal1 >>
rect 7688 16320 7694 16372
rect 7746 16360 7752 16372
rect 15508 16360 15514 16372
rect 7746 16332 15514 16360
rect 7746 16320 7752 16332
rect 15508 16320 15514 16332
rect 15566 16320 15572 16372
rect 38 16066 8870 16088
rect 38 16014 1394 16066
rect 1446 16014 1458 16066
rect 1510 16014 1522 16066
rect 1574 16014 1586 16066
rect 1638 16014 4352 16066
rect 4404 16014 4416 16066
rect 4468 16014 4480 16066
rect 4532 16014 4544 16066
rect 4596 16014 7309 16066
rect 7361 16014 7373 16066
rect 7425 16014 7437 16066
rect 7489 16014 7501 16066
rect 7553 16014 8870 16066
rect 38 15992 8870 16014
rect 7136 15612 7142 15624
rect 7097 15584 7142 15612
rect 7136 15572 7142 15584
rect 7194 15572 7200 15624
rect 38 15522 8870 15544
rect 38 15470 2873 15522
rect 2925 15470 2937 15522
rect 2989 15470 3001 15522
rect 3053 15470 3065 15522
rect 3117 15470 5830 15522
rect 5882 15470 5894 15522
rect 5946 15470 5958 15522
rect 6010 15470 6022 15522
rect 6074 15470 8870 15522
rect 38 15448 8870 15470
rect 4836 15232 4842 15284
rect 4894 15272 4900 15284
rect 7507 15275 7565 15281
rect 7507 15272 7519 15275
rect 4894 15244 7519 15272
rect 4894 15232 4900 15244
rect 7507 15241 7519 15244
rect 7553 15241 7565 15275
rect 7507 15235 7565 15241
rect 7691 15071 7749 15077
rect 7691 15037 7703 15071
rect 7737 15068 7749 15071
rect 7780 15068 7786 15080
rect 7737 15040 7786 15068
rect 7737 15037 7749 15040
rect 7691 15031 7749 15037
rect 7780 15028 7786 15040
rect 7838 15028 7844 15080
rect 38 14978 8870 15000
rect 38 14926 1394 14978
rect 1446 14926 1458 14978
rect 1510 14926 1522 14978
rect 1574 14926 1586 14978
rect 1638 14926 4352 14978
rect 4404 14926 4416 14978
rect 4468 14926 4480 14978
rect 4532 14926 4544 14978
rect 4596 14926 7309 14978
rect 7361 14926 7373 14978
rect 7425 14926 7437 14978
rect 7489 14926 7501 14978
rect 7553 14926 8870 14978
rect 38 14904 8870 14926
rect 1708 14620 1714 14672
rect 1766 14660 1772 14672
rect 6311 14663 6369 14669
rect 6311 14660 6323 14663
rect 1766 14632 6323 14660
rect 1766 14620 1772 14632
rect 6311 14629 6323 14632
rect 6357 14629 6369 14663
rect 6311 14623 6369 14629
rect 7415 14663 7473 14669
rect 7415 14629 7427 14663
rect 7461 14629 7473 14663
rect 7415 14623 7473 14629
rect 1892 14552 1898 14604
rect 1950 14592 1956 14604
rect 7430 14592 7458 14623
rect 1950 14564 7458 14592
rect 1950 14552 1956 14564
rect 4744 14484 4750 14536
rect 4802 14524 4808 14536
rect 6495 14527 6553 14533
rect 6495 14524 6507 14527
rect 4802 14496 6507 14524
rect 4802 14484 4808 14496
rect 6495 14493 6507 14496
rect 6541 14493 6553 14527
rect 7596 14524 7602 14536
rect 7557 14496 7602 14524
rect 6495 14487 6553 14493
rect 7596 14484 7602 14496
rect 7654 14484 7660 14536
rect 38 14434 8870 14456
rect 38 14382 2873 14434
rect 2925 14382 2937 14434
rect 2989 14382 3001 14434
rect 3053 14382 3065 14434
rect 3117 14382 5830 14434
rect 5882 14382 5894 14434
rect 5946 14382 5958 14434
rect 6010 14382 6022 14434
rect 6074 14382 8870 14434
rect 38 14360 8870 14382
rect 6219 14187 6277 14193
rect 6219 14153 6231 14187
rect 6265 14184 6277 14187
rect 7136 14184 7142 14196
rect 6265 14156 7142 14184
rect 6265 14153 6277 14156
rect 6219 14147 6277 14153
rect 7136 14144 7142 14156
rect 7194 14144 7200 14196
rect 7323 14187 7381 14193
rect 7323 14153 7335 14187
rect 7369 14153 7381 14187
rect 7323 14147 7381 14153
rect 6584 14076 6590 14128
rect 6642 14116 6648 14128
rect 7338 14116 7366 14147
rect 7688 14116 7694 14128
rect 6642 14088 7366 14116
rect 7649 14088 7694 14116
rect 6642 14076 6648 14088
rect 7688 14076 7694 14088
rect 7746 14076 7752 14128
rect 38 13890 8870 13912
rect 38 13838 1394 13890
rect 1446 13838 1458 13890
rect 1510 13838 1522 13890
rect 1574 13838 1586 13890
rect 1638 13838 4352 13890
rect 4404 13838 4416 13890
rect 4468 13838 4480 13890
rect 4532 13838 4544 13890
rect 4596 13838 7309 13890
rect 7361 13838 7373 13890
rect 7425 13838 7437 13890
rect 7489 13838 7501 13890
rect 7553 13838 8870 13890
rect 38 13816 8870 13838
rect 3364 13668 3370 13720
rect 3422 13708 3428 13720
rect 4747 13711 4805 13717
rect 4747 13708 4759 13711
rect 3422 13680 4759 13708
rect 3422 13668 3428 13680
rect 4747 13677 4759 13680
rect 4793 13677 4805 13711
rect 4747 13671 4805 13677
rect 15508 13640 15514 13652
rect 4670 13612 15514 13640
rect 4670 13584 4698 13612
rect 15508 13600 15514 13612
rect 15566 13600 15572 13652
rect 4652 13572 4658 13584
rect 4613 13544 4658 13572
rect 4652 13532 4658 13544
rect 4710 13532 4716 13584
rect 5664 13572 5670 13584
rect 5625 13544 5670 13572
rect 5664 13532 5670 13544
rect 5722 13532 5728 13584
rect 7228 13532 7234 13584
rect 7286 13572 7292 13584
rect 7691 13575 7749 13581
rect 7691 13572 7703 13575
rect 7286 13544 7703 13572
rect 7286 13532 7292 13544
rect 7691 13541 7703 13544
rect 7737 13541 7749 13575
rect 7691 13535 7749 13541
rect 1800 13464 1806 13516
rect 1858 13504 1864 13516
rect 5943 13507 6001 13513
rect 1858 13476 5894 13504
rect 1858 13464 1864 13476
rect 5866 13436 5894 13476
rect 5943 13473 5955 13507
rect 5989 13504 6001 13507
rect 6216 13504 6222 13516
rect 5989 13476 6222 13504
rect 5989 13473 6001 13476
rect 5943 13467 6001 13473
rect 6216 13464 6222 13476
rect 6274 13464 6280 13516
rect 6418 13436 6446 13490
rect 5866 13408 6446 13436
rect 38 13346 8870 13368
rect 38 13294 2873 13346
rect 2925 13294 2937 13346
rect 2989 13294 3001 13346
rect 3053 13294 3065 13346
rect 3117 13294 5830 13346
rect 5882 13294 5894 13346
rect 5946 13294 5958 13346
rect 6010 13294 6022 13346
rect 6074 13294 8870 13346
rect 38 13272 8870 13294
rect 4747 13235 4805 13241
rect 4747 13201 4759 13235
rect 4793 13232 4805 13235
rect 4836 13232 4842 13244
rect 4793 13204 4842 13232
rect 4793 13201 4805 13204
rect 4747 13195 4805 13201
rect 4836 13192 4842 13204
rect 4894 13192 4900 13244
rect 6492 13124 6498 13176
rect 6550 13124 6556 13176
rect 3824 13056 3830 13108
rect 3882 13096 3888 13108
rect 4195 13099 4253 13105
rect 4195 13096 4207 13099
rect 3882 13068 4207 13096
rect 3882 13056 3888 13068
rect 4195 13065 4207 13068
rect 4241 13065 4253 13099
rect 4195 13059 4253 13065
rect 4563 13099 4621 13105
rect 4563 13065 4575 13099
rect 4609 13065 4621 13099
rect 4563 13059 4621 13065
rect 4100 12988 4106 13040
rect 4158 13028 4164 13040
rect 4578 13028 4606 13059
rect 4158 13000 4606 13028
rect 4158 12988 4164 13000
rect 5664 12988 5670 13040
rect 5722 13028 5728 13040
rect 5759 13031 5817 13037
rect 5759 13028 5771 13031
rect 5722 13000 5771 13028
rect 5722 12988 5728 13000
rect 5759 12997 5771 13000
rect 5805 12997 5817 13031
rect 5759 12991 5817 12997
rect 6035 13031 6093 13037
rect 6035 12997 6047 13031
rect 6081 13028 6093 13031
rect 6124 13028 6130 13040
rect 6081 13000 6130 13028
rect 6081 12997 6093 13000
rect 6035 12991 6093 12997
rect 6124 12988 6130 13000
rect 6182 12988 6188 13040
rect 6400 12988 6406 13040
rect 6458 13028 6464 13040
rect 7783 13031 7841 13037
rect 7783 13028 7795 13031
rect 6458 13000 7795 13028
rect 6458 12988 6464 13000
rect 7783 12997 7795 13000
rect 7829 12997 7841 13031
rect 7783 12991 7841 12997
rect 2628 12852 2634 12904
rect 2686 12892 2692 12904
rect 4011 12895 4069 12901
rect 4011 12892 4023 12895
rect 2686 12864 4023 12892
rect 2686 12852 2692 12864
rect 4011 12861 4023 12864
rect 4057 12892 4069 12895
rect 4192 12892 4198 12904
rect 4057 12864 4198 12892
rect 4057 12861 4069 12864
rect 4011 12855 4069 12861
rect 4192 12852 4198 12864
rect 4250 12852 4256 12904
rect 38 12802 8870 12824
rect 38 12750 1394 12802
rect 1446 12750 1458 12802
rect 1510 12750 1522 12802
rect 1574 12750 1586 12802
rect 1638 12750 4352 12802
rect 4404 12750 4416 12802
rect 4468 12750 4480 12802
rect 4532 12750 4544 12802
rect 4596 12750 7309 12802
rect 7361 12750 7373 12802
rect 7425 12750 7437 12802
rect 7489 12750 7501 12802
rect 7553 12750 8870 12802
rect 38 12728 8870 12750
rect 4836 12552 4842 12564
rect 3198 12524 4842 12552
rect 2076 12444 2082 12496
rect 2134 12484 2140 12496
rect 3198 12493 3226 12524
rect 4836 12512 4842 12524
rect 4894 12512 4900 12564
rect 5943 12555 6001 12561
rect 5943 12521 5955 12555
rect 5989 12552 6001 12555
rect 6492 12552 6498 12564
rect 5989 12524 6498 12552
rect 5989 12521 6001 12524
rect 5943 12515 6001 12521
rect 6492 12512 6498 12524
rect 6550 12512 6556 12564
rect 6676 12512 6682 12564
rect 6734 12552 6740 12564
rect 7691 12555 7749 12561
rect 7691 12552 7703 12555
rect 6734 12524 7703 12552
rect 6734 12512 6740 12524
rect 7691 12521 7703 12524
rect 7737 12521 7749 12555
rect 7691 12515 7749 12521
rect 3183 12487 3241 12493
rect 3183 12484 3195 12487
rect 2134 12456 3195 12484
rect 2134 12444 2140 12456
rect 3183 12453 3195 12456
rect 3229 12453 3241 12487
rect 3183 12447 3241 12453
rect 4192 12444 4198 12496
rect 4250 12484 4256 12496
rect 4471 12487 4529 12493
rect 4471 12484 4483 12487
rect 4250 12456 4483 12484
rect 4250 12444 4256 12456
rect 4471 12453 4483 12456
rect 4517 12484 4529 12487
rect 5664 12484 5670 12496
rect 4517 12456 5670 12484
rect 4517 12453 4529 12456
rect 4471 12447 4529 12453
rect 5664 12444 5670 12456
rect 5722 12444 5728 12496
rect 4287 12419 4345 12425
rect 4287 12385 4299 12419
rect 4333 12416 4345 12419
rect 4652 12416 4658 12428
rect 4333 12388 4658 12416
rect 4333 12385 4345 12388
rect 4287 12379 4345 12385
rect 4652 12376 4658 12388
rect 4710 12376 4716 12428
rect 3367 12351 3425 12357
rect 3367 12317 3379 12351
rect 3413 12348 3425 12351
rect 3640 12348 3646 12360
rect 3413 12320 3646 12348
rect 3413 12317 3425 12320
rect 3367 12311 3425 12317
rect 3640 12308 3646 12320
rect 3698 12308 3704 12360
rect 4100 12308 4106 12360
rect 4158 12348 4164 12360
rect 4563 12351 4621 12357
rect 4563 12348 4575 12351
rect 4158 12320 4575 12348
rect 4158 12308 4164 12320
rect 4563 12317 4575 12320
rect 4609 12317 4621 12351
rect 4563 12311 4621 12317
rect 6308 12308 6314 12360
rect 6366 12348 6372 12360
rect 6418 12348 6446 12402
rect 6366 12320 6446 12348
rect 6366 12308 6372 12320
rect 38 12258 8870 12280
rect 38 12206 2873 12258
rect 2925 12206 2937 12258
rect 2989 12206 3001 12258
rect 3053 12206 3065 12258
rect 3117 12206 5830 12258
rect 5882 12206 5894 12258
rect 5946 12206 5958 12258
rect 6010 12206 6022 12258
rect 6074 12206 8870 12258
rect 38 12184 8870 12206
rect 7044 12144 7050 12156
rect 3106 12116 7050 12144
rect 3106 12085 3134 12116
rect 7044 12104 7050 12116
rect 7102 12104 7108 12156
rect 3091 12079 3149 12085
rect 3091 12045 3103 12079
rect 3137 12045 3149 12079
rect 4744 12076 4750 12088
rect 4316 12048 4750 12076
rect 3091 12039 3149 12045
rect 4744 12036 4750 12048
rect 4802 12036 4808 12088
rect 5020 12036 5026 12088
rect 5078 12076 5084 12088
rect 5078 12048 6524 12076
rect 5078 12036 5084 12048
rect 5664 11968 5670 12020
rect 5722 12008 5728 12020
rect 5759 12011 5817 12017
rect 5759 12008 5771 12011
rect 5722 11980 5771 12008
rect 5722 11968 5728 11980
rect 5759 11977 5771 11980
rect 5805 11977 5817 12011
rect 5759 11971 5817 11977
rect 2628 11900 2634 11952
rect 2686 11940 2692 11952
rect 2815 11943 2873 11949
rect 2815 11940 2827 11943
rect 2686 11912 2827 11940
rect 2686 11900 2692 11912
rect 2815 11909 2827 11912
rect 2861 11909 2873 11943
rect 4836 11940 4842 11952
rect 4797 11912 4842 11940
rect 2815 11903 2873 11909
rect 4836 11900 4842 11912
rect 4894 11900 4900 11952
rect 6035 11943 6093 11949
rect 6035 11909 6047 11943
rect 6081 11940 6093 11943
rect 7783 11943 7841 11949
rect 6081 11912 7090 11940
rect 6081 11909 6093 11912
rect 6035 11903 6093 11909
rect 7062 11804 7090 11912
rect 7783 11909 7795 11943
rect 7829 11909 7841 11943
rect 7783 11903 7841 11909
rect 7136 11832 7142 11884
rect 7194 11872 7200 11884
rect 7798 11872 7826 11903
rect 7194 11844 7826 11872
rect 7194 11832 7200 11844
rect 7967 11807 8025 11813
rect 7967 11804 7979 11807
rect 7062 11776 7979 11804
rect 7967 11773 7979 11776
rect 8013 11804 8025 11807
rect 15692 11804 15698 11816
rect 8013 11776 15698 11804
rect 8013 11773 8025 11776
rect 7967 11767 8025 11773
rect 15692 11764 15698 11776
rect 15750 11764 15756 11816
rect 38 11714 8870 11736
rect 38 11662 1394 11714
rect 1446 11662 1458 11714
rect 1510 11662 1522 11714
rect 1574 11662 1586 11714
rect 1638 11662 4352 11714
rect 4404 11662 4416 11714
rect 4468 11662 4480 11714
rect 4532 11662 4544 11714
rect 4596 11662 7309 11714
rect 7361 11662 7373 11714
rect 7425 11662 7437 11714
rect 7489 11662 7501 11714
rect 7553 11662 8870 11714
rect 38 11640 8870 11662
rect 6584 11600 6590 11612
rect 4486 11572 6590 11600
rect 3548 11464 3554 11476
rect 2094 11436 3554 11464
rect 2094 11408 2122 11436
rect 3548 11424 3554 11436
rect 3606 11424 3612 11476
rect 4486 11473 4514 11572
rect 6584 11560 6590 11572
rect 6642 11560 6648 11612
rect 4471 11467 4529 11473
rect 4471 11433 4483 11467
rect 4517 11433 4529 11467
rect 4471 11427 4529 11433
rect 4836 11424 4842 11476
rect 4894 11464 4900 11476
rect 5943 11467 6001 11473
rect 5943 11464 5955 11467
rect 4894 11436 5955 11464
rect 4894 11424 4900 11436
rect 5943 11433 5955 11436
rect 5989 11464 6001 11467
rect 9252 11464 9258 11476
rect 5989 11436 9258 11464
rect 5989 11433 6001 11436
rect 5943 11427 6001 11433
rect 9252 11424 9258 11436
rect 9310 11424 9316 11476
rect 604 11356 610 11408
rect 662 11396 668 11408
rect 1803 11399 1861 11405
rect 1803 11396 1815 11399
rect 662 11368 1815 11396
rect 662 11356 668 11368
rect 1803 11365 1815 11368
rect 1849 11396 1861 11399
rect 2076 11396 2082 11408
rect 1849 11368 2082 11396
rect 1849 11365 1861 11368
rect 1803 11359 1861 11365
rect 2076 11356 2082 11368
rect 2134 11356 2140 11408
rect 2999 11399 3057 11405
rect 2999 11365 3011 11399
rect 3045 11365 3057 11399
rect 2999 11359 3057 11365
rect 4379 11399 4437 11405
rect 4379 11365 4391 11399
rect 4425 11365 4437 11399
rect 4379 11359 4437 11365
rect 4747 11399 4805 11405
rect 4747 11365 4759 11399
rect 4793 11365 4805 11399
rect 4747 11359 4805 11365
rect 696 11288 702 11340
rect 754 11328 760 11340
rect 3014 11328 3042 11359
rect 754 11300 3042 11328
rect 754 11288 760 11300
rect 1984 11260 1990 11272
rect 1945 11232 1990 11260
rect 1984 11220 1990 11232
rect 2042 11220 2048 11272
rect 3180 11260 3186 11272
rect 3141 11232 3186 11260
rect 3180 11220 3186 11232
rect 3238 11220 3244 11272
rect 4394 11260 4422 11359
rect 4762 11328 4790 11359
rect 5572 11356 5578 11408
rect 5630 11396 5636 11408
rect 5667 11399 5725 11405
rect 5667 11396 5679 11399
rect 5630 11368 5679 11396
rect 5630 11356 5636 11368
rect 5667 11365 5679 11368
rect 5713 11365 5725 11399
rect 5667 11359 5725 11365
rect 4836 11328 4842 11340
rect 4762 11300 4842 11328
rect 4836 11288 4842 11300
rect 4894 11288 4900 11340
rect 4928 11288 4934 11340
rect 4986 11328 4992 11340
rect 7688 11328 7694 11340
rect 4986 11300 6432 11328
rect 7649 11300 7694 11328
rect 4986 11288 4992 11300
rect 7688 11288 7694 11300
rect 7746 11288 7752 11340
rect 7872 11260 7878 11272
rect 4394 11232 7878 11260
rect 7872 11220 7878 11232
rect 7930 11220 7936 11272
rect 38 11170 8870 11192
rect 38 11118 2873 11170
rect 2925 11118 2937 11170
rect 2989 11118 3001 11170
rect 3053 11118 3065 11170
rect 3117 11118 5830 11170
rect 5882 11118 5894 11170
rect 5946 11118 5958 11170
rect 6010 11118 6022 11170
rect 6074 11118 8870 11170
rect 38 11096 8870 11118
rect 788 11016 794 11068
rect 846 11056 852 11068
rect 1892 11056 1898 11068
rect 846 11028 1898 11056
rect 846 11016 852 11028
rect 1892 11016 1898 11028
rect 1950 11016 1956 11068
rect 1984 11016 1990 11068
rect 2042 11056 2048 11068
rect 2042 11028 6538 11056
rect 2042 11016 2048 11028
rect 2720 10948 2726 11000
rect 2778 10988 2784 11000
rect 4839 10991 4897 10997
rect 2778 10960 3580 10988
rect 2778 10948 2784 10960
rect 4839 10957 4851 10991
rect 4885 10988 4897 10991
rect 6035 10991 6093 10997
rect 6035 10988 6047 10991
rect 4885 10960 6047 10988
rect 4885 10957 4897 10960
rect 4839 10951 4897 10957
rect 6035 10957 6047 10960
rect 6081 10988 6093 10991
rect 6124 10988 6130 11000
rect 6081 10960 6130 10988
rect 6081 10957 6093 10960
rect 6035 10951 6093 10957
rect 6124 10948 6130 10960
rect 6182 10948 6188 11000
rect 6510 10974 6538 11028
rect 604 10920 610 10932
rect 565 10892 610 10920
rect 604 10880 610 10892
rect 662 10880 668 10932
rect 1708 10880 1714 10932
rect 1766 10920 1772 10932
rect 1766 10892 1811 10920
rect 1766 10880 1772 10892
rect 2628 10812 2634 10864
rect 2686 10852 2692 10864
rect 2815 10855 2873 10861
rect 2815 10852 2827 10855
rect 2686 10824 2827 10852
rect 2686 10812 2692 10824
rect 2815 10821 2827 10824
rect 2861 10821 2873 10855
rect 4652 10852 4658 10864
rect 2815 10815 2873 10821
rect 2922 10824 4658 10852
rect 791 10787 849 10793
rect 791 10753 803 10787
rect 837 10784 849 10787
rect 2922 10784 2950 10824
rect 4652 10812 4658 10824
rect 4710 10812 4716 10864
rect 5572 10812 5578 10864
rect 5630 10852 5636 10864
rect 5759 10855 5817 10861
rect 5759 10852 5771 10855
rect 5630 10824 5771 10852
rect 5630 10812 5636 10824
rect 5759 10821 5771 10824
rect 5805 10821 5817 10855
rect 5759 10815 5817 10821
rect 7783 10855 7841 10861
rect 7783 10821 7795 10855
rect 7829 10852 7841 10855
rect 15600 10852 15606 10864
rect 7829 10824 15606 10852
rect 7829 10821 7841 10824
rect 7783 10815 7841 10821
rect 15600 10812 15606 10824
rect 15658 10812 15664 10864
rect 837 10756 2950 10784
rect 837 10753 849 10756
rect 791 10747 849 10753
rect 3078 10719 3136 10725
rect 3078 10685 3090 10719
rect 3124 10716 3136 10719
rect 6676 10716 6682 10728
rect 3124 10688 6682 10716
rect 3124 10685 3136 10688
rect 3078 10679 3136 10685
rect 6676 10676 6682 10688
rect 6734 10676 6740 10728
rect 38 10626 8870 10648
rect 38 10574 1394 10626
rect 1446 10574 1458 10626
rect 1510 10574 1522 10626
rect 1574 10574 1586 10626
rect 1638 10574 4352 10626
rect 4404 10574 4416 10626
rect 4468 10574 4480 10626
rect 4532 10574 4544 10626
rect 4596 10574 7309 10626
rect 7361 10574 7373 10626
rect 7425 10574 7437 10626
rect 7489 10574 7501 10626
rect 7553 10574 8870 10626
rect 38 10552 8870 10574
rect 8608 10512 8614 10524
rect 3934 10484 8614 10512
rect 1527 10379 1585 10385
rect 1527 10345 1539 10379
rect 1573 10376 1585 10379
rect 2628 10376 2634 10388
rect 1573 10348 2634 10376
rect 1573 10345 1585 10348
rect 1527 10339 1585 10345
rect 2628 10336 2634 10348
rect 2686 10336 2692 10388
rect 3275 10379 3333 10385
rect 3275 10345 3287 10379
rect 3321 10376 3333 10379
rect 3934 10376 3962 10484
rect 8608 10472 8614 10484
rect 8666 10472 8672 10524
rect 4928 10444 4934 10456
rect 3321 10348 3962 10376
rect 4026 10416 4934 10444
rect 3321 10345 3333 10348
rect 3275 10339 3333 10345
rect 423 10311 481 10317
rect 423 10277 435 10311
rect 469 10308 481 10311
rect 788 10308 794 10320
rect 469 10280 794 10308
rect 469 10277 481 10280
rect 423 10271 481 10277
rect 788 10268 794 10280
rect 846 10268 852 10320
rect 1619 10311 1677 10317
rect 1619 10277 1631 10311
rect 1665 10308 1677 10311
rect 3364 10308 3370 10320
rect 1665 10280 3370 10308
rect 1665 10277 1677 10280
rect 1619 10271 1677 10277
rect 3364 10268 3370 10280
rect 3422 10268 3428 10320
rect 3732 10308 3738 10320
rect 3693 10280 3738 10308
rect 3732 10268 3738 10280
rect 3790 10268 3796 10320
rect 3824 10268 3830 10320
rect 3882 10308 3888 10320
rect 3919 10311 3977 10317
rect 3919 10308 3931 10311
rect 3882 10280 3931 10308
rect 3882 10268 3888 10280
rect 3919 10277 3931 10280
rect 3965 10277 3977 10311
rect 3919 10271 3977 10277
rect 2076 10240 2082 10252
rect 2037 10212 2082 10240
rect 2076 10200 2082 10212
rect 2134 10200 2140 10252
rect 607 10175 665 10181
rect 607 10141 619 10175
rect 653 10172 665 10175
rect 4026 10172 4054 10416
rect 4928 10404 4934 10416
rect 4986 10404 4992 10456
rect 7323 10379 7381 10385
rect 7323 10376 7335 10379
rect 4670 10348 7335 10376
rect 4195 10311 4253 10317
rect 4195 10277 4207 10311
rect 4241 10277 4253 10311
rect 4468 10308 4474 10320
rect 4429 10280 4474 10308
rect 4195 10271 4253 10277
rect 4210 10240 4238 10271
rect 4468 10268 4474 10280
rect 4526 10268 4532 10320
rect 4670 10240 4698 10348
rect 7323 10345 7335 10348
rect 7369 10345 7381 10379
rect 7323 10339 7381 10345
rect 4747 10311 4805 10317
rect 4747 10277 4759 10311
rect 4793 10308 4805 10311
rect 4836 10308 4842 10320
rect 4793 10280 4842 10308
rect 4793 10277 4805 10280
rect 4747 10271 4805 10277
rect 4836 10268 4842 10280
rect 4894 10268 4900 10320
rect 5572 10308 5578 10320
rect 5533 10280 5578 10308
rect 5572 10268 5578 10280
rect 5630 10268 5636 10320
rect 5664 10268 5670 10320
rect 5722 10308 5728 10320
rect 5943 10311 6001 10317
rect 5943 10308 5955 10311
rect 5722 10280 5955 10308
rect 5722 10268 5728 10280
rect 5943 10277 5955 10280
rect 5989 10277 6001 10311
rect 5943 10271 6001 10277
rect 7596 10240 7602 10252
rect 4210 10212 4698 10240
rect 6984 10212 7602 10240
rect 7596 10200 7602 10212
rect 7654 10200 7660 10252
rect 653 10144 4054 10172
rect 653 10141 665 10144
rect 607 10135 665 10141
rect 4468 10132 4474 10184
rect 4526 10172 4532 10184
rect 8608 10172 8614 10184
rect 4526 10144 8614 10172
rect 4526 10132 4532 10144
rect 8608 10132 8614 10144
rect 8666 10132 8672 10184
rect 38 10082 8870 10104
rect 38 10030 2873 10082
rect 2925 10030 2937 10082
rect 2989 10030 3001 10082
rect 3053 10030 3065 10082
rect 3117 10030 5830 10082
rect 5882 10030 5894 10082
rect 5946 10030 5958 10082
rect 6010 10030 6022 10082
rect 6074 10030 8870 10082
rect 38 10008 8870 10030
rect 8902 10008 11414 10036
rect 1708 9928 1714 9980
rect 1766 9968 1772 9980
rect 1895 9971 1953 9977
rect 1895 9968 1907 9971
rect 1766 9940 1907 9968
rect 1766 9928 1772 9940
rect 1895 9937 1907 9940
rect 1941 9937 1953 9971
rect 4100 9968 4106 9980
rect 1895 9931 1953 9937
rect 3106 9940 4106 9968
rect 3106 9900 3134 9940
rect 4100 9928 4106 9940
rect 4158 9928 4164 9980
rect 8700 9928 8706 9980
rect 8758 9968 8764 9980
rect 8902 9968 8930 10008
rect 8758 9940 8930 9968
rect 11386 9968 11414 10008
rect 23788 9968 23794 9980
rect 11386 9940 23794 9968
rect 8758 9928 8764 9940
rect 23788 9928 23794 9940
rect 23846 9928 23852 9980
rect 1726 9872 3134 9900
rect 607 9835 665 9841
rect 607 9801 619 9835
rect 653 9832 665 9835
rect 696 9832 702 9844
rect 653 9804 702 9832
rect 653 9801 665 9804
rect 607 9795 665 9801
rect 696 9792 702 9804
rect 754 9792 760 9844
rect 1726 9841 1754 9872
rect 3180 9860 3186 9912
rect 3238 9900 3244 9912
rect 3238 9872 3580 9900
rect 3238 9860 3244 9872
rect 4652 9860 4658 9912
rect 4710 9900 4716 9912
rect 4710 9872 6524 9900
rect 4710 9860 4716 9872
rect 1711 9835 1769 9841
rect 1711 9801 1723 9835
rect 1757 9801 1769 9835
rect 1711 9795 1769 9801
rect 2628 9792 2634 9844
rect 2686 9832 2692 9844
rect 2815 9835 2873 9841
rect 2815 9832 2827 9835
rect 2686 9804 2827 9832
rect 2686 9792 2692 9804
rect 2815 9801 2827 9804
rect 2861 9801 2873 9835
rect 2815 9795 2873 9801
rect 5572 9792 5578 9844
rect 5630 9832 5636 9844
rect 5759 9835 5817 9841
rect 5759 9832 5771 9835
rect 5630 9804 5771 9832
rect 5630 9792 5636 9804
rect 5759 9801 5771 9804
rect 5805 9801 5817 9835
rect 5759 9795 5817 9801
rect 3091 9767 3149 9773
rect 3091 9733 3103 9767
rect 3137 9764 3149 9767
rect 4100 9764 4106 9776
rect 3137 9736 4106 9764
rect 3137 9733 3149 9736
rect 3091 9727 3149 9733
rect 4100 9724 4106 9736
rect 4158 9724 4164 9776
rect 4744 9724 4750 9776
rect 4802 9764 4808 9776
rect 4839 9767 4897 9773
rect 4839 9764 4851 9767
rect 4802 9736 4851 9764
rect 4802 9724 4808 9736
rect 4839 9733 4851 9736
rect 4885 9764 4897 9767
rect 5664 9764 5670 9776
rect 4885 9736 5670 9764
rect 4885 9733 4897 9736
rect 4839 9727 4897 9733
rect 5664 9724 5670 9736
rect 5722 9724 5728 9776
rect 6035 9767 6093 9773
rect 6035 9733 6047 9767
rect 6081 9764 6093 9767
rect 6676 9764 6682 9776
rect 6081 9736 6682 9764
rect 6081 9733 6093 9736
rect 6035 9727 6093 9733
rect 6676 9724 6682 9736
rect 6734 9724 6740 9776
rect 7783 9767 7841 9773
rect 7783 9733 7795 9767
rect 7829 9764 7841 9767
rect 11460 9764 11466 9776
rect 7829 9736 11466 9764
rect 7829 9733 7841 9736
rect 7783 9727 7841 9733
rect 11460 9724 11466 9736
rect 11518 9724 11524 9776
rect 791 9699 849 9705
rect 791 9665 803 9699
rect 837 9696 849 9699
rect 837 9668 2950 9696
rect 837 9665 849 9668
rect 791 9659 849 9665
rect 2922 9628 2950 9668
rect 5020 9628 5026 9640
rect 2922 9600 5026 9628
rect 5020 9588 5026 9600
rect 5078 9588 5084 9640
rect 38 9538 8870 9560
rect 38 9486 1394 9538
rect 1446 9486 1458 9538
rect 1510 9486 1522 9538
rect 1574 9486 1586 9538
rect 1638 9486 4352 9538
rect 4404 9486 4416 9538
rect 4468 9486 4480 9538
rect 4532 9486 4544 9538
rect 4596 9486 7309 9538
rect 7361 9486 7373 9538
rect 7425 9486 7437 9538
rect 7489 9486 7501 9538
rect 7553 9486 8870 9538
rect 38 9464 8870 9486
rect 4100 9384 4106 9436
rect 4158 9424 4164 9436
rect 5940 9424 5946 9436
rect 4158 9396 5946 9424
rect 4158 9384 4164 9396
rect 5940 9384 5946 9396
rect 5998 9424 6004 9436
rect 7136 9424 7142 9436
rect 5998 9396 7142 9424
rect 5998 9384 6004 9396
rect 7136 9384 7142 9396
rect 7194 9384 7200 9436
rect 3916 9316 3922 9368
rect 3974 9356 3980 9368
rect 5023 9359 5081 9365
rect 5023 9356 5035 9359
rect 3974 9328 5035 9356
rect 3974 9316 3980 9328
rect 5023 9325 5035 9328
rect 5069 9325 5081 9359
rect 5023 9319 5081 9325
rect 11279 9291 11337 9297
rect 11279 9288 11291 9291
rect 3750 9260 11291 9288
rect 512 9180 518 9232
rect 570 9220 576 9232
rect 687 9223 745 9229
rect 687 9220 699 9223
rect 570 9192 699 9220
rect 570 9180 576 9192
rect 687 9189 699 9192
rect 733 9189 745 9223
rect 1800 9220 1806 9232
rect 1761 9192 1806 9220
rect 687 9183 745 9189
rect 1800 9180 1806 9192
rect 1858 9180 1864 9232
rect 3750 9229 3778 9260
rect 11279 9257 11291 9260
rect 11325 9257 11337 9291
rect 11279 9251 11337 9257
rect 11371 9291 11429 9297
rect 11371 9257 11383 9291
rect 11417 9288 11429 9291
rect 15968 9288 15974 9300
rect 11417 9260 15974 9288
rect 11417 9257 11429 9260
rect 11371 9251 11429 9257
rect 15968 9248 15974 9260
rect 16026 9248 16032 9300
rect 3735 9223 3793 9229
rect 3735 9189 3747 9223
rect 3781 9189 3793 9223
rect 5572 9220 5578 9232
rect 5533 9192 5578 9220
rect 3735 9183 3793 9189
rect 5572 9180 5578 9192
rect 5630 9180 5636 9232
rect 5940 9220 5946 9232
rect 5901 9192 5946 9220
rect 5940 9180 5946 9192
rect 5998 9180 6004 9232
rect 7780 9152 7786 9164
rect 2002 9124 5158 9152
rect 6984 9124 7786 9152
rect 880 9084 886 9096
rect 841 9056 886 9084
rect 880 9044 886 9056
rect 938 9044 944 9096
rect 2002 9093 2030 9124
rect 1987 9087 2045 9093
rect 1987 9053 1999 9087
rect 2033 9053 2045 9087
rect 5130 9084 5158 9124
rect 7780 9112 7786 9124
rect 7838 9112 7844 9164
rect 6400 9084 6406 9096
rect 5130 9056 6406 9084
rect 1987 9047 2045 9053
rect 6400 9044 6406 9056
rect 6458 9044 6464 9096
rect 7691 9087 7749 9093
rect 7691 9053 7703 9087
rect 7737 9084 7749 9087
rect 7964 9084 7970 9096
rect 7737 9056 7970 9084
rect 7737 9053 7749 9056
rect 7691 9047 7749 9053
rect 7964 9044 7970 9056
rect 8022 9044 8028 9096
rect 11279 9087 11337 9093
rect 11279 9053 11291 9087
rect 11325 9084 11337 9087
rect 24064 9084 24070 9096
rect 11325 9056 24070 9084
rect 11325 9053 11337 9056
rect 11279 9047 11337 9053
rect 24064 9044 24070 9056
rect 24122 9044 24128 9096
rect 38 8994 8870 9016
rect 38 8942 2873 8994
rect 2925 8942 2937 8994
rect 2989 8942 3001 8994
rect 3053 8942 3065 8994
rect 3117 8942 5830 8994
rect 5882 8942 5894 8994
rect 5946 8942 5958 8994
rect 6010 8942 6022 8994
rect 6074 8942 8870 8994
rect 38 8920 8870 8942
rect 1800 8840 1806 8892
rect 1858 8880 1864 8892
rect 1895 8883 1953 8889
rect 1895 8880 1907 8883
rect 1858 8852 1907 8880
rect 1858 8840 1864 8852
rect 1895 8849 1907 8852
rect 1941 8849 1953 8883
rect 1895 8843 1953 8849
rect 4652 8840 4658 8892
rect 4710 8880 4716 8892
rect 11279 8883 11337 8889
rect 11279 8880 11291 8883
rect 4710 8852 11291 8880
rect 4710 8840 4716 8852
rect 11279 8849 11291 8852
rect 11325 8849 11337 8883
rect 11279 8843 11337 8849
rect 880 8772 886 8824
rect 938 8812 944 8824
rect 6035 8815 6093 8821
rect 6035 8812 6047 8815
rect 938 8784 3580 8812
rect 4854 8784 6047 8812
rect 938 8772 944 8784
rect 604 8744 610 8756
rect 565 8716 610 8744
rect 604 8704 610 8716
rect 662 8744 668 8756
rect 1616 8744 1622 8756
rect 662 8716 1622 8744
rect 662 8704 668 8716
rect 1616 8704 1622 8716
rect 1674 8744 1680 8756
rect 1711 8747 1769 8753
rect 1711 8744 1723 8747
rect 1674 8716 1723 8744
rect 1674 8704 1680 8716
rect 1711 8713 1723 8716
rect 1757 8713 1769 8747
rect 4744 8744 4750 8756
rect 1711 8707 1769 8713
rect 4670 8716 4750 8744
rect 2536 8636 2542 8688
rect 2594 8676 2600 8688
rect 2815 8679 2873 8685
rect 2815 8676 2827 8679
rect 2594 8648 2827 8676
rect 2594 8636 2600 8648
rect 2815 8645 2827 8648
rect 2861 8645 2873 8679
rect 2815 8639 2873 8645
rect 3091 8679 3149 8685
rect 3091 8645 3103 8679
rect 3137 8676 3149 8679
rect 4670 8676 4698 8716
rect 4744 8704 4750 8716
rect 4802 8704 4808 8756
rect 4854 8688 4882 8784
rect 6035 8781 6047 8784
rect 6081 8781 6093 8815
rect 6035 8775 6093 8781
rect 6492 8772 6498 8824
rect 6550 8772 6556 8824
rect 7872 8772 7878 8824
rect 7930 8812 7936 8824
rect 8516 8812 8522 8824
rect 7930 8784 8522 8812
rect 7930 8772 7936 8784
rect 8516 8772 8522 8784
rect 8574 8812 8580 8824
rect 11368 8812 11374 8824
rect 8574 8784 11374 8812
rect 8574 8772 8580 8784
rect 11368 8772 11374 8784
rect 11426 8772 11432 8824
rect 5572 8704 5578 8756
rect 5630 8744 5636 8756
rect 5759 8747 5817 8753
rect 5759 8744 5771 8747
rect 5630 8716 5771 8744
rect 5630 8704 5636 8716
rect 5759 8713 5771 8716
rect 5805 8713 5817 8747
rect 5759 8707 5817 8713
rect 8608 8704 8614 8756
rect 8666 8744 8672 8756
rect 11644 8744 11650 8756
rect 8666 8716 11650 8744
rect 8666 8704 8672 8716
rect 11644 8704 11650 8716
rect 11702 8704 11708 8756
rect 4836 8676 4842 8688
rect 3137 8648 4698 8676
rect 4797 8648 4842 8676
rect 3137 8645 3149 8648
rect 3091 8639 3149 8645
rect 4836 8636 4842 8648
rect 4894 8636 4900 8688
rect 7783 8679 7841 8685
rect 4946 8648 7090 8676
rect 4100 8568 4106 8620
rect 4158 8608 4164 8620
rect 4946 8608 4974 8648
rect 4158 8580 4974 8608
rect 7062 8608 7090 8648
rect 7783 8645 7795 8679
rect 7829 8676 7841 8679
rect 11460 8676 11466 8688
rect 7829 8648 11466 8676
rect 7829 8645 7841 8648
rect 7783 8639 7841 8645
rect 11460 8636 11466 8648
rect 11518 8636 11524 8688
rect 7964 8608 7970 8620
rect 7062 8580 7970 8608
rect 4158 8568 4164 8580
rect 7964 8568 7970 8580
rect 8022 8568 8028 8620
rect 512 8500 518 8552
rect 570 8540 576 8552
rect 791 8543 849 8549
rect 791 8540 803 8543
rect 570 8512 803 8540
rect 570 8500 576 8512
rect 791 8509 803 8512
rect 837 8540 849 8543
rect 1984 8540 1990 8552
rect 837 8512 1990 8540
rect 837 8509 849 8512
rect 791 8503 849 8509
rect 1984 8500 1990 8512
rect 2042 8500 2048 8552
rect 2168 8500 2174 8552
rect 2226 8540 2232 8552
rect 6400 8540 6406 8552
rect 2226 8512 6406 8540
rect 2226 8500 2232 8512
rect 6400 8500 6406 8512
rect 6458 8500 6464 8552
rect 38 8450 8870 8472
rect 38 8398 1394 8450
rect 1446 8398 1458 8450
rect 1510 8398 1522 8450
rect 1574 8398 1586 8450
rect 1638 8398 4352 8450
rect 4404 8398 4416 8450
rect 4468 8398 4480 8450
rect 4532 8398 4544 8450
rect 4596 8398 7309 8450
rect 7361 8398 7373 8450
rect 7425 8398 7437 8450
rect 7489 8398 7501 8450
rect 7553 8398 8870 8450
rect 38 8376 8870 8398
rect 1987 8339 2045 8345
rect 1987 8305 1999 8339
rect 2033 8336 2045 8339
rect 2168 8336 2174 8348
rect 2033 8308 2174 8336
rect 2033 8305 2045 8308
rect 1987 8299 2045 8305
rect 2168 8296 2174 8308
rect 2226 8296 2232 8348
rect 8332 8296 8338 8348
rect 8390 8336 8396 8348
rect 8608 8336 8614 8348
rect 8390 8308 8614 8336
rect 8390 8296 8396 8308
rect 8608 8296 8614 8308
rect 8666 8296 8672 8348
rect 883 8271 941 8277
rect 883 8237 895 8271
rect 929 8268 941 8271
rect 2628 8268 2634 8280
rect 929 8240 2634 8268
rect 929 8237 941 8240
rect 883 8231 941 8237
rect 2628 8228 2634 8240
rect 2686 8228 2692 8280
rect 3364 8228 3370 8280
rect 3422 8268 3428 8280
rect 3732 8268 3738 8280
rect 3422 8240 3738 8268
rect 3422 8228 3428 8240
rect 3732 8228 3738 8240
rect 3790 8268 3796 8280
rect 4100 8268 4106 8280
rect 3790 8240 4106 8268
rect 3790 8228 3796 8240
rect 4100 8228 4106 8240
rect 4158 8228 4164 8280
rect 3272 8200 3278 8212
rect 3233 8172 3278 8200
rect 3272 8160 3278 8172
rect 3330 8160 3336 8212
rect 512 8092 518 8144
rect 570 8132 576 8144
rect 687 8135 745 8141
rect 687 8132 699 8135
rect 570 8104 699 8132
rect 570 8092 576 8104
rect 687 8101 699 8104
rect 733 8101 745 8135
rect 1800 8132 1806 8144
rect 1761 8104 1806 8132
rect 687 8095 745 8101
rect 1800 8092 1806 8104
rect 1858 8092 1864 8144
rect 2999 8135 3057 8141
rect 2999 8101 3011 8135
rect 3045 8101 3057 8135
rect 3732 8132 3738 8144
rect 3693 8104 3738 8132
rect 2999 8095 3057 8101
rect 3014 8064 3042 8095
rect 3732 8092 3738 8104
rect 3790 8092 3796 8144
rect 4008 8132 4014 8144
rect 3969 8104 4014 8132
rect 4008 8092 4014 8104
rect 4066 8092 4072 8144
rect 4118 8141 4146 8228
rect 4652 8200 4658 8212
rect 4613 8172 4658 8200
rect 4652 8160 4658 8172
rect 4710 8160 4716 8212
rect 5572 8200 5578 8212
rect 5533 8172 5578 8200
rect 5572 8160 5578 8172
rect 5630 8160 5636 8212
rect 5943 8203 6001 8209
rect 5943 8169 5955 8203
rect 5989 8200 6001 8203
rect 6216 8200 6222 8212
rect 5989 8172 6222 8200
rect 5989 8169 6001 8172
rect 5943 8163 6001 8169
rect 6216 8160 6222 8172
rect 6274 8160 6280 8212
rect 4103 8135 4161 8141
rect 4103 8101 4115 8135
rect 4149 8101 4161 8135
rect 4103 8095 4161 8101
rect 4563 8135 4621 8141
rect 4563 8101 4575 8135
rect 4609 8132 4621 8135
rect 4928 8132 4934 8144
rect 4609 8104 4934 8132
rect 4609 8101 4621 8104
rect 4563 8095 4621 8101
rect 3364 8064 3370 8076
rect 3014 8036 3370 8064
rect 3364 8024 3370 8036
rect 3422 8024 3428 8076
rect 3091 7999 3149 8005
rect 3091 7965 3103 7999
rect 3137 7996 3149 7999
rect 4578 7996 4606 8095
rect 4928 8092 4934 8104
rect 4986 8092 4992 8144
rect 7596 8064 7602 8076
rect 6984 8036 7602 8064
rect 7596 8024 7602 8036
rect 7654 8024 7660 8076
rect 7691 8067 7749 8073
rect 7691 8033 7703 8067
rect 7737 8064 7749 8067
rect 7872 8064 7878 8076
rect 7737 8036 7878 8064
rect 7737 8033 7749 8036
rect 7691 8027 7749 8033
rect 7872 8024 7878 8036
rect 7930 8024 7936 8076
rect 3137 7968 4606 7996
rect 3137 7965 3149 7968
rect 3091 7959 3149 7965
rect 38 7906 8870 7928
rect 38 7854 2873 7906
rect 2925 7854 2937 7906
rect 2989 7854 3001 7906
rect 3053 7854 3065 7906
rect 3117 7854 5830 7906
rect 5882 7854 5894 7906
rect 5946 7854 5958 7906
rect 6010 7854 6022 7906
rect 6074 7854 8870 7906
rect 38 7832 8870 7854
rect 696 7752 702 7804
rect 754 7792 760 7804
rect 791 7795 849 7801
rect 791 7792 803 7795
rect 754 7764 803 7792
rect 754 7752 760 7764
rect 791 7761 803 7764
rect 837 7761 849 7795
rect 4836 7792 4842 7804
rect 791 7755 849 7761
rect 3106 7764 4842 7792
rect 3106 7733 3134 7764
rect 4836 7752 4842 7764
rect 4894 7752 4900 7804
rect 3091 7727 3149 7733
rect 3091 7693 3103 7727
rect 3137 7693 3149 7727
rect 3091 7687 3149 7693
rect 3364 7684 3370 7736
rect 3422 7724 3428 7736
rect 6035 7727 6093 7733
rect 6035 7724 6047 7727
rect 3422 7696 3580 7724
rect 4854 7696 6047 7724
rect 3422 7684 3428 7696
rect 604 7656 610 7668
rect 565 7628 610 7656
rect 604 7616 610 7628
rect 662 7616 668 7668
rect 1711 7659 1769 7665
rect 1711 7625 1723 7659
rect 1757 7656 1769 7659
rect 1800 7656 1806 7668
rect 1757 7628 1806 7656
rect 1757 7625 1769 7628
rect 1711 7619 1769 7625
rect 1800 7616 1806 7628
rect 1858 7616 1864 7668
rect 2536 7616 2542 7668
rect 2594 7656 2600 7668
rect 2815 7659 2873 7665
rect 2815 7656 2827 7659
rect 2594 7628 2827 7656
rect 2594 7616 2600 7628
rect 2815 7625 2827 7628
rect 2861 7625 2873 7659
rect 2815 7619 2873 7625
rect 3640 7548 3646 7600
rect 3698 7588 3704 7600
rect 3698 7560 4146 7588
rect 3698 7548 3704 7560
rect 4118 7520 4146 7560
rect 4652 7548 4658 7600
rect 4710 7588 4716 7600
rect 4854 7597 4882 7696
rect 6035 7693 6047 7696
rect 6081 7693 6093 7727
rect 6035 7687 6093 7693
rect 5572 7616 5578 7668
rect 5630 7656 5636 7668
rect 5759 7659 5817 7665
rect 5759 7656 5771 7659
rect 5630 7628 5771 7656
rect 5630 7616 5636 7628
rect 5759 7625 5771 7628
rect 5805 7625 5817 7659
rect 5759 7619 5817 7625
rect 4839 7591 4897 7597
rect 4839 7588 4851 7591
rect 4710 7560 4851 7588
rect 4710 7548 4716 7560
rect 4839 7557 4851 7560
rect 4885 7557 4897 7591
rect 7154 7588 7182 7642
rect 4839 7551 4897 7557
rect 5866 7560 7182 7588
rect 7783 7591 7841 7597
rect 5866 7520 5894 7560
rect 7783 7557 7795 7591
rect 7829 7588 7841 7591
rect 11552 7588 11558 7600
rect 7829 7560 11558 7588
rect 7829 7557 7841 7560
rect 7783 7551 7841 7557
rect 11552 7548 11558 7560
rect 11610 7548 11616 7600
rect 4118 7492 5894 7520
rect 1892 7452 1898 7464
rect 1853 7424 1898 7452
rect 1892 7412 1898 7424
rect 1950 7412 1956 7464
rect 3824 7412 3830 7464
rect 3882 7452 3888 7464
rect 4100 7452 4106 7464
rect 3882 7424 4106 7452
rect 3882 7412 3888 7424
rect 4100 7412 4106 7424
rect 4158 7452 4164 7464
rect 11279 7455 11337 7461
rect 11279 7452 11291 7455
rect 4158 7424 11291 7452
rect 4158 7412 4164 7424
rect 11279 7421 11291 7424
rect 11325 7421 11337 7455
rect 11279 7415 11337 7421
rect 38 7362 8870 7384
rect 38 7310 1394 7362
rect 1446 7310 1458 7362
rect 1510 7310 1522 7362
rect 1574 7310 1586 7362
rect 1638 7310 4352 7362
rect 4404 7310 4416 7362
rect 4468 7310 4480 7362
rect 4532 7310 4544 7362
rect 4596 7310 7309 7362
rect 7361 7310 7373 7362
rect 7425 7310 7437 7362
rect 7489 7310 7501 7362
rect 7553 7310 8870 7362
rect 38 7288 8870 7310
rect 2720 7248 2726 7260
rect 2681 7220 2726 7248
rect 2720 7208 2726 7220
rect 2778 7208 2784 7260
rect 3548 7208 3554 7260
rect 3606 7248 3612 7260
rect 4192 7248 4198 7260
rect 3606 7220 4198 7248
rect 3606 7208 3612 7220
rect 4192 7208 4198 7220
rect 4250 7248 4256 7260
rect 4563 7251 4621 7257
rect 4563 7248 4575 7251
rect 4250 7220 4575 7248
rect 4250 7208 4256 7220
rect 4563 7217 4575 7220
rect 4609 7217 4621 7251
rect 4563 7211 4621 7217
rect 1800 7140 1806 7192
rect 1858 7140 1864 7192
rect 1987 7183 2045 7189
rect 1987 7149 1999 7183
rect 2033 7180 2045 7183
rect 4836 7180 4842 7192
rect 2033 7152 4842 7180
rect 2033 7149 2045 7152
rect 1987 7143 2045 7149
rect 4836 7140 4842 7152
rect 4894 7140 4900 7192
rect 11279 7183 11337 7189
rect 11279 7149 11291 7183
rect 11325 7180 11337 7183
rect 23788 7180 23794 7192
rect 11325 7152 23794 7180
rect 11325 7149 11337 7152
rect 11279 7143 11337 7149
rect 23788 7140 23794 7152
rect 23846 7140 23852 7192
rect 1818 7112 1846 7140
rect 3643 7115 3701 7121
rect 1818 7084 2582 7112
rect 699 7047 757 7053
rect 699 7013 711 7047
rect 745 7044 757 7047
rect 788 7044 794 7056
rect 745 7016 794 7044
rect 745 7013 757 7016
rect 699 7007 757 7013
rect 788 7004 794 7016
rect 846 7004 852 7056
rect 1803 7047 1861 7053
rect 1803 7013 1815 7047
rect 1849 7044 1861 7047
rect 1984 7044 1990 7056
rect 1849 7016 1990 7044
rect 1849 7013 1861 7016
rect 1803 7007 1861 7013
rect 1984 7004 1990 7016
rect 2042 7004 2048 7056
rect 2554 7053 2582 7084
rect 3643 7081 3655 7115
rect 3689 7112 3701 7115
rect 3732 7112 3738 7124
rect 3689 7084 3738 7112
rect 3689 7081 3701 7084
rect 3643 7075 3701 7081
rect 3732 7072 3738 7084
rect 3790 7072 3796 7124
rect 7872 7112 7878 7124
rect 3934 7084 7878 7112
rect 2539 7047 2597 7053
rect 2539 7013 2551 7047
rect 2585 7013 2597 7047
rect 3548 7044 3554 7056
rect 3509 7016 3554 7044
rect 2539 7007 2597 7013
rect 3548 7004 3554 7016
rect 3606 7004 3612 7056
rect 3934 7053 3962 7084
rect 7872 7072 7878 7084
rect 7930 7072 7936 7124
rect 3919 7047 3977 7053
rect 3919 7013 3931 7047
rect 3965 7013 3977 7047
rect 4100 7044 4106 7056
rect 4061 7016 4106 7044
rect 3919 7007 3977 7013
rect 4100 7004 4106 7016
rect 4158 7004 4164 7056
rect 4379 7047 4437 7053
rect 4379 7013 4391 7047
rect 4425 7013 4437 7047
rect 4379 7007 4437 7013
rect 3180 6936 3186 6988
rect 3238 6976 3244 6988
rect 4287 6979 4345 6985
rect 4287 6976 4299 6979
rect 3238 6948 4299 6976
rect 3238 6936 3244 6948
rect 4287 6945 4299 6948
rect 4333 6945 4345 6979
rect 4287 6939 4345 6945
rect 880 6908 886 6920
rect 841 6880 886 6908
rect 880 6868 886 6880
rect 938 6868 944 6920
rect 4394 6908 4422 7007
rect 5572 7004 5578 7056
rect 5630 7044 5636 7056
rect 5667 7047 5725 7053
rect 5667 7044 5679 7047
rect 5630 7016 5679 7044
rect 5630 7004 5636 7016
rect 5667 7013 5679 7016
rect 5713 7013 5725 7047
rect 5667 7007 5725 7013
rect 5943 6979 6001 6985
rect 5943 6945 5955 6979
rect 5989 6976 6001 6979
rect 6216 6976 6222 6988
rect 5989 6948 6222 6976
rect 5989 6945 6001 6948
rect 5943 6939 6001 6945
rect 6216 6936 6222 6948
rect 6274 6936 6280 6988
rect 6400 6936 6406 6988
rect 6458 6936 6464 6988
rect 7691 6979 7749 6985
rect 7691 6945 7703 6979
rect 7737 6976 7749 6979
rect 11368 6976 11374 6988
rect 7737 6948 11374 6976
rect 7737 6945 7749 6948
rect 7691 6939 7749 6945
rect 11368 6936 11374 6948
rect 11426 6936 11432 6988
rect 6768 6908 6774 6920
rect 4394 6880 6774 6908
rect 6768 6868 6774 6880
rect 6826 6868 6832 6920
rect 38 6818 8870 6840
rect 38 6766 2873 6818
rect 2925 6766 2937 6818
rect 2989 6766 3001 6818
rect 3053 6766 3065 6818
rect 3117 6766 5830 6818
rect 5882 6766 5894 6818
rect 5946 6766 5958 6818
rect 6010 6766 6022 6818
rect 6074 6766 8870 6818
rect 38 6744 8870 6766
rect 880 6664 886 6716
rect 938 6704 944 6716
rect 938 6676 4422 6704
rect 938 6664 944 6676
rect 696 6596 702 6648
rect 754 6636 760 6648
rect 754 6608 1754 6636
rect 754 6596 760 6608
rect 1726 6580 1754 6608
rect 2628 6596 2634 6648
rect 2686 6636 2692 6648
rect 4394 6636 4422 6676
rect 2686 6608 3580 6636
rect 4394 6608 6524 6636
rect 2686 6596 2692 6608
rect 1708 6528 1714 6580
rect 1766 6568 1772 6580
rect 1766 6540 1811 6568
rect 1766 6528 1772 6540
rect 2536 6528 2542 6580
rect 2594 6568 2600 6580
rect 2815 6571 2873 6577
rect 2815 6568 2827 6571
rect 2594 6540 2827 6568
rect 2594 6528 2600 6540
rect 2815 6537 2827 6540
rect 2861 6537 2873 6571
rect 2815 6531 2873 6537
rect 5572 6528 5578 6580
rect 5630 6568 5636 6580
rect 5759 6571 5817 6577
rect 5759 6568 5771 6571
rect 5630 6540 5771 6568
rect 5630 6528 5636 6540
rect 5759 6537 5771 6540
rect 5805 6537 5817 6571
rect 5759 6531 5817 6537
rect 7688 6528 7694 6580
rect 7746 6568 7752 6580
rect 11368 6568 11374 6580
rect 7746 6540 11374 6568
rect 7746 6528 7752 6540
rect 11368 6528 11374 6540
rect 11426 6528 11432 6580
rect 3091 6503 3149 6509
rect 3091 6469 3103 6503
rect 3137 6500 3149 6503
rect 4652 6500 4658 6512
rect 3137 6472 4658 6500
rect 3137 6469 3149 6472
rect 3091 6463 3149 6469
rect 4652 6460 4658 6472
rect 4710 6460 4716 6512
rect 4839 6503 4897 6509
rect 4839 6469 4851 6503
rect 4885 6469 4897 6503
rect 4839 6463 4897 6469
rect 6035 6503 6093 6509
rect 6035 6469 6047 6503
rect 6081 6500 6093 6503
rect 6676 6500 6682 6512
rect 6081 6472 6682 6500
rect 6081 6469 6093 6472
rect 6035 6463 6093 6469
rect 1895 6367 1953 6373
rect 1895 6333 1907 6367
rect 1941 6364 1953 6367
rect 4652 6364 4658 6376
rect 1941 6336 4658 6364
rect 1941 6333 1953 6336
rect 1895 6327 1953 6333
rect 4652 6324 4658 6336
rect 4710 6324 4716 6376
rect 4854 6364 4882 6463
rect 6676 6460 6682 6472
rect 6734 6460 6740 6512
rect 6768 6460 6774 6512
rect 6826 6500 6832 6512
rect 7783 6503 7841 6509
rect 7783 6500 7795 6503
rect 6826 6472 7795 6500
rect 6826 6460 6832 6472
rect 7783 6469 7795 6472
rect 7829 6500 7841 6503
rect 11460 6500 11466 6512
rect 7829 6472 11466 6500
rect 7829 6469 7841 6472
rect 7783 6463 7841 6469
rect 11460 6460 11466 6472
rect 11518 6460 11524 6512
rect 6216 6364 6222 6376
rect 4854 6336 6222 6364
rect 6216 6324 6222 6336
rect 6274 6324 6280 6376
rect 38 6274 8870 6296
rect 38 6222 1394 6274
rect 1446 6222 1458 6274
rect 1510 6222 1522 6274
rect 1574 6222 1586 6274
rect 1638 6222 4352 6274
rect 4404 6222 4416 6274
rect 4468 6222 4480 6274
rect 4532 6222 4544 6274
rect 4596 6222 7309 6274
rect 7361 6222 7373 6274
rect 7425 6222 7437 6274
rect 7489 6222 7501 6274
rect 7553 6222 8870 6274
rect 38 6200 8870 6222
rect 1987 6163 2045 6169
rect 1987 6129 1999 6163
rect 2033 6160 2045 6163
rect 3180 6160 3186 6172
rect 2033 6132 3186 6160
rect 2033 6129 2045 6132
rect 1987 6123 2045 6129
rect 3180 6120 3186 6132
rect 3238 6120 3244 6172
rect 3364 6160 3370 6172
rect 3325 6132 3370 6160
rect 3364 6120 3370 6132
rect 3422 6120 3428 6172
rect 4008 6120 4014 6172
rect 4066 6160 4072 6172
rect 4563 6163 4621 6169
rect 4563 6160 4575 6163
rect 4066 6132 4575 6160
rect 4066 6120 4072 6132
rect 4563 6129 4575 6132
rect 4609 6129 4621 6163
rect 7688 6160 7694 6172
rect 4563 6123 4621 6129
rect 5774 6132 7694 6160
rect 5774 6092 5802 6132
rect 7688 6120 7694 6132
rect 7746 6120 7752 6172
rect 1910 6064 5802 6092
rect 1910 5965 1938 6064
rect 4928 5984 4934 6036
rect 4986 6024 4992 6036
rect 5943 6027 6001 6033
rect 5943 6024 5955 6027
rect 4986 5996 5955 6024
rect 4986 5984 4992 5996
rect 5943 5993 5955 5996
rect 5989 6024 6001 6027
rect 7688 6024 7694 6036
rect 5989 5996 7694 6024
rect 5989 5993 6001 5996
rect 5943 5987 6001 5993
rect 7688 5984 7694 5996
rect 7746 5984 7752 6036
rect 1895 5959 1953 5965
rect 1895 5925 1907 5959
rect 1941 5925 1953 5959
rect 1895 5919 1953 5925
rect 1984 5916 1990 5968
rect 2042 5956 2048 5968
rect 3183 5959 3241 5965
rect 3183 5956 3195 5959
rect 2042 5928 3195 5956
rect 2042 5916 2048 5928
rect 3183 5925 3195 5928
rect 3229 5956 3241 5959
rect 3548 5956 3554 5968
rect 3229 5928 3554 5956
rect 3229 5925 3241 5928
rect 3183 5919 3241 5925
rect 3548 5916 3554 5928
rect 3606 5916 3612 5968
rect 4192 5916 4198 5968
rect 4250 5956 4256 5968
rect 4287 5959 4345 5965
rect 4287 5956 4299 5959
rect 4250 5928 4299 5956
rect 4250 5916 4256 5928
rect 4287 5925 4299 5928
rect 4333 5925 4345 5959
rect 4287 5919 4345 5925
rect 4471 5959 4529 5965
rect 4471 5925 4483 5959
rect 4517 5956 4529 5959
rect 5296 5956 5302 5968
rect 4517 5928 5302 5956
rect 4517 5925 4529 5928
rect 4471 5919 4529 5925
rect 5296 5916 5302 5928
rect 5354 5916 5360 5968
rect 5572 5916 5578 5968
rect 5630 5956 5636 5968
rect 5667 5959 5725 5965
rect 5667 5956 5679 5959
rect 5630 5928 5679 5956
rect 5630 5916 5636 5928
rect 5667 5925 5679 5928
rect 5713 5925 5725 5959
rect 5667 5919 5725 5925
rect 7044 5916 7050 5968
rect 7102 5916 7108 5968
rect 7691 5891 7749 5897
rect 7691 5857 7703 5891
rect 7737 5888 7749 5891
rect 11552 5888 11558 5900
rect 7737 5860 11558 5888
rect 7737 5857 7749 5860
rect 7691 5851 7749 5857
rect 11552 5848 11558 5860
rect 11610 5848 11616 5900
rect 38 5730 8870 5752
rect 38 5678 2873 5730
rect 2925 5678 2937 5730
rect 2989 5678 3001 5730
rect 3053 5678 3065 5730
rect 3117 5678 5830 5730
rect 5882 5678 5894 5730
rect 5946 5678 5958 5730
rect 6010 5678 6022 5730
rect 6074 5678 8870 5730
rect 38 5656 8870 5678
rect 1892 5508 1898 5560
rect 1950 5548 1956 5560
rect 4839 5551 4897 5557
rect 1950 5520 3580 5548
rect 1950 5508 1956 5520
rect 4839 5517 4851 5551
rect 4885 5548 4897 5551
rect 5940 5548 5946 5560
rect 4885 5520 5946 5548
rect 4885 5517 4897 5520
rect 4839 5511 4897 5517
rect 5940 5508 5946 5520
rect 5998 5508 6004 5560
rect 6308 5508 6314 5560
rect 6366 5548 6372 5560
rect 6366 5520 6524 5548
rect 6366 5508 6372 5520
rect 2536 5440 2542 5492
rect 2594 5480 2600 5492
rect 2815 5483 2873 5489
rect 2815 5480 2827 5483
rect 2594 5452 2827 5480
rect 2594 5440 2600 5452
rect 2815 5449 2827 5452
rect 2861 5449 2873 5483
rect 4928 5480 4934 5492
rect 2815 5443 2873 5449
rect 4762 5452 4934 5480
rect 2830 5276 2858 5443
rect 3091 5415 3149 5421
rect 3091 5381 3103 5415
rect 3137 5412 3149 5415
rect 4762 5412 4790 5452
rect 4928 5440 4934 5452
rect 4986 5440 4992 5492
rect 5572 5440 5578 5492
rect 5630 5480 5636 5492
rect 5759 5483 5817 5489
rect 5759 5480 5771 5483
rect 5630 5452 5771 5480
rect 5630 5440 5636 5452
rect 5759 5449 5771 5452
rect 5805 5449 5817 5483
rect 5759 5443 5817 5449
rect 3137 5384 4790 5412
rect 6035 5415 6093 5421
rect 3137 5381 3149 5384
rect 3091 5375 3149 5381
rect 6035 5381 6047 5415
rect 6081 5412 6093 5415
rect 6124 5412 6130 5424
rect 6081 5384 6130 5412
rect 6081 5381 6093 5384
rect 6035 5375 6093 5381
rect 6124 5372 6130 5384
rect 6182 5372 6188 5424
rect 7780 5412 7786 5424
rect 7741 5384 7786 5412
rect 7780 5372 7786 5384
rect 7838 5372 7844 5424
rect 3732 5276 3738 5288
rect 2830 5248 3738 5276
rect 3732 5236 3738 5248
rect 3790 5236 3796 5288
rect 38 5186 8870 5208
rect 38 5134 1394 5186
rect 1446 5134 1458 5186
rect 1510 5134 1522 5186
rect 1574 5134 1586 5186
rect 1638 5134 4352 5186
rect 4404 5134 4416 5186
rect 4468 5134 4480 5186
rect 4532 5134 4544 5186
rect 4596 5134 7309 5186
rect 7361 5134 7373 5186
rect 7425 5134 7437 5186
rect 7489 5134 7501 5186
rect 7553 5134 8870 5186
rect 38 5112 8870 5134
rect 3643 5075 3701 5081
rect 3643 5041 3655 5075
rect 3689 5072 3701 5075
rect 6492 5072 6498 5084
rect 3689 5044 6498 5072
rect 3689 5041 3701 5044
rect 3643 5035 3701 5041
rect 6492 5032 6498 5044
rect 6550 5032 6556 5084
rect 7872 5032 7878 5084
rect 7930 5072 7936 5084
rect 11368 5072 11374 5084
rect 7930 5044 11374 5072
rect 7930 5032 7936 5044
rect 11368 5032 11374 5044
rect 11426 5032 11432 5084
rect 3640 4936 3646 4948
rect 3474 4908 3646 4936
rect 3474 4877 3502 4908
rect 3640 4896 3646 4908
rect 3698 4896 3704 4948
rect 5572 4896 5578 4948
rect 5630 4936 5636 4948
rect 5667 4939 5725 4945
rect 5667 4936 5679 4939
rect 5630 4908 5679 4936
rect 5630 4896 5636 4908
rect 5667 4905 5679 4908
rect 5713 4905 5725 4939
rect 5940 4936 5946 4948
rect 5853 4908 5946 4936
rect 5667 4899 5725 4905
rect 5940 4896 5946 4908
rect 5998 4936 6004 4948
rect 6584 4936 6590 4948
rect 5998 4908 6590 4936
rect 5998 4896 6004 4908
rect 6584 4896 6590 4908
rect 6642 4896 6648 4948
rect 3459 4871 3517 4877
rect 3459 4837 3471 4871
rect 3505 4837 3517 4871
rect 3459 4831 3517 4837
rect 3548 4828 3554 4880
rect 3606 4868 3612 4880
rect 4563 4871 4621 4877
rect 4563 4868 4575 4871
rect 3606 4840 4575 4868
rect 3606 4828 3612 4840
rect 4563 4837 4575 4840
rect 4609 4837 4621 4871
rect 4563 4831 4621 4837
rect 4652 4760 4658 4812
rect 4710 4800 4716 4812
rect 7691 4803 7749 4809
rect 4710 4772 4882 4800
rect 4710 4760 4716 4772
rect 4744 4732 4750 4744
rect 4705 4704 4750 4732
rect 4744 4692 4750 4704
rect 4802 4692 4808 4744
rect 4854 4732 4882 4772
rect 6418 4732 6446 4786
rect 7691 4769 7703 4803
rect 7737 4800 7749 4803
rect 7737 4772 11414 4800
rect 7737 4769 7749 4772
rect 7691 4763 7749 4769
rect 11386 4744 11414 4772
rect 4854 4704 6446 4732
rect 11368 4692 11374 4744
rect 11426 4692 11432 4744
rect 38 4642 8870 4664
rect 38 4590 2873 4642
rect 2925 4590 2937 4642
rect 2989 4590 3001 4642
rect 3053 4590 3065 4642
rect 3117 4590 5830 4642
rect 5882 4590 5894 4642
rect 5946 4590 5958 4642
rect 6010 4590 6022 4642
rect 6074 4590 8870 4642
rect 38 4568 8870 4590
rect 3732 4528 3738 4540
rect 3693 4500 3738 4528
rect 3732 4488 3738 4500
rect 3790 4488 3796 4540
rect 6400 4528 6406 4540
rect 4670 4500 6406 4528
rect 788 4420 794 4472
rect 846 4460 852 4472
rect 846 4432 4606 4460
rect 846 4420 852 4432
rect 4578 4404 4606 4432
rect 3916 4392 3922 4404
rect 3877 4364 3922 4392
rect 3916 4352 3922 4364
rect 3974 4352 3980 4404
rect 4560 4392 4566 4404
rect 4473 4364 4566 4392
rect 4560 4352 4566 4364
rect 4618 4352 4624 4404
rect 4670 4256 4698 4500
rect 6400 4488 6406 4500
rect 6458 4488 6464 4540
rect 4744 4420 4750 4472
rect 4802 4460 4808 4472
rect 4802 4432 6524 4460
rect 4802 4420 4808 4432
rect 5759 4327 5817 4333
rect 5759 4293 5771 4327
rect 5805 4293 5817 4327
rect 5759 4287 5817 4293
rect 4747 4259 4805 4265
rect 4747 4256 4759 4259
rect 4670 4228 4759 4256
rect 4747 4225 4759 4228
rect 4793 4225 4805 4259
rect 4747 4219 4805 4225
rect 3732 4148 3738 4200
rect 3790 4188 3796 4200
rect 5664 4188 5670 4200
rect 3790 4160 5670 4188
rect 3790 4148 3796 4160
rect 5664 4148 5670 4160
rect 5722 4188 5728 4200
rect 5774 4188 5802 4287
rect 6124 4284 6130 4336
rect 6182 4324 6188 4336
rect 7783 4327 7841 4333
rect 7783 4324 7795 4327
rect 6182 4296 7795 4324
rect 6182 4284 6188 4296
rect 7783 4293 7795 4296
rect 7829 4293 7841 4327
rect 7783 4287 7841 4293
rect 5722 4160 5802 4188
rect 6022 4191 6080 4197
rect 5722 4148 5728 4160
rect 6022 4157 6034 4191
rect 6068 4188 6080 4191
rect 6216 4188 6222 4200
rect 6068 4160 6222 4188
rect 6068 4157 6080 4160
rect 6022 4151 6080 4157
rect 6216 4148 6222 4160
rect 6274 4148 6280 4200
rect 38 4098 8870 4120
rect 38 4046 1394 4098
rect 1446 4046 1458 4098
rect 1510 4046 1522 4098
rect 1574 4046 1586 4098
rect 1638 4046 4352 4098
rect 4404 4046 4416 4098
rect 4468 4046 4480 4098
rect 4532 4046 4544 4098
rect 4596 4046 7309 4098
rect 7361 4046 7373 4098
rect 7425 4046 7437 4098
rect 7489 4046 7501 4098
rect 7553 4046 8870 4098
rect 38 4024 8870 4046
rect 5930 3987 5988 3993
rect 5930 3953 5942 3987
rect 5976 3984 5988 3987
rect 6124 3984 6130 3996
rect 5976 3956 6130 3984
rect 5976 3953 5988 3956
rect 5930 3947 5988 3953
rect 6124 3944 6130 3956
rect 6182 3944 6188 3996
rect 5664 3848 5670 3860
rect 5625 3820 5670 3848
rect 5664 3808 5670 3820
rect 5722 3808 5728 3860
rect 7688 3848 7694 3860
rect 7649 3820 7694 3848
rect 7688 3808 7694 3820
rect 7746 3808 7752 3860
rect 4836 3672 4842 3724
rect 4894 3712 4900 3724
rect 4894 3684 6432 3712
rect 4894 3672 4900 3684
rect 38 3554 8870 3576
rect 38 3502 2873 3554
rect 2925 3502 2937 3554
rect 2989 3502 3001 3554
rect 3053 3502 3065 3554
rect 3117 3502 5830 3554
rect 5882 3502 5894 3554
rect 5946 3502 5958 3554
rect 6010 3502 6022 3554
rect 6074 3502 8870 3554
rect 38 3480 8870 3502
rect 6308 3440 6314 3452
rect 6269 3412 6314 3440
rect 6308 3400 6314 3412
rect 6366 3400 6372 3452
rect 1708 3264 1714 3316
rect 1766 3304 1772 3316
rect 6124 3304 6130 3316
rect 1766 3276 6130 3304
rect 1766 3264 1772 3276
rect 6124 3264 6130 3276
rect 6182 3264 6188 3316
rect 7323 3307 7381 3313
rect 7323 3273 7335 3307
rect 7369 3304 7381 3307
rect 8516 3304 8522 3316
rect 7369 3276 8522 3304
rect 7369 3273 7381 3276
rect 7323 3267 7381 3273
rect 8516 3264 8522 3276
rect 8574 3264 8580 3316
rect 7231 3239 7289 3245
rect 7231 3205 7243 3239
rect 7277 3236 7289 3239
rect 7964 3236 7970 3248
rect 7277 3208 7970 3236
rect 7277 3205 7289 3208
rect 7231 3199 7289 3205
rect 7964 3196 7970 3208
rect 8022 3196 8028 3248
rect 7507 3103 7565 3109
rect 7507 3069 7519 3103
rect 7553 3100 7565 3103
rect 15692 3100 15698 3112
rect 7553 3072 15698 3100
rect 7553 3069 7565 3072
rect 7507 3063 7565 3069
rect 15692 3060 15698 3072
rect 15750 3060 15756 3112
rect 38 3010 8870 3032
rect 38 2958 1394 3010
rect 1446 2958 1458 3010
rect 1510 2958 1522 3010
rect 1574 2958 1586 3010
rect 1638 2958 4352 3010
rect 4404 2958 4416 3010
rect 4468 2958 4480 3010
rect 4532 2958 4544 3010
rect 4596 2958 7309 3010
rect 7361 2958 7373 3010
rect 7425 2958 7437 3010
rect 7489 2958 7501 3010
rect 7553 2958 8870 3010
rect 38 2936 8870 2958
rect 7044 2856 7050 2908
rect 7102 2896 7108 2908
rect 7599 2899 7657 2905
rect 7599 2896 7611 2899
rect 7102 2868 7611 2896
rect 7102 2856 7108 2868
rect 7599 2865 7611 2868
rect 7645 2865 7657 2899
rect 7599 2859 7657 2865
rect 6124 2652 6130 2704
rect 6182 2692 6188 2704
rect 7415 2695 7473 2701
rect 7415 2692 7427 2695
rect 6182 2664 7427 2692
rect 6182 2652 6188 2664
rect 7415 2661 7427 2664
rect 7461 2661 7473 2695
rect 7415 2655 7473 2661
rect 38 2466 8870 2488
rect 38 2414 2873 2466
rect 2925 2414 2937 2466
rect 2989 2414 3001 2466
rect 3053 2414 3065 2466
rect 3117 2414 5830 2466
rect 5882 2414 5894 2466
rect 5946 2414 5958 2466
rect 6010 2414 6022 2466
rect 6074 2414 8870 2466
rect 38 2392 8870 2414
rect 5296 2312 5302 2364
rect 5354 2352 5360 2364
rect 15600 2352 15606 2364
rect 5354 2324 15606 2352
rect 5354 2312 5360 2324
rect 15600 2312 15606 2324
rect 15658 2312 15664 2364
rect 7780 2244 7786 2296
rect 7838 2284 7844 2296
rect 15508 2284 15514 2296
rect 7838 2256 15514 2284
rect 7838 2244 7844 2256
rect 15508 2244 15514 2256
rect 15566 2244 15572 2296
rect 4652 2176 4658 2228
rect 4710 2216 4716 2228
rect 7507 2219 7565 2225
rect 7507 2216 7519 2219
rect 4710 2188 7519 2216
rect 4710 2176 4716 2188
rect 7507 2185 7519 2188
rect 7553 2185 7565 2219
rect 7507 2179 7565 2185
rect 7596 2040 7602 2092
rect 7654 2080 7660 2092
rect 7691 2083 7749 2089
rect 7691 2080 7703 2083
rect 7654 2052 7703 2080
rect 7654 2040 7660 2052
rect 7691 2049 7703 2052
rect 7737 2049 7749 2083
rect 7691 2043 7749 2049
rect 38 1922 8870 1944
rect 38 1870 1394 1922
rect 1446 1870 1458 1922
rect 1510 1870 1522 1922
rect 1574 1870 1586 1922
rect 1638 1870 4352 1922
rect 4404 1870 4416 1922
rect 4468 1870 4480 1922
rect 4532 1870 4544 1922
rect 4596 1870 7309 1922
rect 7361 1870 7373 1922
rect 7425 1870 7437 1922
rect 7489 1870 7501 1922
rect 7553 1870 8870 1922
rect 38 1848 8870 1870
<< via1 >>
rect 7694 16320 7746 16372
rect 15514 16320 15566 16372
rect 1394 16014 1446 16066
rect 1458 16014 1510 16066
rect 1522 16014 1574 16066
rect 1586 16014 1638 16066
rect 4352 16014 4404 16066
rect 4416 16014 4468 16066
rect 4480 16014 4532 16066
rect 4544 16014 4596 16066
rect 7309 16014 7361 16066
rect 7373 16014 7425 16066
rect 7437 16014 7489 16066
rect 7501 16014 7553 16066
rect 7142 15615 7194 15624
rect 7142 15581 7151 15615
rect 7151 15581 7185 15615
rect 7185 15581 7194 15615
rect 7142 15572 7194 15581
rect 2873 15470 2925 15522
rect 2937 15470 2989 15522
rect 3001 15470 3053 15522
rect 3065 15470 3117 15522
rect 5830 15470 5882 15522
rect 5894 15470 5946 15522
rect 5958 15470 6010 15522
rect 6022 15470 6074 15522
rect 4842 15232 4894 15284
rect 7786 15028 7838 15080
rect 1394 14926 1446 14978
rect 1458 14926 1510 14978
rect 1522 14926 1574 14978
rect 1586 14926 1638 14978
rect 4352 14926 4404 14978
rect 4416 14926 4468 14978
rect 4480 14926 4532 14978
rect 4544 14926 4596 14978
rect 7309 14926 7361 14978
rect 7373 14926 7425 14978
rect 7437 14926 7489 14978
rect 7501 14926 7553 14978
rect 1714 14620 1766 14672
rect 1898 14552 1950 14604
rect 4750 14484 4802 14536
rect 7602 14527 7654 14536
rect 7602 14493 7611 14527
rect 7611 14493 7645 14527
rect 7645 14493 7654 14527
rect 7602 14484 7654 14493
rect 2873 14382 2925 14434
rect 2937 14382 2989 14434
rect 3001 14382 3053 14434
rect 3065 14382 3117 14434
rect 5830 14382 5882 14434
rect 5894 14382 5946 14434
rect 5958 14382 6010 14434
rect 6022 14382 6074 14434
rect 7142 14144 7194 14196
rect 6590 14076 6642 14128
rect 7694 14119 7746 14128
rect 7694 14085 7703 14119
rect 7703 14085 7737 14119
rect 7737 14085 7746 14119
rect 7694 14076 7746 14085
rect 1394 13838 1446 13890
rect 1458 13838 1510 13890
rect 1522 13838 1574 13890
rect 1586 13838 1638 13890
rect 4352 13838 4404 13890
rect 4416 13838 4468 13890
rect 4480 13838 4532 13890
rect 4544 13838 4596 13890
rect 7309 13838 7361 13890
rect 7373 13838 7425 13890
rect 7437 13838 7489 13890
rect 7501 13838 7553 13890
rect 3370 13668 3422 13720
rect 15514 13600 15566 13652
rect 4658 13575 4710 13584
rect 4658 13541 4667 13575
rect 4667 13541 4701 13575
rect 4701 13541 4710 13575
rect 4658 13532 4710 13541
rect 5670 13575 5722 13584
rect 5670 13541 5679 13575
rect 5679 13541 5713 13575
rect 5713 13541 5722 13575
rect 5670 13532 5722 13541
rect 7234 13532 7286 13584
rect 1806 13464 1858 13516
rect 6222 13464 6274 13516
rect 2873 13294 2925 13346
rect 2937 13294 2989 13346
rect 3001 13294 3053 13346
rect 3065 13294 3117 13346
rect 5830 13294 5882 13346
rect 5894 13294 5946 13346
rect 5958 13294 6010 13346
rect 6022 13294 6074 13346
rect 4842 13192 4894 13244
rect 6498 13124 6550 13176
rect 3830 13056 3882 13108
rect 4106 12988 4158 13040
rect 5670 12988 5722 13040
rect 6130 12988 6182 13040
rect 6406 12988 6458 13040
rect 2634 12852 2686 12904
rect 4198 12852 4250 12904
rect 1394 12750 1446 12802
rect 1458 12750 1510 12802
rect 1522 12750 1574 12802
rect 1586 12750 1638 12802
rect 4352 12750 4404 12802
rect 4416 12750 4468 12802
rect 4480 12750 4532 12802
rect 4544 12750 4596 12802
rect 7309 12750 7361 12802
rect 7373 12750 7425 12802
rect 7437 12750 7489 12802
rect 7501 12750 7553 12802
rect 2082 12444 2134 12496
rect 4842 12512 4894 12564
rect 6498 12512 6550 12564
rect 6682 12512 6734 12564
rect 4198 12444 4250 12496
rect 5670 12487 5722 12496
rect 5670 12453 5679 12487
rect 5679 12453 5713 12487
rect 5713 12453 5722 12487
rect 5670 12444 5722 12453
rect 4658 12376 4710 12428
rect 3646 12308 3698 12360
rect 4106 12308 4158 12360
rect 6314 12308 6366 12360
rect 2873 12206 2925 12258
rect 2937 12206 2989 12258
rect 3001 12206 3053 12258
rect 3065 12206 3117 12258
rect 5830 12206 5882 12258
rect 5894 12206 5946 12258
rect 5958 12206 6010 12258
rect 6022 12206 6074 12258
rect 7050 12104 7102 12156
rect 4750 12036 4802 12088
rect 5026 12036 5078 12088
rect 5670 11968 5722 12020
rect 2634 11900 2686 11952
rect 4842 11943 4894 11952
rect 4842 11909 4851 11943
rect 4851 11909 4885 11943
rect 4885 11909 4894 11943
rect 4842 11900 4894 11909
rect 7142 11832 7194 11884
rect 15698 11764 15750 11816
rect 1394 11662 1446 11714
rect 1458 11662 1510 11714
rect 1522 11662 1574 11714
rect 1586 11662 1638 11714
rect 4352 11662 4404 11714
rect 4416 11662 4468 11714
rect 4480 11662 4532 11714
rect 4544 11662 4596 11714
rect 7309 11662 7361 11714
rect 7373 11662 7425 11714
rect 7437 11662 7489 11714
rect 7501 11662 7553 11714
rect 3554 11424 3606 11476
rect 6590 11560 6642 11612
rect 4842 11424 4894 11476
rect 9258 11424 9310 11476
rect 610 11356 662 11408
rect 2082 11356 2134 11408
rect 702 11288 754 11340
rect 1990 11263 2042 11272
rect 1990 11229 1999 11263
rect 1999 11229 2033 11263
rect 2033 11229 2042 11263
rect 1990 11220 2042 11229
rect 3186 11263 3238 11272
rect 3186 11229 3195 11263
rect 3195 11229 3229 11263
rect 3229 11229 3238 11263
rect 3186 11220 3238 11229
rect 5578 11356 5630 11408
rect 4842 11288 4894 11340
rect 4934 11288 4986 11340
rect 7694 11331 7746 11340
rect 7694 11297 7703 11331
rect 7703 11297 7737 11331
rect 7737 11297 7746 11331
rect 7694 11288 7746 11297
rect 7878 11220 7930 11272
rect 2873 11118 2925 11170
rect 2937 11118 2989 11170
rect 3001 11118 3053 11170
rect 3065 11118 3117 11170
rect 5830 11118 5882 11170
rect 5894 11118 5946 11170
rect 5958 11118 6010 11170
rect 6022 11118 6074 11170
rect 794 11016 846 11068
rect 1898 11059 1950 11068
rect 1898 11025 1907 11059
rect 1907 11025 1941 11059
rect 1941 11025 1950 11059
rect 1898 11016 1950 11025
rect 1990 11016 2042 11068
rect 2726 10948 2778 11000
rect 6130 10948 6182 11000
rect 610 10923 662 10932
rect 610 10889 619 10923
rect 619 10889 653 10923
rect 653 10889 662 10923
rect 610 10880 662 10889
rect 1714 10923 1766 10932
rect 1714 10889 1723 10923
rect 1723 10889 1757 10923
rect 1757 10889 1766 10923
rect 1714 10880 1766 10889
rect 2634 10812 2686 10864
rect 4658 10812 4710 10864
rect 5578 10812 5630 10864
rect 15606 10812 15658 10864
rect 6682 10676 6734 10728
rect 1394 10574 1446 10626
rect 1458 10574 1510 10626
rect 1522 10574 1574 10626
rect 1586 10574 1638 10626
rect 4352 10574 4404 10626
rect 4416 10574 4468 10626
rect 4480 10574 4532 10626
rect 4544 10574 4596 10626
rect 7309 10574 7361 10626
rect 7373 10574 7425 10626
rect 7437 10574 7489 10626
rect 7501 10574 7553 10626
rect 2634 10336 2686 10388
rect 8614 10472 8666 10524
rect 794 10268 846 10320
rect 3370 10268 3422 10320
rect 3738 10311 3790 10320
rect 3738 10277 3747 10311
rect 3747 10277 3781 10311
rect 3781 10277 3790 10311
rect 3738 10268 3790 10277
rect 3830 10268 3882 10320
rect 2082 10243 2134 10252
rect 2082 10209 2091 10243
rect 2091 10209 2125 10243
rect 2125 10209 2134 10243
rect 2082 10200 2134 10209
rect 4934 10404 4986 10456
rect 4474 10311 4526 10320
rect 4474 10277 4483 10311
rect 4483 10277 4517 10311
rect 4517 10277 4526 10311
rect 4474 10268 4526 10277
rect 4842 10268 4894 10320
rect 5578 10311 5630 10320
rect 5578 10277 5587 10311
rect 5587 10277 5621 10311
rect 5621 10277 5630 10311
rect 5578 10268 5630 10277
rect 5670 10268 5722 10320
rect 7602 10200 7654 10252
rect 4474 10132 4526 10184
rect 8614 10132 8666 10184
rect 2873 10030 2925 10082
rect 2937 10030 2989 10082
rect 3001 10030 3053 10082
rect 3065 10030 3117 10082
rect 5830 10030 5882 10082
rect 5894 10030 5946 10082
rect 5958 10030 6010 10082
rect 6022 10030 6074 10082
rect 1714 9928 1766 9980
rect 4106 9928 4158 9980
rect 8706 9928 8758 9980
rect 23794 9928 23846 9980
rect 702 9792 754 9844
rect 3186 9860 3238 9912
rect 4658 9860 4710 9912
rect 2634 9792 2686 9844
rect 5578 9792 5630 9844
rect 4106 9724 4158 9776
rect 4750 9724 4802 9776
rect 5670 9724 5722 9776
rect 6682 9724 6734 9776
rect 11466 9724 11518 9776
rect 5026 9588 5078 9640
rect 1394 9486 1446 9538
rect 1458 9486 1510 9538
rect 1522 9486 1574 9538
rect 1586 9486 1638 9538
rect 4352 9486 4404 9538
rect 4416 9486 4468 9538
rect 4480 9486 4532 9538
rect 4544 9486 4596 9538
rect 7309 9486 7361 9538
rect 7373 9486 7425 9538
rect 7437 9486 7489 9538
rect 7501 9486 7553 9538
rect 4106 9384 4158 9436
rect 5946 9384 5998 9436
rect 7142 9384 7194 9436
rect 3922 9316 3974 9368
rect 518 9180 570 9232
rect 1806 9223 1858 9232
rect 1806 9189 1815 9223
rect 1815 9189 1849 9223
rect 1849 9189 1858 9223
rect 1806 9180 1858 9189
rect 15974 9248 16026 9300
rect 5578 9223 5630 9232
rect 5578 9189 5587 9223
rect 5587 9189 5621 9223
rect 5621 9189 5630 9223
rect 5578 9180 5630 9189
rect 5946 9223 5998 9232
rect 5946 9189 5955 9223
rect 5955 9189 5989 9223
rect 5989 9189 5998 9223
rect 5946 9180 5998 9189
rect 886 9087 938 9096
rect 886 9053 895 9087
rect 895 9053 929 9087
rect 929 9053 938 9087
rect 886 9044 938 9053
rect 7786 9112 7838 9164
rect 6406 9044 6458 9096
rect 7970 9044 8022 9096
rect 24070 9044 24122 9096
rect 2873 8942 2925 8994
rect 2937 8942 2989 8994
rect 3001 8942 3053 8994
rect 3065 8942 3117 8994
rect 5830 8942 5882 8994
rect 5894 8942 5946 8994
rect 5958 8942 6010 8994
rect 6022 8942 6074 8994
rect 1806 8840 1858 8892
rect 4658 8840 4710 8892
rect 886 8772 938 8824
rect 610 8747 662 8756
rect 610 8713 619 8747
rect 619 8713 653 8747
rect 653 8713 662 8747
rect 610 8704 662 8713
rect 1622 8704 1674 8756
rect 2542 8636 2594 8688
rect 4750 8704 4802 8756
rect 6498 8772 6550 8824
rect 7878 8772 7930 8824
rect 8522 8772 8574 8824
rect 11374 8772 11426 8824
rect 5578 8704 5630 8756
rect 8614 8704 8666 8756
rect 11650 8704 11702 8756
rect 4842 8679 4894 8688
rect 4842 8645 4851 8679
rect 4851 8645 4885 8679
rect 4885 8645 4894 8679
rect 4842 8636 4894 8645
rect 4106 8568 4158 8620
rect 11466 8636 11518 8688
rect 7970 8568 8022 8620
rect 518 8500 570 8552
rect 1990 8500 2042 8552
rect 2174 8500 2226 8552
rect 6406 8500 6458 8552
rect 1394 8398 1446 8450
rect 1458 8398 1510 8450
rect 1522 8398 1574 8450
rect 1586 8398 1638 8450
rect 4352 8398 4404 8450
rect 4416 8398 4468 8450
rect 4480 8398 4532 8450
rect 4544 8398 4596 8450
rect 7309 8398 7361 8450
rect 7373 8398 7425 8450
rect 7437 8398 7489 8450
rect 7501 8398 7553 8450
rect 2174 8296 2226 8348
rect 8338 8296 8390 8348
rect 8614 8296 8666 8348
rect 2634 8228 2686 8280
rect 3370 8228 3422 8280
rect 3738 8228 3790 8280
rect 4106 8228 4158 8280
rect 3278 8203 3330 8212
rect 3278 8169 3287 8203
rect 3287 8169 3321 8203
rect 3321 8169 3330 8203
rect 3278 8160 3330 8169
rect 518 8092 570 8144
rect 1806 8135 1858 8144
rect 1806 8101 1815 8135
rect 1815 8101 1849 8135
rect 1849 8101 1858 8135
rect 1806 8092 1858 8101
rect 3738 8135 3790 8144
rect 3738 8101 3747 8135
rect 3747 8101 3781 8135
rect 3781 8101 3790 8135
rect 3738 8092 3790 8101
rect 4014 8135 4066 8144
rect 4014 8101 4023 8135
rect 4023 8101 4057 8135
rect 4057 8101 4066 8135
rect 4014 8092 4066 8101
rect 4658 8203 4710 8212
rect 4658 8169 4667 8203
rect 4667 8169 4701 8203
rect 4701 8169 4710 8203
rect 4658 8160 4710 8169
rect 5578 8203 5630 8212
rect 5578 8169 5587 8203
rect 5587 8169 5621 8203
rect 5621 8169 5630 8203
rect 5578 8160 5630 8169
rect 6222 8160 6274 8212
rect 3370 8024 3422 8076
rect 4934 8092 4986 8144
rect 7602 8024 7654 8076
rect 7878 8024 7930 8076
rect 2873 7854 2925 7906
rect 2937 7854 2989 7906
rect 3001 7854 3053 7906
rect 3065 7854 3117 7906
rect 5830 7854 5882 7906
rect 5894 7854 5946 7906
rect 5958 7854 6010 7906
rect 6022 7854 6074 7906
rect 702 7752 754 7804
rect 4842 7752 4894 7804
rect 3370 7684 3422 7736
rect 610 7659 662 7668
rect 610 7625 619 7659
rect 619 7625 653 7659
rect 653 7625 662 7659
rect 610 7616 662 7625
rect 1806 7616 1858 7668
rect 2542 7616 2594 7668
rect 3646 7548 3698 7600
rect 4658 7548 4710 7600
rect 5578 7616 5630 7668
rect 11558 7548 11610 7600
rect 1898 7455 1950 7464
rect 1898 7421 1907 7455
rect 1907 7421 1941 7455
rect 1941 7421 1950 7455
rect 1898 7412 1950 7421
rect 3830 7412 3882 7464
rect 4106 7412 4158 7464
rect 1394 7310 1446 7362
rect 1458 7310 1510 7362
rect 1522 7310 1574 7362
rect 1586 7310 1638 7362
rect 4352 7310 4404 7362
rect 4416 7310 4468 7362
rect 4480 7310 4532 7362
rect 4544 7310 4596 7362
rect 7309 7310 7361 7362
rect 7373 7310 7425 7362
rect 7437 7310 7489 7362
rect 7501 7310 7553 7362
rect 2726 7251 2778 7260
rect 2726 7217 2735 7251
rect 2735 7217 2769 7251
rect 2769 7217 2778 7251
rect 2726 7208 2778 7217
rect 3554 7208 3606 7260
rect 4198 7208 4250 7260
rect 1806 7140 1858 7192
rect 4842 7140 4894 7192
rect 23794 7140 23846 7192
rect 794 7004 846 7056
rect 1990 7004 2042 7056
rect 3738 7072 3790 7124
rect 3554 7047 3606 7056
rect 3554 7013 3563 7047
rect 3563 7013 3597 7047
rect 3597 7013 3606 7047
rect 3554 7004 3606 7013
rect 7878 7072 7930 7124
rect 4106 7047 4158 7056
rect 4106 7013 4115 7047
rect 4115 7013 4149 7047
rect 4149 7013 4158 7047
rect 4106 7004 4158 7013
rect 3186 6936 3238 6988
rect 886 6911 938 6920
rect 886 6877 895 6911
rect 895 6877 929 6911
rect 929 6877 938 6911
rect 886 6868 938 6877
rect 5578 7004 5630 7056
rect 6222 6936 6274 6988
rect 6406 6936 6458 6988
rect 11374 6936 11426 6988
rect 6774 6868 6826 6920
rect 2873 6766 2925 6818
rect 2937 6766 2989 6818
rect 3001 6766 3053 6818
rect 3065 6766 3117 6818
rect 5830 6766 5882 6818
rect 5894 6766 5946 6818
rect 5958 6766 6010 6818
rect 6022 6766 6074 6818
rect 886 6664 938 6716
rect 702 6596 754 6648
rect 2634 6596 2686 6648
rect 1714 6571 1766 6580
rect 1714 6537 1723 6571
rect 1723 6537 1757 6571
rect 1757 6537 1766 6571
rect 1714 6528 1766 6537
rect 2542 6528 2594 6580
rect 5578 6528 5630 6580
rect 7694 6528 7746 6580
rect 11374 6528 11426 6580
rect 4658 6460 4710 6512
rect 4658 6324 4710 6376
rect 6682 6460 6734 6512
rect 6774 6460 6826 6512
rect 11466 6460 11518 6512
rect 6222 6324 6274 6376
rect 1394 6222 1446 6274
rect 1458 6222 1510 6274
rect 1522 6222 1574 6274
rect 1586 6222 1638 6274
rect 4352 6222 4404 6274
rect 4416 6222 4468 6274
rect 4480 6222 4532 6274
rect 4544 6222 4596 6274
rect 7309 6222 7361 6274
rect 7373 6222 7425 6274
rect 7437 6222 7489 6274
rect 7501 6222 7553 6274
rect 3186 6120 3238 6172
rect 3370 6163 3422 6172
rect 3370 6129 3379 6163
rect 3379 6129 3413 6163
rect 3413 6129 3422 6163
rect 3370 6120 3422 6129
rect 4014 6120 4066 6172
rect 7694 6120 7746 6172
rect 4934 5984 4986 6036
rect 7694 5984 7746 6036
rect 1990 5916 2042 5968
rect 3554 5916 3606 5968
rect 4198 5916 4250 5968
rect 5302 5916 5354 5968
rect 5578 5916 5630 5968
rect 7050 5916 7102 5968
rect 11558 5848 11610 5900
rect 2873 5678 2925 5730
rect 2937 5678 2989 5730
rect 3001 5678 3053 5730
rect 3065 5678 3117 5730
rect 5830 5678 5882 5730
rect 5894 5678 5946 5730
rect 5958 5678 6010 5730
rect 6022 5678 6074 5730
rect 1898 5508 1950 5560
rect 5946 5508 5998 5560
rect 6314 5508 6366 5560
rect 2542 5440 2594 5492
rect 4934 5440 4986 5492
rect 5578 5440 5630 5492
rect 6130 5372 6182 5424
rect 7786 5415 7838 5424
rect 7786 5381 7795 5415
rect 7795 5381 7829 5415
rect 7829 5381 7838 5415
rect 7786 5372 7838 5381
rect 3738 5236 3790 5288
rect 1394 5134 1446 5186
rect 1458 5134 1510 5186
rect 1522 5134 1574 5186
rect 1586 5134 1638 5186
rect 4352 5134 4404 5186
rect 4416 5134 4468 5186
rect 4480 5134 4532 5186
rect 4544 5134 4596 5186
rect 7309 5134 7361 5186
rect 7373 5134 7425 5186
rect 7437 5134 7489 5186
rect 7501 5134 7553 5186
rect 6498 5032 6550 5084
rect 7878 5032 7930 5084
rect 11374 5032 11426 5084
rect 3646 4896 3698 4948
rect 5578 4896 5630 4948
rect 5946 4939 5998 4948
rect 5946 4905 5955 4939
rect 5955 4905 5989 4939
rect 5989 4905 5998 4939
rect 5946 4896 5998 4905
rect 6590 4896 6642 4948
rect 3554 4828 3606 4880
rect 4658 4760 4710 4812
rect 4750 4735 4802 4744
rect 4750 4701 4759 4735
rect 4759 4701 4793 4735
rect 4793 4701 4802 4735
rect 4750 4692 4802 4701
rect 11374 4692 11426 4744
rect 2873 4590 2925 4642
rect 2937 4590 2989 4642
rect 3001 4590 3053 4642
rect 3065 4590 3117 4642
rect 5830 4590 5882 4642
rect 5894 4590 5946 4642
rect 5958 4590 6010 4642
rect 6022 4590 6074 4642
rect 3738 4531 3790 4540
rect 3738 4497 3747 4531
rect 3747 4497 3781 4531
rect 3781 4497 3790 4531
rect 3738 4488 3790 4497
rect 794 4420 846 4472
rect 3922 4395 3974 4404
rect 3922 4361 3931 4395
rect 3931 4361 3965 4395
rect 3965 4361 3974 4395
rect 3922 4352 3974 4361
rect 4566 4395 4618 4404
rect 4566 4361 4575 4395
rect 4575 4361 4609 4395
rect 4609 4361 4618 4395
rect 4566 4352 4618 4361
rect 6406 4488 6458 4540
rect 4750 4420 4802 4472
rect 3738 4148 3790 4200
rect 5670 4148 5722 4200
rect 6130 4284 6182 4336
rect 6222 4148 6274 4200
rect 1394 4046 1446 4098
rect 1458 4046 1510 4098
rect 1522 4046 1574 4098
rect 1586 4046 1638 4098
rect 4352 4046 4404 4098
rect 4416 4046 4468 4098
rect 4480 4046 4532 4098
rect 4544 4046 4596 4098
rect 7309 4046 7361 4098
rect 7373 4046 7425 4098
rect 7437 4046 7489 4098
rect 7501 4046 7553 4098
rect 6130 3944 6182 3996
rect 5670 3851 5722 3860
rect 5670 3817 5679 3851
rect 5679 3817 5713 3851
rect 5713 3817 5722 3851
rect 5670 3808 5722 3817
rect 7694 3851 7746 3860
rect 7694 3817 7703 3851
rect 7703 3817 7737 3851
rect 7737 3817 7746 3851
rect 7694 3808 7746 3817
rect 4842 3672 4894 3724
rect 2873 3502 2925 3554
rect 2937 3502 2989 3554
rect 3001 3502 3053 3554
rect 3065 3502 3117 3554
rect 5830 3502 5882 3554
rect 5894 3502 5946 3554
rect 5958 3502 6010 3554
rect 6022 3502 6074 3554
rect 6314 3443 6366 3452
rect 6314 3409 6323 3443
rect 6323 3409 6357 3443
rect 6357 3409 6366 3443
rect 6314 3400 6366 3409
rect 1714 3264 1766 3316
rect 6130 3307 6182 3316
rect 6130 3273 6139 3307
rect 6139 3273 6173 3307
rect 6173 3273 6182 3307
rect 6130 3264 6182 3273
rect 8522 3264 8574 3316
rect 7970 3196 8022 3248
rect 15698 3060 15750 3112
rect 1394 2958 1446 3010
rect 1458 2958 1510 3010
rect 1522 2958 1574 3010
rect 1586 2958 1638 3010
rect 4352 2958 4404 3010
rect 4416 2958 4468 3010
rect 4480 2958 4532 3010
rect 4544 2958 4596 3010
rect 7309 2958 7361 3010
rect 7373 2958 7425 3010
rect 7437 2958 7489 3010
rect 7501 2958 7553 3010
rect 7050 2856 7102 2908
rect 6130 2652 6182 2704
rect 2873 2414 2925 2466
rect 2937 2414 2989 2466
rect 3001 2414 3053 2466
rect 3065 2414 3117 2466
rect 5830 2414 5882 2466
rect 5894 2414 5946 2466
rect 5958 2414 6010 2466
rect 6022 2414 6074 2466
rect 5302 2312 5354 2364
rect 15606 2312 15658 2364
rect 7786 2244 7838 2296
rect 15514 2244 15566 2296
rect 4658 2176 4710 2228
rect 7602 2040 7654 2092
rect 1394 1870 1446 1922
rect 1458 1870 1510 1922
rect 1522 1870 1574 1922
rect 1586 1870 1638 1922
rect 4352 1870 4404 1922
rect 4416 1870 4468 1922
rect 4480 1870 4532 1922
rect 4544 1870 4596 1922
rect 7309 1870 7361 1922
rect 7373 1870 7425 1922
rect 7437 1870 7489 1922
rect 7501 1870 7553 1922
<< metal2 >>
rect 24068 18312 24124 18321
rect 24068 18247 24124 18256
rect 23792 17496 23848 17505
rect 23792 17431 23848 17440
rect 15512 16680 15568 16689
rect 15512 16615 15568 16624
rect 15526 16378 15554 16615
rect 7694 16372 7746 16378
rect 7694 16314 7746 16320
rect 15514 16372 15566 16378
rect 15514 16314 15566 16320
rect 1368 16068 1664 16088
rect 1424 16066 1448 16068
rect 1504 16066 1528 16068
rect 1584 16066 1608 16068
rect 1446 16014 1448 16066
rect 1510 16014 1522 16066
rect 1584 16014 1586 16066
rect 1424 16012 1448 16014
rect 1504 16012 1528 16014
rect 1584 16012 1608 16014
rect 1368 15992 1664 16012
rect 4326 16068 4622 16088
rect 4382 16066 4406 16068
rect 4462 16066 4486 16068
rect 4542 16066 4566 16068
rect 4404 16014 4406 16066
rect 4468 16014 4480 16066
rect 4542 16014 4544 16066
rect 4382 16012 4406 16014
rect 4462 16012 4486 16014
rect 4542 16012 4566 16014
rect 4326 15992 4622 16012
rect 7283 16068 7579 16088
rect 7339 16066 7363 16068
rect 7419 16066 7443 16068
rect 7499 16066 7523 16068
rect 7361 16014 7363 16066
rect 7425 16014 7437 16066
rect 7499 16014 7501 16066
rect 7339 16012 7363 16014
rect 7419 16012 7443 16014
rect 7499 16012 7523 16014
rect 7283 15992 7579 16012
rect 7142 15624 7194 15630
rect 7142 15566 7194 15572
rect 2847 15524 3143 15544
rect 2903 15522 2927 15524
rect 2983 15522 3007 15524
rect 3063 15522 3087 15524
rect 2925 15470 2927 15522
rect 2989 15470 3001 15522
rect 3063 15470 3065 15522
rect 2903 15468 2927 15470
rect 2983 15468 3007 15470
rect 3063 15468 3087 15470
rect 2847 15448 3143 15468
rect 5804 15524 6100 15544
rect 5860 15522 5884 15524
rect 5940 15522 5964 15524
rect 6020 15522 6044 15524
rect 5882 15470 5884 15522
rect 5946 15470 5958 15522
rect 6020 15470 6022 15522
rect 5860 15468 5884 15470
rect 5940 15468 5964 15470
rect 6020 15468 6044 15470
rect 5804 15448 6100 15468
rect 4842 15284 4894 15290
rect 4842 15226 4894 15232
rect 1368 14980 1664 15000
rect 1424 14978 1448 14980
rect 1504 14978 1528 14980
rect 1584 14978 1608 14980
rect 1446 14926 1448 14978
rect 1510 14926 1522 14978
rect 1584 14926 1586 14978
rect 1424 14924 1448 14926
rect 1504 14924 1528 14926
rect 1584 14924 1608 14926
rect 1368 14904 1664 14924
rect 4326 14980 4622 15000
rect 4382 14978 4406 14980
rect 4462 14978 4486 14980
rect 4542 14978 4566 14980
rect 4404 14926 4406 14978
rect 4468 14926 4480 14978
rect 4542 14926 4544 14978
rect 4382 14924 4406 14926
rect 4462 14924 4486 14926
rect 4542 14924 4566 14926
rect 4326 14904 4622 14924
rect 1714 14672 1766 14678
rect 1714 14614 1766 14620
rect 1368 13892 1664 13912
rect 1424 13890 1448 13892
rect 1504 13890 1528 13892
rect 1584 13890 1608 13892
rect 1446 13838 1448 13890
rect 1510 13838 1522 13890
rect 1584 13838 1586 13890
rect 1424 13836 1448 13838
rect 1504 13836 1528 13838
rect 1584 13836 1608 13838
rect 1368 13816 1664 13836
rect 1368 12804 1664 12824
rect 1424 12802 1448 12804
rect 1504 12802 1528 12804
rect 1584 12802 1608 12804
rect 1446 12750 1448 12802
rect 1510 12750 1522 12802
rect 1584 12750 1586 12802
rect 1424 12748 1448 12750
rect 1504 12748 1528 12750
rect 1584 12748 1608 12750
rect 1368 12728 1664 12748
rect 1368 11716 1664 11736
rect 1424 11714 1448 11716
rect 1504 11714 1528 11716
rect 1584 11714 1608 11716
rect 1446 11662 1448 11714
rect 1510 11662 1522 11714
rect 1584 11662 1586 11714
rect 1424 11660 1448 11662
rect 1504 11660 1528 11662
rect 1584 11660 1608 11662
rect 1368 11640 1664 11660
rect 610 11408 662 11414
rect 610 11350 662 11356
rect 622 10938 650 11350
rect 702 11340 754 11346
rect 702 11282 754 11288
rect 610 10932 662 10938
rect 610 10874 662 10880
rect 714 9850 742 11282
rect 794 11068 846 11074
rect 794 11010 846 11016
rect 806 10326 834 11010
rect 1726 10938 1754 14614
rect 1898 14604 1950 14610
rect 1898 14546 1950 14552
rect 1806 13516 1858 13522
rect 1806 13458 1858 13464
rect 1714 10932 1766 10938
rect 1714 10874 1766 10880
rect 1368 10628 1664 10648
rect 1424 10626 1448 10628
rect 1504 10626 1528 10628
rect 1584 10626 1608 10628
rect 1446 10574 1448 10626
rect 1510 10574 1522 10626
rect 1584 10574 1586 10626
rect 1424 10572 1448 10574
rect 1504 10572 1528 10574
rect 1584 10572 1608 10574
rect 1368 10552 1664 10572
rect 794 10320 846 10326
rect 794 10262 846 10268
rect 702 9844 754 9850
rect 702 9786 754 9792
rect 518 9232 570 9238
rect 518 9174 570 9180
rect 530 8558 558 9174
rect 610 8756 662 8762
rect 610 8698 662 8704
rect 518 8552 570 8558
rect 518 8494 570 8500
rect 530 8150 558 8494
rect 518 8144 570 8150
rect 518 8086 570 8092
rect 622 7674 650 8698
rect 714 7810 742 9786
rect 702 7804 754 7810
rect 702 7746 754 7752
rect 610 7668 662 7674
rect 610 7610 662 7616
rect 714 6654 742 7746
rect 806 7062 834 10262
rect 1726 9986 1754 10874
rect 1714 9980 1766 9986
rect 1714 9922 1766 9928
rect 1368 9540 1664 9560
rect 1424 9538 1448 9540
rect 1504 9538 1528 9540
rect 1584 9538 1608 9540
rect 1446 9486 1448 9538
rect 1510 9486 1522 9538
rect 1584 9486 1586 9538
rect 1424 9484 1448 9486
rect 1504 9484 1528 9486
rect 1584 9484 1608 9486
rect 1368 9464 1664 9484
rect 1726 9322 1754 9922
rect 1634 9294 1754 9322
rect 886 9096 938 9102
rect 886 9038 938 9044
rect 898 8830 926 9038
rect 886 8824 938 8830
rect 886 8766 938 8772
rect 1634 8762 1662 9294
rect 1818 9238 1846 13458
rect 1910 11074 1938 14546
rect 4750 14536 4802 14542
rect 4750 14478 4802 14484
rect 2847 14436 3143 14456
rect 2903 14434 2927 14436
rect 2983 14434 3007 14436
rect 3063 14434 3087 14436
rect 2925 14382 2927 14434
rect 2989 14382 3001 14434
rect 3063 14382 3065 14434
rect 2903 14380 2927 14382
rect 2983 14380 3007 14382
rect 3063 14380 3087 14382
rect 2847 14360 3143 14380
rect 4326 13892 4622 13912
rect 4382 13890 4406 13892
rect 4462 13890 4486 13892
rect 4542 13890 4566 13892
rect 4404 13838 4406 13890
rect 4468 13838 4480 13890
rect 4542 13838 4544 13890
rect 4382 13836 4406 13838
rect 4462 13836 4486 13838
rect 4542 13836 4566 13838
rect 4326 13816 4622 13836
rect 3370 13720 3422 13726
rect 3370 13662 3422 13668
rect 2847 13348 3143 13368
rect 2903 13346 2927 13348
rect 2983 13346 3007 13348
rect 3063 13346 3087 13348
rect 2925 13294 2927 13346
rect 2989 13294 3001 13346
rect 3063 13294 3065 13346
rect 2903 13292 2927 13294
rect 2983 13292 3007 13294
rect 3063 13292 3087 13294
rect 2847 13272 3143 13292
rect 2634 12904 2686 12910
rect 2634 12846 2686 12852
rect 2082 12496 2134 12502
rect 2082 12438 2134 12444
rect 2094 11414 2122 12438
rect 2646 11958 2674 12846
rect 2847 12260 3143 12280
rect 2903 12258 2927 12260
rect 2983 12258 3007 12260
rect 3063 12258 3087 12260
rect 2925 12206 2927 12258
rect 2989 12206 3001 12258
rect 3063 12206 3065 12258
rect 2903 12204 2927 12206
rect 2983 12204 3007 12206
rect 3063 12204 3087 12206
rect 2847 12184 3143 12204
rect 2634 11952 2686 11958
rect 2634 11894 2686 11900
rect 2082 11408 2134 11414
rect 2082 11350 2134 11356
rect 1990 11272 2042 11278
rect 1990 11214 2042 11220
rect 2002 11074 2030 11214
rect 1898 11068 1950 11074
rect 1898 11010 1950 11016
rect 1990 11068 2042 11074
rect 1990 11010 2042 11016
rect 2646 10870 2674 11894
rect 3186 11272 3238 11278
rect 3186 11214 3238 11220
rect 2847 11172 3143 11192
rect 2903 11170 2927 11172
rect 2983 11170 3007 11172
rect 3063 11170 3087 11172
rect 2925 11118 2927 11170
rect 2989 11118 3001 11170
rect 3063 11118 3065 11170
rect 2903 11116 2927 11118
rect 2983 11116 3007 11118
rect 3063 11116 3087 11118
rect 2847 11096 3143 11116
rect 2726 11000 2778 11006
rect 2726 10942 2778 10948
rect 2634 10864 2686 10870
rect 2634 10806 2686 10812
rect 2646 10394 2674 10806
rect 2634 10388 2686 10394
rect 2634 10330 2686 10336
rect 2080 10288 2136 10297
rect 2080 10223 2082 10232
rect 2134 10223 2136 10232
rect 2082 10194 2134 10200
rect 2646 9850 2674 10330
rect 2634 9844 2686 9850
rect 2634 9786 2686 9792
rect 1806 9232 1858 9238
rect 1806 9174 1858 9180
rect 1818 8898 1846 9174
rect 1806 8892 1858 8898
rect 1806 8834 1858 8840
rect 1622 8756 1674 8762
rect 1622 8698 1674 8704
rect 1368 8452 1664 8472
rect 1424 8450 1448 8452
rect 1504 8450 1528 8452
rect 1584 8450 1608 8452
rect 1446 8398 1448 8450
rect 1510 8398 1522 8450
rect 1584 8398 1586 8450
rect 1424 8396 1448 8398
rect 1504 8396 1528 8398
rect 1584 8396 1608 8398
rect 1368 8376 1664 8396
rect 1818 8150 1846 8834
rect 2542 8688 2594 8694
rect 2542 8630 2594 8636
rect 1990 8552 2042 8558
rect 1990 8494 2042 8500
rect 2174 8552 2226 8558
rect 2174 8494 2226 8500
rect 1806 8144 1858 8150
rect 1806 8086 1858 8092
rect 1818 7674 1846 8086
rect 1806 7668 1858 7674
rect 1806 7610 1858 7616
rect 1368 7364 1664 7384
rect 1424 7362 1448 7364
rect 1504 7362 1528 7364
rect 1584 7362 1608 7364
rect 1446 7310 1448 7362
rect 1510 7310 1522 7362
rect 1584 7310 1586 7362
rect 1424 7308 1448 7310
rect 1504 7308 1528 7310
rect 1584 7308 1608 7310
rect 1368 7288 1664 7308
rect 1818 7198 1846 7610
rect 1898 7464 1950 7470
rect 1898 7406 1950 7412
rect 1806 7192 1858 7198
rect 1806 7134 1858 7140
rect 794 7056 846 7062
rect 794 6998 846 7004
rect 702 6648 754 6654
rect 702 6590 754 6596
rect 806 4478 834 6998
rect 886 6920 938 6926
rect 886 6862 938 6868
rect 898 6722 926 6862
rect 886 6716 938 6722
rect 886 6658 938 6664
rect 1714 6580 1766 6586
rect 1714 6522 1766 6528
rect 1368 6276 1664 6296
rect 1424 6274 1448 6276
rect 1504 6274 1528 6276
rect 1584 6274 1608 6276
rect 1446 6222 1448 6274
rect 1510 6222 1522 6274
rect 1584 6222 1586 6274
rect 1424 6220 1448 6222
rect 1504 6220 1528 6222
rect 1584 6220 1608 6222
rect 1368 6200 1664 6220
rect 1368 5188 1664 5208
rect 1424 5186 1448 5188
rect 1504 5186 1528 5188
rect 1584 5186 1608 5188
rect 1446 5134 1448 5186
rect 1510 5134 1522 5186
rect 1584 5134 1586 5186
rect 1424 5132 1448 5134
rect 1504 5132 1528 5134
rect 1584 5132 1608 5134
rect 1368 5112 1664 5132
rect 794 4472 846 4478
rect 794 4414 846 4420
rect 1368 4100 1664 4120
rect 1424 4098 1448 4100
rect 1504 4098 1528 4100
rect 1584 4098 1608 4100
rect 1446 4046 1448 4098
rect 1510 4046 1522 4098
rect 1584 4046 1586 4098
rect 1424 4044 1448 4046
rect 1504 4044 1528 4046
rect 1584 4044 1608 4046
rect 1368 4024 1664 4044
rect 1726 3322 1754 6522
rect 1910 5566 1938 7406
rect 2002 7062 2030 8494
rect 2186 8354 2214 8494
rect 2174 8348 2226 8354
rect 2174 8290 2226 8296
rect 2554 7674 2582 8630
rect 2634 8280 2686 8286
rect 2634 8222 2686 8228
rect 2542 7668 2594 7674
rect 2542 7610 2594 7616
rect 1990 7056 2042 7062
rect 1990 6998 2042 7004
rect 2002 5974 2030 6998
rect 2554 6586 2582 7610
rect 2646 6654 2674 8222
rect 2738 7266 2766 10942
rect 2847 10084 3143 10104
rect 2903 10082 2927 10084
rect 2983 10082 3007 10084
rect 3063 10082 3087 10084
rect 2925 10030 2927 10082
rect 2989 10030 3001 10082
rect 3063 10030 3065 10082
rect 2903 10028 2927 10030
rect 2983 10028 3007 10030
rect 3063 10028 3087 10030
rect 2847 10008 3143 10028
rect 3198 9918 3226 11214
rect 3382 10326 3410 13662
rect 4658 13584 4710 13590
rect 4658 13526 4710 13532
rect 3830 13108 3882 13114
rect 3830 13050 3882 13056
rect 3646 12360 3698 12366
rect 3646 12302 3698 12308
rect 3554 11476 3606 11482
rect 3554 11418 3606 11424
rect 3370 10320 3422 10326
rect 3370 10262 3422 10268
rect 3186 9912 3238 9918
rect 3186 9854 3238 9860
rect 2847 8996 3143 9016
rect 2903 8994 2927 8996
rect 2983 8994 3007 8996
rect 3063 8994 3087 8996
rect 2925 8942 2927 8994
rect 2989 8942 3001 8994
rect 3063 8942 3065 8994
rect 2903 8940 2927 8942
rect 2983 8940 3007 8942
rect 3063 8940 3087 8942
rect 2847 8920 3143 8940
rect 3370 8280 3422 8286
rect 3276 8248 3332 8257
rect 3370 8222 3422 8228
rect 3276 8183 3278 8192
rect 3330 8183 3332 8192
rect 3278 8154 3330 8160
rect 3382 8082 3410 8222
rect 3370 8076 3422 8082
rect 3370 8018 3422 8024
rect 2847 7908 3143 7928
rect 2903 7906 2927 7908
rect 2983 7906 3007 7908
rect 3063 7906 3087 7908
rect 2925 7854 2927 7906
rect 2989 7854 3001 7906
rect 3063 7854 3065 7906
rect 2903 7852 2927 7854
rect 2983 7852 3007 7854
rect 3063 7852 3087 7854
rect 2847 7832 3143 7852
rect 3370 7736 3422 7742
rect 3370 7678 3422 7684
rect 2726 7260 2778 7266
rect 2726 7202 2778 7208
rect 3186 6988 3238 6994
rect 3186 6930 3238 6936
rect 2847 6820 3143 6840
rect 2903 6818 2927 6820
rect 2983 6818 3007 6820
rect 3063 6818 3087 6820
rect 2925 6766 2927 6818
rect 2989 6766 3001 6818
rect 3063 6766 3065 6818
rect 2903 6764 2927 6766
rect 2983 6764 3007 6766
rect 3063 6764 3087 6766
rect 2847 6744 3143 6764
rect 2634 6648 2686 6654
rect 2634 6590 2686 6596
rect 2542 6580 2594 6586
rect 2542 6522 2594 6528
rect 1990 5968 2042 5974
rect 1990 5910 2042 5916
rect 1898 5560 1950 5566
rect 1898 5502 1950 5508
rect 2554 5498 2582 6522
rect 3198 6178 3226 6930
rect 3382 6178 3410 7678
rect 3566 7452 3594 11418
rect 3658 7606 3686 12302
rect 3842 11260 3870 13050
rect 4106 13040 4158 13046
rect 4106 12982 4158 12988
rect 4118 12366 4146 12982
rect 4198 12904 4250 12910
rect 4198 12846 4250 12852
rect 4210 12502 4238 12846
rect 4326 12804 4622 12824
rect 4382 12802 4406 12804
rect 4462 12802 4486 12804
rect 4542 12802 4566 12804
rect 4404 12750 4406 12802
rect 4468 12750 4480 12802
rect 4542 12750 4544 12802
rect 4382 12748 4406 12750
rect 4462 12748 4486 12750
rect 4542 12748 4566 12750
rect 4326 12728 4622 12748
rect 4198 12496 4250 12502
rect 4198 12438 4250 12444
rect 4670 12434 4698 13526
rect 4658 12428 4710 12434
rect 4658 12370 4710 12376
rect 4106 12360 4158 12366
rect 4106 12302 4158 12308
rect 3842 11232 3962 11260
rect 3738 10320 3790 10326
rect 3738 10262 3790 10268
rect 3830 10320 3882 10326
rect 3830 10262 3882 10268
rect 3750 8286 3778 10262
rect 3738 8280 3790 8286
rect 3738 8222 3790 8228
rect 3738 8144 3790 8150
rect 3738 8086 3790 8092
rect 3646 7600 3698 7606
rect 3646 7542 3698 7548
rect 3566 7424 3686 7452
rect 3554 7260 3606 7266
rect 3554 7202 3606 7208
rect 3566 7062 3594 7202
rect 3554 7056 3606 7062
rect 3554 6998 3606 7004
rect 3186 6172 3238 6178
rect 3186 6114 3238 6120
rect 3370 6172 3422 6178
rect 3370 6114 3422 6120
rect 3554 5968 3606 5974
rect 3554 5910 3606 5916
rect 2847 5732 3143 5752
rect 2903 5730 2927 5732
rect 2983 5730 3007 5732
rect 3063 5730 3087 5732
rect 2925 5678 2927 5730
rect 2989 5678 3001 5730
rect 3063 5678 3065 5730
rect 2903 5676 2927 5678
rect 2983 5676 3007 5678
rect 3063 5676 3087 5678
rect 2847 5656 3143 5676
rect 2542 5492 2594 5498
rect 2542 5434 2594 5440
rect 3566 4886 3594 5910
rect 3658 4954 3686 7424
rect 3750 7130 3778 8086
rect 3842 7470 3870 10262
rect 3934 9374 3962 11232
rect 4118 9986 4146 12302
rect 4762 12094 4790 14478
rect 4854 13250 4882 15226
rect 5804 14436 6100 14456
rect 5860 14434 5884 14436
rect 5940 14434 5964 14436
rect 6020 14434 6044 14436
rect 5882 14382 5884 14434
rect 5946 14382 5958 14434
rect 6020 14382 6022 14434
rect 5860 14380 5884 14382
rect 5940 14380 5964 14382
rect 6020 14380 6044 14382
rect 5804 14360 6100 14380
rect 7154 14202 7182 15566
rect 7283 14980 7579 15000
rect 7339 14978 7363 14980
rect 7419 14978 7443 14980
rect 7499 14978 7523 14980
rect 7361 14926 7363 14978
rect 7425 14926 7437 14978
rect 7499 14926 7501 14978
rect 7339 14924 7363 14926
rect 7419 14924 7443 14926
rect 7499 14924 7523 14926
rect 7283 14904 7579 14924
rect 7602 14536 7654 14542
rect 7602 14478 7654 14484
rect 7142 14196 7194 14202
rect 7142 14138 7194 14144
rect 6590 14128 6642 14134
rect 6590 14070 6642 14076
rect 5670 13584 5722 13590
rect 5670 13526 5722 13532
rect 4842 13244 4894 13250
rect 4842 13186 4894 13192
rect 4854 12570 4882 13186
rect 5682 13046 5710 13526
rect 6222 13516 6274 13522
rect 6222 13458 6274 13464
rect 5804 13348 6100 13368
rect 5860 13346 5884 13348
rect 5940 13346 5964 13348
rect 6020 13346 6044 13348
rect 5882 13294 5884 13346
rect 5946 13294 5958 13346
rect 6020 13294 6022 13346
rect 5860 13292 5884 13294
rect 5940 13292 5964 13294
rect 6020 13292 6044 13294
rect 5804 13272 6100 13292
rect 5670 13040 5722 13046
rect 5670 12982 5722 12988
rect 6130 13040 6182 13046
rect 6130 12982 6182 12988
rect 6234 13028 6262 13458
rect 6498 13176 6550 13182
rect 6498 13118 6550 13124
rect 6406 13040 6458 13046
rect 6234 13000 6406 13028
rect 4842 12564 4894 12570
rect 4842 12506 4894 12512
rect 5682 12502 5710 12982
rect 5670 12496 5722 12502
rect 5670 12438 5722 12444
rect 4750 12088 4802 12094
rect 4750 12030 4802 12036
rect 5026 12088 5078 12094
rect 5026 12030 5078 12036
rect 4842 11952 4894 11958
rect 4842 11894 4894 11900
rect 4326 11716 4622 11736
rect 4382 11714 4406 11716
rect 4462 11714 4486 11716
rect 4542 11714 4566 11716
rect 4404 11662 4406 11714
rect 4468 11662 4480 11714
rect 4542 11662 4544 11714
rect 4382 11660 4406 11662
rect 4462 11660 4486 11662
rect 4542 11660 4566 11662
rect 4326 11640 4622 11660
rect 4854 11482 4882 11894
rect 4842 11476 4894 11482
rect 4842 11418 4894 11424
rect 4842 11340 4894 11346
rect 4842 11282 4894 11288
rect 4934 11340 4986 11346
rect 4934 11282 4986 11288
rect 4658 10864 4710 10870
rect 4658 10806 4710 10812
rect 4326 10628 4622 10648
rect 4382 10626 4406 10628
rect 4462 10626 4486 10628
rect 4542 10626 4566 10628
rect 4404 10574 4406 10626
rect 4468 10574 4480 10626
rect 4542 10574 4544 10626
rect 4382 10572 4406 10574
rect 4462 10572 4486 10574
rect 4542 10572 4566 10574
rect 4326 10552 4622 10572
rect 4474 10320 4526 10326
rect 4474 10262 4526 10268
rect 4486 10190 4514 10262
rect 4474 10184 4526 10190
rect 4474 10126 4526 10132
rect 4106 9980 4158 9986
rect 4106 9922 4158 9928
rect 4670 9918 4698 10806
rect 4854 10326 4882 11282
rect 4946 10462 4974 11282
rect 4934 10456 4986 10462
rect 4934 10398 4986 10404
rect 4842 10320 4894 10326
rect 4842 10262 4894 10268
rect 4658 9912 4710 9918
rect 4658 9854 4710 9860
rect 4106 9776 4158 9782
rect 4106 9718 4158 9724
rect 4750 9776 4802 9782
rect 4750 9718 4802 9724
rect 4118 9442 4146 9718
rect 4326 9540 4622 9560
rect 4382 9538 4406 9540
rect 4462 9538 4486 9540
rect 4542 9538 4566 9540
rect 4404 9486 4406 9538
rect 4468 9486 4480 9538
rect 4542 9486 4544 9538
rect 4382 9484 4406 9486
rect 4462 9484 4486 9486
rect 4542 9484 4566 9486
rect 4326 9464 4622 9484
rect 4106 9436 4158 9442
rect 4106 9378 4158 9384
rect 3922 9368 3974 9374
rect 3922 9310 3974 9316
rect 3830 7464 3882 7470
rect 3830 7406 3882 7412
rect 3738 7124 3790 7130
rect 3738 7066 3790 7072
rect 3738 5288 3790 5294
rect 3738 5230 3790 5236
rect 3646 4948 3698 4954
rect 3646 4890 3698 4896
rect 3554 4880 3606 4886
rect 3554 4822 3606 4828
rect 2847 4644 3143 4664
rect 2903 4642 2927 4644
rect 2983 4642 3007 4644
rect 3063 4642 3087 4644
rect 2925 4590 2927 4642
rect 2989 4590 3001 4642
rect 3063 4590 3065 4642
rect 2903 4588 2927 4590
rect 2983 4588 3007 4590
rect 3063 4588 3087 4590
rect 2847 4568 3143 4588
rect 3750 4546 3778 5230
rect 3738 4540 3790 4546
rect 3738 4482 3790 4488
rect 3750 4206 3778 4482
rect 3934 4410 3962 9310
rect 4658 8892 4710 8898
rect 4658 8834 4710 8840
rect 4106 8620 4158 8626
rect 4106 8562 4158 8568
rect 4118 8286 4146 8562
rect 4326 8452 4622 8472
rect 4382 8450 4406 8452
rect 4462 8450 4486 8452
rect 4542 8450 4566 8452
rect 4404 8398 4406 8450
rect 4468 8398 4480 8450
rect 4542 8398 4544 8450
rect 4382 8396 4406 8398
rect 4462 8396 4486 8398
rect 4542 8396 4566 8398
rect 4326 8376 4622 8396
rect 4106 8280 4158 8286
rect 4106 8222 4158 8228
rect 4670 8218 4698 8834
rect 4762 8762 4790 9718
rect 4854 8778 4882 10262
rect 5038 9646 5066 12030
rect 5682 12026 5710 12438
rect 5804 12260 6100 12280
rect 5860 12258 5884 12260
rect 5940 12258 5964 12260
rect 6020 12258 6044 12260
rect 5882 12206 5884 12258
rect 5946 12206 5958 12258
rect 6020 12206 6022 12258
rect 5860 12204 5884 12206
rect 5940 12204 5964 12206
rect 6020 12204 6044 12206
rect 5804 12184 6100 12204
rect 5670 12020 5722 12026
rect 5670 11962 5722 11968
rect 5578 11408 5630 11414
rect 5578 11350 5630 11356
rect 5590 10870 5618 11350
rect 5804 11172 6100 11192
rect 5860 11170 5884 11172
rect 5940 11170 5964 11172
rect 6020 11170 6044 11172
rect 5882 11118 5884 11170
rect 5946 11118 5958 11170
rect 6020 11118 6022 11170
rect 5860 11116 5884 11118
rect 5940 11116 5964 11118
rect 6020 11116 6044 11118
rect 5804 11096 6100 11116
rect 6142 11006 6170 12982
rect 6130 11000 6182 11006
rect 6130 10942 6182 10948
rect 5578 10864 5630 10870
rect 5578 10806 5630 10812
rect 5590 10326 5618 10806
rect 5578 10320 5630 10326
rect 5576 10288 5578 10297
rect 5670 10320 5722 10326
rect 5630 10288 5632 10297
rect 5670 10262 5722 10268
rect 5576 10223 5632 10232
rect 5590 9850 5618 10223
rect 5578 9844 5630 9850
rect 5578 9786 5630 9792
rect 5026 9640 5078 9646
rect 5026 9582 5078 9588
rect 5590 9238 5618 9786
rect 5682 9782 5710 10262
rect 5804 10084 6100 10104
rect 5860 10082 5884 10084
rect 5940 10082 5964 10084
rect 6020 10082 6044 10084
rect 5882 10030 5884 10082
rect 5946 10030 5958 10082
rect 6020 10030 6022 10082
rect 5860 10028 5884 10030
rect 5940 10028 5964 10030
rect 6020 10028 6044 10030
rect 5804 10008 6100 10028
rect 5670 9776 5722 9782
rect 5670 9718 5722 9724
rect 5946 9436 5998 9442
rect 5946 9378 5998 9384
rect 5958 9238 5986 9378
rect 5578 9232 5630 9238
rect 5578 9174 5630 9180
rect 5946 9232 5998 9238
rect 5946 9174 5998 9180
rect 4750 8756 4802 8762
rect 4854 8750 4974 8778
rect 5590 8762 5618 9174
rect 5804 8996 6100 9016
rect 5860 8994 5884 8996
rect 5940 8994 5964 8996
rect 6020 8994 6044 8996
rect 5882 8942 5884 8994
rect 5946 8942 5958 8994
rect 6020 8942 6022 8994
rect 5860 8940 5884 8942
rect 5940 8940 5964 8942
rect 6020 8940 6044 8942
rect 5804 8920 6100 8940
rect 4750 8698 4802 8704
rect 4842 8688 4894 8694
rect 4842 8630 4894 8636
rect 4658 8212 4710 8218
rect 4658 8154 4710 8160
rect 4014 8144 4066 8150
rect 4014 8086 4066 8092
rect 4026 6178 4054 8086
rect 4854 7810 4882 8630
rect 4946 8150 4974 8750
rect 5578 8756 5630 8762
rect 5578 8698 5630 8704
rect 5590 8218 5618 8698
rect 6234 8218 6262 13000
rect 6406 12982 6458 12988
rect 6510 12722 6538 13118
rect 6418 12694 6538 12722
rect 6314 12360 6366 12366
rect 6314 12302 6366 12308
rect 6326 8540 6354 12302
rect 6418 9102 6446 12694
rect 6498 12564 6550 12570
rect 6498 12506 6550 12512
rect 6406 9096 6458 9102
rect 6406 9038 6458 9044
rect 6510 8914 6538 12506
rect 6602 11618 6630 14070
rect 7283 13892 7579 13912
rect 7339 13890 7363 13892
rect 7419 13890 7443 13892
rect 7499 13890 7523 13892
rect 7361 13838 7363 13890
rect 7425 13838 7437 13890
rect 7499 13838 7501 13890
rect 7339 13836 7363 13838
rect 7419 13836 7443 13838
rect 7499 13836 7523 13838
rect 7283 13816 7579 13836
rect 7234 13584 7286 13590
rect 7062 13544 7234 13572
rect 6682 12564 6734 12570
rect 6682 12506 6734 12512
rect 6590 11612 6642 11618
rect 6590 11554 6642 11560
rect 6694 10734 6722 12506
rect 7062 12162 7090 13544
rect 7234 13526 7286 13532
rect 7283 12804 7579 12824
rect 7339 12802 7363 12804
rect 7419 12802 7443 12804
rect 7499 12802 7523 12804
rect 7361 12750 7363 12802
rect 7425 12750 7437 12802
rect 7499 12750 7501 12802
rect 7339 12748 7363 12750
rect 7419 12748 7443 12750
rect 7499 12748 7523 12750
rect 7283 12728 7579 12748
rect 7050 12156 7102 12162
rect 7050 12098 7102 12104
rect 6682 10728 6734 10734
rect 6682 10670 6734 10676
rect 6694 9782 6722 10670
rect 6682 9776 6734 9782
rect 6682 9718 6734 9724
rect 7062 9594 7090 12098
rect 7142 11884 7194 11890
rect 7142 11826 7194 11832
rect 6694 9566 7090 9594
rect 6510 8886 6630 8914
rect 6498 8824 6550 8830
rect 6498 8766 6550 8772
rect 6406 8552 6458 8558
rect 6326 8512 6406 8540
rect 6406 8494 6458 8500
rect 5578 8212 5630 8218
rect 5578 8154 5630 8160
rect 6222 8212 6274 8218
rect 6222 8154 6274 8160
rect 4934 8144 4986 8150
rect 4934 8086 4986 8092
rect 4842 7804 4894 7810
rect 4842 7746 4894 7752
rect 5590 7674 5618 8154
rect 5804 7908 6100 7928
rect 5860 7906 5884 7908
rect 5940 7906 5964 7908
rect 6020 7906 6044 7908
rect 5882 7854 5884 7906
rect 5946 7854 5958 7906
rect 6020 7854 6022 7906
rect 5860 7852 5884 7854
rect 5940 7852 5964 7854
rect 6020 7852 6044 7854
rect 5804 7832 6100 7852
rect 5578 7668 5630 7674
rect 5578 7610 5630 7616
rect 4658 7600 4710 7606
rect 4658 7542 4710 7548
rect 4106 7464 4158 7470
rect 4106 7406 4158 7412
rect 4118 7062 4146 7406
rect 4326 7364 4622 7384
rect 4382 7362 4406 7364
rect 4462 7362 4486 7364
rect 4542 7362 4566 7364
rect 4404 7310 4406 7362
rect 4468 7310 4480 7362
rect 4542 7310 4544 7362
rect 4382 7308 4406 7310
rect 4462 7308 4486 7310
rect 4542 7308 4566 7310
rect 4326 7288 4622 7308
rect 4198 7260 4250 7266
rect 4198 7202 4250 7208
rect 4106 7056 4158 7062
rect 4106 6998 4158 7004
rect 4014 6172 4066 6178
rect 4014 6114 4066 6120
rect 4210 5974 4238 7202
rect 4670 6518 4698 7542
rect 4842 7192 4894 7198
rect 4842 7134 4894 7140
rect 4658 6512 4710 6518
rect 4658 6454 4710 6460
rect 4658 6376 4710 6382
rect 4658 6318 4710 6324
rect 4326 6276 4622 6296
rect 4382 6274 4406 6276
rect 4462 6274 4486 6276
rect 4542 6274 4566 6276
rect 4404 6222 4406 6274
rect 4468 6222 4480 6274
rect 4542 6222 4544 6274
rect 4382 6220 4406 6222
rect 4462 6220 4486 6222
rect 4542 6220 4566 6222
rect 4326 6200 4622 6220
rect 4198 5968 4250 5974
rect 4198 5910 4250 5916
rect 4326 5188 4622 5208
rect 4382 5186 4406 5188
rect 4462 5186 4486 5188
rect 4542 5186 4566 5188
rect 4404 5134 4406 5186
rect 4468 5134 4480 5186
rect 4542 5134 4544 5186
rect 4382 5132 4406 5134
rect 4462 5132 4486 5134
rect 4542 5132 4566 5134
rect 4326 5112 4622 5132
rect 4670 4818 4698 6318
rect 4658 4812 4710 4818
rect 4658 4754 4710 4760
rect 4750 4744 4802 4750
rect 4750 4686 4802 4692
rect 4762 4478 4790 4686
rect 4750 4472 4802 4478
rect 4750 4414 4802 4420
rect 3922 4404 3974 4410
rect 3922 4346 3974 4352
rect 4566 4404 4618 4410
rect 4566 4346 4618 4352
rect 4578 4290 4606 4346
rect 4578 4262 4698 4290
rect 3738 4200 3790 4206
rect 3738 4142 3790 4148
rect 4326 4100 4622 4120
rect 4382 4098 4406 4100
rect 4462 4098 4486 4100
rect 4542 4098 4566 4100
rect 4404 4046 4406 4098
rect 4468 4046 4480 4098
rect 4542 4046 4544 4098
rect 4382 4044 4406 4046
rect 4462 4044 4486 4046
rect 4542 4044 4566 4046
rect 4326 4024 4622 4044
rect 2847 3556 3143 3576
rect 2903 3554 2927 3556
rect 2983 3554 3007 3556
rect 3063 3554 3087 3556
rect 2925 3502 2927 3554
rect 2989 3502 3001 3554
rect 3063 3502 3065 3554
rect 2903 3500 2927 3502
rect 2983 3500 3007 3502
rect 3063 3500 3087 3502
rect 2847 3480 3143 3500
rect 1714 3316 1766 3322
rect 1714 3258 1766 3264
rect 1368 3012 1664 3032
rect 1424 3010 1448 3012
rect 1504 3010 1528 3012
rect 1584 3010 1608 3012
rect 1446 2958 1448 3010
rect 1510 2958 1522 3010
rect 1584 2958 1586 3010
rect 1424 2956 1448 2958
rect 1504 2956 1528 2958
rect 1584 2956 1608 2958
rect 1368 2936 1664 2956
rect 4326 3012 4622 3032
rect 4382 3010 4406 3012
rect 4462 3010 4486 3012
rect 4542 3010 4566 3012
rect 4404 2958 4406 3010
rect 4468 2958 4480 3010
rect 4542 2958 4544 3010
rect 4382 2956 4406 2958
rect 4462 2956 4486 2958
rect 4542 2956 4566 2958
rect 4326 2936 4622 2956
rect 2847 2468 3143 2488
rect 2903 2466 2927 2468
rect 2983 2466 3007 2468
rect 3063 2466 3087 2468
rect 2925 2414 2927 2466
rect 2989 2414 3001 2466
rect 3063 2414 3065 2466
rect 2903 2412 2927 2414
rect 2983 2412 3007 2414
rect 3063 2412 3087 2414
rect 2847 2392 3143 2412
rect 4670 2234 4698 4262
rect 4854 3730 4882 7134
rect 5590 7062 5618 7610
rect 5578 7056 5630 7062
rect 5578 6998 5630 7004
rect 5590 6586 5618 6998
rect 6222 6988 6274 6994
rect 6222 6930 6274 6936
rect 6406 6988 6458 6994
rect 6406 6930 6458 6936
rect 5804 6820 6100 6840
rect 5860 6818 5884 6820
rect 5940 6818 5964 6820
rect 6020 6818 6044 6820
rect 5882 6766 5884 6818
rect 5946 6766 5958 6818
rect 6020 6766 6022 6818
rect 5860 6764 5884 6766
rect 5940 6764 5964 6766
rect 6020 6764 6044 6766
rect 5804 6744 6100 6764
rect 5578 6580 5630 6586
rect 5578 6522 5630 6528
rect 4934 6036 4986 6042
rect 4934 5978 4986 5984
rect 4946 5498 4974 5978
rect 5590 5974 5618 6522
rect 6234 6382 6262 6930
rect 6222 6376 6274 6382
rect 6222 6318 6274 6324
rect 5302 5968 5354 5974
rect 5302 5910 5354 5916
rect 5578 5968 5630 5974
rect 5578 5910 5630 5916
rect 4934 5492 4986 5498
rect 4934 5434 4986 5440
rect 4842 3724 4894 3730
rect 4842 3666 4894 3672
rect 5314 2370 5342 5910
rect 5590 5498 5618 5910
rect 5804 5732 6100 5752
rect 5860 5730 5884 5732
rect 5940 5730 5964 5732
rect 6020 5730 6044 5732
rect 5882 5678 5884 5730
rect 5946 5678 5958 5730
rect 6020 5678 6022 5730
rect 5860 5676 5884 5678
rect 5940 5676 5964 5678
rect 6020 5676 6044 5678
rect 5804 5656 6100 5676
rect 5946 5560 5998 5566
rect 5946 5502 5998 5508
rect 5578 5492 5630 5498
rect 5578 5434 5630 5440
rect 5590 4954 5618 5434
rect 5958 4954 5986 5502
rect 6130 5424 6182 5430
rect 6130 5366 6182 5372
rect 5578 4948 5630 4954
rect 5578 4890 5630 4896
rect 5946 4948 5998 4954
rect 5946 4890 5998 4896
rect 5804 4644 6100 4664
rect 5860 4642 5884 4644
rect 5940 4642 5964 4644
rect 6020 4642 6044 4644
rect 5882 4590 5884 4642
rect 5946 4590 5958 4642
rect 6020 4590 6022 4642
rect 5860 4588 5884 4590
rect 5940 4588 5964 4590
rect 6020 4588 6044 4590
rect 5804 4568 6100 4588
rect 6142 4342 6170 5366
rect 6130 4336 6182 4342
rect 6130 4278 6182 4284
rect 5670 4200 5722 4206
rect 5670 4142 5722 4148
rect 5682 3866 5710 4142
rect 6142 4002 6170 4278
rect 6234 4206 6262 6318
rect 6314 5560 6366 5566
rect 6314 5502 6366 5508
rect 6222 4200 6274 4206
rect 6222 4142 6274 4148
rect 6130 3996 6182 4002
rect 6130 3938 6182 3944
rect 5670 3860 5722 3866
rect 5670 3802 5722 3808
rect 5804 3556 6100 3576
rect 5860 3554 5884 3556
rect 5940 3554 5964 3556
rect 6020 3554 6044 3556
rect 5882 3502 5884 3554
rect 5946 3502 5958 3554
rect 6020 3502 6022 3554
rect 5860 3500 5884 3502
rect 5940 3500 5964 3502
rect 6020 3500 6044 3502
rect 5804 3480 6100 3500
rect 6326 3458 6354 5502
rect 6418 4546 6446 6930
rect 6510 5090 6538 8766
rect 6498 5084 6550 5090
rect 6498 5026 6550 5032
rect 6602 4954 6630 8886
rect 6694 6518 6722 9566
rect 7154 9442 7182 11826
rect 7283 11716 7579 11736
rect 7339 11714 7363 11716
rect 7419 11714 7443 11716
rect 7499 11714 7523 11716
rect 7361 11662 7363 11714
rect 7425 11662 7437 11714
rect 7499 11662 7501 11714
rect 7339 11660 7363 11662
rect 7419 11660 7443 11662
rect 7499 11660 7523 11662
rect 7283 11640 7579 11660
rect 7283 10628 7579 10648
rect 7339 10626 7363 10628
rect 7419 10626 7443 10628
rect 7499 10626 7523 10628
rect 7361 10574 7363 10626
rect 7425 10574 7437 10626
rect 7499 10574 7501 10626
rect 7339 10572 7363 10574
rect 7419 10572 7443 10574
rect 7499 10572 7523 10574
rect 7283 10552 7579 10572
rect 7614 10258 7642 14478
rect 7706 14134 7734 16314
rect 9256 15864 9312 15873
rect 9256 15799 9312 15808
rect 7786 15080 7838 15086
rect 7786 15022 7838 15028
rect 7694 14128 7746 14134
rect 7694 14070 7746 14076
rect 7694 11340 7746 11346
rect 7694 11282 7746 11288
rect 7602 10252 7654 10258
rect 7602 10194 7654 10200
rect 7283 9540 7579 9560
rect 7339 9538 7363 9540
rect 7419 9538 7443 9540
rect 7499 9538 7523 9540
rect 7361 9486 7363 9538
rect 7425 9486 7437 9538
rect 7499 9486 7501 9538
rect 7339 9484 7363 9486
rect 7419 9484 7443 9486
rect 7499 9484 7523 9486
rect 7283 9464 7579 9484
rect 7142 9436 7194 9442
rect 7142 9378 7194 9384
rect 7283 8452 7579 8472
rect 7339 8450 7363 8452
rect 7419 8450 7443 8452
rect 7499 8450 7523 8452
rect 7361 8398 7363 8450
rect 7425 8398 7437 8450
rect 7499 8398 7501 8450
rect 7339 8396 7363 8398
rect 7419 8396 7443 8398
rect 7499 8396 7523 8398
rect 7283 8376 7579 8396
rect 7602 8076 7654 8082
rect 7602 8018 7654 8024
rect 7283 7364 7579 7384
rect 7339 7362 7363 7364
rect 7419 7362 7443 7364
rect 7499 7362 7523 7364
rect 7361 7310 7363 7362
rect 7425 7310 7437 7362
rect 7499 7310 7501 7362
rect 7339 7308 7363 7310
rect 7419 7308 7443 7310
rect 7499 7308 7523 7310
rect 7283 7288 7579 7308
rect 6774 6920 6826 6926
rect 6774 6862 6826 6868
rect 6786 6518 6814 6862
rect 6682 6512 6734 6518
rect 6682 6454 6734 6460
rect 6774 6512 6826 6518
rect 6774 6454 6826 6460
rect 7283 6276 7579 6296
rect 7339 6274 7363 6276
rect 7419 6274 7443 6276
rect 7499 6274 7523 6276
rect 7361 6222 7363 6274
rect 7425 6222 7437 6274
rect 7499 6222 7501 6274
rect 7339 6220 7363 6222
rect 7419 6220 7443 6222
rect 7499 6220 7523 6222
rect 7283 6200 7579 6220
rect 7050 5968 7102 5974
rect 7050 5910 7102 5916
rect 6590 4948 6642 4954
rect 6590 4890 6642 4896
rect 6406 4540 6458 4546
rect 6406 4482 6458 4488
rect 6314 3452 6366 3458
rect 6314 3394 6366 3400
rect 6130 3316 6182 3322
rect 6130 3258 6182 3264
rect 6142 2710 6170 3258
rect 7062 2914 7090 5910
rect 7283 5188 7579 5208
rect 7339 5186 7363 5188
rect 7419 5186 7443 5188
rect 7499 5186 7523 5188
rect 7361 5134 7363 5186
rect 7425 5134 7437 5186
rect 7499 5134 7501 5186
rect 7339 5132 7363 5134
rect 7419 5132 7443 5134
rect 7499 5132 7523 5134
rect 7283 5112 7579 5132
rect 7283 4100 7579 4120
rect 7339 4098 7363 4100
rect 7419 4098 7443 4100
rect 7499 4098 7523 4100
rect 7361 4046 7363 4098
rect 7425 4046 7437 4098
rect 7499 4046 7501 4098
rect 7339 4044 7363 4046
rect 7419 4044 7443 4046
rect 7499 4044 7523 4046
rect 7283 4024 7579 4044
rect 7283 3012 7579 3032
rect 7339 3010 7363 3012
rect 7419 3010 7443 3012
rect 7499 3010 7523 3012
rect 7361 2958 7363 3010
rect 7425 2958 7437 3010
rect 7499 2958 7501 3010
rect 7339 2956 7363 2958
rect 7419 2956 7443 2958
rect 7499 2956 7523 2958
rect 7283 2936 7579 2956
rect 7050 2908 7102 2914
rect 7050 2850 7102 2856
rect 6130 2704 6182 2710
rect 6130 2646 6182 2652
rect 5804 2468 6100 2488
rect 5860 2466 5884 2468
rect 5940 2466 5964 2468
rect 6020 2466 6044 2468
rect 5882 2414 5884 2466
rect 5946 2414 5958 2466
rect 6020 2414 6022 2466
rect 5860 2412 5884 2414
rect 5940 2412 5964 2414
rect 6020 2412 6044 2414
rect 5804 2392 6100 2412
rect 5302 2364 5354 2370
rect 5302 2306 5354 2312
rect 4658 2228 4710 2234
rect 4658 2170 4710 2176
rect 7614 2098 7642 8018
rect 7706 6586 7734 11282
rect 7798 9170 7826 15022
rect 9270 11482 9298 15799
rect 15696 15048 15752 15057
rect 15696 14983 15752 14992
rect 15514 13652 15566 13658
rect 15514 13594 15566 13600
rect 15526 13561 15554 13594
rect 15512 13552 15568 13561
rect 15512 13487 15568 13496
rect 15604 12736 15660 12745
rect 15604 12671 15660 12680
rect 11464 11920 11520 11929
rect 11464 11855 11520 11864
rect 9258 11476 9310 11482
rect 9258 11418 9310 11424
rect 7878 11272 7930 11278
rect 7878 11214 7930 11220
rect 7786 9164 7838 9170
rect 7786 9106 7838 9112
rect 7890 8830 7918 11214
rect 8704 11104 8760 11113
rect 8704 11039 8760 11048
rect 8614 10524 8666 10530
rect 8614 10466 8666 10472
rect 8626 10410 8654 10466
rect 8718 10410 8746 11039
rect 8626 10382 8746 10410
rect 8626 10246 8746 10274
rect 8626 10190 8654 10246
rect 8614 10184 8666 10190
rect 8614 10126 8666 10132
rect 8718 9986 8746 10246
rect 8706 9980 8758 9986
rect 8706 9922 8758 9928
rect 11478 9782 11506 11855
rect 15618 10870 15646 12671
rect 15710 11822 15738 14983
rect 15972 14368 16028 14377
rect 15972 14303 16028 14312
rect 15698 11816 15750 11822
rect 15698 11758 15750 11764
rect 15606 10864 15658 10870
rect 15606 10806 15658 10812
rect 11648 10288 11704 10297
rect 11648 10223 11704 10232
rect 11466 9776 11518 9782
rect 11466 9718 11518 9724
rect 11556 9608 11612 9617
rect 11556 9543 11612 9552
rect 7970 9096 8022 9102
rect 7970 9038 8022 9044
rect 7878 8824 7930 8830
rect 7878 8766 7930 8772
rect 7982 8626 8010 9038
rect 8522 8824 8574 8830
rect 11374 8824 11426 8830
rect 8522 8766 8574 8772
rect 11372 8792 11374 8801
rect 11426 8792 11428 8801
rect 7970 8620 8022 8626
rect 7970 8562 8022 8568
rect 7878 8076 7930 8082
rect 7878 8018 7930 8024
rect 7890 7130 7918 8018
rect 7878 7124 7930 7130
rect 7878 7066 7930 7072
rect 7694 6580 7746 6586
rect 7694 6522 7746 6528
rect 7706 6178 7734 6522
rect 7694 6172 7746 6178
rect 7694 6114 7746 6120
rect 7694 6036 7746 6042
rect 7694 5978 7746 5984
rect 7706 3866 7734 5978
rect 7786 5424 7838 5430
rect 7786 5366 7838 5372
rect 7694 3860 7746 3866
rect 7694 3802 7746 3808
rect 7798 2302 7826 5366
rect 7890 5090 7918 7066
rect 7878 5084 7930 5090
rect 7878 5026 7930 5032
rect 7982 3254 8010 8562
rect 8338 8348 8390 8354
rect 8338 8290 8390 8296
rect 8350 8257 8378 8290
rect 8336 8248 8392 8257
rect 8336 8183 8392 8192
rect 8534 3322 8562 8766
rect 8614 8756 8666 8762
rect 11372 8727 11428 8736
rect 8614 8698 8666 8704
rect 8626 8354 8654 8698
rect 11466 8688 11518 8694
rect 11466 8630 11518 8636
rect 8614 8348 8666 8354
rect 8614 8290 8666 8296
rect 11372 7976 11428 7985
rect 11372 7911 11428 7920
rect 11386 6994 11414 7911
rect 11478 7169 11506 8630
rect 11570 7606 11598 9543
rect 11662 8762 11690 10223
rect 15986 9306 16014 14303
rect 23806 9986 23834 17431
rect 23794 9980 23846 9986
rect 23794 9922 23846 9928
rect 15974 9300 16026 9306
rect 15974 9242 16026 9248
rect 24082 9102 24110 18247
rect 24070 9096 24122 9102
rect 24070 9038 24122 9044
rect 11650 8756 11702 8762
rect 11650 8698 11702 8704
rect 11558 7600 11610 7606
rect 11558 7542 11610 7548
rect 23794 7192 23846 7198
rect 11464 7160 11520 7169
rect 23794 7134 23846 7140
rect 11464 7095 11520 7104
rect 11374 6988 11426 6994
rect 11374 6930 11426 6936
rect 11374 6580 11426 6586
rect 11374 6522 11426 6528
rect 11386 6353 11414 6522
rect 11466 6512 11518 6518
rect 11466 6454 11518 6460
rect 11372 6344 11428 6353
rect 11372 6279 11428 6288
rect 11478 5537 11506 6454
rect 11558 5900 11610 5906
rect 11558 5842 11610 5848
rect 11464 5528 11520 5537
rect 11464 5463 11520 5472
rect 11374 5084 11426 5090
rect 11374 5026 11426 5032
rect 11386 4857 11414 5026
rect 11372 4848 11428 4857
rect 11372 4783 11428 4792
rect 11374 4744 11426 4750
rect 11374 4686 11426 4692
rect 8522 3316 8574 3322
rect 8522 3258 8574 3264
rect 7970 3248 8022 3254
rect 11386 3225 11414 4686
rect 11570 4041 11598 5842
rect 11556 4032 11612 4041
rect 11556 3967 11612 3976
rect 7970 3190 8022 3196
rect 11372 3216 11428 3225
rect 11372 3151 11428 3160
rect 15698 3112 15750 3118
rect 15698 3054 15750 3060
rect 15512 2400 15568 2409
rect 15512 2335 15568 2344
rect 15606 2364 15658 2370
rect 15526 2302 15554 2335
rect 15606 2306 15658 2312
rect 7786 2296 7838 2302
rect 7786 2238 7838 2244
rect 15514 2296 15566 2302
rect 15514 2238 15566 2244
rect 7602 2092 7654 2098
rect 7602 2034 7654 2040
rect 1368 1924 1664 1944
rect 1424 1922 1448 1924
rect 1504 1922 1528 1924
rect 1584 1922 1608 1924
rect 1446 1870 1448 1922
rect 1510 1870 1522 1922
rect 1584 1870 1586 1922
rect 1424 1868 1448 1870
rect 1504 1868 1528 1870
rect 1584 1868 1608 1870
rect 1368 1848 1664 1868
rect 4326 1924 4622 1944
rect 4382 1922 4406 1924
rect 4462 1922 4486 1924
rect 4542 1922 4566 1924
rect 4404 1870 4406 1922
rect 4468 1870 4480 1922
rect 4542 1870 4544 1922
rect 4382 1868 4406 1870
rect 4462 1868 4486 1870
rect 4542 1868 4566 1870
rect 4326 1848 4622 1868
rect 7283 1924 7579 1944
rect 7339 1922 7363 1924
rect 7419 1922 7443 1924
rect 7499 1922 7523 1924
rect 7361 1870 7363 1922
rect 7425 1870 7437 1922
rect 7499 1870 7501 1922
rect 7339 1868 7363 1870
rect 7419 1868 7443 1870
rect 7499 1868 7523 1870
rect 7283 1848 7579 1868
rect 15618 1593 15646 2306
rect 15604 1584 15660 1593
rect 15604 1519 15660 1528
rect 15710 97 15738 3054
rect 23806 777 23834 7134
rect 23792 768 23848 777
rect 23792 703 23848 712
rect 15696 88 15752 97
rect 15696 23 15752 32
<< via2 >>
rect 24068 18256 24124 18312
rect 23792 17440 23848 17496
rect 15512 16624 15568 16680
rect 1368 16066 1424 16068
rect 1448 16066 1504 16068
rect 1528 16066 1584 16068
rect 1608 16066 1664 16068
rect 1368 16014 1394 16066
rect 1394 16014 1424 16066
rect 1448 16014 1458 16066
rect 1458 16014 1504 16066
rect 1528 16014 1574 16066
rect 1574 16014 1584 16066
rect 1608 16014 1638 16066
rect 1638 16014 1664 16066
rect 1368 16012 1424 16014
rect 1448 16012 1504 16014
rect 1528 16012 1584 16014
rect 1608 16012 1664 16014
rect 4326 16066 4382 16068
rect 4406 16066 4462 16068
rect 4486 16066 4542 16068
rect 4566 16066 4622 16068
rect 4326 16014 4352 16066
rect 4352 16014 4382 16066
rect 4406 16014 4416 16066
rect 4416 16014 4462 16066
rect 4486 16014 4532 16066
rect 4532 16014 4542 16066
rect 4566 16014 4596 16066
rect 4596 16014 4622 16066
rect 4326 16012 4382 16014
rect 4406 16012 4462 16014
rect 4486 16012 4542 16014
rect 4566 16012 4622 16014
rect 7283 16066 7339 16068
rect 7363 16066 7419 16068
rect 7443 16066 7499 16068
rect 7523 16066 7579 16068
rect 7283 16014 7309 16066
rect 7309 16014 7339 16066
rect 7363 16014 7373 16066
rect 7373 16014 7419 16066
rect 7443 16014 7489 16066
rect 7489 16014 7499 16066
rect 7523 16014 7553 16066
rect 7553 16014 7579 16066
rect 7283 16012 7339 16014
rect 7363 16012 7419 16014
rect 7443 16012 7499 16014
rect 7523 16012 7579 16014
rect 2847 15522 2903 15524
rect 2927 15522 2983 15524
rect 3007 15522 3063 15524
rect 3087 15522 3143 15524
rect 2847 15470 2873 15522
rect 2873 15470 2903 15522
rect 2927 15470 2937 15522
rect 2937 15470 2983 15522
rect 3007 15470 3053 15522
rect 3053 15470 3063 15522
rect 3087 15470 3117 15522
rect 3117 15470 3143 15522
rect 2847 15468 2903 15470
rect 2927 15468 2983 15470
rect 3007 15468 3063 15470
rect 3087 15468 3143 15470
rect 5804 15522 5860 15524
rect 5884 15522 5940 15524
rect 5964 15522 6020 15524
rect 6044 15522 6100 15524
rect 5804 15470 5830 15522
rect 5830 15470 5860 15522
rect 5884 15470 5894 15522
rect 5894 15470 5940 15522
rect 5964 15470 6010 15522
rect 6010 15470 6020 15522
rect 6044 15470 6074 15522
rect 6074 15470 6100 15522
rect 5804 15468 5860 15470
rect 5884 15468 5940 15470
rect 5964 15468 6020 15470
rect 6044 15468 6100 15470
rect 1368 14978 1424 14980
rect 1448 14978 1504 14980
rect 1528 14978 1584 14980
rect 1608 14978 1664 14980
rect 1368 14926 1394 14978
rect 1394 14926 1424 14978
rect 1448 14926 1458 14978
rect 1458 14926 1504 14978
rect 1528 14926 1574 14978
rect 1574 14926 1584 14978
rect 1608 14926 1638 14978
rect 1638 14926 1664 14978
rect 1368 14924 1424 14926
rect 1448 14924 1504 14926
rect 1528 14924 1584 14926
rect 1608 14924 1664 14926
rect 4326 14978 4382 14980
rect 4406 14978 4462 14980
rect 4486 14978 4542 14980
rect 4566 14978 4622 14980
rect 4326 14926 4352 14978
rect 4352 14926 4382 14978
rect 4406 14926 4416 14978
rect 4416 14926 4462 14978
rect 4486 14926 4532 14978
rect 4532 14926 4542 14978
rect 4566 14926 4596 14978
rect 4596 14926 4622 14978
rect 4326 14924 4382 14926
rect 4406 14924 4462 14926
rect 4486 14924 4542 14926
rect 4566 14924 4622 14926
rect 1368 13890 1424 13892
rect 1448 13890 1504 13892
rect 1528 13890 1584 13892
rect 1608 13890 1664 13892
rect 1368 13838 1394 13890
rect 1394 13838 1424 13890
rect 1448 13838 1458 13890
rect 1458 13838 1504 13890
rect 1528 13838 1574 13890
rect 1574 13838 1584 13890
rect 1608 13838 1638 13890
rect 1638 13838 1664 13890
rect 1368 13836 1424 13838
rect 1448 13836 1504 13838
rect 1528 13836 1584 13838
rect 1608 13836 1664 13838
rect 1368 12802 1424 12804
rect 1448 12802 1504 12804
rect 1528 12802 1584 12804
rect 1608 12802 1664 12804
rect 1368 12750 1394 12802
rect 1394 12750 1424 12802
rect 1448 12750 1458 12802
rect 1458 12750 1504 12802
rect 1528 12750 1574 12802
rect 1574 12750 1584 12802
rect 1608 12750 1638 12802
rect 1638 12750 1664 12802
rect 1368 12748 1424 12750
rect 1448 12748 1504 12750
rect 1528 12748 1584 12750
rect 1608 12748 1664 12750
rect 1368 11714 1424 11716
rect 1448 11714 1504 11716
rect 1528 11714 1584 11716
rect 1608 11714 1664 11716
rect 1368 11662 1394 11714
rect 1394 11662 1424 11714
rect 1448 11662 1458 11714
rect 1458 11662 1504 11714
rect 1528 11662 1574 11714
rect 1574 11662 1584 11714
rect 1608 11662 1638 11714
rect 1638 11662 1664 11714
rect 1368 11660 1424 11662
rect 1448 11660 1504 11662
rect 1528 11660 1584 11662
rect 1608 11660 1664 11662
rect 1368 10626 1424 10628
rect 1448 10626 1504 10628
rect 1528 10626 1584 10628
rect 1608 10626 1664 10628
rect 1368 10574 1394 10626
rect 1394 10574 1424 10626
rect 1448 10574 1458 10626
rect 1458 10574 1504 10626
rect 1528 10574 1574 10626
rect 1574 10574 1584 10626
rect 1608 10574 1638 10626
rect 1638 10574 1664 10626
rect 1368 10572 1424 10574
rect 1448 10572 1504 10574
rect 1528 10572 1584 10574
rect 1608 10572 1664 10574
rect 1368 9538 1424 9540
rect 1448 9538 1504 9540
rect 1528 9538 1584 9540
rect 1608 9538 1664 9540
rect 1368 9486 1394 9538
rect 1394 9486 1424 9538
rect 1448 9486 1458 9538
rect 1458 9486 1504 9538
rect 1528 9486 1574 9538
rect 1574 9486 1584 9538
rect 1608 9486 1638 9538
rect 1638 9486 1664 9538
rect 1368 9484 1424 9486
rect 1448 9484 1504 9486
rect 1528 9484 1584 9486
rect 1608 9484 1664 9486
rect 2847 14434 2903 14436
rect 2927 14434 2983 14436
rect 3007 14434 3063 14436
rect 3087 14434 3143 14436
rect 2847 14382 2873 14434
rect 2873 14382 2903 14434
rect 2927 14382 2937 14434
rect 2937 14382 2983 14434
rect 3007 14382 3053 14434
rect 3053 14382 3063 14434
rect 3087 14382 3117 14434
rect 3117 14382 3143 14434
rect 2847 14380 2903 14382
rect 2927 14380 2983 14382
rect 3007 14380 3063 14382
rect 3087 14380 3143 14382
rect 4326 13890 4382 13892
rect 4406 13890 4462 13892
rect 4486 13890 4542 13892
rect 4566 13890 4622 13892
rect 4326 13838 4352 13890
rect 4352 13838 4382 13890
rect 4406 13838 4416 13890
rect 4416 13838 4462 13890
rect 4486 13838 4532 13890
rect 4532 13838 4542 13890
rect 4566 13838 4596 13890
rect 4596 13838 4622 13890
rect 4326 13836 4382 13838
rect 4406 13836 4462 13838
rect 4486 13836 4542 13838
rect 4566 13836 4622 13838
rect 2847 13346 2903 13348
rect 2927 13346 2983 13348
rect 3007 13346 3063 13348
rect 3087 13346 3143 13348
rect 2847 13294 2873 13346
rect 2873 13294 2903 13346
rect 2927 13294 2937 13346
rect 2937 13294 2983 13346
rect 3007 13294 3053 13346
rect 3053 13294 3063 13346
rect 3087 13294 3117 13346
rect 3117 13294 3143 13346
rect 2847 13292 2903 13294
rect 2927 13292 2983 13294
rect 3007 13292 3063 13294
rect 3087 13292 3143 13294
rect 2847 12258 2903 12260
rect 2927 12258 2983 12260
rect 3007 12258 3063 12260
rect 3087 12258 3143 12260
rect 2847 12206 2873 12258
rect 2873 12206 2903 12258
rect 2927 12206 2937 12258
rect 2937 12206 2983 12258
rect 3007 12206 3053 12258
rect 3053 12206 3063 12258
rect 3087 12206 3117 12258
rect 3117 12206 3143 12258
rect 2847 12204 2903 12206
rect 2927 12204 2983 12206
rect 3007 12204 3063 12206
rect 3087 12204 3143 12206
rect 2847 11170 2903 11172
rect 2927 11170 2983 11172
rect 3007 11170 3063 11172
rect 3087 11170 3143 11172
rect 2847 11118 2873 11170
rect 2873 11118 2903 11170
rect 2927 11118 2937 11170
rect 2937 11118 2983 11170
rect 3007 11118 3053 11170
rect 3053 11118 3063 11170
rect 3087 11118 3117 11170
rect 3117 11118 3143 11170
rect 2847 11116 2903 11118
rect 2927 11116 2983 11118
rect 3007 11116 3063 11118
rect 3087 11116 3143 11118
rect 2080 10252 2136 10288
rect 2080 10232 2082 10252
rect 2082 10232 2134 10252
rect 2134 10232 2136 10252
rect 1368 8450 1424 8452
rect 1448 8450 1504 8452
rect 1528 8450 1584 8452
rect 1608 8450 1664 8452
rect 1368 8398 1394 8450
rect 1394 8398 1424 8450
rect 1448 8398 1458 8450
rect 1458 8398 1504 8450
rect 1528 8398 1574 8450
rect 1574 8398 1584 8450
rect 1608 8398 1638 8450
rect 1638 8398 1664 8450
rect 1368 8396 1424 8398
rect 1448 8396 1504 8398
rect 1528 8396 1584 8398
rect 1608 8396 1664 8398
rect 1368 7362 1424 7364
rect 1448 7362 1504 7364
rect 1528 7362 1584 7364
rect 1608 7362 1664 7364
rect 1368 7310 1394 7362
rect 1394 7310 1424 7362
rect 1448 7310 1458 7362
rect 1458 7310 1504 7362
rect 1528 7310 1574 7362
rect 1574 7310 1584 7362
rect 1608 7310 1638 7362
rect 1638 7310 1664 7362
rect 1368 7308 1424 7310
rect 1448 7308 1504 7310
rect 1528 7308 1584 7310
rect 1608 7308 1664 7310
rect 1368 6274 1424 6276
rect 1448 6274 1504 6276
rect 1528 6274 1584 6276
rect 1608 6274 1664 6276
rect 1368 6222 1394 6274
rect 1394 6222 1424 6274
rect 1448 6222 1458 6274
rect 1458 6222 1504 6274
rect 1528 6222 1574 6274
rect 1574 6222 1584 6274
rect 1608 6222 1638 6274
rect 1638 6222 1664 6274
rect 1368 6220 1424 6222
rect 1448 6220 1504 6222
rect 1528 6220 1584 6222
rect 1608 6220 1664 6222
rect 1368 5186 1424 5188
rect 1448 5186 1504 5188
rect 1528 5186 1584 5188
rect 1608 5186 1664 5188
rect 1368 5134 1394 5186
rect 1394 5134 1424 5186
rect 1448 5134 1458 5186
rect 1458 5134 1504 5186
rect 1528 5134 1574 5186
rect 1574 5134 1584 5186
rect 1608 5134 1638 5186
rect 1638 5134 1664 5186
rect 1368 5132 1424 5134
rect 1448 5132 1504 5134
rect 1528 5132 1584 5134
rect 1608 5132 1664 5134
rect 1368 4098 1424 4100
rect 1448 4098 1504 4100
rect 1528 4098 1584 4100
rect 1608 4098 1664 4100
rect 1368 4046 1394 4098
rect 1394 4046 1424 4098
rect 1448 4046 1458 4098
rect 1458 4046 1504 4098
rect 1528 4046 1574 4098
rect 1574 4046 1584 4098
rect 1608 4046 1638 4098
rect 1638 4046 1664 4098
rect 1368 4044 1424 4046
rect 1448 4044 1504 4046
rect 1528 4044 1584 4046
rect 1608 4044 1664 4046
rect 2847 10082 2903 10084
rect 2927 10082 2983 10084
rect 3007 10082 3063 10084
rect 3087 10082 3143 10084
rect 2847 10030 2873 10082
rect 2873 10030 2903 10082
rect 2927 10030 2937 10082
rect 2937 10030 2983 10082
rect 3007 10030 3053 10082
rect 3053 10030 3063 10082
rect 3087 10030 3117 10082
rect 3117 10030 3143 10082
rect 2847 10028 2903 10030
rect 2927 10028 2983 10030
rect 3007 10028 3063 10030
rect 3087 10028 3143 10030
rect 2847 8994 2903 8996
rect 2927 8994 2983 8996
rect 3007 8994 3063 8996
rect 3087 8994 3143 8996
rect 2847 8942 2873 8994
rect 2873 8942 2903 8994
rect 2927 8942 2937 8994
rect 2937 8942 2983 8994
rect 3007 8942 3053 8994
rect 3053 8942 3063 8994
rect 3087 8942 3117 8994
rect 3117 8942 3143 8994
rect 2847 8940 2903 8942
rect 2927 8940 2983 8942
rect 3007 8940 3063 8942
rect 3087 8940 3143 8942
rect 3276 8212 3332 8248
rect 3276 8192 3278 8212
rect 3278 8192 3330 8212
rect 3330 8192 3332 8212
rect 2847 7906 2903 7908
rect 2927 7906 2983 7908
rect 3007 7906 3063 7908
rect 3087 7906 3143 7908
rect 2847 7854 2873 7906
rect 2873 7854 2903 7906
rect 2927 7854 2937 7906
rect 2937 7854 2983 7906
rect 3007 7854 3053 7906
rect 3053 7854 3063 7906
rect 3087 7854 3117 7906
rect 3117 7854 3143 7906
rect 2847 7852 2903 7854
rect 2927 7852 2983 7854
rect 3007 7852 3063 7854
rect 3087 7852 3143 7854
rect 2847 6818 2903 6820
rect 2927 6818 2983 6820
rect 3007 6818 3063 6820
rect 3087 6818 3143 6820
rect 2847 6766 2873 6818
rect 2873 6766 2903 6818
rect 2927 6766 2937 6818
rect 2937 6766 2983 6818
rect 3007 6766 3053 6818
rect 3053 6766 3063 6818
rect 3087 6766 3117 6818
rect 3117 6766 3143 6818
rect 2847 6764 2903 6766
rect 2927 6764 2983 6766
rect 3007 6764 3063 6766
rect 3087 6764 3143 6766
rect 4326 12802 4382 12804
rect 4406 12802 4462 12804
rect 4486 12802 4542 12804
rect 4566 12802 4622 12804
rect 4326 12750 4352 12802
rect 4352 12750 4382 12802
rect 4406 12750 4416 12802
rect 4416 12750 4462 12802
rect 4486 12750 4532 12802
rect 4532 12750 4542 12802
rect 4566 12750 4596 12802
rect 4596 12750 4622 12802
rect 4326 12748 4382 12750
rect 4406 12748 4462 12750
rect 4486 12748 4542 12750
rect 4566 12748 4622 12750
rect 2847 5730 2903 5732
rect 2927 5730 2983 5732
rect 3007 5730 3063 5732
rect 3087 5730 3143 5732
rect 2847 5678 2873 5730
rect 2873 5678 2903 5730
rect 2927 5678 2937 5730
rect 2937 5678 2983 5730
rect 3007 5678 3053 5730
rect 3053 5678 3063 5730
rect 3087 5678 3117 5730
rect 3117 5678 3143 5730
rect 2847 5676 2903 5678
rect 2927 5676 2983 5678
rect 3007 5676 3063 5678
rect 3087 5676 3143 5678
rect 5804 14434 5860 14436
rect 5884 14434 5940 14436
rect 5964 14434 6020 14436
rect 6044 14434 6100 14436
rect 5804 14382 5830 14434
rect 5830 14382 5860 14434
rect 5884 14382 5894 14434
rect 5894 14382 5940 14434
rect 5964 14382 6010 14434
rect 6010 14382 6020 14434
rect 6044 14382 6074 14434
rect 6074 14382 6100 14434
rect 5804 14380 5860 14382
rect 5884 14380 5940 14382
rect 5964 14380 6020 14382
rect 6044 14380 6100 14382
rect 7283 14978 7339 14980
rect 7363 14978 7419 14980
rect 7443 14978 7499 14980
rect 7523 14978 7579 14980
rect 7283 14926 7309 14978
rect 7309 14926 7339 14978
rect 7363 14926 7373 14978
rect 7373 14926 7419 14978
rect 7443 14926 7489 14978
rect 7489 14926 7499 14978
rect 7523 14926 7553 14978
rect 7553 14926 7579 14978
rect 7283 14924 7339 14926
rect 7363 14924 7419 14926
rect 7443 14924 7499 14926
rect 7523 14924 7579 14926
rect 5804 13346 5860 13348
rect 5884 13346 5940 13348
rect 5964 13346 6020 13348
rect 6044 13346 6100 13348
rect 5804 13294 5830 13346
rect 5830 13294 5860 13346
rect 5884 13294 5894 13346
rect 5894 13294 5940 13346
rect 5964 13294 6010 13346
rect 6010 13294 6020 13346
rect 6044 13294 6074 13346
rect 6074 13294 6100 13346
rect 5804 13292 5860 13294
rect 5884 13292 5940 13294
rect 5964 13292 6020 13294
rect 6044 13292 6100 13294
rect 4326 11714 4382 11716
rect 4406 11714 4462 11716
rect 4486 11714 4542 11716
rect 4566 11714 4622 11716
rect 4326 11662 4352 11714
rect 4352 11662 4382 11714
rect 4406 11662 4416 11714
rect 4416 11662 4462 11714
rect 4486 11662 4532 11714
rect 4532 11662 4542 11714
rect 4566 11662 4596 11714
rect 4596 11662 4622 11714
rect 4326 11660 4382 11662
rect 4406 11660 4462 11662
rect 4486 11660 4542 11662
rect 4566 11660 4622 11662
rect 4326 10626 4382 10628
rect 4406 10626 4462 10628
rect 4486 10626 4542 10628
rect 4566 10626 4622 10628
rect 4326 10574 4352 10626
rect 4352 10574 4382 10626
rect 4406 10574 4416 10626
rect 4416 10574 4462 10626
rect 4486 10574 4532 10626
rect 4532 10574 4542 10626
rect 4566 10574 4596 10626
rect 4596 10574 4622 10626
rect 4326 10572 4382 10574
rect 4406 10572 4462 10574
rect 4486 10572 4542 10574
rect 4566 10572 4622 10574
rect 4326 9538 4382 9540
rect 4406 9538 4462 9540
rect 4486 9538 4542 9540
rect 4566 9538 4622 9540
rect 4326 9486 4352 9538
rect 4352 9486 4382 9538
rect 4406 9486 4416 9538
rect 4416 9486 4462 9538
rect 4486 9486 4532 9538
rect 4532 9486 4542 9538
rect 4566 9486 4596 9538
rect 4596 9486 4622 9538
rect 4326 9484 4382 9486
rect 4406 9484 4462 9486
rect 4486 9484 4542 9486
rect 4566 9484 4622 9486
rect 2847 4642 2903 4644
rect 2927 4642 2983 4644
rect 3007 4642 3063 4644
rect 3087 4642 3143 4644
rect 2847 4590 2873 4642
rect 2873 4590 2903 4642
rect 2927 4590 2937 4642
rect 2937 4590 2983 4642
rect 3007 4590 3053 4642
rect 3053 4590 3063 4642
rect 3087 4590 3117 4642
rect 3117 4590 3143 4642
rect 2847 4588 2903 4590
rect 2927 4588 2983 4590
rect 3007 4588 3063 4590
rect 3087 4588 3143 4590
rect 4326 8450 4382 8452
rect 4406 8450 4462 8452
rect 4486 8450 4542 8452
rect 4566 8450 4622 8452
rect 4326 8398 4352 8450
rect 4352 8398 4382 8450
rect 4406 8398 4416 8450
rect 4416 8398 4462 8450
rect 4486 8398 4532 8450
rect 4532 8398 4542 8450
rect 4566 8398 4596 8450
rect 4596 8398 4622 8450
rect 4326 8396 4382 8398
rect 4406 8396 4462 8398
rect 4486 8396 4542 8398
rect 4566 8396 4622 8398
rect 5804 12258 5860 12260
rect 5884 12258 5940 12260
rect 5964 12258 6020 12260
rect 6044 12258 6100 12260
rect 5804 12206 5830 12258
rect 5830 12206 5860 12258
rect 5884 12206 5894 12258
rect 5894 12206 5940 12258
rect 5964 12206 6010 12258
rect 6010 12206 6020 12258
rect 6044 12206 6074 12258
rect 6074 12206 6100 12258
rect 5804 12204 5860 12206
rect 5884 12204 5940 12206
rect 5964 12204 6020 12206
rect 6044 12204 6100 12206
rect 5804 11170 5860 11172
rect 5884 11170 5940 11172
rect 5964 11170 6020 11172
rect 6044 11170 6100 11172
rect 5804 11118 5830 11170
rect 5830 11118 5860 11170
rect 5884 11118 5894 11170
rect 5894 11118 5940 11170
rect 5964 11118 6010 11170
rect 6010 11118 6020 11170
rect 6044 11118 6074 11170
rect 6074 11118 6100 11170
rect 5804 11116 5860 11118
rect 5884 11116 5940 11118
rect 5964 11116 6020 11118
rect 6044 11116 6100 11118
rect 5576 10268 5578 10288
rect 5578 10268 5630 10288
rect 5630 10268 5632 10288
rect 5576 10232 5632 10268
rect 5804 10082 5860 10084
rect 5884 10082 5940 10084
rect 5964 10082 6020 10084
rect 6044 10082 6100 10084
rect 5804 10030 5830 10082
rect 5830 10030 5860 10082
rect 5884 10030 5894 10082
rect 5894 10030 5940 10082
rect 5964 10030 6010 10082
rect 6010 10030 6020 10082
rect 6044 10030 6074 10082
rect 6074 10030 6100 10082
rect 5804 10028 5860 10030
rect 5884 10028 5940 10030
rect 5964 10028 6020 10030
rect 6044 10028 6100 10030
rect 5804 8994 5860 8996
rect 5884 8994 5940 8996
rect 5964 8994 6020 8996
rect 6044 8994 6100 8996
rect 5804 8942 5830 8994
rect 5830 8942 5860 8994
rect 5884 8942 5894 8994
rect 5894 8942 5940 8994
rect 5964 8942 6010 8994
rect 6010 8942 6020 8994
rect 6044 8942 6074 8994
rect 6074 8942 6100 8994
rect 5804 8940 5860 8942
rect 5884 8940 5940 8942
rect 5964 8940 6020 8942
rect 6044 8940 6100 8942
rect 7283 13890 7339 13892
rect 7363 13890 7419 13892
rect 7443 13890 7499 13892
rect 7523 13890 7579 13892
rect 7283 13838 7309 13890
rect 7309 13838 7339 13890
rect 7363 13838 7373 13890
rect 7373 13838 7419 13890
rect 7443 13838 7489 13890
rect 7489 13838 7499 13890
rect 7523 13838 7553 13890
rect 7553 13838 7579 13890
rect 7283 13836 7339 13838
rect 7363 13836 7419 13838
rect 7443 13836 7499 13838
rect 7523 13836 7579 13838
rect 7283 12802 7339 12804
rect 7363 12802 7419 12804
rect 7443 12802 7499 12804
rect 7523 12802 7579 12804
rect 7283 12750 7309 12802
rect 7309 12750 7339 12802
rect 7363 12750 7373 12802
rect 7373 12750 7419 12802
rect 7443 12750 7489 12802
rect 7489 12750 7499 12802
rect 7523 12750 7553 12802
rect 7553 12750 7579 12802
rect 7283 12748 7339 12750
rect 7363 12748 7419 12750
rect 7443 12748 7499 12750
rect 7523 12748 7579 12750
rect 5804 7906 5860 7908
rect 5884 7906 5940 7908
rect 5964 7906 6020 7908
rect 6044 7906 6100 7908
rect 5804 7854 5830 7906
rect 5830 7854 5860 7906
rect 5884 7854 5894 7906
rect 5894 7854 5940 7906
rect 5964 7854 6010 7906
rect 6010 7854 6020 7906
rect 6044 7854 6074 7906
rect 6074 7854 6100 7906
rect 5804 7852 5860 7854
rect 5884 7852 5940 7854
rect 5964 7852 6020 7854
rect 6044 7852 6100 7854
rect 4326 7362 4382 7364
rect 4406 7362 4462 7364
rect 4486 7362 4542 7364
rect 4566 7362 4622 7364
rect 4326 7310 4352 7362
rect 4352 7310 4382 7362
rect 4406 7310 4416 7362
rect 4416 7310 4462 7362
rect 4486 7310 4532 7362
rect 4532 7310 4542 7362
rect 4566 7310 4596 7362
rect 4596 7310 4622 7362
rect 4326 7308 4382 7310
rect 4406 7308 4462 7310
rect 4486 7308 4542 7310
rect 4566 7308 4622 7310
rect 4326 6274 4382 6276
rect 4406 6274 4462 6276
rect 4486 6274 4542 6276
rect 4566 6274 4622 6276
rect 4326 6222 4352 6274
rect 4352 6222 4382 6274
rect 4406 6222 4416 6274
rect 4416 6222 4462 6274
rect 4486 6222 4532 6274
rect 4532 6222 4542 6274
rect 4566 6222 4596 6274
rect 4596 6222 4622 6274
rect 4326 6220 4382 6222
rect 4406 6220 4462 6222
rect 4486 6220 4542 6222
rect 4566 6220 4622 6222
rect 4326 5186 4382 5188
rect 4406 5186 4462 5188
rect 4486 5186 4542 5188
rect 4566 5186 4622 5188
rect 4326 5134 4352 5186
rect 4352 5134 4382 5186
rect 4406 5134 4416 5186
rect 4416 5134 4462 5186
rect 4486 5134 4532 5186
rect 4532 5134 4542 5186
rect 4566 5134 4596 5186
rect 4596 5134 4622 5186
rect 4326 5132 4382 5134
rect 4406 5132 4462 5134
rect 4486 5132 4542 5134
rect 4566 5132 4622 5134
rect 4326 4098 4382 4100
rect 4406 4098 4462 4100
rect 4486 4098 4542 4100
rect 4566 4098 4622 4100
rect 4326 4046 4352 4098
rect 4352 4046 4382 4098
rect 4406 4046 4416 4098
rect 4416 4046 4462 4098
rect 4486 4046 4532 4098
rect 4532 4046 4542 4098
rect 4566 4046 4596 4098
rect 4596 4046 4622 4098
rect 4326 4044 4382 4046
rect 4406 4044 4462 4046
rect 4486 4044 4542 4046
rect 4566 4044 4622 4046
rect 2847 3554 2903 3556
rect 2927 3554 2983 3556
rect 3007 3554 3063 3556
rect 3087 3554 3143 3556
rect 2847 3502 2873 3554
rect 2873 3502 2903 3554
rect 2927 3502 2937 3554
rect 2937 3502 2983 3554
rect 3007 3502 3053 3554
rect 3053 3502 3063 3554
rect 3087 3502 3117 3554
rect 3117 3502 3143 3554
rect 2847 3500 2903 3502
rect 2927 3500 2983 3502
rect 3007 3500 3063 3502
rect 3087 3500 3143 3502
rect 1368 3010 1424 3012
rect 1448 3010 1504 3012
rect 1528 3010 1584 3012
rect 1608 3010 1664 3012
rect 1368 2958 1394 3010
rect 1394 2958 1424 3010
rect 1448 2958 1458 3010
rect 1458 2958 1504 3010
rect 1528 2958 1574 3010
rect 1574 2958 1584 3010
rect 1608 2958 1638 3010
rect 1638 2958 1664 3010
rect 1368 2956 1424 2958
rect 1448 2956 1504 2958
rect 1528 2956 1584 2958
rect 1608 2956 1664 2958
rect 4326 3010 4382 3012
rect 4406 3010 4462 3012
rect 4486 3010 4542 3012
rect 4566 3010 4622 3012
rect 4326 2958 4352 3010
rect 4352 2958 4382 3010
rect 4406 2958 4416 3010
rect 4416 2958 4462 3010
rect 4486 2958 4532 3010
rect 4532 2958 4542 3010
rect 4566 2958 4596 3010
rect 4596 2958 4622 3010
rect 4326 2956 4382 2958
rect 4406 2956 4462 2958
rect 4486 2956 4542 2958
rect 4566 2956 4622 2958
rect 2847 2466 2903 2468
rect 2927 2466 2983 2468
rect 3007 2466 3063 2468
rect 3087 2466 3143 2468
rect 2847 2414 2873 2466
rect 2873 2414 2903 2466
rect 2927 2414 2937 2466
rect 2937 2414 2983 2466
rect 3007 2414 3053 2466
rect 3053 2414 3063 2466
rect 3087 2414 3117 2466
rect 3117 2414 3143 2466
rect 2847 2412 2903 2414
rect 2927 2412 2983 2414
rect 3007 2412 3063 2414
rect 3087 2412 3143 2414
rect 5804 6818 5860 6820
rect 5884 6818 5940 6820
rect 5964 6818 6020 6820
rect 6044 6818 6100 6820
rect 5804 6766 5830 6818
rect 5830 6766 5860 6818
rect 5884 6766 5894 6818
rect 5894 6766 5940 6818
rect 5964 6766 6010 6818
rect 6010 6766 6020 6818
rect 6044 6766 6074 6818
rect 6074 6766 6100 6818
rect 5804 6764 5860 6766
rect 5884 6764 5940 6766
rect 5964 6764 6020 6766
rect 6044 6764 6100 6766
rect 5804 5730 5860 5732
rect 5884 5730 5940 5732
rect 5964 5730 6020 5732
rect 6044 5730 6100 5732
rect 5804 5678 5830 5730
rect 5830 5678 5860 5730
rect 5884 5678 5894 5730
rect 5894 5678 5940 5730
rect 5964 5678 6010 5730
rect 6010 5678 6020 5730
rect 6044 5678 6074 5730
rect 6074 5678 6100 5730
rect 5804 5676 5860 5678
rect 5884 5676 5940 5678
rect 5964 5676 6020 5678
rect 6044 5676 6100 5678
rect 5804 4642 5860 4644
rect 5884 4642 5940 4644
rect 5964 4642 6020 4644
rect 6044 4642 6100 4644
rect 5804 4590 5830 4642
rect 5830 4590 5860 4642
rect 5884 4590 5894 4642
rect 5894 4590 5940 4642
rect 5964 4590 6010 4642
rect 6010 4590 6020 4642
rect 6044 4590 6074 4642
rect 6074 4590 6100 4642
rect 5804 4588 5860 4590
rect 5884 4588 5940 4590
rect 5964 4588 6020 4590
rect 6044 4588 6100 4590
rect 5804 3554 5860 3556
rect 5884 3554 5940 3556
rect 5964 3554 6020 3556
rect 6044 3554 6100 3556
rect 5804 3502 5830 3554
rect 5830 3502 5860 3554
rect 5884 3502 5894 3554
rect 5894 3502 5940 3554
rect 5964 3502 6010 3554
rect 6010 3502 6020 3554
rect 6044 3502 6074 3554
rect 6074 3502 6100 3554
rect 5804 3500 5860 3502
rect 5884 3500 5940 3502
rect 5964 3500 6020 3502
rect 6044 3500 6100 3502
rect 7283 11714 7339 11716
rect 7363 11714 7419 11716
rect 7443 11714 7499 11716
rect 7523 11714 7579 11716
rect 7283 11662 7309 11714
rect 7309 11662 7339 11714
rect 7363 11662 7373 11714
rect 7373 11662 7419 11714
rect 7443 11662 7489 11714
rect 7489 11662 7499 11714
rect 7523 11662 7553 11714
rect 7553 11662 7579 11714
rect 7283 11660 7339 11662
rect 7363 11660 7419 11662
rect 7443 11660 7499 11662
rect 7523 11660 7579 11662
rect 7283 10626 7339 10628
rect 7363 10626 7419 10628
rect 7443 10626 7499 10628
rect 7523 10626 7579 10628
rect 7283 10574 7309 10626
rect 7309 10574 7339 10626
rect 7363 10574 7373 10626
rect 7373 10574 7419 10626
rect 7443 10574 7489 10626
rect 7489 10574 7499 10626
rect 7523 10574 7553 10626
rect 7553 10574 7579 10626
rect 7283 10572 7339 10574
rect 7363 10572 7419 10574
rect 7443 10572 7499 10574
rect 7523 10572 7579 10574
rect 9256 15808 9312 15864
rect 7283 9538 7339 9540
rect 7363 9538 7419 9540
rect 7443 9538 7499 9540
rect 7523 9538 7579 9540
rect 7283 9486 7309 9538
rect 7309 9486 7339 9538
rect 7363 9486 7373 9538
rect 7373 9486 7419 9538
rect 7443 9486 7489 9538
rect 7489 9486 7499 9538
rect 7523 9486 7553 9538
rect 7553 9486 7579 9538
rect 7283 9484 7339 9486
rect 7363 9484 7419 9486
rect 7443 9484 7499 9486
rect 7523 9484 7579 9486
rect 7283 8450 7339 8452
rect 7363 8450 7419 8452
rect 7443 8450 7499 8452
rect 7523 8450 7579 8452
rect 7283 8398 7309 8450
rect 7309 8398 7339 8450
rect 7363 8398 7373 8450
rect 7373 8398 7419 8450
rect 7443 8398 7489 8450
rect 7489 8398 7499 8450
rect 7523 8398 7553 8450
rect 7553 8398 7579 8450
rect 7283 8396 7339 8398
rect 7363 8396 7419 8398
rect 7443 8396 7499 8398
rect 7523 8396 7579 8398
rect 7283 7362 7339 7364
rect 7363 7362 7419 7364
rect 7443 7362 7499 7364
rect 7523 7362 7579 7364
rect 7283 7310 7309 7362
rect 7309 7310 7339 7362
rect 7363 7310 7373 7362
rect 7373 7310 7419 7362
rect 7443 7310 7489 7362
rect 7489 7310 7499 7362
rect 7523 7310 7553 7362
rect 7553 7310 7579 7362
rect 7283 7308 7339 7310
rect 7363 7308 7419 7310
rect 7443 7308 7499 7310
rect 7523 7308 7579 7310
rect 7283 6274 7339 6276
rect 7363 6274 7419 6276
rect 7443 6274 7499 6276
rect 7523 6274 7579 6276
rect 7283 6222 7309 6274
rect 7309 6222 7339 6274
rect 7363 6222 7373 6274
rect 7373 6222 7419 6274
rect 7443 6222 7489 6274
rect 7489 6222 7499 6274
rect 7523 6222 7553 6274
rect 7553 6222 7579 6274
rect 7283 6220 7339 6222
rect 7363 6220 7419 6222
rect 7443 6220 7499 6222
rect 7523 6220 7579 6222
rect 7283 5186 7339 5188
rect 7363 5186 7419 5188
rect 7443 5186 7499 5188
rect 7523 5186 7579 5188
rect 7283 5134 7309 5186
rect 7309 5134 7339 5186
rect 7363 5134 7373 5186
rect 7373 5134 7419 5186
rect 7443 5134 7489 5186
rect 7489 5134 7499 5186
rect 7523 5134 7553 5186
rect 7553 5134 7579 5186
rect 7283 5132 7339 5134
rect 7363 5132 7419 5134
rect 7443 5132 7499 5134
rect 7523 5132 7579 5134
rect 7283 4098 7339 4100
rect 7363 4098 7419 4100
rect 7443 4098 7499 4100
rect 7523 4098 7579 4100
rect 7283 4046 7309 4098
rect 7309 4046 7339 4098
rect 7363 4046 7373 4098
rect 7373 4046 7419 4098
rect 7443 4046 7489 4098
rect 7489 4046 7499 4098
rect 7523 4046 7553 4098
rect 7553 4046 7579 4098
rect 7283 4044 7339 4046
rect 7363 4044 7419 4046
rect 7443 4044 7499 4046
rect 7523 4044 7579 4046
rect 7283 3010 7339 3012
rect 7363 3010 7419 3012
rect 7443 3010 7499 3012
rect 7523 3010 7579 3012
rect 7283 2958 7309 3010
rect 7309 2958 7339 3010
rect 7363 2958 7373 3010
rect 7373 2958 7419 3010
rect 7443 2958 7489 3010
rect 7489 2958 7499 3010
rect 7523 2958 7553 3010
rect 7553 2958 7579 3010
rect 7283 2956 7339 2958
rect 7363 2956 7419 2958
rect 7443 2956 7499 2958
rect 7523 2956 7579 2958
rect 5804 2466 5860 2468
rect 5884 2466 5940 2468
rect 5964 2466 6020 2468
rect 6044 2466 6100 2468
rect 5804 2414 5830 2466
rect 5830 2414 5860 2466
rect 5884 2414 5894 2466
rect 5894 2414 5940 2466
rect 5964 2414 6010 2466
rect 6010 2414 6020 2466
rect 6044 2414 6074 2466
rect 6074 2414 6100 2466
rect 5804 2412 5860 2414
rect 5884 2412 5940 2414
rect 5964 2412 6020 2414
rect 6044 2412 6100 2414
rect 15696 14992 15752 15048
rect 15512 13496 15568 13552
rect 15604 12680 15660 12736
rect 11464 11864 11520 11920
rect 8704 11048 8760 11104
rect 15972 14312 16028 14368
rect 11648 10232 11704 10288
rect 11556 9552 11612 9608
rect 11372 8772 11374 8792
rect 11374 8772 11426 8792
rect 11426 8772 11428 8792
rect 8336 8192 8392 8248
rect 11372 8736 11428 8772
rect 11372 7920 11428 7976
rect 11464 7104 11520 7160
rect 11372 6288 11428 6344
rect 11464 5472 11520 5528
rect 11372 4792 11428 4848
rect 11556 3976 11612 4032
rect 11372 3160 11428 3216
rect 15512 2344 15568 2400
rect 1368 1922 1424 1924
rect 1448 1922 1504 1924
rect 1528 1922 1584 1924
rect 1608 1922 1664 1924
rect 1368 1870 1394 1922
rect 1394 1870 1424 1922
rect 1448 1870 1458 1922
rect 1458 1870 1504 1922
rect 1528 1870 1574 1922
rect 1574 1870 1584 1922
rect 1608 1870 1638 1922
rect 1638 1870 1664 1922
rect 1368 1868 1424 1870
rect 1448 1868 1504 1870
rect 1528 1868 1584 1870
rect 1608 1868 1664 1870
rect 4326 1922 4382 1924
rect 4406 1922 4462 1924
rect 4486 1922 4542 1924
rect 4566 1922 4622 1924
rect 4326 1870 4352 1922
rect 4352 1870 4382 1922
rect 4406 1870 4416 1922
rect 4416 1870 4462 1922
rect 4486 1870 4532 1922
rect 4532 1870 4542 1922
rect 4566 1870 4596 1922
rect 4596 1870 4622 1922
rect 4326 1868 4382 1870
rect 4406 1868 4462 1870
rect 4486 1868 4542 1870
rect 4566 1868 4622 1870
rect 7283 1922 7339 1924
rect 7363 1922 7419 1924
rect 7443 1922 7499 1924
rect 7523 1922 7579 1924
rect 7283 1870 7309 1922
rect 7309 1870 7339 1922
rect 7363 1870 7373 1922
rect 7373 1870 7419 1922
rect 7443 1870 7489 1922
rect 7489 1870 7499 1922
rect 7523 1870 7553 1922
rect 7553 1870 7579 1922
rect 7283 1868 7339 1870
rect 7363 1868 7419 1870
rect 7443 1868 7499 1870
rect 7523 1868 7579 1870
rect 15604 1528 15660 1584
rect 23792 712 23848 768
rect 15696 32 15752 88
<< metal3 >>
rect 9934 18312 33934 18344
rect 9934 18256 24068 18312
rect 24124 18256 33934 18312
rect 9934 18224 33934 18256
rect 9934 17496 33934 17528
rect 9934 17440 23792 17496
rect 23848 17440 33934 17496
rect 9934 17408 33934 17440
rect 9934 16680 33934 16712
rect 9934 16624 15512 16680
rect 15568 16624 33934 16680
rect 9934 16592 33934 16624
rect 1356 16072 1676 16073
rect 1356 16008 1364 16072
rect 1428 16008 1444 16072
rect 1508 16008 1524 16072
rect 1588 16008 1604 16072
rect 1668 16008 1676 16072
rect 1356 16007 1676 16008
rect 4314 16072 4634 16073
rect 4314 16008 4322 16072
rect 4386 16008 4402 16072
rect 4466 16008 4482 16072
rect 4546 16008 4562 16072
rect 4626 16008 4634 16072
rect 4314 16007 4634 16008
rect 7271 16072 7591 16073
rect 7271 16008 7279 16072
rect 7343 16008 7359 16072
rect 7423 16008 7439 16072
rect 7503 16008 7519 16072
rect 7583 16008 7591 16072
rect 7271 16007 7591 16008
rect 9251 15866 9317 15869
rect 9934 15866 33934 15896
rect 9251 15864 33934 15866
rect 9251 15808 9256 15864
rect 9312 15808 33934 15864
rect 9251 15806 33934 15808
rect 9251 15803 9317 15806
rect 9934 15776 33934 15806
rect 2835 15528 3155 15529
rect 2835 15464 2843 15528
rect 2907 15464 2923 15528
rect 2987 15464 3003 15528
rect 3067 15464 3083 15528
rect 3147 15464 3155 15528
rect 2835 15463 3155 15464
rect 5792 15528 6112 15529
rect 5792 15464 5800 15528
rect 5864 15464 5880 15528
rect 5944 15464 5960 15528
rect 6024 15464 6040 15528
rect 6104 15464 6112 15528
rect 5792 15463 6112 15464
rect 9934 15048 33934 15080
rect 9934 14992 15696 15048
rect 15752 14992 33934 15048
rect 1356 14984 1676 14985
rect 1356 14920 1364 14984
rect 1428 14920 1444 14984
rect 1508 14920 1524 14984
rect 1588 14920 1604 14984
rect 1668 14920 1676 14984
rect 1356 14919 1676 14920
rect 4314 14984 4634 14985
rect 4314 14920 4322 14984
rect 4386 14920 4402 14984
rect 4466 14920 4482 14984
rect 4546 14920 4562 14984
rect 4626 14920 4634 14984
rect 4314 14919 4634 14920
rect 7271 14984 7591 14985
rect 7271 14920 7279 14984
rect 7343 14920 7359 14984
rect 7423 14920 7439 14984
rect 7503 14920 7519 14984
rect 7583 14920 7591 14984
rect 9934 14960 33934 14992
rect 7271 14919 7591 14920
rect 2835 14440 3155 14441
rect 2835 14376 2843 14440
rect 2907 14376 2923 14440
rect 2987 14376 3003 14440
rect 3067 14376 3083 14440
rect 3147 14376 3155 14440
rect 2835 14375 3155 14376
rect 5792 14440 6112 14441
rect 5792 14376 5800 14440
rect 5864 14376 5880 14440
rect 5944 14376 5960 14440
rect 6024 14376 6040 14440
rect 6104 14376 6112 14440
rect 5792 14375 6112 14376
rect 9934 14368 33934 14400
rect 9934 14312 15972 14368
rect 16028 14312 33934 14368
rect 9934 14280 33934 14312
rect 1356 13896 1676 13897
rect 1356 13832 1364 13896
rect 1428 13832 1444 13896
rect 1508 13832 1524 13896
rect 1588 13832 1604 13896
rect 1668 13832 1676 13896
rect 1356 13831 1676 13832
rect 4314 13896 4634 13897
rect 4314 13832 4322 13896
rect 4386 13832 4402 13896
rect 4466 13832 4482 13896
rect 4546 13832 4562 13896
rect 4626 13832 4634 13896
rect 4314 13831 4634 13832
rect 7271 13896 7591 13897
rect 7271 13832 7279 13896
rect 7343 13832 7359 13896
rect 7423 13832 7439 13896
rect 7503 13832 7519 13896
rect 7583 13832 7591 13896
rect 7271 13831 7591 13832
rect 9934 13552 33934 13584
rect 9934 13496 15512 13552
rect 15568 13496 33934 13552
rect 9934 13464 33934 13496
rect 2835 13352 3155 13353
rect 2835 13288 2843 13352
rect 2907 13288 2923 13352
rect 2987 13288 3003 13352
rect 3067 13288 3083 13352
rect 3147 13288 3155 13352
rect 2835 13287 3155 13288
rect 5792 13352 6112 13353
rect 5792 13288 5800 13352
rect 5864 13288 5880 13352
rect 5944 13288 5960 13352
rect 6024 13288 6040 13352
rect 6104 13288 6112 13352
rect 5792 13287 6112 13288
rect 1356 12808 1676 12809
rect 1356 12744 1364 12808
rect 1428 12744 1444 12808
rect 1508 12744 1524 12808
rect 1588 12744 1604 12808
rect 1668 12744 1676 12808
rect 1356 12743 1676 12744
rect 4314 12808 4634 12809
rect 4314 12744 4322 12808
rect 4386 12744 4402 12808
rect 4466 12744 4482 12808
rect 4546 12744 4562 12808
rect 4626 12744 4634 12808
rect 4314 12743 4634 12744
rect 7271 12808 7591 12809
rect 7271 12744 7279 12808
rect 7343 12744 7359 12808
rect 7423 12744 7439 12808
rect 7503 12744 7519 12808
rect 7583 12744 7591 12808
rect 7271 12743 7591 12744
rect 9934 12736 33934 12768
rect 9934 12680 15604 12736
rect 15660 12680 33934 12736
rect 9934 12648 33934 12680
rect 2835 12264 3155 12265
rect 2835 12200 2843 12264
rect 2907 12200 2923 12264
rect 2987 12200 3003 12264
rect 3067 12200 3083 12264
rect 3147 12200 3155 12264
rect 2835 12199 3155 12200
rect 5792 12264 6112 12265
rect 5792 12200 5800 12264
rect 5864 12200 5880 12264
rect 5944 12200 5960 12264
rect 6024 12200 6040 12264
rect 6104 12200 6112 12264
rect 5792 12199 6112 12200
rect 9934 11920 33934 11952
rect 9934 11864 11464 11920
rect 11520 11864 33934 11920
rect 9934 11832 33934 11864
rect 1356 11720 1676 11721
rect 1356 11656 1364 11720
rect 1428 11656 1444 11720
rect 1508 11656 1524 11720
rect 1588 11656 1604 11720
rect 1668 11656 1676 11720
rect 1356 11655 1676 11656
rect 4314 11720 4634 11721
rect 4314 11656 4322 11720
rect 4386 11656 4402 11720
rect 4466 11656 4482 11720
rect 4546 11656 4562 11720
rect 4626 11656 4634 11720
rect 4314 11655 4634 11656
rect 7271 11720 7591 11721
rect 7271 11656 7279 11720
rect 7343 11656 7359 11720
rect 7423 11656 7439 11720
rect 7503 11656 7519 11720
rect 7583 11656 7591 11720
rect 7271 11655 7591 11656
rect 2835 11176 3155 11177
rect 2835 11112 2843 11176
rect 2907 11112 2923 11176
rect 2987 11112 3003 11176
rect 3067 11112 3083 11176
rect 3147 11112 3155 11176
rect 2835 11111 3155 11112
rect 5792 11176 6112 11177
rect 5792 11112 5800 11176
rect 5864 11112 5880 11176
rect 5944 11112 5960 11176
rect 6024 11112 6040 11176
rect 6104 11112 6112 11176
rect 5792 11111 6112 11112
rect 8699 11106 8765 11109
rect 9934 11106 33934 11136
rect 8699 11104 33934 11106
rect 8699 11048 8704 11104
rect 8760 11048 33934 11104
rect 8699 11046 33934 11048
rect 8699 11043 8765 11046
rect 9934 11016 33934 11046
rect 1356 10632 1676 10633
rect 1356 10568 1364 10632
rect 1428 10568 1444 10632
rect 1508 10568 1524 10632
rect 1588 10568 1604 10632
rect 1668 10568 1676 10632
rect 1356 10567 1676 10568
rect 4314 10632 4634 10633
rect 4314 10568 4322 10632
rect 4386 10568 4402 10632
rect 4466 10568 4482 10632
rect 4546 10568 4562 10632
rect 4626 10568 4634 10632
rect 4314 10567 4634 10568
rect 7271 10632 7591 10633
rect 7271 10568 7279 10632
rect 7343 10568 7359 10632
rect 7423 10568 7439 10632
rect 7503 10568 7519 10632
rect 7583 10568 7591 10632
rect 7271 10567 7591 10568
rect 2075 10290 2141 10293
rect 5571 10290 5637 10293
rect 2075 10288 5637 10290
rect 2075 10232 2080 10288
rect 2136 10232 5576 10288
rect 5632 10232 5637 10288
rect 2075 10230 5637 10232
rect 2075 10227 2141 10230
rect 5571 10227 5637 10230
rect 9934 10288 33934 10320
rect 9934 10232 11648 10288
rect 11704 10232 33934 10288
rect 9934 10200 33934 10232
rect 2835 10088 3155 10089
rect 2835 10024 2843 10088
rect 2907 10024 2923 10088
rect 2987 10024 3003 10088
rect 3067 10024 3083 10088
rect 3147 10024 3155 10088
rect 2835 10023 3155 10024
rect 5792 10088 6112 10089
rect 5792 10024 5800 10088
rect 5864 10024 5880 10088
rect 5944 10024 5960 10088
rect 6024 10024 6040 10088
rect 6104 10024 6112 10088
rect 5792 10023 6112 10024
rect 9934 9608 33934 9640
rect 9934 9552 11556 9608
rect 11612 9552 33934 9608
rect 1356 9544 1676 9545
rect 1356 9480 1364 9544
rect 1428 9480 1444 9544
rect 1508 9480 1524 9544
rect 1588 9480 1604 9544
rect 1668 9480 1676 9544
rect 1356 9479 1676 9480
rect 4314 9544 4634 9545
rect 4314 9480 4322 9544
rect 4386 9480 4402 9544
rect 4466 9480 4482 9544
rect 4546 9480 4562 9544
rect 4626 9480 4634 9544
rect 4314 9479 4634 9480
rect 7271 9544 7591 9545
rect 7271 9480 7279 9544
rect 7343 9480 7359 9544
rect 7423 9480 7439 9544
rect 7503 9480 7519 9544
rect 7583 9480 7591 9544
rect 9934 9520 33934 9552
rect 7271 9479 7591 9480
rect 2835 9000 3155 9001
rect 2835 8936 2843 9000
rect 2907 8936 2923 9000
rect 2987 8936 3003 9000
rect 3067 8936 3083 9000
rect 3147 8936 3155 9000
rect 2835 8935 3155 8936
rect 5792 9000 6112 9001
rect 5792 8936 5800 9000
rect 5864 8936 5880 9000
rect 5944 8936 5960 9000
rect 6024 8936 6040 9000
rect 6104 8936 6112 9000
rect 5792 8935 6112 8936
rect 9934 8792 33934 8824
rect 9934 8736 11372 8792
rect 11428 8736 33934 8792
rect 9934 8704 33934 8736
rect 1356 8456 1676 8457
rect 1356 8392 1364 8456
rect 1428 8392 1444 8456
rect 1508 8392 1524 8456
rect 1588 8392 1604 8456
rect 1668 8392 1676 8456
rect 1356 8391 1676 8392
rect 4314 8456 4634 8457
rect 4314 8392 4322 8456
rect 4386 8392 4402 8456
rect 4466 8392 4482 8456
rect 4546 8392 4562 8456
rect 4626 8392 4634 8456
rect 4314 8391 4634 8392
rect 7271 8456 7591 8457
rect 7271 8392 7279 8456
rect 7343 8392 7359 8456
rect 7423 8392 7439 8456
rect 7503 8392 7519 8456
rect 7583 8392 7591 8456
rect 7271 8391 7591 8392
rect 3271 8250 3337 8253
rect 8331 8250 8397 8253
rect 3271 8248 8397 8250
rect 3271 8192 3276 8248
rect 3332 8192 8336 8248
rect 8392 8192 8397 8248
rect 3271 8190 8397 8192
rect 3271 8187 3337 8190
rect 8331 8187 8397 8190
rect 9934 7976 33934 8008
rect 9934 7920 11372 7976
rect 11428 7920 33934 7976
rect 2835 7912 3155 7913
rect 2835 7848 2843 7912
rect 2907 7848 2923 7912
rect 2987 7848 3003 7912
rect 3067 7848 3083 7912
rect 3147 7848 3155 7912
rect 2835 7847 3155 7848
rect 5792 7912 6112 7913
rect 5792 7848 5800 7912
rect 5864 7848 5880 7912
rect 5944 7848 5960 7912
rect 6024 7848 6040 7912
rect 6104 7848 6112 7912
rect 9934 7888 33934 7920
rect 5792 7847 6112 7848
rect 1356 7368 1676 7369
rect 1356 7304 1364 7368
rect 1428 7304 1444 7368
rect 1508 7304 1524 7368
rect 1588 7304 1604 7368
rect 1668 7304 1676 7368
rect 1356 7303 1676 7304
rect 4314 7368 4634 7369
rect 4314 7304 4322 7368
rect 4386 7304 4402 7368
rect 4466 7304 4482 7368
rect 4546 7304 4562 7368
rect 4626 7304 4634 7368
rect 4314 7303 4634 7304
rect 7271 7368 7591 7369
rect 7271 7304 7279 7368
rect 7343 7304 7359 7368
rect 7423 7304 7439 7368
rect 7503 7304 7519 7368
rect 7583 7304 7591 7368
rect 7271 7303 7591 7304
rect 9934 7160 33934 7192
rect 9934 7104 11464 7160
rect 11520 7104 33934 7160
rect 9934 7072 33934 7104
rect 2835 6824 3155 6825
rect 2835 6760 2843 6824
rect 2907 6760 2923 6824
rect 2987 6760 3003 6824
rect 3067 6760 3083 6824
rect 3147 6760 3155 6824
rect 2835 6759 3155 6760
rect 5792 6824 6112 6825
rect 5792 6760 5800 6824
rect 5864 6760 5880 6824
rect 5944 6760 5960 6824
rect 6024 6760 6040 6824
rect 6104 6760 6112 6824
rect 5792 6759 6112 6760
rect 9934 6344 33934 6376
rect 9934 6288 11372 6344
rect 11428 6288 33934 6344
rect 1356 6280 1676 6281
rect 1356 6216 1364 6280
rect 1428 6216 1444 6280
rect 1508 6216 1524 6280
rect 1588 6216 1604 6280
rect 1668 6216 1676 6280
rect 1356 6215 1676 6216
rect 4314 6280 4634 6281
rect 4314 6216 4322 6280
rect 4386 6216 4402 6280
rect 4466 6216 4482 6280
rect 4546 6216 4562 6280
rect 4626 6216 4634 6280
rect 4314 6215 4634 6216
rect 7271 6280 7591 6281
rect 7271 6216 7279 6280
rect 7343 6216 7359 6280
rect 7423 6216 7439 6280
rect 7503 6216 7519 6280
rect 7583 6216 7591 6280
rect 9934 6256 33934 6288
rect 7271 6215 7591 6216
rect 2835 5736 3155 5737
rect 2835 5672 2843 5736
rect 2907 5672 2923 5736
rect 2987 5672 3003 5736
rect 3067 5672 3083 5736
rect 3147 5672 3155 5736
rect 2835 5671 3155 5672
rect 5792 5736 6112 5737
rect 5792 5672 5800 5736
rect 5864 5672 5880 5736
rect 5944 5672 5960 5736
rect 6024 5672 6040 5736
rect 6104 5672 6112 5736
rect 5792 5671 6112 5672
rect 9934 5528 33934 5560
rect 9934 5472 11464 5528
rect 11520 5472 33934 5528
rect 9934 5440 33934 5472
rect 1356 5192 1676 5193
rect 1356 5128 1364 5192
rect 1428 5128 1444 5192
rect 1508 5128 1524 5192
rect 1588 5128 1604 5192
rect 1668 5128 1676 5192
rect 1356 5127 1676 5128
rect 4314 5192 4634 5193
rect 4314 5128 4322 5192
rect 4386 5128 4402 5192
rect 4466 5128 4482 5192
rect 4546 5128 4562 5192
rect 4626 5128 4634 5192
rect 4314 5127 4634 5128
rect 7271 5192 7591 5193
rect 7271 5128 7279 5192
rect 7343 5128 7359 5192
rect 7423 5128 7439 5192
rect 7503 5128 7519 5192
rect 7583 5128 7591 5192
rect 7271 5127 7591 5128
rect 9934 4848 33934 4880
rect 9934 4792 11372 4848
rect 11428 4792 33934 4848
rect 9934 4760 33934 4792
rect 2835 4648 3155 4649
rect 2835 4584 2843 4648
rect 2907 4584 2923 4648
rect 2987 4584 3003 4648
rect 3067 4584 3083 4648
rect 3147 4584 3155 4648
rect 2835 4583 3155 4584
rect 5792 4648 6112 4649
rect 5792 4584 5800 4648
rect 5864 4584 5880 4648
rect 5944 4584 5960 4648
rect 6024 4584 6040 4648
rect 6104 4584 6112 4648
rect 5792 4583 6112 4584
rect 1356 4104 1676 4105
rect 1356 4040 1364 4104
rect 1428 4040 1444 4104
rect 1508 4040 1524 4104
rect 1588 4040 1604 4104
rect 1668 4040 1676 4104
rect 1356 4039 1676 4040
rect 4314 4104 4634 4105
rect 4314 4040 4322 4104
rect 4386 4040 4402 4104
rect 4466 4040 4482 4104
rect 4546 4040 4562 4104
rect 4626 4040 4634 4104
rect 4314 4039 4634 4040
rect 7271 4104 7591 4105
rect 7271 4040 7279 4104
rect 7343 4040 7359 4104
rect 7423 4040 7439 4104
rect 7503 4040 7519 4104
rect 7583 4040 7591 4104
rect 7271 4039 7591 4040
rect 9934 4032 33934 4064
rect 9934 3976 11556 4032
rect 11612 3976 33934 4032
rect 9934 3944 33934 3976
rect 2835 3560 3155 3561
rect 2835 3496 2843 3560
rect 2907 3496 2923 3560
rect 2987 3496 3003 3560
rect 3067 3496 3083 3560
rect 3147 3496 3155 3560
rect 2835 3495 3155 3496
rect 5792 3560 6112 3561
rect 5792 3496 5800 3560
rect 5864 3496 5880 3560
rect 5944 3496 5960 3560
rect 6024 3496 6040 3560
rect 6104 3496 6112 3560
rect 5792 3495 6112 3496
rect 9934 3216 33934 3248
rect 9934 3160 11372 3216
rect 11428 3160 33934 3216
rect 9934 3128 33934 3160
rect 1356 3016 1676 3017
rect 1356 2952 1364 3016
rect 1428 2952 1444 3016
rect 1508 2952 1524 3016
rect 1588 2952 1604 3016
rect 1668 2952 1676 3016
rect 1356 2951 1676 2952
rect 4314 3016 4634 3017
rect 4314 2952 4322 3016
rect 4386 2952 4402 3016
rect 4466 2952 4482 3016
rect 4546 2952 4562 3016
rect 4626 2952 4634 3016
rect 4314 2951 4634 2952
rect 7271 3016 7591 3017
rect 7271 2952 7279 3016
rect 7343 2952 7359 3016
rect 7423 2952 7439 3016
rect 7503 2952 7519 3016
rect 7583 2952 7591 3016
rect 7271 2951 7591 2952
rect 2835 2472 3155 2473
rect 2835 2408 2843 2472
rect 2907 2408 2923 2472
rect 2987 2408 3003 2472
rect 3067 2408 3083 2472
rect 3147 2408 3155 2472
rect 2835 2407 3155 2408
rect 5792 2472 6112 2473
rect 5792 2408 5800 2472
rect 5864 2408 5880 2472
rect 5944 2408 5960 2472
rect 6024 2408 6040 2472
rect 6104 2408 6112 2472
rect 5792 2407 6112 2408
rect 9934 2400 33934 2432
rect 9934 2344 15512 2400
rect 15568 2344 33934 2400
rect 9934 2312 33934 2344
rect 1356 1928 1676 1929
rect 1356 1864 1364 1928
rect 1428 1864 1444 1928
rect 1508 1864 1524 1928
rect 1588 1864 1604 1928
rect 1668 1864 1676 1928
rect 1356 1863 1676 1864
rect 4314 1928 4634 1929
rect 4314 1864 4322 1928
rect 4386 1864 4402 1928
rect 4466 1864 4482 1928
rect 4546 1864 4562 1928
rect 4626 1864 4634 1928
rect 4314 1863 4634 1864
rect 7271 1928 7591 1929
rect 7271 1864 7279 1928
rect 7343 1864 7359 1928
rect 7423 1864 7439 1928
rect 7503 1864 7519 1928
rect 7583 1864 7591 1928
rect 7271 1863 7591 1864
rect 9934 1584 33934 1616
rect 9934 1528 15604 1584
rect 15660 1528 33934 1584
rect 9934 1496 33934 1528
rect 9934 768 33934 800
rect 9934 712 23792 768
rect 23848 712 33934 768
rect 9934 680 33934 712
rect 9934 88 33934 120
rect 9934 32 15696 88
rect 15752 32 33934 88
rect 9934 0 33934 32
<< via3 >>
rect 1364 16068 1428 16072
rect 1364 16012 1368 16068
rect 1368 16012 1424 16068
rect 1424 16012 1428 16068
rect 1364 16008 1428 16012
rect 1444 16068 1508 16072
rect 1444 16012 1448 16068
rect 1448 16012 1504 16068
rect 1504 16012 1508 16068
rect 1444 16008 1508 16012
rect 1524 16068 1588 16072
rect 1524 16012 1528 16068
rect 1528 16012 1584 16068
rect 1584 16012 1588 16068
rect 1524 16008 1588 16012
rect 1604 16068 1668 16072
rect 1604 16012 1608 16068
rect 1608 16012 1664 16068
rect 1664 16012 1668 16068
rect 1604 16008 1668 16012
rect 4322 16068 4386 16072
rect 4322 16012 4326 16068
rect 4326 16012 4382 16068
rect 4382 16012 4386 16068
rect 4322 16008 4386 16012
rect 4402 16068 4466 16072
rect 4402 16012 4406 16068
rect 4406 16012 4462 16068
rect 4462 16012 4466 16068
rect 4402 16008 4466 16012
rect 4482 16068 4546 16072
rect 4482 16012 4486 16068
rect 4486 16012 4542 16068
rect 4542 16012 4546 16068
rect 4482 16008 4546 16012
rect 4562 16068 4626 16072
rect 4562 16012 4566 16068
rect 4566 16012 4622 16068
rect 4622 16012 4626 16068
rect 4562 16008 4626 16012
rect 7279 16068 7343 16072
rect 7279 16012 7283 16068
rect 7283 16012 7339 16068
rect 7339 16012 7343 16068
rect 7279 16008 7343 16012
rect 7359 16068 7423 16072
rect 7359 16012 7363 16068
rect 7363 16012 7419 16068
rect 7419 16012 7423 16068
rect 7359 16008 7423 16012
rect 7439 16068 7503 16072
rect 7439 16012 7443 16068
rect 7443 16012 7499 16068
rect 7499 16012 7503 16068
rect 7439 16008 7503 16012
rect 7519 16068 7583 16072
rect 7519 16012 7523 16068
rect 7523 16012 7579 16068
rect 7579 16012 7583 16068
rect 7519 16008 7583 16012
rect 2843 15524 2907 15528
rect 2843 15468 2847 15524
rect 2847 15468 2903 15524
rect 2903 15468 2907 15524
rect 2843 15464 2907 15468
rect 2923 15524 2987 15528
rect 2923 15468 2927 15524
rect 2927 15468 2983 15524
rect 2983 15468 2987 15524
rect 2923 15464 2987 15468
rect 3003 15524 3067 15528
rect 3003 15468 3007 15524
rect 3007 15468 3063 15524
rect 3063 15468 3067 15524
rect 3003 15464 3067 15468
rect 3083 15524 3147 15528
rect 3083 15468 3087 15524
rect 3087 15468 3143 15524
rect 3143 15468 3147 15524
rect 3083 15464 3147 15468
rect 5800 15524 5864 15528
rect 5800 15468 5804 15524
rect 5804 15468 5860 15524
rect 5860 15468 5864 15524
rect 5800 15464 5864 15468
rect 5880 15524 5944 15528
rect 5880 15468 5884 15524
rect 5884 15468 5940 15524
rect 5940 15468 5944 15524
rect 5880 15464 5944 15468
rect 5960 15524 6024 15528
rect 5960 15468 5964 15524
rect 5964 15468 6020 15524
rect 6020 15468 6024 15524
rect 5960 15464 6024 15468
rect 6040 15524 6104 15528
rect 6040 15468 6044 15524
rect 6044 15468 6100 15524
rect 6100 15468 6104 15524
rect 6040 15464 6104 15468
rect 1364 14980 1428 14984
rect 1364 14924 1368 14980
rect 1368 14924 1424 14980
rect 1424 14924 1428 14980
rect 1364 14920 1428 14924
rect 1444 14980 1508 14984
rect 1444 14924 1448 14980
rect 1448 14924 1504 14980
rect 1504 14924 1508 14980
rect 1444 14920 1508 14924
rect 1524 14980 1588 14984
rect 1524 14924 1528 14980
rect 1528 14924 1584 14980
rect 1584 14924 1588 14980
rect 1524 14920 1588 14924
rect 1604 14980 1668 14984
rect 1604 14924 1608 14980
rect 1608 14924 1664 14980
rect 1664 14924 1668 14980
rect 1604 14920 1668 14924
rect 4322 14980 4386 14984
rect 4322 14924 4326 14980
rect 4326 14924 4382 14980
rect 4382 14924 4386 14980
rect 4322 14920 4386 14924
rect 4402 14980 4466 14984
rect 4402 14924 4406 14980
rect 4406 14924 4462 14980
rect 4462 14924 4466 14980
rect 4402 14920 4466 14924
rect 4482 14980 4546 14984
rect 4482 14924 4486 14980
rect 4486 14924 4542 14980
rect 4542 14924 4546 14980
rect 4482 14920 4546 14924
rect 4562 14980 4626 14984
rect 4562 14924 4566 14980
rect 4566 14924 4622 14980
rect 4622 14924 4626 14980
rect 4562 14920 4626 14924
rect 7279 14980 7343 14984
rect 7279 14924 7283 14980
rect 7283 14924 7339 14980
rect 7339 14924 7343 14980
rect 7279 14920 7343 14924
rect 7359 14980 7423 14984
rect 7359 14924 7363 14980
rect 7363 14924 7419 14980
rect 7419 14924 7423 14980
rect 7359 14920 7423 14924
rect 7439 14980 7503 14984
rect 7439 14924 7443 14980
rect 7443 14924 7499 14980
rect 7499 14924 7503 14980
rect 7439 14920 7503 14924
rect 7519 14980 7583 14984
rect 7519 14924 7523 14980
rect 7523 14924 7579 14980
rect 7579 14924 7583 14980
rect 7519 14920 7583 14924
rect 2843 14436 2907 14440
rect 2843 14380 2847 14436
rect 2847 14380 2903 14436
rect 2903 14380 2907 14436
rect 2843 14376 2907 14380
rect 2923 14436 2987 14440
rect 2923 14380 2927 14436
rect 2927 14380 2983 14436
rect 2983 14380 2987 14436
rect 2923 14376 2987 14380
rect 3003 14436 3067 14440
rect 3003 14380 3007 14436
rect 3007 14380 3063 14436
rect 3063 14380 3067 14436
rect 3003 14376 3067 14380
rect 3083 14436 3147 14440
rect 3083 14380 3087 14436
rect 3087 14380 3143 14436
rect 3143 14380 3147 14436
rect 3083 14376 3147 14380
rect 5800 14436 5864 14440
rect 5800 14380 5804 14436
rect 5804 14380 5860 14436
rect 5860 14380 5864 14436
rect 5800 14376 5864 14380
rect 5880 14436 5944 14440
rect 5880 14380 5884 14436
rect 5884 14380 5940 14436
rect 5940 14380 5944 14436
rect 5880 14376 5944 14380
rect 5960 14436 6024 14440
rect 5960 14380 5964 14436
rect 5964 14380 6020 14436
rect 6020 14380 6024 14436
rect 5960 14376 6024 14380
rect 6040 14436 6104 14440
rect 6040 14380 6044 14436
rect 6044 14380 6100 14436
rect 6100 14380 6104 14436
rect 6040 14376 6104 14380
rect 1364 13892 1428 13896
rect 1364 13836 1368 13892
rect 1368 13836 1424 13892
rect 1424 13836 1428 13892
rect 1364 13832 1428 13836
rect 1444 13892 1508 13896
rect 1444 13836 1448 13892
rect 1448 13836 1504 13892
rect 1504 13836 1508 13892
rect 1444 13832 1508 13836
rect 1524 13892 1588 13896
rect 1524 13836 1528 13892
rect 1528 13836 1584 13892
rect 1584 13836 1588 13892
rect 1524 13832 1588 13836
rect 1604 13892 1668 13896
rect 1604 13836 1608 13892
rect 1608 13836 1664 13892
rect 1664 13836 1668 13892
rect 1604 13832 1668 13836
rect 4322 13892 4386 13896
rect 4322 13836 4326 13892
rect 4326 13836 4382 13892
rect 4382 13836 4386 13892
rect 4322 13832 4386 13836
rect 4402 13892 4466 13896
rect 4402 13836 4406 13892
rect 4406 13836 4462 13892
rect 4462 13836 4466 13892
rect 4402 13832 4466 13836
rect 4482 13892 4546 13896
rect 4482 13836 4486 13892
rect 4486 13836 4542 13892
rect 4542 13836 4546 13892
rect 4482 13832 4546 13836
rect 4562 13892 4626 13896
rect 4562 13836 4566 13892
rect 4566 13836 4622 13892
rect 4622 13836 4626 13892
rect 4562 13832 4626 13836
rect 7279 13892 7343 13896
rect 7279 13836 7283 13892
rect 7283 13836 7339 13892
rect 7339 13836 7343 13892
rect 7279 13832 7343 13836
rect 7359 13892 7423 13896
rect 7359 13836 7363 13892
rect 7363 13836 7419 13892
rect 7419 13836 7423 13892
rect 7359 13832 7423 13836
rect 7439 13892 7503 13896
rect 7439 13836 7443 13892
rect 7443 13836 7499 13892
rect 7499 13836 7503 13892
rect 7439 13832 7503 13836
rect 7519 13892 7583 13896
rect 7519 13836 7523 13892
rect 7523 13836 7579 13892
rect 7579 13836 7583 13892
rect 7519 13832 7583 13836
rect 2843 13348 2907 13352
rect 2843 13292 2847 13348
rect 2847 13292 2903 13348
rect 2903 13292 2907 13348
rect 2843 13288 2907 13292
rect 2923 13348 2987 13352
rect 2923 13292 2927 13348
rect 2927 13292 2983 13348
rect 2983 13292 2987 13348
rect 2923 13288 2987 13292
rect 3003 13348 3067 13352
rect 3003 13292 3007 13348
rect 3007 13292 3063 13348
rect 3063 13292 3067 13348
rect 3003 13288 3067 13292
rect 3083 13348 3147 13352
rect 3083 13292 3087 13348
rect 3087 13292 3143 13348
rect 3143 13292 3147 13348
rect 3083 13288 3147 13292
rect 5800 13348 5864 13352
rect 5800 13292 5804 13348
rect 5804 13292 5860 13348
rect 5860 13292 5864 13348
rect 5800 13288 5864 13292
rect 5880 13348 5944 13352
rect 5880 13292 5884 13348
rect 5884 13292 5940 13348
rect 5940 13292 5944 13348
rect 5880 13288 5944 13292
rect 5960 13348 6024 13352
rect 5960 13292 5964 13348
rect 5964 13292 6020 13348
rect 6020 13292 6024 13348
rect 5960 13288 6024 13292
rect 6040 13348 6104 13352
rect 6040 13292 6044 13348
rect 6044 13292 6100 13348
rect 6100 13292 6104 13348
rect 6040 13288 6104 13292
rect 1364 12804 1428 12808
rect 1364 12748 1368 12804
rect 1368 12748 1424 12804
rect 1424 12748 1428 12804
rect 1364 12744 1428 12748
rect 1444 12804 1508 12808
rect 1444 12748 1448 12804
rect 1448 12748 1504 12804
rect 1504 12748 1508 12804
rect 1444 12744 1508 12748
rect 1524 12804 1588 12808
rect 1524 12748 1528 12804
rect 1528 12748 1584 12804
rect 1584 12748 1588 12804
rect 1524 12744 1588 12748
rect 1604 12804 1668 12808
rect 1604 12748 1608 12804
rect 1608 12748 1664 12804
rect 1664 12748 1668 12804
rect 1604 12744 1668 12748
rect 4322 12804 4386 12808
rect 4322 12748 4326 12804
rect 4326 12748 4382 12804
rect 4382 12748 4386 12804
rect 4322 12744 4386 12748
rect 4402 12804 4466 12808
rect 4402 12748 4406 12804
rect 4406 12748 4462 12804
rect 4462 12748 4466 12804
rect 4402 12744 4466 12748
rect 4482 12804 4546 12808
rect 4482 12748 4486 12804
rect 4486 12748 4542 12804
rect 4542 12748 4546 12804
rect 4482 12744 4546 12748
rect 4562 12804 4626 12808
rect 4562 12748 4566 12804
rect 4566 12748 4622 12804
rect 4622 12748 4626 12804
rect 4562 12744 4626 12748
rect 7279 12804 7343 12808
rect 7279 12748 7283 12804
rect 7283 12748 7339 12804
rect 7339 12748 7343 12804
rect 7279 12744 7343 12748
rect 7359 12804 7423 12808
rect 7359 12748 7363 12804
rect 7363 12748 7419 12804
rect 7419 12748 7423 12804
rect 7359 12744 7423 12748
rect 7439 12804 7503 12808
rect 7439 12748 7443 12804
rect 7443 12748 7499 12804
rect 7499 12748 7503 12804
rect 7439 12744 7503 12748
rect 7519 12804 7583 12808
rect 7519 12748 7523 12804
rect 7523 12748 7579 12804
rect 7579 12748 7583 12804
rect 7519 12744 7583 12748
rect 2843 12260 2907 12264
rect 2843 12204 2847 12260
rect 2847 12204 2903 12260
rect 2903 12204 2907 12260
rect 2843 12200 2907 12204
rect 2923 12260 2987 12264
rect 2923 12204 2927 12260
rect 2927 12204 2983 12260
rect 2983 12204 2987 12260
rect 2923 12200 2987 12204
rect 3003 12260 3067 12264
rect 3003 12204 3007 12260
rect 3007 12204 3063 12260
rect 3063 12204 3067 12260
rect 3003 12200 3067 12204
rect 3083 12260 3147 12264
rect 3083 12204 3087 12260
rect 3087 12204 3143 12260
rect 3143 12204 3147 12260
rect 3083 12200 3147 12204
rect 5800 12260 5864 12264
rect 5800 12204 5804 12260
rect 5804 12204 5860 12260
rect 5860 12204 5864 12260
rect 5800 12200 5864 12204
rect 5880 12260 5944 12264
rect 5880 12204 5884 12260
rect 5884 12204 5940 12260
rect 5940 12204 5944 12260
rect 5880 12200 5944 12204
rect 5960 12260 6024 12264
rect 5960 12204 5964 12260
rect 5964 12204 6020 12260
rect 6020 12204 6024 12260
rect 5960 12200 6024 12204
rect 6040 12260 6104 12264
rect 6040 12204 6044 12260
rect 6044 12204 6100 12260
rect 6100 12204 6104 12260
rect 6040 12200 6104 12204
rect 1364 11716 1428 11720
rect 1364 11660 1368 11716
rect 1368 11660 1424 11716
rect 1424 11660 1428 11716
rect 1364 11656 1428 11660
rect 1444 11716 1508 11720
rect 1444 11660 1448 11716
rect 1448 11660 1504 11716
rect 1504 11660 1508 11716
rect 1444 11656 1508 11660
rect 1524 11716 1588 11720
rect 1524 11660 1528 11716
rect 1528 11660 1584 11716
rect 1584 11660 1588 11716
rect 1524 11656 1588 11660
rect 1604 11716 1668 11720
rect 1604 11660 1608 11716
rect 1608 11660 1664 11716
rect 1664 11660 1668 11716
rect 1604 11656 1668 11660
rect 4322 11716 4386 11720
rect 4322 11660 4326 11716
rect 4326 11660 4382 11716
rect 4382 11660 4386 11716
rect 4322 11656 4386 11660
rect 4402 11716 4466 11720
rect 4402 11660 4406 11716
rect 4406 11660 4462 11716
rect 4462 11660 4466 11716
rect 4402 11656 4466 11660
rect 4482 11716 4546 11720
rect 4482 11660 4486 11716
rect 4486 11660 4542 11716
rect 4542 11660 4546 11716
rect 4482 11656 4546 11660
rect 4562 11716 4626 11720
rect 4562 11660 4566 11716
rect 4566 11660 4622 11716
rect 4622 11660 4626 11716
rect 4562 11656 4626 11660
rect 7279 11716 7343 11720
rect 7279 11660 7283 11716
rect 7283 11660 7339 11716
rect 7339 11660 7343 11716
rect 7279 11656 7343 11660
rect 7359 11716 7423 11720
rect 7359 11660 7363 11716
rect 7363 11660 7419 11716
rect 7419 11660 7423 11716
rect 7359 11656 7423 11660
rect 7439 11716 7503 11720
rect 7439 11660 7443 11716
rect 7443 11660 7499 11716
rect 7499 11660 7503 11716
rect 7439 11656 7503 11660
rect 7519 11716 7583 11720
rect 7519 11660 7523 11716
rect 7523 11660 7579 11716
rect 7579 11660 7583 11716
rect 7519 11656 7583 11660
rect 2843 11172 2907 11176
rect 2843 11116 2847 11172
rect 2847 11116 2903 11172
rect 2903 11116 2907 11172
rect 2843 11112 2907 11116
rect 2923 11172 2987 11176
rect 2923 11116 2927 11172
rect 2927 11116 2983 11172
rect 2983 11116 2987 11172
rect 2923 11112 2987 11116
rect 3003 11172 3067 11176
rect 3003 11116 3007 11172
rect 3007 11116 3063 11172
rect 3063 11116 3067 11172
rect 3003 11112 3067 11116
rect 3083 11172 3147 11176
rect 3083 11116 3087 11172
rect 3087 11116 3143 11172
rect 3143 11116 3147 11172
rect 3083 11112 3147 11116
rect 5800 11172 5864 11176
rect 5800 11116 5804 11172
rect 5804 11116 5860 11172
rect 5860 11116 5864 11172
rect 5800 11112 5864 11116
rect 5880 11172 5944 11176
rect 5880 11116 5884 11172
rect 5884 11116 5940 11172
rect 5940 11116 5944 11172
rect 5880 11112 5944 11116
rect 5960 11172 6024 11176
rect 5960 11116 5964 11172
rect 5964 11116 6020 11172
rect 6020 11116 6024 11172
rect 5960 11112 6024 11116
rect 6040 11172 6104 11176
rect 6040 11116 6044 11172
rect 6044 11116 6100 11172
rect 6100 11116 6104 11172
rect 6040 11112 6104 11116
rect 1364 10628 1428 10632
rect 1364 10572 1368 10628
rect 1368 10572 1424 10628
rect 1424 10572 1428 10628
rect 1364 10568 1428 10572
rect 1444 10628 1508 10632
rect 1444 10572 1448 10628
rect 1448 10572 1504 10628
rect 1504 10572 1508 10628
rect 1444 10568 1508 10572
rect 1524 10628 1588 10632
rect 1524 10572 1528 10628
rect 1528 10572 1584 10628
rect 1584 10572 1588 10628
rect 1524 10568 1588 10572
rect 1604 10628 1668 10632
rect 1604 10572 1608 10628
rect 1608 10572 1664 10628
rect 1664 10572 1668 10628
rect 1604 10568 1668 10572
rect 4322 10628 4386 10632
rect 4322 10572 4326 10628
rect 4326 10572 4382 10628
rect 4382 10572 4386 10628
rect 4322 10568 4386 10572
rect 4402 10628 4466 10632
rect 4402 10572 4406 10628
rect 4406 10572 4462 10628
rect 4462 10572 4466 10628
rect 4402 10568 4466 10572
rect 4482 10628 4546 10632
rect 4482 10572 4486 10628
rect 4486 10572 4542 10628
rect 4542 10572 4546 10628
rect 4482 10568 4546 10572
rect 4562 10628 4626 10632
rect 4562 10572 4566 10628
rect 4566 10572 4622 10628
rect 4622 10572 4626 10628
rect 4562 10568 4626 10572
rect 7279 10628 7343 10632
rect 7279 10572 7283 10628
rect 7283 10572 7339 10628
rect 7339 10572 7343 10628
rect 7279 10568 7343 10572
rect 7359 10628 7423 10632
rect 7359 10572 7363 10628
rect 7363 10572 7419 10628
rect 7419 10572 7423 10628
rect 7359 10568 7423 10572
rect 7439 10628 7503 10632
rect 7439 10572 7443 10628
rect 7443 10572 7499 10628
rect 7499 10572 7503 10628
rect 7439 10568 7503 10572
rect 7519 10628 7583 10632
rect 7519 10572 7523 10628
rect 7523 10572 7579 10628
rect 7579 10572 7583 10628
rect 7519 10568 7583 10572
rect 2843 10084 2907 10088
rect 2843 10028 2847 10084
rect 2847 10028 2903 10084
rect 2903 10028 2907 10084
rect 2843 10024 2907 10028
rect 2923 10084 2987 10088
rect 2923 10028 2927 10084
rect 2927 10028 2983 10084
rect 2983 10028 2987 10084
rect 2923 10024 2987 10028
rect 3003 10084 3067 10088
rect 3003 10028 3007 10084
rect 3007 10028 3063 10084
rect 3063 10028 3067 10084
rect 3003 10024 3067 10028
rect 3083 10084 3147 10088
rect 3083 10028 3087 10084
rect 3087 10028 3143 10084
rect 3143 10028 3147 10084
rect 3083 10024 3147 10028
rect 5800 10084 5864 10088
rect 5800 10028 5804 10084
rect 5804 10028 5860 10084
rect 5860 10028 5864 10084
rect 5800 10024 5864 10028
rect 5880 10084 5944 10088
rect 5880 10028 5884 10084
rect 5884 10028 5940 10084
rect 5940 10028 5944 10084
rect 5880 10024 5944 10028
rect 5960 10084 6024 10088
rect 5960 10028 5964 10084
rect 5964 10028 6020 10084
rect 6020 10028 6024 10084
rect 5960 10024 6024 10028
rect 6040 10084 6104 10088
rect 6040 10028 6044 10084
rect 6044 10028 6100 10084
rect 6100 10028 6104 10084
rect 6040 10024 6104 10028
rect 1364 9540 1428 9544
rect 1364 9484 1368 9540
rect 1368 9484 1424 9540
rect 1424 9484 1428 9540
rect 1364 9480 1428 9484
rect 1444 9540 1508 9544
rect 1444 9484 1448 9540
rect 1448 9484 1504 9540
rect 1504 9484 1508 9540
rect 1444 9480 1508 9484
rect 1524 9540 1588 9544
rect 1524 9484 1528 9540
rect 1528 9484 1584 9540
rect 1584 9484 1588 9540
rect 1524 9480 1588 9484
rect 1604 9540 1668 9544
rect 1604 9484 1608 9540
rect 1608 9484 1664 9540
rect 1664 9484 1668 9540
rect 1604 9480 1668 9484
rect 4322 9540 4386 9544
rect 4322 9484 4326 9540
rect 4326 9484 4382 9540
rect 4382 9484 4386 9540
rect 4322 9480 4386 9484
rect 4402 9540 4466 9544
rect 4402 9484 4406 9540
rect 4406 9484 4462 9540
rect 4462 9484 4466 9540
rect 4402 9480 4466 9484
rect 4482 9540 4546 9544
rect 4482 9484 4486 9540
rect 4486 9484 4542 9540
rect 4542 9484 4546 9540
rect 4482 9480 4546 9484
rect 4562 9540 4626 9544
rect 4562 9484 4566 9540
rect 4566 9484 4622 9540
rect 4622 9484 4626 9540
rect 4562 9480 4626 9484
rect 7279 9540 7343 9544
rect 7279 9484 7283 9540
rect 7283 9484 7339 9540
rect 7339 9484 7343 9540
rect 7279 9480 7343 9484
rect 7359 9540 7423 9544
rect 7359 9484 7363 9540
rect 7363 9484 7419 9540
rect 7419 9484 7423 9540
rect 7359 9480 7423 9484
rect 7439 9540 7503 9544
rect 7439 9484 7443 9540
rect 7443 9484 7499 9540
rect 7499 9484 7503 9540
rect 7439 9480 7503 9484
rect 7519 9540 7583 9544
rect 7519 9484 7523 9540
rect 7523 9484 7579 9540
rect 7579 9484 7583 9540
rect 7519 9480 7583 9484
rect 2843 8996 2907 9000
rect 2843 8940 2847 8996
rect 2847 8940 2903 8996
rect 2903 8940 2907 8996
rect 2843 8936 2907 8940
rect 2923 8996 2987 9000
rect 2923 8940 2927 8996
rect 2927 8940 2983 8996
rect 2983 8940 2987 8996
rect 2923 8936 2987 8940
rect 3003 8996 3067 9000
rect 3003 8940 3007 8996
rect 3007 8940 3063 8996
rect 3063 8940 3067 8996
rect 3003 8936 3067 8940
rect 3083 8996 3147 9000
rect 3083 8940 3087 8996
rect 3087 8940 3143 8996
rect 3143 8940 3147 8996
rect 3083 8936 3147 8940
rect 5800 8996 5864 9000
rect 5800 8940 5804 8996
rect 5804 8940 5860 8996
rect 5860 8940 5864 8996
rect 5800 8936 5864 8940
rect 5880 8996 5944 9000
rect 5880 8940 5884 8996
rect 5884 8940 5940 8996
rect 5940 8940 5944 8996
rect 5880 8936 5944 8940
rect 5960 8996 6024 9000
rect 5960 8940 5964 8996
rect 5964 8940 6020 8996
rect 6020 8940 6024 8996
rect 5960 8936 6024 8940
rect 6040 8996 6104 9000
rect 6040 8940 6044 8996
rect 6044 8940 6100 8996
rect 6100 8940 6104 8996
rect 6040 8936 6104 8940
rect 1364 8452 1428 8456
rect 1364 8396 1368 8452
rect 1368 8396 1424 8452
rect 1424 8396 1428 8452
rect 1364 8392 1428 8396
rect 1444 8452 1508 8456
rect 1444 8396 1448 8452
rect 1448 8396 1504 8452
rect 1504 8396 1508 8452
rect 1444 8392 1508 8396
rect 1524 8452 1588 8456
rect 1524 8396 1528 8452
rect 1528 8396 1584 8452
rect 1584 8396 1588 8452
rect 1524 8392 1588 8396
rect 1604 8452 1668 8456
rect 1604 8396 1608 8452
rect 1608 8396 1664 8452
rect 1664 8396 1668 8452
rect 1604 8392 1668 8396
rect 4322 8452 4386 8456
rect 4322 8396 4326 8452
rect 4326 8396 4382 8452
rect 4382 8396 4386 8452
rect 4322 8392 4386 8396
rect 4402 8452 4466 8456
rect 4402 8396 4406 8452
rect 4406 8396 4462 8452
rect 4462 8396 4466 8452
rect 4402 8392 4466 8396
rect 4482 8452 4546 8456
rect 4482 8396 4486 8452
rect 4486 8396 4542 8452
rect 4542 8396 4546 8452
rect 4482 8392 4546 8396
rect 4562 8452 4626 8456
rect 4562 8396 4566 8452
rect 4566 8396 4622 8452
rect 4622 8396 4626 8452
rect 4562 8392 4626 8396
rect 7279 8452 7343 8456
rect 7279 8396 7283 8452
rect 7283 8396 7339 8452
rect 7339 8396 7343 8452
rect 7279 8392 7343 8396
rect 7359 8452 7423 8456
rect 7359 8396 7363 8452
rect 7363 8396 7419 8452
rect 7419 8396 7423 8452
rect 7359 8392 7423 8396
rect 7439 8452 7503 8456
rect 7439 8396 7443 8452
rect 7443 8396 7499 8452
rect 7499 8396 7503 8452
rect 7439 8392 7503 8396
rect 7519 8452 7583 8456
rect 7519 8396 7523 8452
rect 7523 8396 7579 8452
rect 7579 8396 7583 8452
rect 7519 8392 7583 8396
rect 2843 7908 2907 7912
rect 2843 7852 2847 7908
rect 2847 7852 2903 7908
rect 2903 7852 2907 7908
rect 2843 7848 2907 7852
rect 2923 7908 2987 7912
rect 2923 7852 2927 7908
rect 2927 7852 2983 7908
rect 2983 7852 2987 7908
rect 2923 7848 2987 7852
rect 3003 7908 3067 7912
rect 3003 7852 3007 7908
rect 3007 7852 3063 7908
rect 3063 7852 3067 7908
rect 3003 7848 3067 7852
rect 3083 7908 3147 7912
rect 3083 7852 3087 7908
rect 3087 7852 3143 7908
rect 3143 7852 3147 7908
rect 3083 7848 3147 7852
rect 5800 7908 5864 7912
rect 5800 7852 5804 7908
rect 5804 7852 5860 7908
rect 5860 7852 5864 7908
rect 5800 7848 5864 7852
rect 5880 7908 5944 7912
rect 5880 7852 5884 7908
rect 5884 7852 5940 7908
rect 5940 7852 5944 7908
rect 5880 7848 5944 7852
rect 5960 7908 6024 7912
rect 5960 7852 5964 7908
rect 5964 7852 6020 7908
rect 6020 7852 6024 7908
rect 5960 7848 6024 7852
rect 6040 7908 6104 7912
rect 6040 7852 6044 7908
rect 6044 7852 6100 7908
rect 6100 7852 6104 7908
rect 6040 7848 6104 7852
rect 1364 7364 1428 7368
rect 1364 7308 1368 7364
rect 1368 7308 1424 7364
rect 1424 7308 1428 7364
rect 1364 7304 1428 7308
rect 1444 7364 1508 7368
rect 1444 7308 1448 7364
rect 1448 7308 1504 7364
rect 1504 7308 1508 7364
rect 1444 7304 1508 7308
rect 1524 7364 1588 7368
rect 1524 7308 1528 7364
rect 1528 7308 1584 7364
rect 1584 7308 1588 7364
rect 1524 7304 1588 7308
rect 1604 7364 1668 7368
rect 1604 7308 1608 7364
rect 1608 7308 1664 7364
rect 1664 7308 1668 7364
rect 1604 7304 1668 7308
rect 4322 7364 4386 7368
rect 4322 7308 4326 7364
rect 4326 7308 4382 7364
rect 4382 7308 4386 7364
rect 4322 7304 4386 7308
rect 4402 7364 4466 7368
rect 4402 7308 4406 7364
rect 4406 7308 4462 7364
rect 4462 7308 4466 7364
rect 4402 7304 4466 7308
rect 4482 7364 4546 7368
rect 4482 7308 4486 7364
rect 4486 7308 4542 7364
rect 4542 7308 4546 7364
rect 4482 7304 4546 7308
rect 4562 7364 4626 7368
rect 4562 7308 4566 7364
rect 4566 7308 4622 7364
rect 4622 7308 4626 7364
rect 4562 7304 4626 7308
rect 7279 7364 7343 7368
rect 7279 7308 7283 7364
rect 7283 7308 7339 7364
rect 7339 7308 7343 7364
rect 7279 7304 7343 7308
rect 7359 7364 7423 7368
rect 7359 7308 7363 7364
rect 7363 7308 7419 7364
rect 7419 7308 7423 7364
rect 7359 7304 7423 7308
rect 7439 7364 7503 7368
rect 7439 7308 7443 7364
rect 7443 7308 7499 7364
rect 7499 7308 7503 7364
rect 7439 7304 7503 7308
rect 7519 7364 7583 7368
rect 7519 7308 7523 7364
rect 7523 7308 7579 7364
rect 7579 7308 7583 7364
rect 7519 7304 7583 7308
rect 2843 6820 2907 6824
rect 2843 6764 2847 6820
rect 2847 6764 2903 6820
rect 2903 6764 2907 6820
rect 2843 6760 2907 6764
rect 2923 6820 2987 6824
rect 2923 6764 2927 6820
rect 2927 6764 2983 6820
rect 2983 6764 2987 6820
rect 2923 6760 2987 6764
rect 3003 6820 3067 6824
rect 3003 6764 3007 6820
rect 3007 6764 3063 6820
rect 3063 6764 3067 6820
rect 3003 6760 3067 6764
rect 3083 6820 3147 6824
rect 3083 6764 3087 6820
rect 3087 6764 3143 6820
rect 3143 6764 3147 6820
rect 3083 6760 3147 6764
rect 5800 6820 5864 6824
rect 5800 6764 5804 6820
rect 5804 6764 5860 6820
rect 5860 6764 5864 6820
rect 5800 6760 5864 6764
rect 5880 6820 5944 6824
rect 5880 6764 5884 6820
rect 5884 6764 5940 6820
rect 5940 6764 5944 6820
rect 5880 6760 5944 6764
rect 5960 6820 6024 6824
rect 5960 6764 5964 6820
rect 5964 6764 6020 6820
rect 6020 6764 6024 6820
rect 5960 6760 6024 6764
rect 6040 6820 6104 6824
rect 6040 6764 6044 6820
rect 6044 6764 6100 6820
rect 6100 6764 6104 6820
rect 6040 6760 6104 6764
rect 1364 6276 1428 6280
rect 1364 6220 1368 6276
rect 1368 6220 1424 6276
rect 1424 6220 1428 6276
rect 1364 6216 1428 6220
rect 1444 6276 1508 6280
rect 1444 6220 1448 6276
rect 1448 6220 1504 6276
rect 1504 6220 1508 6276
rect 1444 6216 1508 6220
rect 1524 6276 1588 6280
rect 1524 6220 1528 6276
rect 1528 6220 1584 6276
rect 1584 6220 1588 6276
rect 1524 6216 1588 6220
rect 1604 6276 1668 6280
rect 1604 6220 1608 6276
rect 1608 6220 1664 6276
rect 1664 6220 1668 6276
rect 1604 6216 1668 6220
rect 4322 6276 4386 6280
rect 4322 6220 4326 6276
rect 4326 6220 4382 6276
rect 4382 6220 4386 6276
rect 4322 6216 4386 6220
rect 4402 6276 4466 6280
rect 4402 6220 4406 6276
rect 4406 6220 4462 6276
rect 4462 6220 4466 6276
rect 4402 6216 4466 6220
rect 4482 6276 4546 6280
rect 4482 6220 4486 6276
rect 4486 6220 4542 6276
rect 4542 6220 4546 6276
rect 4482 6216 4546 6220
rect 4562 6276 4626 6280
rect 4562 6220 4566 6276
rect 4566 6220 4622 6276
rect 4622 6220 4626 6276
rect 4562 6216 4626 6220
rect 7279 6276 7343 6280
rect 7279 6220 7283 6276
rect 7283 6220 7339 6276
rect 7339 6220 7343 6276
rect 7279 6216 7343 6220
rect 7359 6276 7423 6280
rect 7359 6220 7363 6276
rect 7363 6220 7419 6276
rect 7419 6220 7423 6276
rect 7359 6216 7423 6220
rect 7439 6276 7503 6280
rect 7439 6220 7443 6276
rect 7443 6220 7499 6276
rect 7499 6220 7503 6276
rect 7439 6216 7503 6220
rect 7519 6276 7583 6280
rect 7519 6220 7523 6276
rect 7523 6220 7579 6276
rect 7579 6220 7583 6276
rect 7519 6216 7583 6220
rect 2843 5732 2907 5736
rect 2843 5676 2847 5732
rect 2847 5676 2903 5732
rect 2903 5676 2907 5732
rect 2843 5672 2907 5676
rect 2923 5732 2987 5736
rect 2923 5676 2927 5732
rect 2927 5676 2983 5732
rect 2983 5676 2987 5732
rect 2923 5672 2987 5676
rect 3003 5732 3067 5736
rect 3003 5676 3007 5732
rect 3007 5676 3063 5732
rect 3063 5676 3067 5732
rect 3003 5672 3067 5676
rect 3083 5732 3147 5736
rect 3083 5676 3087 5732
rect 3087 5676 3143 5732
rect 3143 5676 3147 5732
rect 3083 5672 3147 5676
rect 5800 5732 5864 5736
rect 5800 5676 5804 5732
rect 5804 5676 5860 5732
rect 5860 5676 5864 5732
rect 5800 5672 5864 5676
rect 5880 5732 5944 5736
rect 5880 5676 5884 5732
rect 5884 5676 5940 5732
rect 5940 5676 5944 5732
rect 5880 5672 5944 5676
rect 5960 5732 6024 5736
rect 5960 5676 5964 5732
rect 5964 5676 6020 5732
rect 6020 5676 6024 5732
rect 5960 5672 6024 5676
rect 6040 5732 6104 5736
rect 6040 5676 6044 5732
rect 6044 5676 6100 5732
rect 6100 5676 6104 5732
rect 6040 5672 6104 5676
rect 1364 5188 1428 5192
rect 1364 5132 1368 5188
rect 1368 5132 1424 5188
rect 1424 5132 1428 5188
rect 1364 5128 1428 5132
rect 1444 5188 1508 5192
rect 1444 5132 1448 5188
rect 1448 5132 1504 5188
rect 1504 5132 1508 5188
rect 1444 5128 1508 5132
rect 1524 5188 1588 5192
rect 1524 5132 1528 5188
rect 1528 5132 1584 5188
rect 1584 5132 1588 5188
rect 1524 5128 1588 5132
rect 1604 5188 1668 5192
rect 1604 5132 1608 5188
rect 1608 5132 1664 5188
rect 1664 5132 1668 5188
rect 1604 5128 1668 5132
rect 4322 5188 4386 5192
rect 4322 5132 4326 5188
rect 4326 5132 4382 5188
rect 4382 5132 4386 5188
rect 4322 5128 4386 5132
rect 4402 5188 4466 5192
rect 4402 5132 4406 5188
rect 4406 5132 4462 5188
rect 4462 5132 4466 5188
rect 4402 5128 4466 5132
rect 4482 5188 4546 5192
rect 4482 5132 4486 5188
rect 4486 5132 4542 5188
rect 4542 5132 4546 5188
rect 4482 5128 4546 5132
rect 4562 5188 4626 5192
rect 4562 5132 4566 5188
rect 4566 5132 4622 5188
rect 4622 5132 4626 5188
rect 4562 5128 4626 5132
rect 7279 5188 7343 5192
rect 7279 5132 7283 5188
rect 7283 5132 7339 5188
rect 7339 5132 7343 5188
rect 7279 5128 7343 5132
rect 7359 5188 7423 5192
rect 7359 5132 7363 5188
rect 7363 5132 7419 5188
rect 7419 5132 7423 5188
rect 7359 5128 7423 5132
rect 7439 5188 7503 5192
rect 7439 5132 7443 5188
rect 7443 5132 7499 5188
rect 7499 5132 7503 5188
rect 7439 5128 7503 5132
rect 7519 5188 7583 5192
rect 7519 5132 7523 5188
rect 7523 5132 7579 5188
rect 7579 5132 7583 5188
rect 7519 5128 7583 5132
rect 2843 4644 2907 4648
rect 2843 4588 2847 4644
rect 2847 4588 2903 4644
rect 2903 4588 2907 4644
rect 2843 4584 2907 4588
rect 2923 4644 2987 4648
rect 2923 4588 2927 4644
rect 2927 4588 2983 4644
rect 2983 4588 2987 4644
rect 2923 4584 2987 4588
rect 3003 4644 3067 4648
rect 3003 4588 3007 4644
rect 3007 4588 3063 4644
rect 3063 4588 3067 4644
rect 3003 4584 3067 4588
rect 3083 4644 3147 4648
rect 3083 4588 3087 4644
rect 3087 4588 3143 4644
rect 3143 4588 3147 4644
rect 3083 4584 3147 4588
rect 5800 4644 5864 4648
rect 5800 4588 5804 4644
rect 5804 4588 5860 4644
rect 5860 4588 5864 4644
rect 5800 4584 5864 4588
rect 5880 4644 5944 4648
rect 5880 4588 5884 4644
rect 5884 4588 5940 4644
rect 5940 4588 5944 4644
rect 5880 4584 5944 4588
rect 5960 4644 6024 4648
rect 5960 4588 5964 4644
rect 5964 4588 6020 4644
rect 6020 4588 6024 4644
rect 5960 4584 6024 4588
rect 6040 4644 6104 4648
rect 6040 4588 6044 4644
rect 6044 4588 6100 4644
rect 6100 4588 6104 4644
rect 6040 4584 6104 4588
rect 1364 4100 1428 4104
rect 1364 4044 1368 4100
rect 1368 4044 1424 4100
rect 1424 4044 1428 4100
rect 1364 4040 1428 4044
rect 1444 4100 1508 4104
rect 1444 4044 1448 4100
rect 1448 4044 1504 4100
rect 1504 4044 1508 4100
rect 1444 4040 1508 4044
rect 1524 4100 1588 4104
rect 1524 4044 1528 4100
rect 1528 4044 1584 4100
rect 1584 4044 1588 4100
rect 1524 4040 1588 4044
rect 1604 4100 1668 4104
rect 1604 4044 1608 4100
rect 1608 4044 1664 4100
rect 1664 4044 1668 4100
rect 1604 4040 1668 4044
rect 4322 4100 4386 4104
rect 4322 4044 4326 4100
rect 4326 4044 4382 4100
rect 4382 4044 4386 4100
rect 4322 4040 4386 4044
rect 4402 4100 4466 4104
rect 4402 4044 4406 4100
rect 4406 4044 4462 4100
rect 4462 4044 4466 4100
rect 4402 4040 4466 4044
rect 4482 4100 4546 4104
rect 4482 4044 4486 4100
rect 4486 4044 4542 4100
rect 4542 4044 4546 4100
rect 4482 4040 4546 4044
rect 4562 4100 4626 4104
rect 4562 4044 4566 4100
rect 4566 4044 4622 4100
rect 4622 4044 4626 4100
rect 4562 4040 4626 4044
rect 7279 4100 7343 4104
rect 7279 4044 7283 4100
rect 7283 4044 7339 4100
rect 7339 4044 7343 4100
rect 7279 4040 7343 4044
rect 7359 4100 7423 4104
rect 7359 4044 7363 4100
rect 7363 4044 7419 4100
rect 7419 4044 7423 4100
rect 7359 4040 7423 4044
rect 7439 4100 7503 4104
rect 7439 4044 7443 4100
rect 7443 4044 7499 4100
rect 7499 4044 7503 4100
rect 7439 4040 7503 4044
rect 7519 4100 7583 4104
rect 7519 4044 7523 4100
rect 7523 4044 7579 4100
rect 7579 4044 7583 4100
rect 7519 4040 7583 4044
rect 2843 3556 2907 3560
rect 2843 3500 2847 3556
rect 2847 3500 2903 3556
rect 2903 3500 2907 3556
rect 2843 3496 2907 3500
rect 2923 3556 2987 3560
rect 2923 3500 2927 3556
rect 2927 3500 2983 3556
rect 2983 3500 2987 3556
rect 2923 3496 2987 3500
rect 3003 3556 3067 3560
rect 3003 3500 3007 3556
rect 3007 3500 3063 3556
rect 3063 3500 3067 3556
rect 3003 3496 3067 3500
rect 3083 3556 3147 3560
rect 3083 3500 3087 3556
rect 3087 3500 3143 3556
rect 3143 3500 3147 3556
rect 3083 3496 3147 3500
rect 5800 3556 5864 3560
rect 5800 3500 5804 3556
rect 5804 3500 5860 3556
rect 5860 3500 5864 3556
rect 5800 3496 5864 3500
rect 5880 3556 5944 3560
rect 5880 3500 5884 3556
rect 5884 3500 5940 3556
rect 5940 3500 5944 3556
rect 5880 3496 5944 3500
rect 5960 3556 6024 3560
rect 5960 3500 5964 3556
rect 5964 3500 6020 3556
rect 6020 3500 6024 3556
rect 5960 3496 6024 3500
rect 6040 3556 6104 3560
rect 6040 3500 6044 3556
rect 6044 3500 6100 3556
rect 6100 3500 6104 3556
rect 6040 3496 6104 3500
rect 1364 3012 1428 3016
rect 1364 2956 1368 3012
rect 1368 2956 1424 3012
rect 1424 2956 1428 3012
rect 1364 2952 1428 2956
rect 1444 3012 1508 3016
rect 1444 2956 1448 3012
rect 1448 2956 1504 3012
rect 1504 2956 1508 3012
rect 1444 2952 1508 2956
rect 1524 3012 1588 3016
rect 1524 2956 1528 3012
rect 1528 2956 1584 3012
rect 1584 2956 1588 3012
rect 1524 2952 1588 2956
rect 1604 3012 1668 3016
rect 1604 2956 1608 3012
rect 1608 2956 1664 3012
rect 1664 2956 1668 3012
rect 1604 2952 1668 2956
rect 4322 3012 4386 3016
rect 4322 2956 4326 3012
rect 4326 2956 4382 3012
rect 4382 2956 4386 3012
rect 4322 2952 4386 2956
rect 4402 3012 4466 3016
rect 4402 2956 4406 3012
rect 4406 2956 4462 3012
rect 4462 2956 4466 3012
rect 4402 2952 4466 2956
rect 4482 3012 4546 3016
rect 4482 2956 4486 3012
rect 4486 2956 4542 3012
rect 4542 2956 4546 3012
rect 4482 2952 4546 2956
rect 4562 3012 4626 3016
rect 4562 2956 4566 3012
rect 4566 2956 4622 3012
rect 4622 2956 4626 3012
rect 4562 2952 4626 2956
rect 7279 3012 7343 3016
rect 7279 2956 7283 3012
rect 7283 2956 7339 3012
rect 7339 2956 7343 3012
rect 7279 2952 7343 2956
rect 7359 3012 7423 3016
rect 7359 2956 7363 3012
rect 7363 2956 7419 3012
rect 7419 2956 7423 3012
rect 7359 2952 7423 2956
rect 7439 3012 7503 3016
rect 7439 2956 7443 3012
rect 7443 2956 7499 3012
rect 7499 2956 7503 3012
rect 7439 2952 7503 2956
rect 7519 3012 7583 3016
rect 7519 2956 7523 3012
rect 7523 2956 7579 3012
rect 7579 2956 7583 3012
rect 7519 2952 7583 2956
rect 2843 2468 2907 2472
rect 2843 2412 2847 2468
rect 2847 2412 2903 2468
rect 2903 2412 2907 2468
rect 2843 2408 2907 2412
rect 2923 2468 2987 2472
rect 2923 2412 2927 2468
rect 2927 2412 2983 2468
rect 2983 2412 2987 2468
rect 2923 2408 2987 2412
rect 3003 2468 3067 2472
rect 3003 2412 3007 2468
rect 3007 2412 3063 2468
rect 3063 2412 3067 2468
rect 3003 2408 3067 2412
rect 3083 2468 3147 2472
rect 3083 2412 3087 2468
rect 3087 2412 3143 2468
rect 3143 2412 3147 2468
rect 3083 2408 3147 2412
rect 5800 2468 5864 2472
rect 5800 2412 5804 2468
rect 5804 2412 5860 2468
rect 5860 2412 5864 2468
rect 5800 2408 5864 2412
rect 5880 2468 5944 2472
rect 5880 2412 5884 2468
rect 5884 2412 5940 2468
rect 5940 2412 5944 2468
rect 5880 2408 5944 2412
rect 5960 2468 6024 2472
rect 5960 2412 5964 2468
rect 5964 2412 6020 2468
rect 6020 2412 6024 2468
rect 5960 2408 6024 2412
rect 6040 2468 6104 2472
rect 6040 2412 6044 2468
rect 6044 2412 6100 2468
rect 6100 2412 6104 2468
rect 6040 2408 6104 2412
rect 1364 1924 1428 1928
rect 1364 1868 1368 1924
rect 1368 1868 1424 1924
rect 1424 1868 1428 1924
rect 1364 1864 1428 1868
rect 1444 1924 1508 1928
rect 1444 1868 1448 1924
rect 1448 1868 1504 1924
rect 1504 1868 1508 1924
rect 1444 1864 1508 1868
rect 1524 1924 1588 1928
rect 1524 1868 1528 1924
rect 1528 1868 1584 1924
rect 1584 1868 1588 1924
rect 1524 1864 1588 1868
rect 1604 1924 1668 1928
rect 1604 1868 1608 1924
rect 1608 1868 1664 1924
rect 1664 1868 1668 1924
rect 1604 1864 1668 1868
rect 4322 1924 4386 1928
rect 4322 1868 4326 1924
rect 4326 1868 4382 1924
rect 4382 1868 4386 1924
rect 4322 1864 4386 1868
rect 4402 1924 4466 1928
rect 4402 1868 4406 1924
rect 4406 1868 4462 1924
rect 4462 1868 4466 1924
rect 4402 1864 4466 1868
rect 4482 1924 4546 1928
rect 4482 1868 4486 1924
rect 4486 1868 4542 1924
rect 4542 1868 4546 1924
rect 4482 1864 4546 1868
rect 4562 1924 4626 1928
rect 4562 1868 4566 1924
rect 4566 1868 4622 1924
rect 4622 1868 4626 1924
rect 4562 1864 4626 1868
rect 7279 1924 7343 1928
rect 7279 1868 7283 1924
rect 7283 1868 7339 1924
rect 7339 1868 7343 1924
rect 7279 1864 7343 1868
rect 7359 1924 7423 1928
rect 7359 1868 7363 1924
rect 7363 1868 7419 1924
rect 7419 1868 7423 1924
rect 7359 1864 7423 1868
rect 7439 1924 7503 1928
rect 7439 1868 7443 1924
rect 7443 1868 7499 1924
rect 7499 1868 7503 1924
rect 7439 1864 7503 1868
rect 7519 1924 7583 1928
rect 7519 1868 7523 1924
rect 7523 1868 7579 1924
rect 7579 1868 7583 1924
rect 7519 1864 7583 1868
<< metal4 >>
rect 1356 16072 1676 16088
rect 1356 16008 1364 16072
rect 1428 16008 1444 16072
rect 1508 16008 1524 16072
rect 1588 16008 1604 16072
rect 1668 16008 1676 16072
rect 1356 14984 1676 16008
rect 1356 14920 1364 14984
rect 1428 14920 1444 14984
rect 1508 14920 1524 14984
rect 1588 14920 1604 14984
rect 1668 14920 1676 14984
rect 1356 14172 1676 14920
rect 1356 13936 1398 14172
rect 1634 13936 1676 14172
rect 1356 13896 1676 13936
rect 1356 13832 1364 13896
rect 1428 13832 1444 13896
rect 1508 13832 1524 13896
rect 1588 13832 1604 13896
rect 1668 13832 1676 13896
rect 1356 12808 1676 13832
rect 1356 12744 1364 12808
rect 1428 12744 1444 12808
rect 1508 12744 1524 12808
rect 1588 12744 1604 12808
rect 1668 12744 1676 12808
rect 1356 11720 1676 12744
rect 1356 11656 1364 11720
rect 1428 11656 1444 11720
rect 1508 11656 1524 11720
rect 1588 11656 1604 11720
rect 1668 11656 1676 11720
rect 1356 10632 1676 11656
rect 1356 10568 1364 10632
rect 1428 10568 1444 10632
rect 1508 10568 1524 10632
rect 1588 10568 1604 10632
rect 1668 10568 1676 10632
rect 1356 9544 1676 10568
rect 1356 9480 1364 9544
rect 1428 9480 1444 9544
rect 1508 9480 1524 9544
rect 1588 9480 1604 9544
rect 1668 9480 1676 9544
rect 1356 9290 1676 9480
rect 1356 9054 1398 9290
rect 1634 9054 1676 9290
rect 1356 8456 1676 9054
rect 1356 8392 1364 8456
rect 1428 8392 1444 8456
rect 1508 8392 1524 8456
rect 1588 8392 1604 8456
rect 1668 8392 1676 8456
rect 1356 7368 1676 8392
rect 1356 7304 1364 7368
rect 1428 7304 1444 7368
rect 1508 7304 1524 7368
rect 1588 7304 1604 7368
rect 1668 7304 1676 7368
rect 1356 6280 1676 7304
rect 1356 6216 1364 6280
rect 1428 6216 1444 6280
rect 1508 6216 1524 6280
rect 1588 6216 1604 6280
rect 1668 6216 1676 6280
rect 1356 5192 1676 6216
rect 1356 5128 1364 5192
rect 1428 5128 1444 5192
rect 1508 5128 1524 5192
rect 1588 5128 1604 5192
rect 1668 5128 1676 5192
rect 1356 4407 1676 5128
rect 1356 4171 1398 4407
rect 1634 4171 1676 4407
rect 1356 4104 1676 4171
rect 1356 4040 1364 4104
rect 1428 4040 1444 4104
rect 1508 4040 1524 4104
rect 1588 4040 1604 4104
rect 1668 4040 1676 4104
rect 1356 3016 1676 4040
rect 1356 2952 1364 3016
rect 1428 2952 1444 3016
rect 1508 2952 1524 3016
rect 1588 2952 1604 3016
rect 1668 2952 1676 3016
rect 1356 1928 1676 2952
rect 1356 1864 1364 1928
rect 1428 1864 1444 1928
rect 1508 1864 1524 1928
rect 1588 1864 1604 1928
rect 1668 1864 1676 1928
rect 1356 1848 1676 1864
rect 2835 15528 3155 16088
rect 2835 15464 2843 15528
rect 2907 15464 2923 15528
rect 2987 15464 3003 15528
rect 3067 15464 3083 15528
rect 3147 15464 3155 15528
rect 2835 14440 3155 15464
rect 2835 14376 2843 14440
rect 2907 14376 2923 14440
rect 2987 14376 3003 14440
rect 3067 14376 3083 14440
rect 3147 14376 3155 14440
rect 2835 13352 3155 14376
rect 2835 13288 2843 13352
rect 2907 13288 2923 13352
rect 2987 13288 3003 13352
rect 3067 13288 3083 13352
rect 3147 13288 3155 13352
rect 2835 12264 3155 13288
rect 2835 12200 2843 12264
rect 2907 12200 2923 12264
rect 2987 12200 3003 12264
rect 3067 12200 3083 12264
rect 3147 12200 3155 12264
rect 2835 11731 3155 12200
rect 2835 11495 2877 11731
rect 3113 11495 3155 11731
rect 2835 11176 3155 11495
rect 2835 11112 2843 11176
rect 2907 11112 2923 11176
rect 2987 11112 3003 11176
rect 3067 11112 3083 11176
rect 3147 11112 3155 11176
rect 2835 10088 3155 11112
rect 2835 10024 2843 10088
rect 2907 10024 2923 10088
rect 2987 10024 3003 10088
rect 3067 10024 3083 10088
rect 3147 10024 3155 10088
rect 2835 9000 3155 10024
rect 2835 8936 2843 9000
rect 2907 8936 2923 9000
rect 2987 8936 3003 9000
rect 3067 8936 3083 9000
rect 3147 8936 3155 9000
rect 2835 7912 3155 8936
rect 2835 7848 2843 7912
rect 2907 7848 2923 7912
rect 2987 7848 3003 7912
rect 3067 7848 3083 7912
rect 3147 7848 3155 7912
rect 2835 6848 3155 7848
rect 2835 6824 2877 6848
rect 3113 6824 3155 6848
rect 2835 6760 2843 6824
rect 3147 6760 3155 6824
rect 2835 6612 2877 6760
rect 3113 6612 3155 6760
rect 2835 5736 3155 6612
rect 2835 5672 2843 5736
rect 2907 5672 2923 5736
rect 2987 5672 3003 5736
rect 3067 5672 3083 5736
rect 3147 5672 3155 5736
rect 2835 4648 3155 5672
rect 2835 4584 2843 4648
rect 2907 4584 2923 4648
rect 2987 4584 3003 4648
rect 3067 4584 3083 4648
rect 3147 4584 3155 4648
rect 2835 3560 3155 4584
rect 2835 3496 2843 3560
rect 2907 3496 2923 3560
rect 2987 3496 3003 3560
rect 3067 3496 3083 3560
rect 3147 3496 3155 3560
rect 2835 2472 3155 3496
rect 2835 2408 2843 2472
rect 2907 2408 2923 2472
rect 2987 2408 3003 2472
rect 3067 2408 3083 2472
rect 3147 2408 3155 2472
rect 2835 1848 3155 2408
rect 4314 16072 4634 16088
rect 4314 16008 4322 16072
rect 4386 16008 4402 16072
rect 4466 16008 4482 16072
rect 4546 16008 4562 16072
rect 4626 16008 4634 16072
rect 4314 14984 4634 16008
rect 4314 14920 4322 14984
rect 4386 14920 4402 14984
rect 4466 14920 4482 14984
rect 4546 14920 4562 14984
rect 4626 14920 4634 14984
rect 4314 14172 4634 14920
rect 4314 13936 4356 14172
rect 4592 13936 4634 14172
rect 4314 13896 4634 13936
rect 4314 13832 4322 13896
rect 4386 13832 4402 13896
rect 4466 13832 4482 13896
rect 4546 13832 4562 13896
rect 4626 13832 4634 13896
rect 4314 12808 4634 13832
rect 4314 12744 4322 12808
rect 4386 12744 4402 12808
rect 4466 12744 4482 12808
rect 4546 12744 4562 12808
rect 4626 12744 4634 12808
rect 4314 11720 4634 12744
rect 4314 11656 4322 11720
rect 4386 11656 4402 11720
rect 4466 11656 4482 11720
rect 4546 11656 4562 11720
rect 4626 11656 4634 11720
rect 4314 10632 4634 11656
rect 4314 10568 4322 10632
rect 4386 10568 4402 10632
rect 4466 10568 4482 10632
rect 4546 10568 4562 10632
rect 4626 10568 4634 10632
rect 4314 9544 4634 10568
rect 4314 9480 4322 9544
rect 4386 9480 4402 9544
rect 4466 9480 4482 9544
rect 4546 9480 4562 9544
rect 4626 9480 4634 9544
rect 4314 9290 4634 9480
rect 4314 9054 4356 9290
rect 4592 9054 4634 9290
rect 4314 8456 4634 9054
rect 4314 8392 4322 8456
rect 4386 8392 4402 8456
rect 4466 8392 4482 8456
rect 4546 8392 4562 8456
rect 4626 8392 4634 8456
rect 4314 7368 4634 8392
rect 4314 7304 4322 7368
rect 4386 7304 4402 7368
rect 4466 7304 4482 7368
rect 4546 7304 4562 7368
rect 4626 7304 4634 7368
rect 4314 6280 4634 7304
rect 4314 6216 4322 6280
rect 4386 6216 4402 6280
rect 4466 6216 4482 6280
rect 4546 6216 4562 6280
rect 4626 6216 4634 6280
rect 4314 5192 4634 6216
rect 4314 5128 4322 5192
rect 4386 5128 4402 5192
rect 4466 5128 4482 5192
rect 4546 5128 4562 5192
rect 4626 5128 4634 5192
rect 4314 4407 4634 5128
rect 4314 4171 4356 4407
rect 4592 4171 4634 4407
rect 4314 4104 4634 4171
rect 4314 4040 4322 4104
rect 4386 4040 4402 4104
rect 4466 4040 4482 4104
rect 4546 4040 4562 4104
rect 4626 4040 4634 4104
rect 4314 3016 4634 4040
rect 4314 2952 4322 3016
rect 4386 2952 4402 3016
rect 4466 2952 4482 3016
rect 4546 2952 4562 3016
rect 4626 2952 4634 3016
rect 4314 1928 4634 2952
rect 4314 1864 4322 1928
rect 4386 1864 4402 1928
rect 4466 1864 4482 1928
rect 4546 1864 4562 1928
rect 4626 1864 4634 1928
rect 4314 1848 4634 1864
rect 5792 15528 6112 16088
rect 5792 15464 5800 15528
rect 5864 15464 5880 15528
rect 5944 15464 5960 15528
rect 6024 15464 6040 15528
rect 6104 15464 6112 15528
rect 5792 14440 6112 15464
rect 5792 14376 5800 14440
rect 5864 14376 5880 14440
rect 5944 14376 5960 14440
rect 6024 14376 6040 14440
rect 6104 14376 6112 14440
rect 5792 13352 6112 14376
rect 5792 13288 5800 13352
rect 5864 13288 5880 13352
rect 5944 13288 5960 13352
rect 6024 13288 6040 13352
rect 6104 13288 6112 13352
rect 5792 12264 6112 13288
rect 5792 12200 5800 12264
rect 5864 12200 5880 12264
rect 5944 12200 5960 12264
rect 6024 12200 6040 12264
rect 6104 12200 6112 12264
rect 5792 11731 6112 12200
rect 5792 11495 5834 11731
rect 6070 11495 6112 11731
rect 5792 11176 6112 11495
rect 5792 11112 5800 11176
rect 5864 11112 5880 11176
rect 5944 11112 5960 11176
rect 6024 11112 6040 11176
rect 6104 11112 6112 11176
rect 5792 10088 6112 11112
rect 5792 10024 5800 10088
rect 5864 10024 5880 10088
rect 5944 10024 5960 10088
rect 6024 10024 6040 10088
rect 6104 10024 6112 10088
rect 5792 9000 6112 10024
rect 5792 8936 5800 9000
rect 5864 8936 5880 9000
rect 5944 8936 5960 9000
rect 6024 8936 6040 9000
rect 6104 8936 6112 9000
rect 5792 7912 6112 8936
rect 5792 7848 5800 7912
rect 5864 7848 5880 7912
rect 5944 7848 5960 7912
rect 6024 7848 6040 7912
rect 6104 7848 6112 7912
rect 5792 6848 6112 7848
rect 5792 6824 5834 6848
rect 6070 6824 6112 6848
rect 5792 6760 5800 6824
rect 6104 6760 6112 6824
rect 5792 6612 5834 6760
rect 6070 6612 6112 6760
rect 5792 5736 6112 6612
rect 5792 5672 5800 5736
rect 5864 5672 5880 5736
rect 5944 5672 5960 5736
rect 6024 5672 6040 5736
rect 6104 5672 6112 5736
rect 5792 4648 6112 5672
rect 5792 4584 5800 4648
rect 5864 4584 5880 4648
rect 5944 4584 5960 4648
rect 6024 4584 6040 4648
rect 6104 4584 6112 4648
rect 5792 3560 6112 4584
rect 5792 3496 5800 3560
rect 5864 3496 5880 3560
rect 5944 3496 5960 3560
rect 6024 3496 6040 3560
rect 6104 3496 6112 3560
rect 5792 2472 6112 3496
rect 5792 2408 5800 2472
rect 5864 2408 5880 2472
rect 5944 2408 5960 2472
rect 6024 2408 6040 2472
rect 6104 2408 6112 2472
rect 5792 1848 6112 2408
rect 7271 16072 7591 16088
rect 7271 16008 7279 16072
rect 7343 16008 7359 16072
rect 7423 16008 7439 16072
rect 7503 16008 7519 16072
rect 7583 16008 7591 16072
rect 7271 14984 7591 16008
rect 7271 14920 7279 14984
rect 7343 14920 7359 14984
rect 7423 14920 7439 14984
rect 7503 14920 7519 14984
rect 7583 14920 7591 14984
rect 7271 14172 7591 14920
rect 7271 13936 7313 14172
rect 7549 13936 7591 14172
rect 7271 13896 7591 13936
rect 7271 13832 7279 13896
rect 7343 13832 7359 13896
rect 7423 13832 7439 13896
rect 7503 13832 7519 13896
rect 7583 13832 7591 13896
rect 7271 12808 7591 13832
rect 7271 12744 7279 12808
rect 7343 12744 7359 12808
rect 7423 12744 7439 12808
rect 7503 12744 7519 12808
rect 7583 12744 7591 12808
rect 7271 11720 7591 12744
rect 7271 11656 7279 11720
rect 7343 11656 7359 11720
rect 7423 11656 7439 11720
rect 7503 11656 7519 11720
rect 7583 11656 7591 11720
rect 7271 10632 7591 11656
rect 7271 10568 7279 10632
rect 7343 10568 7359 10632
rect 7423 10568 7439 10632
rect 7503 10568 7519 10632
rect 7583 10568 7591 10632
rect 7271 9544 7591 10568
rect 7271 9480 7279 9544
rect 7343 9480 7359 9544
rect 7423 9480 7439 9544
rect 7503 9480 7519 9544
rect 7583 9480 7591 9544
rect 7271 9290 7591 9480
rect 7271 9054 7313 9290
rect 7549 9054 7591 9290
rect 7271 8456 7591 9054
rect 7271 8392 7279 8456
rect 7343 8392 7359 8456
rect 7423 8392 7439 8456
rect 7503 8392 7519 8456
rect 7583 8392 7591 8456
rect 7271 7368 7591 8392
rect 7271 7304 7279 7368
rect 7343 7304 7359 7368
rect 7423 7304 7439 7368
rect 7503 7304 7519 7368
rect 7583 7304 7591 7368
rect 7271 6280 7591 7304
rect 7271 6216 7279 6280
rect 7343 6216 7359 6280
rect 7423 6216 7439 6280
rect 7503 6216 7519 6280
rect 7583 6216 7591 6280
rect 7271 5192 7591 6216
rect 7271 5128 7279 5192
rect 7343 5128 7359 5192
rect 7423 5128 7439 5192
rect 7503 5128 7519 5192
rect 7583 5128 7591 5192
rect 7271 4407 7591 5128
rect 7271 4171 7313 4407
rect 7549 4171 7591 4407
rect 7271 4104 7591 4171
rect 7271 4040 7279 4104
rect 7343 4040 7359 4104
rect 7423 4040 7439 4104
rect 7503 4040 7519 4104
rect 7583 4040 7591 4104
rect 7271 3016 7591 4040
rect 7271 2952 7279 3016
rect 7343 2952 7359 3016
rect 7423 2952 7439 3016
rect 7503 2952 7519 3016
rect 7583 2952 7591 3016
rect 7271 1928 7591 2952
rect 7271 1864 7279 1928
rect 7343 1864 7359 1928
rect 7423 1864 7439 1928
rect 7503 1864 7519 1928
rect 7583 1864 7591 1928
rect 7271 1848 7591 1864
<< via4 >>
rect 1398 13936 1634 14172
rect 1398 9054 1634 9290
rect 1398 4171 1634 4407
rect 2877 11495 3113 11731
rect 2877 6824 3113 6848
rect 2877 6760 2907 6824
rect 2907 6760 2923 6824
rect 2923 6760 2987 6824
rect 2987 6760 3003 6824
rect 3003 6760 3067 6824
rect 3067 6760 3083 6824
rect 3083 6760 3113 6824
rect 2877 6612 3113 6760
rect 4356 13936 4592 14172
rect 4356 9054 4592 9290
rect 4356 4171 4592 4407
rect 5834 11495 6070 11731
rect 5834 6824 6070 6848
rect 5834 6760 5864 6824
rect 5864 6760 5880 6824
rect 5880 6760 5944 6824
rect 5944 6760 5960 6824
rect 5960 6760 6024 6824
rect 6024 6760 6040 6824
rect 6040 6760 6070 6824
rect 5834 6612 6070 6760
rect 7313 13936 7549 14172
rect 7313 9054 7549 9290
rect 7313 4171 7549 4407
<< metal5 >>
rect 38 14172 8870 14214
rect 38 13936 1398 14172
rect 1634 13936 4356 14172
rect 4592 13936 7313 14172
rect 7549 13936 8870 14172
rect 38 13894 8870 13936
rect 38 11731 8870 11773
rect 38 11495 2877 11731
rect 3113 11495 5834 11731
rect 6070 11495 8870 11731
rect 38 11453 8870 11495
rect 38 9290 8870 9332
rect 38 9054 1398 9290
rect 1634 9054 4356 9290
rect 4592 9054 7313 9290
rect 7549 9054 8870 9290
rect 38 9012 8870 9054
rect 38 6848 8870 6891
rect 38 6612 2877 6848
rect 3113 6612 5834 6848
rect 6070 6612 8870 6848
rect 38 6570 8870 6612
rect 38 4407 8870 4449
rect 38 4171 1398 4407
rect 1634 4171 4356 4407
rect 4592 4171 7313 4407
rect 7549 4171 8870 4407
rect 38 4129 8870 4171
use sky130_fd_sc_hd__conb_1  gpio_logic_high
timestamp 1606789160
transform 1 0 7122 0 1 15496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606789160
transform -1 0 8870 0 1 15496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_75
timestamp 1606789160
transform 1 0 6938 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_80
timestamp 1606789160
transform 1 0 7398 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_92
timestamp 1606789160
transform 1 0 8502 0 1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606789160
transform 1 0 5742 0 1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_56
timestamp 1606789160
transform 1 0 5190 0 1 15496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_63
timestamp 1606789160
transform 1 0 5834 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606789160
transform 1 0 2890 0 1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_27
timestamp 1606789160
transform 1 0 2522 0 1 15496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_32
timestamp 1606789160
transform 1 0 2982 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_44
timestamp 1606789160
transform 1 0 4086 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606789160
transform 1 0 38 0 1 15496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1606789160
transform 1 0 314 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1606789160
transform 1 0 1418 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1606789160
transform 1 0 7490 0 -1 15496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606789160
transform -1 0 8870 0 -1 15496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_80
timestamp 1606789160
transform 1 0 7398 0 -1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1606789160
transform 1 0 7858 0 -1 15496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606789160
transform 1 0 5650 0 -1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_51
timestamp 1606789160
transform 1 0 4730 0 -1 15496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_59
timestamp 1606789160
transform 1 0 5466 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_62
timestamp 1606789160
transform 1 0 5742 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_74
timestamp 1606789160
transform 1 0 6846 0 -1 15496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_27
timestamp 1606789160
transform 1 0 2522 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_39
timestamp 1606789160
transform 1 0 3626 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606789160
transform 1 0 38 0 -1 15496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1606789160
transform 1 0 314 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1606789160
transform 1 0 1418 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1606789160
transform 1 0 7398 0 1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606789160
transform -1 0 8870 0 1 14408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606789160
transform 1 0 8502 0 1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_84
timestamp 1606789160
transform 1 0 7766 0 1 14408
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1606789160
transform 1 0 6294 0 1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_56
timestamp 1606789160
transform 1 0 5190 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_72
timestamp 1606789160
transform 1 0 6662 0 1 14408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606789160
transform 1 0 2890 0 1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_27
timestamp 1606789160
transform 1 0 2522 0 1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_32
timestamp 1606789160
transform 1 0 2982 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_44
timestamp 1606789160
transform 1 0 4086 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606789160
transform 1 0 38 0 1 14408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1606789160
transform 1 0 314 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1606789160
transform 1 0 1418 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606789160
transform -1 0 8870 0 -1 14408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1606789160
transform 1 0 7858 0 -1 14408
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_8  gpio_in_buf
timestamp 1606789160
transform 1 0 6202 0 -1 14408
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606789160
transform 1 0 5650 0 -1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_51
timestamp 1606789160
transform 1 0 4730 0 -1 14408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_59
timestamp 1606789160
transform 1 0 5466 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_62
timestamp 1606789160
transform 1 0 5742 0 -1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_66
timestamp 1606789160
transform 1 0 6110 0 -1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_27
timestamp 1606789160
transform 1 0 2522 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_39
timestamp 1606789160
transform 1 0 3626 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606789160
transform 1 0 38 0 -1 14408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1606789160
transform 1 0 314 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1606789160
transform 1 0 1418 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606789160
transform -1 0 8870 0 1 13320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606789160
transform 1 0 8502 0 1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_84
timestamp 1606789160
transform 1 0 7766 0 1 13320
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _078_
timestamp 1606789160
transform 1 0 4638 0 1 13320
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _106_
timestamp 1606789160
transform 1 0 5650 0 1 13320
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_8  FILLER_21_53
timestamp 1606789160
transform 1 0 4914 0 1 13320
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606789160
transform 1 0 2890 0 1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_27
timestamp 1606789160
transform 1 0 2522 0 1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_32
timestamp 1606789160
transform 1 0 2982 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_44
timestamp 1606789160
transform 1 0 4086 0 1 13320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606789160
transform 1 0 38 0 1 13320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1606789160
transform 1 0 314 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1606789160
transform 1 0 1418 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606789160
transform -1 0 8870 0 1 12232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606789160
transform -1 0 8870 0 -1 13320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606789160
transform 1 0 8502 0 1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_84
timestamp 1606789160
transform 1 0 7766 0 1 12232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_85
timestamp 1606789160
transform 1 0 7858 0 -1 13320
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _103_
timestamp 1606789160
transform 1 0 5650 0 1 12232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _105_
timestamp 1606789160
transform 1 0 5742 0 -1 13320
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606789160
transform 1 0 5650 0 -1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_53
timestamp 1606789160
transform 1 0 4914 0 1 12232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_53
timestamp 1606789160
transform 1 0 4914 0 -1 13320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_27
timestamp 1606789160
transform 1 0 2522 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _039_
timestamp 1606789160
transform 1 0 4270 0 1 12232
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1606789160
transform 1 0 4546 0 -1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_serial_clock
timestamp 1606789160
transform 1 0 3994 0 -1 13320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_38
timestamp 1606789160
transform 1 0 3534 0 1 12232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_39
timestamp 1606789160
transform 1 0 3626 0 -1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_46
timestamp 1606789160
transform 1 0 4270 0 -1 13320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1606789160
transform 1 0 3166 0 1 12232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606789160
transform 1 0 2890 0 1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_27
timestamp 1606789160
transform 1 0 2522 0 1 12232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_32
timestamp 1606789160
transform 1 0 2982 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606789160
transform 1 0 38 0 1 12232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606789160
transform 1 0 38 0 -1 13320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1606789160
transform 1 0 314 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1606789160
transform 1 0 1418 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1606789160
transform 1 0 314 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1606789160
transform 1 0 1418 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606789160
transform -1 0 8870 0 -1 12232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1606789160
transform 1 0 7858 0 -1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_87
timestamp 1606789160
transform 1 0 8042 0 -1 12232
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_4  _095_
timestamp 1606789160
transform 1 0 5742 0 -1 12232
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606789160
transform 1 0 5650 0 -1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_53
timestamp 1606789160
transform 1 0 4914 0 -1 12232
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _107_
timestamp 1606789160
transform 1 0 2798 0 -1 12232
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  FILLER_18_27
timestamp 1606789160
transform 1 0 2522 0 -1 12232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606789160
transform 1 0 38 0 -1 12232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1606789160
transform 1 0 314 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1606789160
transform 1 0 1418 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606789160
transform -1 0 8870 0 1 11144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606789160
transform 1 0 8502 0 1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_84
timestamp 1606789160
transform 1 0 7766 0 1 11144
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _091_
timestamp 1606789160
transform 1 0 5650 0 1 11144
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_8  FILLER_17_53
timestamp 1606789160
transform 1 0 4914 0 1 11144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _053_
timestamp 1606789160
transform 1 0 2982 0 1 11144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _077_
timestamp 1606789160
transform 1 0 4086 0 1 11144
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606789160
transform 1 0 2890 0 1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_36
timestamp 1606789160
transform 1 0 3350 0 1 11144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1606789160
transform 1 0 1786 0 1 11144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606789160
transform 1 0 38 0 1 11144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1606789160
transform 1 0 314 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_15
timestamp 1606789160
transform 1 0 1418 0 1 11144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_23
timestamp 1606789160
transform 1 0 2154 0 1 11144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606789160
transform -1 0 8870 0 -1 11144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_85
timestamp 1606789160
transform 1 0 7858 0 -1 11144
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _085_
timestamp 1606789160
transform 1 0 5742 0 -1 11144
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606789160
transform 1 0 5650 0 -1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_53
timestamp 1606789160
transform 1 0 4914 0 -1 11144
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _104_
timestamp 1606789160
transform 1 0 2798 0 -1 11144
box -38 -48 2154 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1606789160
transform 1 0 1694 0 -1 11144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1606789160
transform 1 0 590 0 -1 11144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606789160
transform 1 0 38 0 -1 11144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1606789160
transform 1 0 314 0 -1 11144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_10
timestamp 1606789160
transform 1 0 958 0 -1 11144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_22
timestamp 1606789160
transform 1 0 2062 0 -1 11144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606789160
transform -1 0 8870 0 1 10056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606789160
transform 1 0 8502 0 1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_84
timestamp 1606789160
transform 1 0 7766 0 1 10056
box -38 -48 774 592
use sky130_fd_sc_hd__dfstp_4  _088_
timestamp 1606789160
transform 1 0 5558 0 1 10056
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_8  FILLER_15_52
timestamp 1606789160
transform 1 0 4822 0 1 10056
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_4  _071_
timestamp 1606789160
transform 1 0 3258 0 1 10056
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606789160
transform 1 0 2890 0 1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_32
timestamp 1606789160
transform 1 0 2982 0 1 10056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1606789160
transform 1 0 406 0 1 10056
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _079_
timestamp 1606789160
transform 1 0 1510 0 1 10056
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606789160
transform 1 0 38 0 1 10056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1606789160
transform 1 0 314 0 1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_8
timestamp 1606789160
transform 1 0 774 0 1 10056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_23
timestamp 1606789160
transform 1 0 2154 0 1 10056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606789160
transform -1 0 8870 0 1 8968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606789160
transform -1 0 8870 0 -1 10056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606789160
transform 1 0 8502 0 1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_84
timestamp 1606789160
transform 1 0 7766 0 1 8968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_85
timestamp 1606789160
transform 1 0 7858 0 -1 10056
box -38 -48 774 592
use sky130_fd_sc_hd__dfstp_4  _082_
timestamp 1606789160
transform 1 0 5558 0 1 8968
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrtp_4  _084_
timestamp 1606789160
transform 1 0 5742 0 -1 10056
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606789160
transform 1 0 5650 0 -1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_53
timestamp 1606789160
transform 1 0 4914 0 -1 10056
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _096_
timestamp 1606789160
transform 1 0 2798 0 -1 10056
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606789160
transform 1 0 2890 0 1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock
timestamp 1606789160
transform 1 0 3718 0 1 8968
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_13_32
timestamp 1606789160
transform 1 0 2982 0 1 8968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _040_
timestamp 1606789160
transform 1 0 1694 0 -1 10056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _042_
timestamp 1606789160
transform 1 0 1786 0 1 8968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_23
timestamp 1606789160
transform 1 0 2154 0 1 8968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_22
timestamp 1606789160
transform 1 0 2062 0 -1 10056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_11
timestamp 1606789160
transform 1 0 1050 0 1 8968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_10
timestamp 1606789160
transform 1 0 958 0 -1 10056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _051_
timestamp 1606789160
transform 1 0 682 0 1 8968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _054_
timestamp 1606789160
transform 1 0 590 0 -1 10056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606789160
transform 1 0 38 0 1 8968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606789160
transform 1 0 38 0 -1 10056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1606789160
transform 1 0 314 0 1 8968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1606789160
transform 1 0 314 0 -1 10056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606789160
transform -1 0 8870 0 -1 8968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 1606789160
transform 1 0 7858 0 -1 8968
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _083_
timestamp 1606789160
transform 1 0 5742 0 -1 8968
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606789160
transform 1 0 5650 0 -1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_53
timestamp 1606789160
transform 1 0 4914 0 -1 8968
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _097_
timestamp 1606789160
transform 1 0 2798 0 -1 8968
box -38 -48 2154 592
use sky130_fd_sc_hd__buf_2  _041_
timestamp 1606789160
transform 1 0 1694 0 -1 8968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _046_
timestamp 1606789160
transform 1 0 590 0 -1 8968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606789160
transform 1 0 38 0 -1 8968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 1606789160
transform 1 0 314 0 -1 8968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_10
timestamp 1606789160
transform 1 0 958 0 -1 8968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_22
timestamp 1606789160
transform 1 0 2062 0 -1 8968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606789160
transform -1 0 8870 0 1 7880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606789160
transform 1 0 8502 0 1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_84
timestamp 1606789160
transform 1 0 7766 0 1 7880
box -38 -48 774 592
use sky130_fd_sc_hd__dfstp_4  _089_
timestamp 1606789160
transform 1 0 5558 0 1 7880
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_8  FILLER_11_52
timestamp 1606789160
transform 1 0 4822 0 1 7880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _070_
timestamp 1606789160
transform 1 0 2982 0 1 7880
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_4  _076_
timestamp 1606789160
transform 1 0 3258 0 1 7880
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606789160
transform 1 0 2890 0 1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _044_
timestamp 1606789160
transform 1 0 1786 0 1 7880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _049_
timestamp 1606789160
transform 1 0 682 0 1 7880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606789160
transform 1 0 38 0 1 7880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1606789160
transform 1 0 314 0 1 7880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_11
timestamp 1606789160
transform 1 0 1050 0 1 7880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_23
timestamp 1606789160
transform 1 0 2154 0 1 7880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606789160
transform -1 0 8870 0 -1 7880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1606789160
transform 1 0 7858 0 -1 7880
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _086_
timestamp 1606789160
transform 1 0 5742 0 -1 7880
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606789160
transform 1 0 5650 0 -1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_53
timestamp 1606789160
transform 1 0 4914 0 -1 7880
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _098_
timestamp 1606789160
transform 1 0 2798 0 -1 7880
box -38 -48 2154 592
use sky130_fd_sc_hd__buf_2  _045_
timestamp 1606789160
transform 1 0 1694 0 -1 7880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _052_
timestamp 1606789160
transform 1 0 590 0 -1 7880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606789160
transform 1 0 38 0 -1 7880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1606789160
transform 1 0 314 0 -1 7880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_10
timestamp 1606789160
transform 1 0 958 0 -1 7880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_22
timestamp 1606789160
transform 1 0 2062 0 -1 7880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606789160
transform -1 0 8870 0 1 6792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606789160
transform 1 0 8502 0 1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_84
timestamp 1606789160
transform 1 0 7766 0 1 6792
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _087_
timestamp 1606789160
transform 1 0 5650 0 1 6792
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_8  FILLER_9_53
timestamp 1606789160
transform 1 0 4914 0 1 6792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _043_
timestamp 1606789160
transform 1 0 2522 0 1 6792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _073_
timestamp 1606789160
transform 1 0 4086 0 1 6792
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _075_
timestamp 1606789160
transform 1 0 3258 0 1 6792
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1606789160
transform 1 0 2890 0 1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_32
timestamp 1606789160
transform 1 0 2982 0 1 6792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _047_
timestamp 1606789160
transform 1 0 1786 0 1 6792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1606789160
transform 1 0 682 0 1 6792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606789160
transform 1 0 38 0 1 6792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1606789160
transform 1 0 314 0 1 6792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_11
timestamp 1606789160
transform 1 0 1050 0 1 6792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_23
timestamp 1606789160
transform 1 0 2154 0 1 6792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606789160
transform -1 0 8870 0 -1 6792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85
timestamp 1606789160
transform 1 0 7858 0 -1 6792
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _090_
timestamp 1606789160
transform 1 0 5742 0 -1 6792
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1606789160
transform 1 0 5650 0 -1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_53
timestamp 1606789160
transform 1 0 4914 0 -1 6792
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _099_
timestamp 1606789160
transform 1 0 2798 0 -1 6792
box -38 -48 2154 592
use sky130_fd_sc_hd__buf_2  _055_
timestamp 1606789160
transform 1 0 1694 0 -1 6792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606789160
transform 1 0 38 0 -1 6792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1606789160
transform 1 0 314 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_15
timestamp 1606789160
transform 1 0 1418 0 -1 6792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_22
timestamp 1606789160
transform 1 0 2062 0 -1 6792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606789160
transform -1 0 8870 0 -1 5704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606789160
transform -1 0 8870 0 1 5704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1606789160
transform 1 0 8502 0 1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_85
timestamp 1606789160
transform 1 0 7858 0 -1 5704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_84
timestamp 1606789160
transform 1 0 7766 0 1 5704
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _092_
timestamp 1606789160
transform 1 0 5742 0 -1 5704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _093_
timestamp 1606789160
transform 1 0 5650 0 1 5704
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1606789160
transform 1 0 5650 0 -1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_53
timestamp 1606789160
transform 1 0 4914 0 -1 5704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_53
timestamp 1606789160
transform 1 0 4914 0 1 5704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _050_
timestamp 1606789160
transform 1 0 3166 0 1 5704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _074_
timestamp 1606789160
transform 1 0 4270 0 1 5704
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_4  _102_
timestamp 1606789160
transform 1 0 2798 0 -1 5704
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1606789160
transform 1 0 2890 0 1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_27
timestamp 1606789160
transform 1 0 2522 0 -1 5704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_32
timestamp 1606789160
transform 1 0 2982 0 1 5704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_38
timestamp 1606789160
transform 1 0 3534 0 1 5704
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _072_
timestamp 1606789160
transform 1 0 1878 0 1 5704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606789160
transform 1 0 38 0 -1 5704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606789160
transform 1 0 38 0 1 5704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1606789160
transform 1 0 314 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1606789160
transform 1 0 1418 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1606789160
transform 1 0 314 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_15
timestamp 1606789160
transform 1 0 1418 0 1 5704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_19
timestamp 1606789160
transform 1 0 1786 0 1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_23
timestamp 1606789160
transform 1 0 2154 0 1 5704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606789160
transform -1 0 8870 0 1 4616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1606789160
transform 1 0 8502 0 1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_84
timestamp 1606789160
transform 1 0 7766 0 1 4616
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _094_
timestamp 1606789160
transform 1 0 5650 0 1 4616
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_8  FILLER_5_53
timestamp 1606789160
transform 1 0 4914 0 1 4616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _048_
timestamp 1606789160
transform 1 0 4546 0 1 4616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1606789160
transform 1 0 3442 0 1 4616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1606789160
transform 1 0 2890 0 1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1606789160
transform 1 0 2522 0 1 4616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_32
timestamp 1606789160
transform 1 0 2982 0 1 4616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_36
timestamp 1606789160
transform 1 0 3350 0 1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_41
timestamp 1606789160
transform 1 0 3810 0 1 4616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606789160
transform 1 0 38 0 1 4616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1606789160
transform 1 0 314 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1606789160
transform 1 0 1418 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606789160
transform -1 0 8870 0 -1 4616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp 1606789160
transform 1 0 7858 0 -1 4616
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _100_
timestamp 1606789160
transform 1 0 5742 0 -1 4616
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1606789160
transform 1 0 5650 0 -1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_53
timestamp 1606789160
transform 1 0 4914 0 -1 4616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1606789160
transform 1 0 4546 0 -1 4616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_serial_clock
timestamp 1606789160
transform 1 0 3718 0 -1 4616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_27
timestamp 1606789160
transform 1 0 2522 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_39
timestamp 1606789160
transform 1 0 3626 0 -1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_43
timestamp 1606789160
transform 1 0 3994 0 -1 4616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606789160
transform 1 0 38 0 -1 4616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1606789160
transform 1 0 314 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1606789160
transform 1 0 1418 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606789160
transform -1 0 8870 0 1 3528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1606789160
transform 1 0 8502 0 1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_84
timestamp 1606789160
transform 1 0 7766 0 1 3528
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _101_
timestamp 1606789160
transform 1 0 5650 0 1 3528
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_3_56
timestamp 1606789160
transform 1 0 5190 0 1 3528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_60
timestamp 1606789160
transform 1 0 5558 0 1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1606789160
transform 1 0 2890 0 1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1606789160
transform 1 0 2522 0 1 3528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_32
timestamp 1606789160
transform 1 0 2982 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1606789160
transform 1 0 4086 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606789160
transform 1 0 38 0 1 3528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1606789160
transform 1 0 314 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1606789160
transform 1 0 1418 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _080_
timestamp 1606789160
transform 1 0 7214 0 -1 3528
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606789160
transform -1 0 8870 0 -1 3528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1606789160
transform 1 0 7858 0 -1 3528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1606789160
transform 1 0 6110 0 -1 3528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1606789160
transform 1 0 5650 0 -1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_51
timestamp 1606789160
transform 1 0 4730 0 -1 3528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_59
timestamp 1606789160
transform 1 0 5466 0 -1 3528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_62
timestamp 1606789160
transform 1 0 5742 0 -1 3528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_70
timestamp 1606789160
transform 1 0 6478 0 -1 3528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_27
timestamp 1606789160
transform 1 0 2522 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_39
timestamp 1606789160
transform 1 0 3626 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606789160
transform 1 0 38 0 -1 3528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1606789160
transform 1 0 314 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1606789160
transform 1 0 1418 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1606789160
transform 1 0 7398 0 1 2440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1606789160
transform 1 0 7490 0 -1 2440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606789160
transform -1 0 8870 0 -1 2440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606789160
transform -1 0 8870 0 1 2440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1606789160
transform 1 0 8502 0 1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75
timestamp 1606789160
transform 1 0 6938 0 -1 2440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1606789160
transform 1 0 7858 0 -1 2440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_84
timestamp 1606789160
transform 1 0 7766 0 1 2440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1606789160
transform 1 0 5742 0 -1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56
timestamp 1606789160
transform 1 0 5190 0 -1 2440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1606789160
transform 1 0 5834 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_56
timestamp 1606789160
transform 1 0 5190 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_68
timestamp 1606789160
transform 1 0 6294 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1606789160
transform 1 0 2890 0 -1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1606789160
transform 1 0 2890 0 1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1606789160
transform 1 0 2522 0 -1 2440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1606789160
transform 1 0 2982 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1606789160
transform 1 0 4086 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1606789160
transform 1 0 2522 0 1 2440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_32
timestamp 1606789160
transform 1 0 2982 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_44
timestamp 1606789160
transform 1 0 4086 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1606789160
transform 1 0 38 0 -1 2440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606789160
transform 1 0 38 0 1 2440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1606789160
transform 1 0 314 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1606789160
transform 1 0 1418 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1606789160
transform 1 0 314 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1606789160
transform 1 0 1418 0 1 2440
box -38 -48 1142 592
<< labels >>
rlabel metal3 s 9934 0 33934 120 4 mgmt_gpio_in
port 1 nsew
rlabel metal3 s 9934 680 33934 800 4 mgmt_gpio_oeb
port 2 nsew
rlabel metal3 s 9934 1496 33934 1616 4 mgmt_gpio_out
port 3 nsew
rlabel metal3 s 9934 2312 33934 2432 4 pad_gpio_ana_en
port 4 nsew
rlabel metal3 s 9934 3128 33934 3248 4 pad_gpio_ana_pol
port 5 nsew
rlabel metal3 s 9934 3944 33934 4064 4 pad_gpio_ana_sel
port 6 nsew
rlabel metal3 s 9934 4760 33934 4880 4 pad_gpio_dm[0]
port 7 nsew
rlabel metal3 s 9934 5440 33934 5560 4 pad_gpio_dm[1]
port 8 nsew
rlabel metal3 s 9934 6256 33934 6376 4 pad_gpio_dm[2]
port 9 nsew
rlabel metal3 s 9934 7072 33934 7192 4 pad_gpio_holdover
port 10 nsew
rlabel metal3 s 9934 7888 33934 8008 4 pad_gpio_ib_mode_sel
port 11 nsew
rlabel metal3 s 9934 8704 33934 8824 4 pad_gpio_in
port 12 nsew
rlabel metal3 s 9934 9520 33934 9640 4 pad_gpio_inenb
port 13 nsew
rlabel metal3 s 9934 10200 33934 10320 4 pad_gpio_out
port 14 nsew
rlabel metal3 s 9934 11016 33934 11136 4 pad_gpio_outenb
port 15 nsew
rlabel metal3 s 9934 11832 33934 11952 4 pad_gpio_slow_sel
port 16 nsew
rlabel metal3 s 9934 12648 33934 12768 4 pad_gpio_vtrip_sel
port 17 nsew
rlabel metal3 s 9934 13464 33934 13584 4 resetn
port 18 nsew
rlabel metal3 s 9934 14280 33934 14400 4 serial_clock
port 19 nsew
rlabel metal3 s 9934 14960 33934 15080 4 serial_data_in
port 20 nsew
rlabel metal3 s 9934 15776 33934 15896 4 serial_data_out
port 21 nsew
rlabel metal3 s 9934 16592 33934 16712 4 user_gpio_in
port 22 nsew
rlabel metal3 s 9934 17408 33934 17528 4 user_gpio_oeb
port 23 nsew
rlabel metal3 s 9934 18224 33934 18344 4 user_gpio_out
port 24 nsew
rlabel metal5 s 38 4129 8870 4449 4 VPWR
port 25 nsew
rlabel metal5 s 38 6571 8870 6891 4 VGND
port 26 nsew
<< properties >>
string FIXED_BBOX 0 0 33934 18344
string GDS_FILE gpio_control_block.gds
string GDS_END 380356
string GDS_START 138912
<< end >>
