magic
tech sky130A
magscale 1 2
timestamp 1611581575
<< locali >>
rect 7573 7191 7607 7497
rect 765 6443 799 6817
rect 6653 4539 6687 4641
<< viali >>
rect 121 11237 155 11271
rect 2789 11169 2823 11203
rect 3157 11169 3191 11203
rect 3709 11169 3743 11203
rect 4445 11169 4479 11203
rect 4997 11169 5031 11203
rect 6377 11169 6411 11203
rect 4353 11101 4387 11135
rect 6469 11101 6503 11135
rect 3341 11033 3375 11067
rect 3525 11033 3559 11067
rect 2973 10965 3007 10999
rect 4629 10965 4663 10999
rect 6653 10761 6687 10795
rect 1593 10625 1627 10659
rect 1961 10625 1995 10659
rect 1685 10557 1719 10591
rect 4077 10557 4111 10591
rect 4445 10557 4479 10591
rect 6561 10557 6595 10591
rect 3709 10489 3743 10523
rect 4721 10489 4755 10523
rect 6469 10489 6503 10523
rect 4261 10421 4295 10455
rect 6377 10217 6411 10251
rect 5549 10149 5583 10183
rect 3709 10081 3743 10115
rect 5733 10081 5767 10115
rect 6285 10081 6319 10115
rect 1225 10013 1259 10047
rect 1501 10013 1535 10047
rect 3249 10013 3283 10047
rect 3341 10013 3375 10047
rect 5089 10013 5123 10047
rect 5825 9877 5859 9911
rect 2237 9537 2271 9571
rect 5917 9537 5951 9571
rect 1869 9469 1903 9503
rect 2697 9469 2731 9503
rect 2973 9469 3007 9503
rect 3157 9469 3191 9503
rect 3433 9469 3467 9503
rect 3709 9469 3743 9503
rect 3893 9469 3927 9503
rect 6009 9469 6043 9503
rect 6377 9469 6411 9503
rect 4169 9401 4203 9435
rect 2053 9333 2087 9367
rect 6193 9333 6227 9367
rect 6469 9333 6503 9367
rect 5641 9129 5675 9163
rect 6009 9129 6043 9163
rect 1961 8993 1995 9027
rect 2145 8993 2179 9027
rect 2329 8993 2363 9027
rect 2697 8993 2731 9027
rect 5089 8993 5123 9027
rect 5457 8993 5491 9027
rect 5825 8993 5859 9027
rect 6285 8993 6319 9027
rect 1409 8925 1443 8959
rect 2789 8925 2823 8959
rect 2973 8925 3007 8959
rect 3249 8925 3283 8959
rect 4997 8925 5031 8959
rect 5273 8857 5307 8891
rect 6377 8789 6411 8823
rect 6653 8585 6687 8619
rect 1225 8449 1259 8483
rect 1501 8449 1535 8483
rect 3341 8381 3375 8415
rect 3985 8381 4019 8415
rect 4353 8381 4387 8415
rect 6469 8381 6503 8415
rect 3249 8313 3283 8347
rect 4629 8313 4663 8347
rect 6377 8313 6411 8347
rect 3525 8245 3559 8279
rect 4169 8245 4203 8279
rect 6101 8041 6135 8075
rect 6377 8041 6411 8075
rect 1501 7973 1535 8007
rect 3341 7905 3375 7939
rect 3893 7905 3927 7939
rect 4353 7905 4387 7939
rect 6193 7905 6227 7939
rect 1225 7837 1259 7871
rect 3249 7837 3283 7871
rect 3985 7837 4019 7871
rect 3709 7769 3743 7803
rect 3525 7701 3559 7735
rect 7573 7497 7607 7531
rect 1593 7361 1627 7395
rect 4169 7361 4203 7395
rect 1317 7293 1351 7327
rect 3433 7293 3467 7327
rect 3893 7293 3927 7327
rect 6193 7293 6227 7327
rect 3341 7225 3375 7259
rect 5917 7225 5951 7259
rect 6009 7225 6043 7259
rect 3617 7157 3651 7191
rect 6285 7157 6319 7191
rect 7573 7157 7607 7191
rect 2973 6885 3007 6919
rect 5825 6885 5859 6919
rect 5917 6885 5951 6919
rect 765 6817 799 6851
rect 1225 6817 1259 6851
rect 3065 6817 3099 6851
rect 5181 6817 5215 6851
rect 3341 6749 3375 6783
rect 5089 6749 5123 6783
rect 6469 6749 6503 6783
rect 5365 6681 5399 6715
rect 765 6409 799 6443
rect 1501 6273 1535 6307
rect 4629 6273 4663 6307
rect 1225 6205 1259 6239
rect 3341 6205 3375 6239
rect 3893 6205 3927 6239
rect 4353 6205 4387 6239
rect 6469 6205 6503 6239
rect 3249 6137 3283 6171
rect 6377 6137 6411 6171
rect 3525 6069 3559 6103
rect 4077 6069 4111 6103
rect 6653 6069 6687 6103
rect 5825 5865 5859 5899
rect 3525 5729 3559 5763
rect 5549 5729 5583 5763
rect 5641 5729 5675 5763
rect 6009 5729 6043 5763
rect 1409 5661 1443 5695
rect 1685 5661 1719 5695
rect 3433 5661 3467 5695
rect 3801 5661 3835 5695
rect 6193 5525 6227 5559
rect 3525 5321 3559 5355
rect 1225 5185 1259 5219
rect 1501 5185 1535 5219
rect 4997 5185 5031 5219
rect 3341 5117 3375 5151
rect 3985 5117 4019 5151
rect 4629 5117 4663 5151
rect 3249 5049 3283 5083
rect 4169 4981 4203 5015
rect 6745 4981 6779 5015
rect 1593 4777 1627 4811
rect 2329 4777 2363 4811
rect 5273 4777 5307 4811
rect 1409 4641 1443 4675
rect 1777 4641 1811 4675
rect 2145 4641 2179 4675
rect 5089 4641 5123 4675
rect 5457 4641 5491 4675
rect 6009 4641 6043 4675
rect 6469 4641 6503 4675
rect 6653 4641 6687 4675
rect 2513 4573 2547 4607
rect 2789 4573 2823 4607
rect 4537 4573 4571 4607
rect 4813 4573 4847 4607
rect 4997 4505 5031 4539
rect 5549 4505 5583 4539
rect 6653 4505 6687 4539
rect 1961 4437 1995 4471
rect 5825 4437 5859 4471
rect 1488 4233 1522 4267
rect 3525 4233 3559 4267
rect 4156 4233 4190 4267
rect 1225 4097 1259 4131
rect 3893 4097 3927 4131
rect 5917 4097 5951 4131
rect 6009 4097 6043 4131
rect 3341 4029 3375 4063
rect 6193 4029 6227 4063
rect 6285 4029 6319 4063
rect 3249 3961 3283 3995
rect 6745 3961 6779 3995
rect 6193 3689 6227 3723
rect 2881 3621 2915 3655
rect 5825 3621 5859 3655
rect 4813 3553 4847 3587
rect 5181 3553 5215 3587
rect 5917 3553 5951 3587
rect 6101 3553 6135 3587
rect 2605 3485 2639 3519
rect 4629 3485 4663 3519
rect 4997 3349 5031 3383
rect 5365 3349 5399 3383
rect 1961 3009 1995 3043
rect 3709 3009 3743 3043
rect 4813 3009 4847 3043
rect 6285 3009 6319 3043
rect 1685 2941 1719 2975
rect 3893 2941 3927 2975
rect 4445 2941 4479 2975
rect 4077 2805 4111 2839
rect 3433 2601 3467 2635
rect 4813 2533 4847 2567
rect 6561 2533 6595 2567
rect 3249 2465 3283 2499
rect 4537 2465 4571 2499
<< metal1 >>
rect 12526 12724 12532 12776
rect 12584 12764 12590 12776
rect 14090 12764 14096 12776
rect 12584 12736 14096 12764
rect 12584 12724 12590 12736
rect 14090 12724 14096 12736
rect 14148 12724 14154 12776
rect 12434 12452 12440 12504
rect 12492 12492 12498 12504
rect 14182 12492 14188 12504
rect 12492 12464 14188 12492
rect 12492 12452 12498 12464
rect 14182 12452 14188 12464
rect 14240 12452 14246 12504
rect -1664 11462 506 11472
rect -1664 11386 -1610 11462
rect -1312 11386 506 11462
rect -1664 11376 506 11386
rect 626 11450 7084 11472
rect 626 11398 3598 11450
rect 3650 11398 3662 11450
rect 3714 11398 3726 11450
rect 3778 11398 3790 11450
rect 3842 11398 7084 11450
rect 626 11376 7084 11398
rect 1946 11296 1952 11348
rect 2004 11336 2010 11348
rect 14182 11336 14188 11348
rect 2004 11308 14188 11336
rect 2004 11296 2010 11308
rect 14182 11296 14188 11308
rect 14240 11296 14246 11348
rect 109 11271 167 11277
rect 109 11237 121 11271
rect 155 11268 167 11271
rect 155 11240 5028 11268
rect 155 11237 167 11240
rect 109 11231 167 11237
rect 2774 11160 2780 11212
rect 2832 11200 2838 11212
rect 3145 11203 3203 11209
rect 3145 11200 3157 11203
rect 2832 11172 3157 11200
rect 2832 11160 2838 11172
rect 3145 11169 3157 11172
rect 3191 11169 3203 11203
rect 3145 11163 3203 11169
rect 3697 11203 3755 11209
rect 3697 11169 3709 11203
rect 3743 11200 3755 11203
rect 3878 11200 3884 11212
rect 3743 11172 3884 11200
rect 3743 11169 3755 11172
rect 3697 11163 3755 11169
rect 3878 11160 3884 11172
rect 3936 11160 3942 11212
rect 4430 11200 4436 11212
rect 4391 11172 4436 11200
rect 4430 11160 4436 11172
rect 4488 11160 4494 11212
rect 5000 11209 5028 11240
rect 4985 11203 5043 11209
rect 4985 11169 4997 11203
rect 5031 11169 5043 11203
rect 6362 11200 6368 11212
rect 6323 11172 6368 11200
rect 4985 11163 5043 11169
rect 6362 11160 6368 11172
rect 6420 11160 6426 11212
rect 13722 11200 13728 11212
rect 6472 11172 13728 11200
rect 4341 11135 4399 11141
rect 4341 11132 4353 11135
rect 2746 11104 4353 11132
rect 1210 10956 1216 11008
rect 1268 10996 1274 11008
rect 2746 10996 2774 11104
rect 3326 11064 3332 11076
rect 3287 11036 3332 11064
rect 3326 11024 3332 11036
rect 3384 11024 3390 11076
rect 3528 11073 3556 11104
rect 4341 11101 4353 11104
rect 4387 11132 4399 11135
rect 5442 11132 5448 11144
rect 4387 11104 5448 11132
rect 4387 11101 4399 11104
rect 4341 11095 4399 11101
rect 5442 11092 5448 11104
rect 5500 11092 5506 11144
rect 6472 11141 6500 11172
rect 13722 11160 13728 11172
rect 13780 11160 13786 11212
rect 6457 11135 6515 11141
rect 6457 11101 6469 11135
rect 6503 11101 6515 11135
rect 6457 11095 6515 11101
rect 6638 11092 6644 11144
rect 6696 11132 6702 11144
rect 14090 11132 14096 11144
rect 6696 11104 14096 11132
rect 6696 11092 6702 11104
rect 14090 11092 14096 11104
rect 14148 11092 14154 11144
rect 3513 11067 3571 11073
rect 3513 11033 3525 11067
rect 3559 11033 3571 11067
rect 3513 11027 3571 11033
rect 2958 10996 2964 11008
rect 1268 10968 2774 10996
rect 2919 10968 2964 10996
rect 1268 10956 1274 10968
rect 2958 10956 2964 10968
rect 3016 10956 3022 11008
rect 4522 10956 4528 11008
rect 4580 10996 4586 11008
rect 4617 10999 4675 11005
rect 4617 10996 4629 10999
rect 4580 10968 4629 10996
rect 4580 10956 4586 10968
rect 4617 10965 4629 10968
rect 4663 10965 4675 10999
rect 4617 10959 4675 10965
rect -1048 10918 522 10928
rect -1048 10842 -950 10918
rect -652 10842 522 10918
rect -1048 10832 522 10842
rect 642 10906 7084 10928
rect 642 10854 2098 10906
rect 2150 10854 2162 10906
rect 2214 10854 2226 10906
rect 2278 10854 2290 10906
rect 2342 10854 5098 10906
rect 5150 10854 5162 10906
rect 5214 10854 5226 10906
rect 5278 10854 5290 10906
rect 5342 10854 7084 10906
rect 642 10832 7084 10854
rect 4430 10752 4436 10804
rect 4488 10792 4494 10804
rect 6641 10795 6699 10801
rect 6641 10792 6653 10795
rect 4488 10764 6653 10792
rect 4488 10752 4494 10764
rect 6641 10761 6653 10764
rect 6687 10761 6699 10795
rect 6641 10755 6699 10761
rect 1581 10659 1639 10665
rect 1581 10625 1593 10659
rect 1627 10656 1639 10659
rect 1946 10656 1952 10668
rect 1627 10628 1952 10656
rect 1627 10625 1639 10628
rect 1581 10619 1639 10625
rect 1946 10616 1952 10628
rect 2004 10616 2010 10668
rect 13262 10616 13268 10668
rect 13320 10656 13326 10668
rect 14090 10656 14096 10668
rect 13320 10628 14096 10656
rect 13320 10616 13326 10628
rect 14090 10616 14096 10628
rect 14148 10616 14154 10668
rect 1210 10548 1216 10600
rect 1268 10588 1274 10600
rect 1673 10591 1731 10597
rect 1673 10588 1685 10591
rect 1268 10560 1685 10588
rect 1268 10548 1274 10560
rect 1673 10557 1685 10560
rect 1719 10557 1731 10591
rect 4062 10588 4068 10600
rect 4023 10560 4068 10588
rect 1673 10551 1731 10557
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 4430 10588 4436 10600
rect 4391 10560 4436 10588
rect 4430 10548 4436 10560
rect 4488 10548 4494 10600
rect 6546 10588 6552 10600
rect 6459 10560 6552 10588
rect 6546 10548 6552 10560
rect 6604 10588 6610 10600
rect 14182 10588 14188 10600
rect 6604 10560 14188 10588
rect 6604 10548 6610 10560
rect 14182 10548 14188 10560
rect 14240 10548 14246 10600
rect 3326 10520 3332 10532
rect 3174 10492 3332 10520
rect 3326 10480 3332 10492
rect 3384 10480 3390 10532
rect 3418 10480 3424 10532
rect 3476 10520 3482 10532
rect 3697 10523 3755 10529
rect 3697 10520 3709 10523
rect 3476 10492 3709 10520
rect 3476 10480 3482 10492
rect 3697 10489 3709 10492
rect 3743 10489 3755 10523
rect 3697 10483 3755 10489
rect 4614 10480 4620 10532
rect 4672 10520 4678 10532
rect 4709 10523 4767 10529
rect 4709 10520 4721 10523
rect 4672 10492 4721 10520
rect 4672 10480 4678 10492
rect 4709 10489 4721 10492
rect 4755 10489 4767 10523
rect 6086 10520 6092 10532
rect 5934 10492 6092 10520
rect 4709 10483 4767 10489
rect 6086 10480 6092 10492
rect 6144 10480 6150 10532
rect 6457 10523 6515 10529
rect 6457 10489 6469 10523
rect 6503 10520 6515 10523
rect 14090 10520 14096 10532
rect 6503 10492 14096 10520
rect 6503 10489 6515 10492
rect 6457 10483 6515 10489
rect 14090 10480 14096 10492
rect 14148 10480 14154 10532
rect 4246 10452 4252 10464
rect 4207 10424 4252 10452
rect 4246 10412 4252 10424
rect 4304 10412 4310 10464
rect 920 10362 7084 10384
rect 920 10310 3598 10362
rect 3650 10310 3662 10362
rect 3714 10310 3726 10362
rect 3778 10310 3790 10362
rect 3842 10310 7084 10362
rect 920 10288 7084 10310
rect 6362 10248 6368 10260
rect 6323 10220 6368 10248
rect 6362 10208 6368 10220
rect 6420 10208 6426 10260
rect 2958 10180 2964 10192
rect 2714 10152 2964 10180
rect 2958 10140 2964 10152
rect 3016 10140 3022 10192
rect 4246 10140 4252 10192
rect 4304 10140 4310 10192
rect 5537 10183 5595 10189
rect 5537 10149 5549 10183
rect 5583 10180 5595 10183
rect 6546 10180 6552 10192
rect 5583 10152 6552 10180
rect 5583 10149 5595 10152
rect 5537 10143 5595 10149
rect 6546 10140 6552 10152
rect 6604 10140 6610 10192
rect 3418 10112 3424 10124
rect 2746 10084 3424 10112
rect 1210 10044 1216 10056
rect 1171 10016 1216 10044
rect 1210 10004 1216 10016
rect 1268 10004 1274 10056
rect 1489 10047 1547 10053
rect 1489 10013 1501 10047
rect 1535 10044 1547 10047
rect 2746 10044 2774 10084
rect 3418 10072 3424 10084
rect 3476 10112 3482 10124
rect 3697 10115 3755 10121
rect 3697 10112 3709 10115
rect 3476 10084 3709 10112
rect 3476 10072 3482 10084
rect 3697 10081 3709 10084
rect 3743 10081 3755 10115
rect 3697 10075 3755 10081
rect 4522 10072 4528 10124
rect 4580 10112 4586 10124
rect 5442 10112 5448 10124
rect 4580 10084 5448 10112
rect 4580 10072 4586 10084
rect 5442 10072 5448 10084
rect 5500 10112 5506 10124
rect 5721 10115 5779 10121
rect 5721 10112 5733 10115
rect 5500 10084 5733 10112
rect 5500 10072 5506 10084
rect 5721 10081 5733 10084
rect 5767 10081 5779 10115
rect 5721 10075 5779 10081
rect 6273 10115 6331 10121
rect 6273 10081 6285 10115
rect 6319 10112 6331 10115
rect 6362 10112 6368 10124
rect 6319 10084 6368 10112
rect 6319 10081 6331 10084
rect 6273 10075 6331 10081
rect 6362 10072 6368 10084
rect 6420 10072 6426 10124
rect 1535 10016 2774 10044
rect 1535 10013 1547 10016
rect 1489 10007 1547 10013
rect 3142 10004 3148 10056
rect 3200 10044 3206 10056
rect 3237 10047 3295 10053
rect 3237 10044 3249 10047
rect 3200 10016 3249 10044
rect 3200 10004 3206 10016
rect 3237 10013 3249 10016
rect 3283 10013 3295 10047
rect 3237 10007 3295 10013
rect 3329 10047 3387 10053
rect 3329 10013 3341 10047
rect 3375 10013 3387 10047
rect 3329 10007 3387 10013
rect 2866 9936 2872 9988
rect 2924 9976 2930 9988
rect 3344 9976 3372 10007
rect 4982 10004 4988 10056
rect 5040 10044 5046 10056
rect 5077 10047 5135 10053
rect 5077 10044 5089 10047
rect 5040 10016 5089 10044
rect 5040 10004 5046 10016
rect 5077 10013 5089 10016
rect 5123 10013 5135 10047
rect 5077 10007 5135 10013
rect 2924 9948 3372 9976
rect 2924 9936 2930 9948
rect 3344 9908 3372 9948
rect 3694 9908 3700 9920
rect 3344 9880 3700 9908
rect 3694 9868 3700 9880
rect 3752 9908 3758 9920
rect 4430 9908 4436 9920
rect 3752 9880 4436 9908
rect 3752 9868 3758 9880
rect 4430 9868 4436 9880
rect 4488 9868 4494 9920
rect 5442 9868 5448 9920
rect 5500 9908 5506 9920
rect 5813 9911 5871 9917
rect 5813 9908 5825 9911
rect 5500 9880 5825 9908
rect 5500 9868 5506 9880
rect 5813 9877 5825 9880
rect 5859 9877 5871 9911
rect 5813 9871 5871 9877
rect 920 9818 7084 9840
rect 920 9766 2098 9818
rect 2150 9766 2162 9818
rect 2214 9766 2226 9818
rect 2278 9766 2290 9818
rect 2342 9766 5098 9818
rect 5150 9766 5162 9818
rect 5214 9766 5226 9818
rect 5278 9766 5290 9818
rect 5342 9766 7084 9818
rect 920 9744 7084 9766
rect 5718 9704 5724 9716
rect 3160 9676 3372 9704
rect 2225 9571 2283 9577
rect 2225 9537 2237 9571
rect 2271 9568 2283 9571
rect 3160 9568 3188 9676
rect 3234 9596 3240 9648
rect 3292 9636 3298 9648
rect 3344 9636 3372 9676
rect 3988 9676 5724 9704
rect 3988 9636 4016 9676
rect 5718 9664 5724 9676
rect 5776 9664 5782 9716
rect 6086 9664 6092 9716
rect 6144 9704 6150 9716
rect 6144 9676 6224 9704
rect 6144 9664 6150 9676
rect 6196 9674 6224 9676
rect 6196 9648 6316 9674
rect 6196 9646 6276 9648
rect 3292 9608 3372 9636
rect 3436 9608 4016 9636
rect 3292 9596 3298 9608
rect 3436 9568 3464 9608
rect 6270 9596 6276 9646
rect 6328 9596 6334 9648
rect 2271 9540 3188 9568
rect 3252 9540 3464 9568
rect 5905 9571 5963 9577
rect 2271 9537 2283 9540
rect 2225 9531 2283 9537
rect 1857 9503 1915 9509
rect 1857 9469 1869 9503
rect 1903 9469 1915 9503
rect 1857 9463 1915 9469
rect 1872 9432 1900 9463
rect 2314 9460 2320 9512
rect 2372 9500 2378 9512
rect 2682 9500 2688 9512
rect 2372 9472 2688 9500
rect 2372 9460 2378 9472
rect 2682 9460 2688 9472
rect 2740 9460 2746 9512
rect 2958 9500 2964 9512
rect 2919 9472 2964 9500
rect 2958 9460 2964 9472
rect 3016 9460 3022 9512
rect 3145 9503 3203 9509
rect 3145 9469 3157 9503
rect 3191 9500 3203 9503
rect 3252 9500 3280 9540
rect 5905 9537 5917 9571
rect 5951 9568 5963 9571
rect 6178 9568 6184 9580
rect 5951 9540 6184 9568
rect 5951 9537 5963 9540
rect 5905 9531 5963 9537
rect 6178 9528 6184 9540
rect 6236 9528 6242 9580
rect 6454 9528 6460 9580
rect 6512 9568 6518 9580
rect 14090 9568 14096 9580
rect 6512 9540 14096 9568
rect 6512 9528 6518 9540
rect 14090 9528 14096 9540
rect 14148 9528 14154 9580
rect 3418 9500 3424 9512
rect 3191 9472 3280 9500
rect 3379 9472 3424 9500
rect 3191 9469 3203 9472
rect 3145 9463 3203 9469
rect 3418 9460 3424 9472
rect 3476 9460 3482 9512
rect 3697 9503 3755 9509
rect 3697 9469 3709 9503
rect 3743 9469 3755 9503
rect 3697 9463 3755 9469
rect 3050 9432 3056 9444
rect 1872 9404 3056 9432
rect 3050 9392 3056 9404
rect 3108 9392 3114 9444
rect 2041 9367 2099 9373
rect 2041 9333 2053 9367
rect 2087 9364 2099 9367
rect 2774 9364 2780 9376
rect 2087 9336 2780 9364
rect 2087 9333 2099 9336
rect 2041 9327 2099 9333
rect 2774 9324 2780 9336
rect 2832 9364 2838 9376
rect 2958 9364 2964 9376
rect 2832 9336 2964 9364
rect 2832 9324 2838 9336
rect 2958 9324 2964 9336
rect 3016 9324 3022 9376
rect 3326 9324 3332 9376
rect 3384 9364 3390 9376
rect 3712 9364 3740 9463
rect 3786 9460 3792 9512
rect 3844 9500 3850 9512
rect 3881 9503 3939 9509
rect 3881 9500 3893 9503
rect 3844 9472 3893 9500
rect 3844 9460 3850 9472
rect 3881 9469 3893 9472
rect 3927 9469 3939 9503
rect 3881 9463 3939 9469
rect 5626 9460 5632 9512
rect 5684 9500 5690 9512
rect 5997 9503 6055 9509
rect 5997 9500 6009 9503
rect 5684 9472 6009 9500
rect 5684 9460 5690 9472
rect 5997 9469 6009 9472
rect 6043 9469 6055 9503
rect 5997 9463 6055 9469
rect 6365 9503 6423 9509
rect 6365 9469 6377 9503
rect 6411 9500 6423 9503
rect 6546 9500 6552 9512
rect 6411 9472 6552 9500
rect 6411 9469 6423 9472
rect 6365 9463 6423 9469
rect 6546 9460 6552 9472
rect 6604 9460 6610 9512
rect 4154 9432 4160 9444
rect 4115 9404 4160 9432
rect 4154 9392 4160 9404
rect 4212 9392 4218 9444
rect 5810 9432 5816 9444
rect 5382 9404 5816 9432
rect 5810 9392 5816 9404
rect 5868 9392 5874 9444
rect 7190 9392 7196 9444
rect 7248 9432 7254 9444
rect 14182 9432 14188 9444
rect 7248 9404 14188 9432
rect 7248 9392 7254 9404
rect 14182 9392 14188 9404
rect 14240 9392 14246 9444
rect 6086 9364 6092 9376
rect 3384 9336 6092 9364
rect 3384 9324 3390 9336
rect 6086 9324 6092 9336
rect 6144 9324 6150 9376
rect 6178 9324 6184 9376
rect 6236 9364 6242 9376
rect 6457 9367 6515 9373
rect 6236 9336 6281 9364
rect 6236 9324 6242 9336
rect 6457 9333 6469 9367
rect 6503 9364 6515 9367
rect 6546 9364 6552 9376
rect 6503 9336 6552 9364
rect 6503 9333 6515 9336
rect 6457 9327 6515 9333
rect 6546 9324 6552 9336
rect 6604 9324 6610 9376
rect 920 9274 7084 9296
rect 920 9222 3598 9274
rect 3650 9222 3662 9274
rect 3714 9222 3726 9274
rect 3778 9222 3790 9274
rect 3842 9222 7084 9274
rect 920 9200 7084 9222
rect 5626 9160 5632 9172
rect 5539 9132 5632 9160
rect 5626 9120 5632 9132
rect 5684 9120 5690 9172
rect 5810 9120 5816 9172
rect 5868 9160 5874 9172
rect 5997 9163 6055 9169
rect 5997 9160 6009 9163
rect 5868 9132 6009 9160
rect 5868 9120 5874 9132
rect 5997 9129 6009 9132
rect 6043 9129 6055 9163
rect 5997 9123 6055 9129
rect 6086 9120 6092 9172
rect 6144 9160 6150 9172
rect 6546 9160 6552 9172
rect 6144 9132 6552 9160
rect 6144 9120 6150 9132
rect 6546 9120 6552 9132
rect 6604 9120 6610 9172
rect 2590 9092 2596 9104
rect 2148 9064 2596 9092
rect 2148 9033 2176 9064
rect 2590 9052 2596 9064
rect 2648 9052 2654 9104
rect 3326 9092 3332 9104
rect 2700 9064 3332 9092
rect 1949 9027 2007 9033
rect 1949 8993 1961 9027
rect 1995 8993 2007 9027
rect 1949 8987 2007 8993
rect 2133 9027 2191 9033
rect 2133 8993 2145 9027
rect 2179 8993 2191 9027
rect 2314 9024 2320 9036
rect 2275 8996 2320 9024
rect 2133 8987 2191 8993
rect 1394 8956 1400 8968
rect 1355 8928 1400 8956
rect 1394 8916 1400 8928
rect 1452 8916 1458 8968
rect 1964 8956 1992 8987
rect 2314 8984 2320 8996
rect 2372 8984 2378 9036
rect 2700 9033 2728 9064
rect 3326 9052 3332 9064
rect 3384 9052 3390 9104
rect 5644 9092 5672 9120
rect 4816 9064 5672 9092
rect 2685 9027 2743 9033
rect 2685 8993 2697 9027
rect 2731 8993 2743 9027
rect 2685 8987 2743 8993
rect 4338 8984 4344 9036
rect 4396 8984 4402 9036
rect 2498 8956 2504 8968
rect 1964 8928 2504 8956
rect 2498 8916 2504 8928
rect 2556 8916 2562 8968
rect 2777 8959 2835 8965
rect 2777 8925 2789 8959
rect 2823 8925 2835 8959
rect 2777 8919 2835 8925
rect 2792 8820 2820 8919
rect 2866 8916 2872 8968
rect 2924 8956 2930 8968
rect 2961 8959 3019 8965
rect 2961 8956 2973 8959
rect 2924 8928 2973 8956
rect 2924 8916 2930 8928
rect 2961 8925 2973 8928
rect 3007 8925 3019 8959
rect 3234 8956 3240 8968
rect 3195 8928 3240 8956
rect 2961 8919 3019 8925
rect 3234 8916 3240 8928
rect 3292 8916 3298 8968
rect 3970 8916 3976 8968
rect 4028 8956 4034 8968
rect 4816 8956 4844 9064
rect 5077 9027 5135 9033
rect 5077 8993 5089 9027
rect 5123 9024 5135 9027
rect 5442 9024 5448 9036
rect 5123 8996 5448 9024
rect 5123 8993 5135 8996
rect 5077 8987 5135 8993
rect 5442 8984 5448 8996
rect 5500 8984 5506 9036
rect 5644 9024 5672 9064
rect 5718 9052 5724 9104
rect 5776 9092 5782 9104
rect 5776 9064 6316 9092
rect 5776 9052 5782 9064
rect 6288 9036 6316 9064
rect 5813 9027 5871 9033
rect 5813 9024 5825 9027
rect 5644 8996 5825 9024
rect 5813 8993 5825 8996
rect 5859 9024 5871 9027
rect 6086 9024 6092 9036
rect 5859 8996 6092 9024
rect 5859 8993 5871 8996
rect 5813 8987 5871 8993
rect 6086 8984 6092 8996
rect 6144 8984 6150 9036
rect 6270 9024 6276 9036
rect 6231 8996 6276 9024
rect 6270 8984 6276 8996
rect 6328 8984 6334 9036
rect 4982 8956 4988 8968
rect 4028 8928 4844 8956
rect 4943 8928 4988 8956
rect 4028 8916 4034 8928
rect 4982 8916 4988 8928
rect 5040 8916 5046 8968
rect 12526 8956 12532 8968
rect 6104 8928 12532 8956
rect 4430 8848 4436 8900
rect 4488 8888 4494 8900
rect 5261 8891 5319 8897
rect 5261 8888 5273 8891
rect 4488 8860 5273 8888
rect 4488 8848 4494 8860
rect 5261 8857 5273 8860
rect 5307 8857 5319 8891
rect 5261 8851 5319 8857
rect 6104 8820 6132 8928
rect 12526 8916 12532 8928
rect 12584 8916 12590 8968
rect 2792 8792 6132 8820
rect 6178 8780 6184 8832
rect 6236 8820 6242 8832
rect 6365 8823 6423 8829
rect 6365 8820 6377 8823
rect 6236 8792 6377 8820
rect 6236 8780 6242 8792
rect 6365 8789 6377 8792
rect 6411 8789 6423 8823
rect 6365 8783 6423 8789
rect 920 8730 7084 8752
rect 920 8678 2098 8730
rect 2150 8678 2162 8730
rect 2214 8678 2226 8730
rect 2278 8678 2290 8730
rect 2342 8678 5098 8730
rect 5150 8678 5162 8730
rect 5214 8678 5226 8730
rect 5278 8678 5290 8730
rect 5342 8678 7084 8730
rect 920 8656 7084 8678
rect 3142 8616 3148 8628
rect 2746 8588 3148 8616
rect 1210 8480 1216 8492
rect 1171 8452 1216 8480
rect 1210 8440 1216 8452
rect 1268 8440 1274 8492
rect 1489 8483 1547 8489
rect 1489 8449 1501 8483
rect 1535 8480 1547 8483
rect 2746 8480 2774 8588
rect 3142 8576 3148 8588
rect 3200 8616 3206 8628
rect 3970 8616 3976 8628
rect 3200 8588 3976 8616
rect 3200 8576 3206 8588
rect 3970 8576 3976 8588
rect 4028 8576 4034 8628
rect 4338 8576 4344 8628
rect 4396 8616 4402 8628
rect 6641 8619 6699 8625
rect 6641 8616 6653 8619
rect 4396 8588 6653 8616
rect 4396 8576 4402 8588
rect 6641 8585 6653 8588
rect 6687 8585 6699 8619
rect 6641 8579 6699 8585
rect 4246 8548 4252 8560
rect 1535 8452 2774 8480
rect 3068 8520 4252 8548
rect 1535 8449 1547 8452
rect 1489 8443 1547 8449
rect 3068 8344 3096 8520
rect 4246 8508 4252 8520
rect 4304 8508 4310 8560
rect 3418 8440 3424 8492
rect 3476 8480 3482 8492
rect 12434 8480 12440 8492
rect 3476 8452 12440 8480
rect 3476 8440 3482 8452
rect 12434 8440 12440 8452
rect 12492 8440 12498 8492
rect 3326 8412 3332 8424
rect 3287 8384 3332 8412
rect 3326 8372 3332 8384
rect 3384 8372 3390 8424
rect 3973 8415 4031 8421
rect 3973 8381 3985 8415
rect 4019 8412 4031 8415
rect 4062 8412 4068 8424
rect 4019 8384 4068 8412
rect 4019 8381 4031 8384
rect 3973 8375 4031 8381
rect 4062 8372 4068 8384
rect 4120 8372 4126 8424
rect 4341 8415 4399 8421
rect 4341 8381 4353 8415
rect 4387 8381 4399 8415
rect 4341 8375 4399 8381
rect 3234 8344 3240 8356
rect 2714 8316 3096 8344
rect 3195 8316 3240 8344
rect 3234 8304 3240 8316
rect 3292 8304 3298 8356
rect 4356 8344 4384 8375
rect 6086 8372 6092 8424
rect 6144 8412 6150 8424
rect 6457 8415 6515 8421
rect 6457 8412 6469 8415
rect 6144 8384 6469 8412
rect 6144 8372 6150 8384
rect 6457 8381 6469 8384
rect 6503 8381 6515 8415
rect 6457 8375 6515 8381
rect 4522 8344 4528 8356
rect 4356 8316 4528 8344
rect 4522 8304 4528 8316
rect 4580 8304 4586 8356
rect 4617 8347 4675 8353
rect 4617 8313 4629 8347
rect 4663 8344 4675 8347
rect 4706 8344 4712 8356
rect 4663 8316 4712 8344
rect 4663 8313 4675 8316
rect 4617 8307 4675 8313
rect 4706 8304 4712 8316
rect 4764 8304 4770 8356
rect 6365 8347 6423 8353
rect 5460 8288 5488 8330
rect 6365 8313 6377 8347
rect 6411 8344 6423 8347
rect 6638 8344 6644 8356
rect 6411 8316 6644 8344
rect 6411 8313 6423 8316
rect 6365 8307 6423 8313
rect 6638 8304 6644 8316
rect 6696 8304 6702 8356
rect 3142 8236 3148 8288
rect 3200 8276 3206 8288
rect 3513 8279 3571 8285
rect 3513 8276 3525 8279
rect 3200 8248 3525 8276
rect 3200 8236 3206 8248
rect 3513 8245 3525 8248
rect 3559 8245 3571 8279
rect 3513 8239 3571 8245
rect 4157 8279 4215 8285
rect 4157 8245 4169 8279
rect 4203 8276 4215 8279
rect 4246 8276 4252 8288
rect 4203 8248 4252 8276
rect 4203 8245 4215 8248
rect 4157 8239 4215 8245
rect 4246 8236 4252 8248
rect 4304 8236 4310 8288
rect 5442 8236 5448 8288
rect 5500 8236 5506 8288
rect 920 8186 7084 8208
rect 920 8134 3598 8186
rect 3650 8134 3662 8186
rect 3714 8134 3726 8186
rect 3778 8134 3790 8186
rect 3842 8134 7084 8186
rect 920 8112 7084 8134
rect 3234 8072 3240 8084
rect 1504 8044 3240 8072
rect 1504 8013 1532 8044
rect 3234 8032 3240 8044
rect 3292 8032 3298 8084
rect 4430 8072 4436 8084
rect 3344 8044 4436 8072
rect 1489 8007 1547 8013
rect 1489 7973 1501 8007
rect 1535 7973 1547 8007
rect 3142 8004 3148 8016
rect 2714 7976 3148 8004
rect 1489 7967 1547 7973
rect 3142 7964 3148 7976
rect 3200 7964 3206 8016
rect 3050 7896 3056 7948
rect 3108 7936 3114 7948
rect 3344 7945 3372 8044
rect 4430 8032 4436 8044
rect 4488 8032 4494 8084
rect 6089 8075 6147 8081
rect 6089 8041 6101 8075
rect 6135 8072 6147 8075
rect 6270 8072 6276 8084
rect 6135 8044 6276 8072
rect 6135 8041 6147 8044
rect 6089 8035 6147 8041
rect 6270 8032 6276 8044
rect 6328 8032 6334 8084
rect 6365 8075 6423 8081
rect 6365 8041 6377 8075
rect 6411 8041 6423 8075
rect 6365 8035 6423 8041
rect 3970 7964 3976 8016
rect 4028 7964 4034 8016
rect 6380 8004 6408 8035
rect 5382 7976 6408 8004
rect 3329 7939 3387 7945
rect 3329 7936 3341 7939
rect 3108 7908 3341 7936
rect 3108 7896 3114 7908
rect 3329 7905 3341 7908
rect 3375 7905 3387 7939
rect 3329 7899 3387 7905
rect 3418 7896 3424 7948
rect 3476 7936 3482 7948
rect 3878 7936 3884 7948
rect 3476 7908 3884 7936
rect 3476 7896 3482 7908
rect 3878 7896 3884 7908
rect 3936 7896 3942 7948
rect 3988 7936 4016 7964
rect 4341 7939 4399 7945
rect 4341 7936 4353 7939
rect 3988 7908 4353 7936
rect 4341 7905 4353 7908
rect 4387 7905 4399 7939
rect 4341 7899 4399 7905
rect 6086 7896 6092 7948
rect 6144 7936 6150 7948
rect 6181 7939 6239 7945
rect 6181 7936 6193 7939
rect 6144 7908 6193 7936
rect 6144 7896 6150 7908
rect 6181 7905 6193 7908
rect 6227 7905 6239 7939
rect 6181 7899 6239 7905
rect 1210 7868 1216 7880
rect 1171 7840 1216 7868
rect 1210 7828 1216 7840
rect 1268 7828 1274 7880
rect 3234 7868 3240 7880
rect 3195 7840 3240 7868
rect 3234 7828 3240 7840
rect 3292 7828 3298 7880
rect 3970 7868 3976 7880
rect 3931 7840 3976 7868
rect 3970 7828 3976 7840
rect 4028 7828 4034 7880
rect 3050 7760 3056 7812
rect 3108 7800 3114 7812
rect 3697 7803 3755 7809
rect 3697 7800 3709 7803
rect 3108 7772 3709 7800
rect 3108 7760 3114 7772
rect 3697 7769 3709 7772
rect 3743 7769 3755 7803
rect 3697 7763 3755 7769
rect 3142 7692 3148 7744
rect 3200 7732 3206 7744
rect 3326 7732 3332 7744
rect 3200 7704 3332 7732
rect 3200 7692 3206 7704
rect 3326 7692 3332 7704
rect 3384 7732 3390 7744
rect 3513 7735 3571 7741
rect 3513 7732 3525 7735
rect 3384 7704 3525 7732
rect 3384 7692 3390 7704
rect 3513 7701 3525 7704
rect 3559 7701 3571 7735
rect 3513 7695 3571 7701
rect 920 7642 7084 7664
rect 920 7590 2098 7642
rect 2150 7590 2162 7642
rect 2214 7590 2226 7642
rect 2278 7590 2290 7642
rect 2342 7590 5098 7642
rect 5150 7590 5162 7642
rect 5214 7590 5226 7642
rect 5278 7590 5290 7642
rect 5342 7590 7084 7642
rect 920 7568 7084 7590
rect 1394 7488 1400 7540
rect 1452 7528 1458 7540
rect 7561 7531 7619 7537
rect 7561 7528 7573 7531
rect 1452 7500 7573 7528
rect 1452 7488 1458 7500
rect 7561 7497 7573 7500
rect 7607 7497 7619 7531
rect 7561 7491 7619 7497
rect 2866 7420 2872 7472
rect 2924 7460 2930 7472
rect 3878 7460 3884 7472
rect 2924 7432 3884 7460
rect 2924 7420 2930 7432
rect 3878 7420 3884 7432
rect 3936 7420 3942 7472
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7392 1639 7395
rect 3234 7392 3240 7404
rect 1627 7364 3240 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 3234 7352 3240 7364
rect 3292 7392 3298 7404
rect 4157 7395 4215 7401
rect 4157 7392 4169 7395
rect 3292 7364 4169 7392
rect 3292 7352 3298 7364
rect 4157 7361 4169 7364
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 1302 7324 1308 7336
rect 1263 7296 1308 7324
rect 1302 7284 1308 7296
rect 1360 7284 1366 7336
rect 3142 7284 3148 7336
rect 3200 7324 3206 7336
rect 3421 7327 3479 7333
rect 3421 7324 3433 7327
rect 3200 7296 3433 7324
rect 3200 7284 3206 7296
rect 3421 7293 3433 7296
rect 3467 7293 3479 7327
rect 3878 7324 3884 7336
rect 3839 7296 3884 7324
rect 3421 7287 3479 7293
rect 3878 7284 3884 7296
rect 3936 7284 3942 7336
rect 6178 7324 6184 7336
rect 6139 7296 6184 7324
rect 6178 7284 6184 7296
rect 6236 7284 6242 7336
rect 3329 7259 3387 7265
rect 2792 7188 2820 7242
rect 3329 7225 3341 7259
rect 3375 7256 3387 7259
rect 4062 7256 4068 7268
rect 3375 7228 4068 7256
rect 3375 7225 3387 7228
rect 3329 7219 3387 7225
rect 4062 7216 4068 7228
rect 4120 7216 4126 7268
rect 4246 7216 4252 7268
rect 4304 7256 4310 7268
rect 5905 7259 5963 7265
rect 4304 7228 4646 7256
rect 4304 7216 4310 7228
rect 5905 7225 5917 7259
rect 5951 7256 5963 7259
rect 5997 7259 6055 7265
rect 5997 7256 6009 7259
rect 5951 7228 6009 7256
rect 5951 7225 5963 7228
rect 5905 7219 5963 7225
rect 5997 7225 6009 7228
rect 6043 7256 6055 7259
rect 14182 7256 14188 7268
rect 6043 7228 14188 7256
rect 6043 7225 6055 7228
rect 5997 7219 6055 7225
rect 14182 7216 14188 7228
rect 14240 7216 14246 7268
rect 3605 7191 3663 7197
rect 3605 7188 3617 7191
rect 2792 7160 3617 7188
rect 3605 7157 3617 7160
rect 3651 7157 3663 7191
rect 6270 7188 6276 7200
rect 6231 7160 6276 7188
rect 3605 7151 3663 7157
rect 6270 7148 6276 7160
rect 6328 7148 6334 7200
rect 7561 7191 7619 7197
rect 7561 7157 7573 7191
rect 7607 7188 7619 7191
rect 14090 7188 14096 7200
rect 7607 7160 14096 7188
rect 7607 7157 7619 7160
rect 7561 7151 7619 7157
rect 14090 7148 14096 7160
rect 14148 7148 14154 7200
rect 920 7098 7084 7120
rect 920 7046 3598 7098
rect 3650 7046 3662 7098
rect 3714 7046 3726 7098
rect 3778 7046 3790 7098
rect 3842 7046 7084 7098
rect 920 7024 7084 7046
rect 3970 6944 3976 6996
rect 4028 6984 4034 6996
rect 4246 6984 4252 6996
rect 4028 6956 4252 6984
rect 4028 6944 4034 6956
rect 4246 6944 4252 6956
rect 4304 6944 4310 6996
rect 6362 6984 6368 6996
rect 5828 6956 6368 6984
rect 2961 6919 3019 6925
rect 2961 6885 2973 6919
rect 3007 6916 3019 6919
rect 3418 6916 3424 6928
rect 3007 6888 3424 6916
rect 3007 6885 3019 6888
rect 2961 6879 3019 6885
rect 3418 6876 3424 6888
rect 3476 6876 3482 6928
rect 3878 6876 3884 6928
rect 3936 6876 3942 6928
rect 5828 6925 5856 6956
rect 6362 6944 6368 6956
rect 6420 6984 6426 6996
rect 14182 6984 14188 6996
rect 6420 6956 14188 6984
rect 6420 6944 6426 6956
rect 14182 6944 14188 6956
rect 14240 6944 14246 6996
rect 5813 6919 5871 6925
rect 5813 6885 5825 6919
rect 5859 6885 5871 6919
rect 5813 6879 5871 6885
rect 5905 6919 5963 6925
rect 5905 6885 5917 6919
rect 5951 6916 5963 6919
rect 6270 6916 6276 6928
rect 5951 6888 6276 6916
rect 5951 6885 5963 6888
rect 5905 6879 5963 6885
rect 6270 6876 6276 6888
rect 6328 6876 6334 6928
rect 753 6851 811 6857
rect 753 6817 765 6851
rect 799 6848 811 6851
rect 1213 6851 1271 6857
rect 1213 6848 1225 6851
rect 799 6820 1225 6848
rect 799 6817 811 6820
rect 753 6811 811 6817
rect 1213 6817 1225 6820
rect 1259 6817 1271 6851
rect 3050 6848 3056 6860
rect 3011 6820 3056 6848
rect 1213 6811 1271 6817
rect 3050 6808 3056 6820
rect 3108 6808 3114 6860
rect 4890 6848 4896 6860
rect 4724 6820 4896 6848
rect 3329 6783 3387 6789
rect 3329 6749 3341 6783
rect 3375 6780 3387 6783
rect 4724 6780 4752 6820
rect 4890 6808 4896 6820
rect 4948 6808 4954 6860
rect 5169 6851 5227 6857
rect 5169 6817 5181 6851
rect 5215 6848 5227 6851
rect 5215 6820 5488 6848
rect 5215 6817 5227 6820
rect 5169 6811 5227 6817
rect 3375 6752 4752 6780
rect 3375 6749 3387 6752
rect 3329 6743 3387 6749
rect 4798 6740 4804 6792
rect 4856 6780 4862 6792
rect 5077 6783 5135 6789
rect 5077 6780 5089 6783
rect 4856 6752 5089 6780
rect 4856 6740 4862 6752
rect 5077 6749 5089 6752
rect 5123 6749 5135 6783
rect 5077 6743 5135 6749
rect 4338 6672 4344 6724
rect 4396 6712 4402 6724
rect 5353 6715 5411 6721
rect 5353 6712 5365 6715
rect 4396 6684 5365 6712
rect 4396 6672 4402 6684
rect 5353 6681 5365 6684
rect 5399 6681 5411 6715
rect 5353 6675 5411 6681
rect 3142 6604 3148 6656
rect 3200 6644 3206 6656
rect 5460 6644 5488 6820
rect 6454 6780 6460 6792
rect 6415 6752 6460 6780
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 3200 6616 5488 6644
rect 3200 6604 3206 6616
rect 920 6554 7084 6576
rect 920 6502 2098 6554
rect 2150 6502 2162 6554
rect 2214 6502 2226 6554
rect 2278 6502 2290 6554
rect 2342 6502 5098 6554
rect 5150 6502 5162 6554
rect 5214 6502 5226 6554
rect 5278 6502 5290 6554
rect 5342 6502 7084 6554
rect 920 6480 7084 6502
rect 753 6443 811 6449
rect 753 6409 765 6443
rect 799 6440 811 6443
rect 13262 6440 13268 6452
rect 799 6412 13268 6440
rect 799 6409 811 6412
rect 753 6403 811 6409
rect 13262 6400 13268 6412
rect 13320 6400 13326 6452
rect 1489 6307 1547 6313
rect 1489 6273 1501 6307
rect 1535 6304 1547 6307
rect 4062 6304 4068 6316
rect 1535 6276 4068 6304
rect 1535 6273 1547 6276
rect 1489 6267 1547 6273
rect 4062 6264 4068 6276
rect 4120 6304 4126 6316
rect 4617 6307 4675 6313
rect 4617 6304 4629 6307
rect 4120 6276 4629 6304
rect 4120 6264 4126 6276
rect 4617 6273 4629 6276
rect 4663 6273 4675 6307
rect 4617 6267 4675 6273
rect 1210 6236 1216 6248
rect 1171 6208 1216 6236
rect 1210 6196 1216 6208
rect 1268 6196 1274 6248
rect 3142 6196 3148 6248
rect 3200 6236 3206 6248
rect 3329 6239 3387 6245
rect 3329 6236 3341 6239
rect 3200 6208 3341 6236
rect 3200 6196 3206 6208
rect 3329 6205 3341 6208
rect 3375 6205 3387 6239
rect 3878 6236 3884 6248
rect 3839 6208 3884 6236
rect 3329 6199 3387 6205
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 4246 6196 4252 6248
rect 4304 6236 4310 6248
rect 4341 6239 4399 6245
rect 4341 6236 4353 6239
rect 4304 6208 4353 6236
rect 4304 6196 4310 6208
rect 4341 6205 4353 6208
rect 4387 6205 4399 6239
rect 4341 6199 4399 6205
rect 6086 6196 6092 6248
rect 6144 6236 6150 6248
rect 6457 6239 6515 6245
rect 6457 6236 6469 6239
rect 6144 6208 6469 6236
rect 6144 6196 6150 6208
rect 6457 6205 6469 6208
rect 6503 6205 6515 6239
rect 6457 6199 6515 6205
rect 2700 6100 2728 6154
rect 2866 6128 2872 6180
rect 2924 6168 2930 6180
rect 3237 6171 3295 6177
rect 3237 6168 3249 6171
rect 2924 6140 3249 6168
rect 2924 6128 2930 6140
rect 3237 6137 3249 6140
rect 3283 6137 3295 6171
rect 6365 6171 6423 6177
rect 3237 6131 3295 6137
rect 3513 6103 3571 6109
rect 3513 6100 3525 6103
rect 2700 6072 3525 6100
rect 3513 6069 3525 6072
rect 3559 6069 3571 6103
rect 4062 6100 4068 6112
rect 4023 6072 4068 6100
rect 3513 6063 3571 6069
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 5828 6100 5856 6154
rect 6365 6137 6377 6171
rect 6411 6168 6423 6171
rect 14090 6168 14096 6180
rect 6411 6140 14096 6168
rect 6411 6137 6423 6140
rect 6365 6131 6423 6137
rect 14090 6128 14096 6140
rect 14148 6128 14154 6180
rect 6641 6103 6699 6109
rect 6641 6100 6653 6103
rect 5828 6072 6653 6100
rect 6641 6069 6653 6072
rect 6687 6069 6699 6103
rect 6641 6063 6699 6069
rect 920 6010 7084 6032
rect 920 5958 3598 6010
rect 3650 5958 3662 6010
rect 3714 5958 3726 6010
rect 3778 5958 3790 6010
rect 3842 5958 7084 6010
rect 920 5936 7084 5958
rect 4614 5856 4620 5908
rect 4672 5896 4678 5908
rect 4672 5868 5120 5896
rect 4672 5856 4678 5868
rect 2406 5788 2412 5840
rect 2464 5788 2470 5840
rect 4062 5788 4068 5840
rect 4120 5828 4126 5840
rect 4120 5800 4278 5828
rect 4120 5788 4126 5800
rect 3050 5720 3056 5772
rect 3108 5760 3114 5772
rect 3513 5763 3571 5769
rect 3513 5760 3525 5763
rect 3108 5732 3525 5760
rect 3108 5720 3114 5732
rect 3513 5729 3525 5732
rect 3559 5729 3571 5763
rect 5092 5760 5120 5868
rect 5534 5856 5540 5908
rect 5592 5896 5598 5908
rect 5813 5899 5871 5905
rect 5813 5896 5825 5899
rect 5592 5868 5825 5896
rect 5592 5856 5598 5868
rect 5813 5865 5825 5868
rect 5859 5896 5871 5899
rect 5859 5868 6040 5896
rect 5859 5865 5871 5868
rect 5813 5859 5871 5865
rect 6012 5769 6040 5868
rect 5537 5763 5595 5769
rect 5537 5760 5549 5763
rect 5092 5732 5549 5760
rect 3513 5723 3571 5729
rect 5537 5729 5549 5732
rect 5583 5729 5595 5763
rect 5537 5723 5595 5729
rect 5629 5763 5687 5769
rect 5629 5729 5641 5763
rect 5675 5729 5687 5763
rect 5629 5723 5687 5729
rect 5997 5763 6055 5769
rect 5997 5729 6009 5763
rect 6043 5760 6055 5763
rect 6086 5760 6092 5772
rect 6043 5732 6092 5760
rect 6043 5729 6055 5732
rect 5997 5723 6055 5729
rect 1302 5652 1308 5704
rect 1360 5692 1366 5704
rect 1397 5695 1455 5701
rect 1397 5692 1409 5695
rect 1360 5664 1409 5692
rect 1360 5652 1366 5664
rect 1397 5661 1409 5664
rect 1443 5692 1455 5695
rect 1670 5692 1676 5704
rect 1443 5664 1532 5692
rect 1631 5664 1676 5692
rect 1443 5661 1455 5664
rect 1397 5655 1455 5661
rect 1504 5556 1532 5664
rect 1670 5652 1676 5664
rect 1728 5652 1734 5704
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5661 3479 5695
rect 3789 5695 3847 5701
rect 3789 5692 3801 5695
rect 3421 5655 3479 5661
rect 3620 5664 3801 5692
rect 3436 5624 3464 5655
rect 3620 5624 3648 5664
rect 3789 5661 3801 5664
rect 3835 5692 3847 5695
rect 4154 5692 4160 5704
rect 3835 5664 4160 5692
rect 3835 5661 3847 5664
rect 3789 5655 3847 5661
rect 4154 5652 4160 5664
rect 4212 5652 4218 5704
rect 4430 5652 4436 5704
rect 4488 5692 4494 5704
rect 5644 5692 5672 5723
rect 6086 5720 6092 5732
rect 6144 5720 6150 5772
rect 4488 5664 5672 5692
rect 4488 5652 4494 5664
rect 3436 5596 3648 5624
rect 4982 5584 4988 5636
rect 5040 5624 5046 5636
rect 14090 5624 14096 5636
rect 5040 5596 14096 5624
rect 5040 5584 5046 5596
rect 14090 5584 14096 5596
rect 14148 5584 14154 5636
rect 3050 5556 3056 5568
rect 1504 5528 3056 5556
rect 3050 5516 3056 5528
rect 3108 5516 3114 5568
rect 6178 5556 6184 5568
rect 6139 5528 6184 5556
rect 6178 5516 6184 5528
rect 6236 5516 6242 5568
rect 920 5466 7084 5488
rect 920 5414 2098 5466
rect 2150 5414 2162 5466
rect 2214 5414 2226 5466
rect 2278 5414 2290 5466
rect 2342 5414 5098 5466
rect 5150 5414 5162 5466
rect 5214 5414 5226 5466
rect 5278 5414 5290 5466
rect 5342 5414 7084 5466
rect 920 5392 7084 5414
rect 3513 5355 3571 5361
rect 3513 5321 3525 5355
rect 3559 5352 3571 5355
rect 3878 5352 3884 5364
rect 3559 5324 3884 5352
rect 3559 5321 3571 5324
rect 3513 5315 3571 5321
rect 3878 5312 3884 5324
rect 3936 5312 3942 5364
rect 1210 5216 1216 5228
rect 1171 5188 1216 5216
rect 1210 5176 1216 5188
rect 1268 5176 1274 5228
rect 1489 5219 1547 5225
rect 1489 5185 1501 5219
rect 1535 5216 1547 5219
rect 2866 5216 2872 5228
rect 1535 5188 2872 5216
rect 1535 5185 1547 5188
rect 1489 5179 1547 5185
rect 2866 5176 2872 5188
rect 2924 5176 2930 5228
rect 4430 5216 4436 5228
rect 3344 5188 4436 5216
rect 3344 5157 3372 5188
rect 4430 5176 4436 5188
rect 4488 5176 4494 5228
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5216 5043 5219
rect 6638 5216 6644 5228
rect 5031 5188 6644 5216
rect 5031 5185 5043 5188
rect 4985 5179 5043 5185
rect 6638 5176 6644 5188
rect 6696 5176 6702 5228
rect 3329 5151 3387 5157
rect 3329 5117 3341 5151
rect 3375 5117 3387 5151
rect 3329 5111 3387 5117
rect 3878 5108 3884 5160
rect 3936 5148 3942 5160
rect 3973 5151 4031 5157
rect 3973 5148 3985 5151
rect 3936 5120 3985 5148
rect 3936 5108 3942 5120
rect 3973 5117 3985 5120
rect 4019 5117 4031 5151
rect 3973 5111 4031 5117
rect 4246 5108 4252 5160
rect 4304 5148 4310 5160
rect 4617 5151 4675 5157
rect 4617 5148 4629 5151
rect 4304 5120 4629 5148
rect 4304 5108 4310 5120
rect 4617 5117 4629 5120
rect 4663 5117 4675 5151
rect 4617 5111 4675 5117
rect 1578 5040 1584 5092
rect 1636 5080 1642 5092
rect 1636 5052 1978 5080
rect 1636 5040 1642 5052
rect 2774 5040 2780 5092
rect 2832 5080 2838 5092
rect 3237 5083 3295 5089
rect 3237 5080 3249 5083
rect 2832 5052 3249 5080
rect 2832 5040 2838 5052
rect 3237 5049 3249 5052
rect 3283 5049 3295 5083
rect 6178 5080 6184 5092
rect 6026 5052 6184 5080
rect 3237 5043 3295 5049
rect 6178 5040 6184 5052
rect 6236 5040 6242 5092
rect 4157 5015 4215 5021
rect 4157 4981 4169 5015
rect 4203 5012 4215 5015
rect 4614 5012 4620 5024
rect 4203 4984 4620 5012
rect 4203 4981 4215 4984
rect 4157 4975 4215 4981
rect 4614 4972 4620 4984
rect 4672 4972 4678 5024
rect 6733 5015 6791 5021
rect 6733 4981 6745 5015
rect 6779 5012 6791 5015
rect 14182 5012 14188 5024
rect 6779 4984 14188 5012
rect 6779 4981 6791 4984
rect 6733 4975 6791 4981
rect 920 4922 7084 4944
rect 920 4870 3598 4922
rect 3650 4870 3662 4922
rect 3714 4870 3726 4922
rect 3778 4870 3790 4922
rect 3842 4870 7084 4922
rect 920 4848 7084 4870
rect 1578 4808 1584 4820
rect 1539 4780 1584 4808
rect 1578 4768 1584 4780
rect 1636 4768 1642 4820
rect 2317 4811 2375 4817
rect 2317 4777 2329 4811
rect 2363 4808 2375 4811
rect 2406 4808 2412 4820
rect 2363 4780 2412 4808
rect 2363 4777 2375 4780
rect 2317 4771 2375 4777
rect 2406 4768 2412 4780
rect 2464 4768 2470 4820
rect 3142 4808 3148 4820
rect 2746 4780 3148 4808
rect 2746 4740 2774 4780
rect 3142 4768 3148 4780
rect 3200 4768 3206 4820
rect 5261 4811 5319 4817
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 5442 4808 5448 4820
rect 5307 4780 5448 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 5442 4768 5448 4780
rect 5500 4768 5506 4820
rect 1412 4712 2774 4740
rect 1412 4681 1440 4712
rect 3510 4700 3516 4752
rect 3568 4700 3574 4752
rect 7116 4740 7144 4984
rect 14182 4972 14188 4984
rect 14240 4972 14246 5024
rect 5460 4712 7144 4740
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4641 1455 4675
rect 1397 4635 1455 4641
rect 1765 4675 1823 4681
rect 1765 4641 1777 4675
rect 1811 4672 1823 4675
rect 2133 4675 2191 4681
rect 2133 4672 2145 4675
rect 1811 4644 2145 4672
rect 1811 4641 1823 4644
rect 1765 4635 1823 4641
rect 2133 4641 2145 4644
rect 2179 4672 2191 4675
rect 2179 4644 2452 4672
rect 2179 4641 2191 4644
rect 2133 4635 2191 4641
rect 1946 4468 1952 4480
rect 1907 4440 1952 4468
rect 1946 4428 1952 4440
rect 2004 4428 2010 4480
rect 2424 4468 2452 4644
rect 4430 4632 4436 4684
rect 4488 4672 4494 4684
rect 5460 4681 5488 4712
rect 5077 4675 5135 4681
rect 5077 4672 5089 4675
rect 4488 4644 5089 4672
rect 4488 4632 4494 4644
rect 5077 4641 5089 4644
rect 5123 4641 5135 4675
rect 5077 4635 5135 4641
rect 5445 4675 5503 4681
rect 5445 4641 5457 4675
rect 5491 4641 5503 4675
rect 5445 4635 5503 4641
rect 5997 4675 6055 4681
rect 5997 4641 6009 4675
rect 6043 4672 6055 4675
rect 6086 4672 6092 4684
rect 6043 4644 6092 4672
rect 6043 4641 6055 4644
rect 5997 4635 6055 4641
rect 6086 4632 6092 4644
rect 6144 4632 6150 4684
rect 6457 4675 6515 4681
rect 6457 4641 6469 4675
rect 6503 4672 6515 4675
rect 6641 4675 6699 4681
rect 6641 4672 6653 4675
rect 6503 4644 6653 4672
rect 6503 4641 6515 4644
rect 6457 4635 6515 4641
rect 6641 4641 6653 4644
rect 6687 4641 6699 4675
rect 6641 4635 6699 4641
rect 2498 4564 2504 4616
rect 2556 4604 2562 4616
rect 2556 4576 2601 4604
rect 2556 4564 2562 4576
rect 2774 4564 2780 4616
rect 2832 4604 2838 4616
rect 4522 4604 4528 4616
rect 2832 4576 2877 4604
rect 4483 4576 4528 4604
rect 2832 4564 2838 4576
rect 4522 4564 4528 4576
rect 4580 4564 4586 4616
rect 4801 4607 4859 4613
rect 4801 4573 4813 4607
rect 4847 4604 4859 4607
rect 12434 4604 12440 4616
rect 4847 4576 12440 4604
rect 4847 4573 4859 4576
rect 4801 4567 4859 4573
rect 12434 4564 12440 4576
rect 12492 4564 12498 4616
rect 4985 4539 5043 4545
rect 4985 4505 4997 4539
rect 5031 4536 5043 4539
rect 5442 4536 5448 4548
rect 5031 4508 5448 4536
rect 5031 4505 5043 4508
rect 4985 4499 5043 4505
rect 5442 4496 5448 4508
rect 5500 4496 5506 4548
rect 5537 4539 5595 4545
rect 5537 4505 5549 4539
rect 5583 4536 5595 4539
rect 6178 4536 6184 4548
rect 5583 4508 6184 4536
rect 5583 4505 5595 4508
rect 5537 4499 5595 4505
rect 6178 4496 6184 4508
rect 6236 4496 6242 4548
rect 6546 4496 6552 4548
rect 6604 4536 6610 4548
rect 6641 4539 6699 4545
rect 6641 4536 6653 4539
rect 6604 4508 6653 4536
rect 6604 4496 6610 4508
rect 6641 4505 6653 4508
rect 6687 4536 6699 4539
rect 14182 4536 14188 4548
rect 6687 4508 14188 4536
rect 6687 4505 6699 4508
rect 6641 4499 6699 4505
rect 14182 4496 14188 4508
rect 14240 4496 14246 4548
rect 3878 4468 3884 4480
rect 2424 4440 3884 4468
rect 3878 4428 3884 4440
rect 3936 4428 3942 4480
rect 5626 4428 5632 4480
rect 5684 4468 5690 4480
rect 5813 4471 5871 4477
rect 5813 4468 5825 4471
rect 5684 4440 5825 4468
rect 5684 4428 5690 4440
rect 5813 4437 5825 4440
rect 5859 4437 5871 4471
rect 5813 4431 5871 4437
rect 920 4378 7084 4400
rect 920 4326 2098 4378
rect 2150 4326 2162 4378
rect 2214 4326 2226 4378
rect 2278 4326 2290 4378
rect 2342 4326 5098 4378
rect 5150 4326 5162 4378
rect 5214 4326 5226 4378
rect 5278 4326 5290 4378
rect 5342 4326 7084 4378
rect 920 4304 7084 4326
rect 1476 4267 1534 4273
rect 1476 4233 1488 4267
rect 1522 4264 1534 4267
rect 2774 4264 2780 4276
rect 1522 4236 2780 4264
rect 1522 4233 1534 4236
rect 1476 4227 1534 4233
rect 2774 4224 2780 4236
rect 2832 4224 2838 4276
rect 3510 4264 3516 4276
rect 3471 4236 3516 4264
rect 3510 4224 3516 4236
rect 3568 4224 3574 4276
rect 4144 4267 4202 4273
rect 4144 4233 4156 4267
rect 4190 4264 4202 4267
rect 4706 4264 4712 4276
rect 4190 4236 4712 4264
rect 4190 4233 4202 4236
rect 4144 4227 4202 4233
rect 4706 4224 4712 4236
rect 4764 4224 4770 4276
rect 5442 4224 5448 4276
rect 5500 4264 5506 4276
rect 13722 4264 13728 4276
rect 5500 4236 13728 4264
rect 5500 4224 5506 4236
rect 13722 4224 13728 4236
rect 13780 4224 13786 4276
rect 14090 4196 14096 4208
rect 6288 4168 14096 4196
rect 1213 4131 1271 4137
rect 1213 4097 1225 4131
rect 1259 4128 1271 4131
rect 3050 4128 3056 4140
rect 1259 4100 3056 4128
rect 1259 4097 1271 4100
rect 1213 4091 1271 4097
rect 3050 4088 3056 4100
rect 3108 4128 3114 4140
rect 3881 4131 3939 4137
rect 3881 4128 3893 4131
rect 3108 4100 3893 4128
rect 3108 4088 3114 4100
rect 3881 4097 3893 4100
rect 3927 4097 3939 4131
rect 3881 4091 3939 4097
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 5905 4131 5963 4137
rect 5905 4128 5917 4131
rect 4948 4100 5917 4128
rect 4948 4088 4954 4100
rect 5905 4097 5917 4100
rect 5951 4097 5963 4131
rect 5905 4091 5963 4097
rect 5994 4088 6000 4140
rect 6052 4128 6058 4140
rect 6052 4100 6097 4128
rect 6052 4088 6058 4100
rect 6288 4072 6316 4168
rect 14090 4156 14096 4168
rect 14148 4156 14154 4208
rect 2958 4020 2964 4072
rect 3016 4060 3022 4072
rect 3326 4060 3332 4072
rect 3016 4032 3332 4060
rect 3016 4020 3022 4032
rect 3326 4020 3332 4032
rect 3384 4020 3390 4072
rect 6178 4060 6184 4072
rect 6139 4032 6184 4060
rect 6178 4020 6184 4032
rect 6236 4020 6242 4072
rect 6270 4020 6276 4072
rect 6328 4060 6334 4072
rect 6328 4032 6421 4060
rect 6328 4020 6334 4032
rect 1946 3952 1952 4004
rect 2004 3952 2010 4004
rect 3237 3995 3295 4001
rect 3237 3961 3249 3995
rect 3283 3961 3295 3995
rect 3237 3955 3295 3961
rect 1670 3884 1676 3936
rect 1728 3924 1734 3936
rect 3252 3924 3280 3955
rect 4614 3952 4620 4004
rect 4672 3952 4678 4004
rect 6086 3952 6092 4004
rect 6144 3992 6150 4004
rect 6733 3995 6791 4001
rect 6733 3992 6745 3995
rect 6144 3964 6745 3992
rect 6144 3952 6150 3964
rect 6733 3961 6745 3964
rect 6779 3961 6791 3995
rect 6733 3955 6791 3961
rect 1728 3896 3280 3924
rect 1728 3884 1734 3896
rect 5994 3884 6000 3936
rect 6052 3924 6058 3936
rect 6362 3924 6368 3936
rect 6052 3896 6368 3924
rect 6052 3884 6058 3896
rect 6362 3884 6368 3896
rect 6420 3884 6426 3936
rect 920 3834 7084 3856
rect 920 3782 3598 3834
rect 3650 3782 3662 3834
rect 3714 3782 3726 3834
rect 3778 3782 3790 3834
rect 3842 3782 7084 3834
rect 920 3760 7084 3782
rect 2590 3680 2596 3732
rect 2648 3720 2654 3732
rect 6181 3723 6239 3729
rect 6181 3720 6193 3723
rect 2648 3692 6193 3720
rect 2648 3680 2654 3692
rect 6181 3689 6193 3692
rect 6227 3689 6239 3723
rect 6181 3683 6239 3689
rect 2866 3652 2872 3664
rect 2827 3624 2872 3652
rect 2866 3612 2872 3624
rect 2924 3612 2930 3664
rect 3418 3612 3424 3664
rect 3476 3612 3482 3664
rect 5813 3655 5871 3661
rect 5813 3621 5825 3655
rect 5859 3652 5871 3655
rect 5859 3624 6132 3652
rect 5859 3621 5871 3624
rect 5813 3615 5871 3621
rect 6104 3596 6132 3624
rect 4801 3587 4859 3593
rect 4801 3553 4813 3587
rect 4847 3584 4859 3587
rect 5169 3587 5227 3593
rect 5169 3584 5181 3587
rect 4847 3556 5181 3584
rect 4847 3553 4859 3556
rect 4801 3547 4859 3553
rect 5169 3553 5181 3556
rect 5215 3584 5227 3587
rect 5534 3584 5540 3596
rect 5215 3556 5540 3584
rect 5215 3553 5227 3556
rect 5169 3547 5227 3553
rect 5534 3544 5540 3556
rect 5592 3544 5598 3596
rect 5902 3584 5908 3596
rect 5863 3556 5908 3584
rect 5902 3544 5908 3556
rect 5960 3544 5966 3596
rect 6086 3584 6092 3596
rect 6047 3556 6092 3584
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 1578 3476 1584 3528
rect 1636 3516 1642 3528
rect 2498 3516 2504 3528
rect 1636 3488 2504 3516
rect 1636 3476 1642 3488
rect 2498 3476 2504 3488
rect 2556 3516 2562 3528
rect 2593 3519 2651 3525
rect 2593 3516 2605 3519
rect 2556 3488 2605 3516
rect 2556 3476 2562 3488
rect 2593 3485 2605 3488
rect 2639 3516 2651 3519
rect 4246 3516 4252 3528
rect 2639 3488 4252 3516
rect 2639 3485 2651 3488
rect 2593 3479 2651 3485
rect 4246 3476 4252 3488
rect 4304 3476 4310 3528
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3516 4675 3519
rect 14090 3516 14096 3528
rect 4663 3488 14096 3516
rect 4663 3485 4675 3488
rect 4617 3479 4675 3485
rect 14090 3476 14096 3488
rect 14148 3476 14154 3528
rect 4982 3380 4988 3392
rect 4943 3352 4988 3380
rect 4982 3340 4988 3352
rect 5040 3340 5046 3392
rect 5353 3383 5411 3389
rect 5353 3349 5365 3383
rect 5399 3380 5411 3383
rect 5534 3380 5540 3392
rect 5399 3352 5540 3380
rect 5399 3349 5411 3352
rect 5353 3343 5411 3349
rect 5534 3340 5540 3352
rect 5592 3340 5598 3392
rect 920 3290 7084 3312
rect 920 3238 2098 3290
rect 2150 3238 2162 3290
rect 2214 3238 2226 3290
rect 2278 3238 2290 3290
rect 2342 3238 5098 3290
rect 5150 3238 5162 3290
rect 5214 3238 5226 3290
rect 5278 3238 5290 3290
rect 5342 3238 7084 3290
rect 920 3216 7084 3238
rect 14274 3176 14280 3188
rect 3712 3148 14280 3176
rect 1670 3068 1676 3120
rect 1728 3068 1734 3120
rect 1688 3040 1716 3068
rect 3712 3049 3740 3148
rect 14274 3136 14280 3148
rect 14332 3136 14338 3188
rect 1949 3043 2007 3049
rect 1949 3040 1961 3043
rect 1688 3012 1961 3040
rect 1949 3009 1961 3012
rect 1995 3009 2007 3043
rect 1949 3003 2007 3009
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3009 3755 3043
rect 4798 3040 4804 3052
rect 4759 3012 4804 3040
rect 3697 3003 3755 3009
rect 4798 3000 4804 3012
rect 4856 3000 4862 3052
rect 6270 3040 6276 3052
rect 4908 3012 6132 3040
rect 6231 3012 6276 3040
rect 1578 2932 1584 2984
rect 1636 2972 1642 2984
rect 1673 2975 1731 2981
rect 1673 2972 1685 2975
rect 1636 2944 1685 2972
rect 1636 2932 1642 2944
rect 1673 2941 1685 2944
rect 1719 2941 1731 2975
rect 1673 2935 1731 2941
rect 3234 2932 3240 2984
rect 3292 2972 3298 2984
rect 3881 2975 3939 2981
rect 3881 2972 3893 2975
rect 3292 2944 3893 2972
rect 3292 2932 3298 2944
rect 3881 2941 3893 2944
rect 3927 2941 3939 2975
rect 3881 2935 3939 2941
rect 4246 2932 4252 2984
rect 4304 2972 4310 2984
rect 4433 2975 4491 2981
rect 4433 2972 4445 2975
rect 4304 2944 4445 2972
rect 4304 2932 4310 2944
rect 4433 2941 4445 2944
rect 4479 2941 4491 2975
rect 4433 2935 4491 2941
rect 4522 2932 4528 2984
rect 4580 2972 4586 2984
rect 4908 2972 4936 3012
rect 4580 2944 4936 2972
rect 6104 2972 6132 3012
rect 6270 3000 6276 3012
rect 6328 3000 6334 3052
rect 14182 2972 14188 2984
rect 6104 2944 14188 2972
rect 4580 2932 4586 2944
rect 14182 2932 14188 2944
rect 14240 2932 14246 2984
rect 3160 2836 3188 2890
rect 5534 2864 5540 2916
rect 5592 2864 5598 2916
rect 4065 2839 4123 2845
rect 4065 2836 4077 2839
rect 3160 2808 4077 2836
rect 4065 2805 4077 2808
rect 4111 2805 4123 2839
rect 4065 2799 4123 2805
rect 920 2746 7084 2768
rect 920 2694 3598 2746
rect 3650 2694 3662 2746
rect 3714 2694 3726 2746
rect 3778 2694 3790 2746
rect 3842 2694 7084 2746
rect 920 2672 7084 2694
rect 3418 2632 3424 2644
rect 3379 2604 3424 2632
rect 3418 2592 3424 2604
rect 3476 2592 3482 2644
rect 4982 2592 4988 2644
rect 5040 2632 5046 2644
rect 5040 2604 5304 2632
rect 5040 2592 5046 2604
rect 4706 2524 4712 2576
rect 4764 2564 4770 2576
rect 4801 2567 4859 2573
rect 4801 2564 4813 2567
rect 4764 2536 4813 2564
rect 4764 2524 4770 2536
rect 4801 2533 4813 2536
rect 4847 2533 4859 2567
rect 5276 2550 5304 2604
rect 6546 2564 6552 2576
rect 6507 2536 6552 2564
rect 4801 2527 4859 2533
rect 6546 2524 6552 2536
rect 6604 2524 6610 2576
rect 3142 2456 3148 2508
rect 3200 2496 3206 2508
rect 3237 2499 3295 2505
rect 3237 2496 3249 2499
rect 3200 2468 3249 2496
rect 3200 2456 3206 2468
rect 3237 2465 3249 2468
rect 3283 2465 3295 2499
rect 3237 2459 3295 2465
rect 4246 2456 4252 2508
rect 4304 2496 4310 2508
rect 4525 2499 4583 2505
rect 4525 2496 4537 2499
rect 4304 2468 4537 2496
rect 4304 2456 4310 2468
rect 4525 2465 4537 2468
rect 4571 2465 4583 2499
rect 4525 2459 4583 2465
rect 920 2202 7084 2224
rect 920 2150 2098 2202
rect 2150 2150 2162 2202
rect 2214 2150 2226 2202
rect 2278 2150 2290 2202
rect 2342 2150 5098 2202
rect 5150 2150 5162 2202
rect 5214 2150 5226 2202
rect 5278 2150 5290 2202
rect 5342 2150 7084 2202
rect 920 2128 7084 2150
rect 6362 1640 6368 1692
rect 6420 1680 6426 1692
rect 14182 1680 14188 1692
rect 6420 1652 14188 1680
rect 6420 1640 6426 1652
rect 14182 1640 14188 1652
rect 14240 1640 14246 1692
rect 6086 1504 6092 1556
rect 6144 1544 6150 1556
rect 14090 1544 14096 1556
rect 6144 1516 14096 1544
rect 6144 1504 6150 1516
rect 14090 1504 14096 1516
rect 14148 1504 14154 1556
rect 12434 1300 12440 1352
rect 12492 1340 12498 1352
rect 14182 1340 14188 1352
rect 12492 1312 14188 1340
rect 12492 1300 12498 1312
rect 14182 1300 14188 1312
rect 14240 1300 14246 1352
rect 6454 144 6460 196
rect 6512 184 6518 196
rect 14274 184 14280 196
rect 6512 156 14280 184
rect 6512 144 6518 156
rect 14274 144 14280 156
rect 14332 144 14338 196
<< via1 >>
rect 12532 12724 12584 12776
rect 14096 12724 14148 12776
rect 12440 12452 12492 12504
rect 14188 12452 14240 12504
rect -1610 11386 -1312 11462
rect 3598 11398 3650 11450
rect 3662 11398 3714 11450
rect 3726 11398 3778 11450
rect 3790 11398 3842 11450
rect 1952 11296 2004 11348
rect 14188 11296 14240 11348
rect 2780 11203 2832 11212
rect 2780 11169 2789 11203
rect 2789 11169 2823 11203
rect 2823 11169 2832 11203
rect 2780 11160 2832 11169
rect 3884 11160 3936 11212
rect 4436 11203 4488 11212
rect 4436 11169 4445 11203
rect 4445 11169 4479 11203
rect 4479 11169 4488 11203
rect 4436 11160 4488 11169
rect 6368 11203 6420 11212
rect 6368 11169 6377 11203
rect 6377 11169 6411 11203
rect 6411 11169 6420 11203
rect 6368 11160 6420 11169
rect 1216 10956 1268 11008
rect 3332 11067 3384 11076
rect 3332 11033 3341 11067
rect 3341 11033 3375 11067
rect 3375 11033 3384 11067
rect 3332 11024 3384 11033
rect 5448 11092 5500 11144
rect 13728 11160 13780 11212
rect 6644 11092 6696 11144
rect 14096 11092 14148 11144
rect 2964 10999 3016 11008
rect 2964 10965 2973 10999
rect 2973 10965 3007 10999
rect 3007 10965 3016 10999
rect 2964 10956 3016 10965
rect 4528 10956 4580 11008
rect -950 10842 -652 10918
rect 2098 10854 2150 10906
rect 2162 10854 2214 10906
rect 2226 10854 2278 10906
rect 2290 10854 2342 10906
rect 5098 10854 5150 10906
rect 5162 10854 5214 10906
rect 5226 10854 5278 10906
rect 5290 10854 5342 10906
rect 4436 10752 4488 10804
rect 1952 10659 2004 10668
rect 1952 10625 1961 10659
rect 1961 10625 1995 10659
rect 1995 10625 2004 10659
rect 1952 10616 2004 10625
rect 13268 10616 13320 10668
rect 14096 10616 14148 10668
rect 1216 10548 1268 10600
rect 4068 10591 4120 10600
rect 4068 10557 4077 10591
rect 4077 10557 4111 10591
rect 4111 10557 4120 10591
rect 4068 10548 4120 10557
rect 4436 10591 4488 10600
rect 4436 10557 4445 10591
rect 4445 10557 4479 10591
rect 4479 10557 4488 10591
rect 4436 10548 4488 10557
rect 6552 10591 6604 10600
rect 6552 10557 6561 10591
rect 6561 10557 6595 10591
rect 6595 10557 6604 10591
rect 6552 10548 6604 10557
rect 14188 10548 14240 10600
rect 3332 10480 3384 10532
rect 3424 10480 3476 10532
rect 4620 10480 4672 10532
rect 6092 10480 6144 10532
rect 14096 10480 14148 10532
rect 4252 10455 4304 10464
rect 4252 10421 4261 10455
rect 4261 10421 4295 10455
rect 4295 10421 4304 10455
rect 4252 10412 4304 10421
rect 3598 10310 3650 10362
rect 3662 10310 3714 10362
rect 3726 10310 3778 10362
rect 3790 10310 3842 10362
rect 6368 10251 6420 10260
rect 6368 10217 6377 10251
rect 6377 10217 6411 10251
rect 6411 10217 6420 10251
rect 6368 10208 6420 10217
rect 2964 10140 3016 10192
rect 4252 10140 4304 10192
rect 6552 10140 6604 10192
rect 1216 10047 1268 10056
rect 1216 10013 1225 10047
rect 1225 10013 1259 10047
rect 1259 10013 1268 10047
rect 1216 10004 1268 10013
rect 3424 10072 3476 10124
rect 4528 10072 4580 10124
rect 5448 10072 5500 10124
rect 6368 10072 6420 10124
rect 3148 10004 3200 10056
rect 2872 9936 2924 9988
rect 4988 10004 5040 10056
rect 3700 9868 3752 9920
rect 4436 9868 4488 9920
rect 5448 9868 5500 9920
rect 2098 9766 2150 9818
rect 2162 9766 2214 9818
rect 2226 9766 2278 9818
rect 2290 9766 2342 9818
rect 5098 9766 5150 9818
rect 5162 9766 5214 9818
rect 5226 9766 5278 9818
rect 5290 9766 5342 9818
rect 3240 9596 3292 9648
rect 5724 9664 5776 9716
rect 6092 9664 6144 9716
rect 6276 9596 6328 9648
rect 2320 9460 2372 9512
rect 2688 9503 2740 9512
rect 2688 9469 2697 9503
rect 2697 9469 2731 9503
rect 2731 9469 2740 9503
rect 2688 9460 2740 9469
rect 2964 9503 3016 9512
rect 2964 9469 2973 9503
rect 2973 9469 3007 9503
rect 3007 9469 3016 9503
rect 2964 9460 3016 9469
rect 6184 9528 6236 9580
rect 6460 9528 6512 9580
rect 14096 9528 14148 9580
rect 3424 9503 3476 9512
rect 3424 9469 3433 9503
rect 3433 9469 3467 9503
rect 3467 9469 3476 9503
rect 3424 9460 3476 9469
rect 3056 9392 3108 9444
rect 2780 9324 2832 9376
rect 2964 9324 3016 9376
rect 3332 9324 3384 9376
rect 3792 9460 3844 9512
rect 5632 9460 5684 9512
rect 6552 9460 6604 9512
rect 4160 9435 4212 9444
rect 4160 9401 4169 9435
rect 4169 9401 4203 9435
rect 4203 9401 4212 9435
rect 4160 9392 4212 9401
rect 5816 9392 5868 9444
rect 7196 9392 7248 9444
rect 14188 9392 14240 9444
rect 6092 9324 6144 9376
rect 6184 9367 6236 9376
rect 6184 9333 6193 9367
rect 6193 9333 6227 9367
rect 6227 9333 6236 9367
rect 6184 9324 6236 9333
rect 6552 9324 6604 9376
rect 3598 9222 3650 9274
rect 3662 9222 3714 9274
rect 3726 9222 3778 9274
rect 3790 9222 3842 9274
rect 5632 9163 5684 9172
rect 5632 9129 5641 9163
rect 5641 9129 5675 9163
rect 5675 9129 5684 9163
rect 5632 9120 5684 9129
rect 5816 9120 5868 9172
rect 6092 9120 6144 9172
rect 6552 9120 6604 9172
rect 2596 9052 2648 9104
rect 2320 9027 2372 9036
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 2320 8993 2329 9027
rect 2329 8993 2363 9027
rect 2363 8993 2372 9027
rect 2320 8984 2372 8993
rect 3332 9052 3384 9104
rect 4344 8984 4396 9036
rect 2504 8916 2556 8968
rect 2872 8916 2924 8968
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 3976 8916 4028 8968
rect 5448 9027 5500 9036
rect 5448 8993 5457 9027
rect 5457 8993 5491 9027
rect 5491 8993 5500 9027
rect 5448 8984 5500 8993
rect 5724 9052 5776 9104
rect 6092 8984 6144 9036
rect 6276 9027 6328 9036
rect 6276 8993 6285 9027
rect 6285 8993 6319 9027
rect 6319 8993 6328 9027
rect 6276 8984 6328 8993
rect 4988 8959 5040 8968
rect 4988 8925 4997 8959
rect 4997 8925 5031 8959
rect 5031 8925 5040 8959
rect 4988 8916 5040 8925
rect 4436 8848 4488 8900
rect 12532 8916 12584 8968
rect 6184 8780 6236 8832
rect 2098 8678 2150 8730
rect 2162 8678 2214 8730
rect 2226 8678 2278 8730
rect 2290 8678 2342 8730
rect 5098 8678 5150 8730
rect 5162 8678 5214 8730
rect 5226 8678 5278 8730
rect 5290 8678 5342 8730
rect 1216 8483 1268 8492
rect 1216 8449 1225 8483
rect 1225 8449 1259 8483
rect 1259 8449 1268 8483
rect 1216 8440 1268 8449
rect 3148 8576 3200 8628
rect 3976 8576 4028 8628
rect 4344 8576 4396 8628
rect 4252 8508 4304 8560
rect 3424 8440 3476 8492
rect 12440 8440 12492 8492
rect 3332 8415 3384 8424
rect 3332 8381 3341 8415
rect 3341 8381 3375 8415
rect 3375 8381 3384 8415
rect 3332 8372 3384 8381
rect 4068 8372 4120 8424
rect 3240 8347 3292 8356
rect 3240 8313 3249 8347
rect 3249 8313 3283 8347
rect 3283 8313 3292 8347
rect 3240 8304 3292 8313
rect 6092 8372 6144 8424
rect 4528 8304 4580 8356
rect 4712 8304 4764 8356
rect 6644 8304 6696 8356
rect 3148 8236 3200 8288
rect 4252 8236 4304 8288
rect 5448 8236 5500 8288
rect 3598 8134 3650 8186
rect 3662 8134 3714 8186
rect 3726 8134 3778 8186
rect 3790 8134 3842 8186
rect 3240 8032 3292 8084
rect 3148 7964 3200 8016
rect 3056 7896 3108 7948
rect 4436 8032 4488 8084
rect 6276 8032 6328 8084
rect 3976 7964 4028 8016
rect 3424 7896 3476 7948
rect 3884 7939 3936 7948
rect 3884 7905 3893 7939
rect 3893 7905 3927 7939
rect 3927 7905 3936 7939
rect 3884 7896 3936 7905
rect 6092 7896 6144 7948
rect 1216 7871 1268 7880
rect 1216 7837 1225 7871
rect 1225 7837 1259 7871
rect 1259 7837 1268 7871
rect 1216 7828 1268 7837
rect 3240 7871 3292 7880
rect 3240 7837 3249 7871
rect 3249 7837 3283 7871
rect 3283 7837 3292 7871
rect 3240 7828 3292 7837
rect 3976 7871 4028 7880
rect 3976 7837 3985 7871
rect 3985 7837 4019 7871
rect 4019 7837 4028 7871
rect 3976 7828 4028 7837
rect 3056 7760 3108 7812
rect 3148 7692 3200 7744
rect 3332 7692 3384 7744
rect 2098 7590 2150 7642
rect 2162 7590 2214 7642
rect 2226 7590 2278 7642
rect 2290 7590 2342 7642
rect 5098 7590 5150 7642
rect 5162 7590 5214 7642
rect 5226 7590 5278 7642
rect 5290 7590 5342 7642
rect 1400 7488 1452 7540
rect 2872 7420 2924 7472
rect 3884 7420 3936 7472
rect 3240 7352 3292 7404
rect 1308 7327 1360 7336
rect 1308 7293 1317 7327
rect 1317 7293 1351 7327
rect 1351 7293 1360 7327
rect 1308 7284 1360 7293
rect 3148 7284 3200 7336
rect 3884 7327 3936 7336
rect 3884 7293 3893 7327
rect 3893 7293 3927 7327
rect 3927 7293 3936 7327
rect 3884 7284 3936 7293
rect 6184 7327 6236 7336
rect 6184 7293 6193 7327
rect 6193 7293 6227 7327
rect 6227 7293 6236 7327
rect 6184 7284 6236 7293
rect 4068 7216 4120 7268
rect 4252 7216 4304 7268
rect 14188 7216 14240 7268
rect 6276 7191 6328 7200
rect 6276 7157 6285 7191
rect 6285 7157 6319 7191
rect 6319 7157 6328 7191
rect 6276 7148 6328 7157
rect 14096 7148 14148 7200
rect 3598 7046 3650 7098
rect 3662 7046 3714 7098
rect 3726 7046 3778 7098
rect 3790 7046 3842 7098
rect 3976 6944 4028 6996
rect 4252 6944 4304 6996
rect 3424 6876 3476 6928
rect 3884 6876 3936 6928
rect 6368 6944 6420 6996
rect 14188 6944 14240 6996
rect 6276 6876 6328 6928
rect 3056 6851 3108 6860
rect 3056 6817 3065 6851
rect 3065 6817 3099 6851
rect 3099 6817 3108 6851
rect 3056 6808 3108 6817
rect 4896 6808 4948 6860
rect 4804 6740 4856 6792
rect 4344 6672 4396 6724
rect 3148 6604 3200 6656
rect 6460 6783 6512 6792
rect 6460 6749 6469 6783
rect 6469 6749 6503 6783
rect 6503 6749 6512 6783
rect 6460 6740 6512 6749
rect 2098 6502 2150 6554
rect 2162 6502 2214 6554
rect 2226 6502 2278 6554
rect 2290 6502 2342 6554
rect 5098 6502 5150 6554
rect 5162 6502 5214 6554
rect 5226 6502 5278 6554
rect 5290 6502 5342 6554
rect 13268 6400 13320 6452
rect 4068 6264 4120 6316
rect 1216 6239 1268 6248
rect 1216 6205 1225 6239
rect 1225 6205 1259 6239
rect 1259 6205 1268 6239
rect 1216 6196 1268 6205
rect 3148 6196 3200 6248
rect 3884 6239 3936 6248
rect 3884 6205 3893 6239
rect 3893 6205 3927 6239
rect 3927 6205 3936 6239
rect 3884 6196 3936 6205
rect 4252 6196 4304 6248
rect 6092 6196 6144 6248
rect 2872 6128 2924 6180
rect 4068 6103 4120 6112
rect 4068 6069 4077 6103
rect 4077 6069 4111 6103
rect 4111 6069 4120 6103
rect 4068 6060 4120 6069
rect 14096 6128 14148 6180
rect 3598 5958 3650 6010
rect 3662 5958 3714 6010
rect 3726 5958 3778 6010
rect 3790 5958 3842 6010
rect 4620 5856 4672 5908
rect 2412 5788 2464 5840
rect 4068 5788 4120 5840
rect 3056 5720 3108 5772
rect 5540 5856 5592 5908
rect 1308 5652 1360 5704
rect 1676 5695 1728 5704
rect 1676 5661 1685 5695
rect 1685 5661 1719 5695
rect 1719 5661 1728 5695
rect 1676 5652 1728 5661
rect 4160 5652 4212 5704
rect 4436 5652 4488 5704
rect 6092 5720 6144 5772
rect 4988 5584 5040 5636
rect 14096 5584 14148 5636
rect 3056 5516 3108 5568
rect 6184 5559 6236 5568
rect 6184 5525 6193 5559
rect 6193 5525 6227 5559
rect 6227 5525 6236 5559
rect 6184 5516 6236 5525
rect 2098 5414 2150 5466
rect 2162 5414 2214 5466
rect 2226 5414 2278 5466
rect 2290 5414 2342 5466
rect 5098 5414 5150 5466
rect 5162 5414 5214 5466
rect 5226 5414 5278 5466
rect 5290 5414 5342 5466
rect 3884 5312 3936 5364
rect 1216 5219 1268 5228
rect 1216 5185 1225 5219
rect 1225 5185 1259 5219
rect 1259 5185 1268 5219
rect 1216 5176 1268 5185
rect 2872 5176 2924 5228
rect 4436 5176 4488 5228
rect 6644 5176 6696 5228
rect 3884 5108 3936 5160
rect 4252 5108 4304 5160
rect 1584 5040 1636 5092
rect 2780 5040 2832 5092
rect 6184 5040 6236 5092
rect 4620 4972 4672 5024
rect 3598 4870 3650 4922
rect 3662 4870 3714 4922
rect 3726 4870 3778 4922
rect 3790 4870 3842 4922
rect 1584 4811 1636 4820
rect 1584 4777 1593 4811
rect 1593 4777 1627 4811
rect 1627 4777 1636 4811
rect 1584 4768 1636 4777
rect 2412 4768 2464 4820
rect 3148 4768 3200 4820
rect 5448 4768 5500 4820
rect 3516 4700 3568 4752
rect 14188 4972 14240 5024
rect 1952 4471 2004 4480
rect 1952 4437 1961 4471
rect 1961 4437 1995 4471
rect 1995 4437 2004 4471
rect 1952 4428 2004 4437
rect 4436 4632 4488 4684
rect 6092 4632 6144 4684
rect 2504 4607 2556 4616
rect 2504 4573 2513 4607
rect 2513 4573 2547 4607
rect 2547 4573 2556 4607
rect 2504 4564 2556 4573
rect 2780 4607 2832 4616
rect 2780 4573 2789 4607
rect 2789 4573 2823 4607
rect 2823 4573 2832 4607
rect 4528 4607 4580 4616
rect 2780 4564 2832 4573
rect 4528 4573 4537 4607
rect 4537 4573 4571 4607
rect 4571 4573 4580 4607
rect 4528 4564 4580 4573
rect 12440 4564 12492 4616
rect 5448 4496 5500 4548
rect 6184 4496 6236 4548
rect 6552 4496 6604 4548
rect 14188 4496 14240 4548
rect 3884 4428 3936 4480
rect 5632 4428 5684 4480
rect 2098 4326 2150 4378
rect 2162 4326 2214 4378
rect 2226 4326 2278 4378
rect 2290 4326 2342 4378
rect 5098 4326 5150 4378
rect 5162 4326 5214 4378
rect 5226 4326 5278 4378
rect 5290 4326 5342 4378
rect 2780 4224 2832 4276
rect 3516 4267 3568 4276
rect 3516 4233 3525 4267
rect 3525 4233 3559 4267
rect 3559 4233 3568 4267
rect 3516 4224 3568 4233
rect 4712 4224 4764 4276
rect 5448 4224 5500 4276
rect 13728 4224 13780 4276
rect 3056 4088 3108 4140
rect 4896 4088 4948 4140
rect 6000 4131 6052 4140
rect 6000 4097 6009 4131
rect 6009 4097 6043 4131
rect 6043 4097 6052 4131
rect 6000 4088 6052 4097
rect 14096 4156 14148 4208
rect 2964 4020 3016 4072
rect 3332 4063 3384 4072
rect 3332 4029 3341 4063
rect 3341 4029 3375 4063
rect 3375 4029 3384 4063
rect 3332 4020 3384 4029
rect 6184 4063 6236 4072
rect 6184 4029 6193 4063
rect 6193 4029 6227 4063
rect 6227 4029 6236 4063
rect 6184 4020 6236 4029
rect 6276 4063 6328 4072
rect 6276 4029 6285 4063
rect 6285 4029 6319 4063
rect 6319 4029 6328 4063
rect 6276 4020 6328 4029
rect 1952 3952 2004 4004
rect 1676 3884 1728 3936
rect 4620 3952 4672 4004
rect 6092 3952 6144 4004
rect 6000 3884 6052 3936
rect 6368 3884 6420 3936
rect 3598 3782 3650 3834
rect 3662 3782 3714 3834
rect 3726 3782 3778 3834
rect 3790 3782 3842 3834
rect 2596 3680 2648 3732
rect 2872 3655 2924 3664
rect 2872 3621 2881 3655
rect 2881 3621 2915 3655
rect 2915 3621 2924 3655
rect 2872 3612 2924 3621
rect 3424 3612 3476 3664
rect 5540 3544 5592 3596
rect 5908 3587 5960 3596
rect 5908 3553 5917 3587
rect 5917 3553 5951 3587
rect 5951 3553 5960 3587
rect 5908 3544 5960 3553
rect 6092 3587 6144 3596
rect 6092 3553 6101 3587
rect 6101 3553 6135 3587
rect 6135 3553 6144 3587
rect 6092 3544 6144 3553
rect 1584 3476 1636 3528
rect 2504 3476 2556 3528
rect 4252 3476 4304 3528
rect 14096 3476 14148 3528
rect 4988 3383 5040 3392
rect 4988 3349 4997 3383
rect 4997 3349 5031 3383
rect 5031 3349 5040 3383
rect 4988 3340 5040 3349
rect 5540 3340 5592 3392
rect 2098 3238 2150 3290
rect 2162 3238 2214 3290
rect 2226 3238 2278 3290
rect 2290 3238 2342 3290
rect 5098 3238 5150 3290
rect 5162 3238 5214 3290
rect 5226 3238 5278 3290
rect 5290 3238 5342 3290
rect 1676 3068 1728 3120
rect 14280 3136 14332 3188
rect 4804 3043 4856 3052
rect 4804 3009 4813 3043
rect 4813 3009 4847 3043
rect 4847 3009 4856 3043
rect 4804 3000 4856 3009
rect 6276 3043 6328 3052
rect 1584 2932 1636 2984
rect 3240 2932 3292 2984
rect 4252 2932 4304 2984
rect 4528 2932 4580 2984
rect 6276 3009 6285 3043
rect 6285 3009 6319 3043
rect 6319 3009 6328 3043
rect 6276 3000 6328 3009
rect 14188 2932 14240 2984
rect 5540 2864 5592 2916
rect 3598 2694 3650 2746
rect 3662 2694 3714 2746
rect 3726 2694 3778 2746
rect 3790 2694 3842 2746
rect 3424 2635 3476 2644
rect 3424 2601 3433 2635
rect 3433 2601 3467 2635
rect 3467 2601 3476 2635
rect 3424 2592 3476 2601
rect 4988 2592 5040 2644
rect 4712 2524 4764 2576
rect 6552 2567 6604 2576
rect 6552 2533 6561 2567
rect 6561 2533 6595 2567
rect 6595 2533 6604 2567
rect 6552 2524 6604 2533
rect 3148 2456 3200 2508
rect 4252 2456 4304 2508
rect 2098 2150 2150 2202
rect 2162 2150 2214 2202
rect 2226 2150 2278 2202
rect 2290 2150 2342 2202
rect 5098 2150 5150 2202
rect 5162 2150 5214 2202
rect 5226 2150 5278 2202
rect 5290 2150 5342 2202
rect 6368 1640 6420 1692
rect 14188 1640 14240 1692
rect 6092 1504 6144 1556
rect 14096 1504 14148 1556
rect 12440 1300 12492 1352
rect 14188 1300 14240 1352
rect 6460 144 6512 196
rect 14280 144 14332 196
<< metal2 >>
rect 14094 13696 14150 13705
rect 14094 13631 14150 13640
rect 14108 12782 14136 13631
rect 14186 13152 14242 13161
rect 14186 13087 14242 13096
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 12440 12504 12492 12510
rect 12440 12446 12492 12452
rect -1620 11462 -1300 11472
rect -1620 11386 -1610 11462
rect -1312 11386 -1300 11462
rect -1620 11376 -1300 11386
rect 3572 11452 3868 11472
rect 3628 11450 3652 11452
rect 3708 11450 3732 11452
rect 3788 11450 3812 11452
rect 3650 11398 3652 11450
rect 3714 11398 3726 11450
rect 3788 11398 3790 11450
rect 3628 11396 3652 11398
rect 3708 11396 3732 11398
rect 3788 11396 3812 11398
rect 3572 11376 3868 11396
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 1216 11008 1268 11014
rect 1216 10950 1268 10956
rect -960 10918 -640 10928
rect -960 10842 -950 10918
rect -652 10842 -640 10918
rect -960 10832 -640 10842
rect 1228 10606 1256 10950
rect 1964 10674 1992 11290
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 4436 11212 4488 11218
rect 4436 11154 4488 11160
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 2072 10908 2368 10928
rect 2128 10906 2152 10908
rect 2208 10906 2232 10908
rect 2288 10906 2312 10908
rect 2150 10854 2152 10906
rect 2214 10854 2226 10906
rect 2288 10854 2290 10906
rect 2128 10852 2152 10854
rect 2208 10852 2232 10854
rect 2288 10852 2312 10854
rect 2072 10832 2368 10852
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 1216 10600 1268 10606
rect 1216 10542 1268 10548
rect 1228 10062 1256 10542
rect 1216 10056 1268 10062
rect 1216 9998 1268 10004
rect 1228 8498 1256 9998
rect 2072 9820 2368 9840
rect 2128 9818 2152 9820
rect 2208 9818 2232 9820
rect 2288 9818 2312 9820
rect 2150 9766 2152 9818
rect 2214 9766 2226 9818
rect 2288 9766 2290 9818
rect 2128 9764 2152 9766
rect 2208 9764 2232 9766
rect 2288 9764 2312 9766
rect 2072 9744 2368 9764
rect 2686 9616 2742 9625
rect 2686 9551 2742 9560
rect 2700 9518 2728 9551
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2332 9042 2360 9454
rect 2792 9382 2820 11154
rect 3332 11076 3384 11082
rect 3332 11018 3384 11024
rect 2964 11008 3016 11014
rect 2964 10950 3016 10956
rect 2976 10198 3004 10950
rect 3344 10538 3372 11018
rect 3332 10532 3384 10538
rect 3332 10474 3384 10480
rect 3424 10532 3476 10538
rect 3424 10474 3476 10480
rect 2964 10192 3016 10198
rect 2964 10134 3016 10140
rect 3436 10130 3464 10474
rect 3572 10364 3868 10384
rect 3628 10362 3652 10364
rect 3708 10362 3732 10364
rect 3788 10362 3812 10364
rect 3650 10310 3652 10362
rect 3714 10310 3726 10362
rect 3788 10310 3790 10362
rect 3628 10308 3652 10310
rect 3708 10308 3732 10310
rect 3788 10308 3812 10310
rect 3572 10288 3868 10308
rect 3424 10124 3476 10130
rect 3424 10066 3476 10072
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 2872 9988 2924 9994
rect 2872 9930 2924 9936
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2596 9104 2648 9110
rect 2596 9046 2648 9052
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 1400 8968 1452 8974
rect 2504 8968 2556 8974
rect 1400 8910 1452 8916
rect 2502 8936 2504 8945
rect 2556 8936 2558 8945
rect 1216 8492 1268 8498
rect 1216 8434 1268 8440
rect 1216 7880 1268 7886
rect 1216 7822 1268 7828
rect 1228 7426 1256 7822
rect 1412 7546 1440 8910
rect 2502 8871 2558 8880
rect 2072 8732 2368 8752
rect 2128 8730 2152 8732
rect 2208 8730 2232 8732
rect 2288 8730 2312 8732
rect 2150 8678 2152 8730
rect 2214 8678 2226 8730
rect 2288 8678 2290 8730
rect 2128 8676 2152 8678
rect 2208 8676 2232 8678
rect 2288 8676 2312 8678
rect 2072 8656 2368 8676
rect 2072 7644 2368 7664
rect 2128 7642 2152 7644
rect 2208 7642 2232 7644
rect 2288 7642 2312 7644
rect 2150 7590 2152 7642
rect 2214 7590 2226 7642
rect 2288 7590 2290 7642
rect 2128 7588 2152 7590
rect 2208 7588 2232 7590
rect 2288 7588 2312 7590
rect 2072 7568 2368 7588
rect 1400 7540 1452 7546
rect 1400 7482 1452 7488
rect 1228 7398 1348 7426
rect 1320 7342 1348 7398
rect 1308 7336 1360 7342
rect 1308 7278 1360 7284
rect 1216 6248 1268 6254
rect 1320 6202 1348 7278
rect 2072 6556 2368 6576
rect 2128 6554 2152 6556
rect 2208 6554 2232 6556
rect 2288 6554 2312 6556
rect 2150 6502 2152 6554
rect 2214 6502 2226 6554
rect 2288 6502 2290 6554
rect 2128 6500 2152 6502
rect 2208 6500 2232 6502
rect 2288 6500 2312 6502
rect 2072 6480 2368 6500
rect 1268 6196 1348 6202
rect 1216 6190 1348 6196
rect 1228 6174 1348 6190
rect 1320 5710 1348 6174
rect 2412 5840 2464 5846
rect 2412 5782 2464 5788
rect 1308 5704 1360 5710
rect 1228 5652 1308 5658
rect 1228 5646 1360 5652
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1228 5630 1348 5646
rect 1228 5234 1256 5630
rect 1216 5228 1268 5234
rect 1216 5170 1268 5176
rect 1584 5092 1636 5098
rect 1584 5034 1636 5040
rect 1596 4826 1624 5034
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 1688 3942 1716 5646
rect 2072 5468 2368 5488
rect 2128 5466 2152 5468
rect 2208 5466 2232 5468
rect 2288 5466 2312 5468
rect 2150 5414 2152 5466
rect 2214 5414 2226 5466
rect 2288 5414 2290 5466
rect 2128 5412 2152 5414
rect 2208 5412 2232 5414
rect 2288 5412 2312 5414
rect 2072 5392 2368 5412
rect 2424 4826 2452 5782
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 1952 4480 2004 4486
rect 1952 4422 2004 4428
rect 1964 4010 1992 4422
rect 2072 4380 2368 4400
rect 2128 4378 2152 4380
rect 2208 4378 2232 4380
rect 2288 4378 2312 4380
rect 2150 4326 2152 4378
rect 2214 4326 2226 4378
rect 2288 4326 2290 4378
rect 2128 4324 2152 4326
rect 2208 4324 2232 4326
rect 2288 4324 2312 4326
rect 2072 4304 2368 4324
rect 1952 4004 2004 4010
rect 1952 3946 2004 3952
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 1596 2990 1624 3470
rect 1688 3126 1716 3878
rect 2516 3534 2544 4558
rect 2608 3738 2636 9046
rect 2884 8974 2912 9930
rect 2964 9512 3016 9518
rect 2962 9480 2964 9489
rect 3016 9480 3018 9489
rect 2962 9415 3018 9424
rect 3056 9444 3108 9450
rect 3056 9386 3108 9392
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2884 7478 2912 8910
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 2872 6180 2924 6186
rect 2872 6122 2924 6128
rect 2884 5234 2912 6122
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2780 5092 2832 5098
rect 2780 5034 2832 5040
rect 2792 4622 2820 5034
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 2792 4282 2820 4558
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 2884 3670 2912 5170
rect 2976 4078 3004 9318
rect 3068 7954 3096 9386
rect 3160 8634 3188 9998
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 3252 9081 3280 9590
rect 3424 9512 3476 9518
rect 3712 9500 3740 9862
rect 3792 9512 3844 9518
rect 3712 9472 3792 9500
rect 3424 9454 3476 9460
rect 3792 9454 3844 9460
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3344 9110 3372 9318
rect 3332 9104 3384 9110
rect 3238 9072 3294 9081
rect 3332 9046 3384 9052
rect 3238 9007 3294 9016
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3252 8362 3280 8910
rect 3436 8498 3464 9454
rect 3572 9276 3868 9296
rect 3628 9274 3652 9276
rect 3708 9274 3732 9276
rect 3788 9274 3812 9276
rect 3650 9222 3652 9274
rect 3714 9222 3726 9274
rect 3788 9222 3790 9274
rect 3628 9220 3652 9222
rect 3708 9220 3732 9222
rect 3788 9220 3812 9222
rect 3572 9200 3868 9220
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 3160 8022 3188 8230
rect 3252 8090 3280 8298
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3148 8016 3200 8022
rect 3148 7958 3200 7964
rect 3056 7948 3108 7954
rect 3056 7890 3108 7896
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3056 7812 3108 7818
rect 3056 7754 3108 7760
rect 3068 6866 3096 7754
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 3160 7342 3188 7686
rect 3252 7410 3280 7822
rect 3344 7750 3372 8366
rect 3572 8188 3868 8208
rect 3628 8186 3652 8188
rect 3708 8186 3732 8188
rect 3788 8186 3812 8188
rect 3650 8134 3652 8186
rect 3714 8134 3726 8186
rect 3788 8134 3790 8186
rect 3628 8132 3652 8134
rect 3708 8132 3732 8134
rect 3788 8132 3812 8134
rect 3572 8112 3868 8132
rect 3896 7954 3924 11154
rect 4448 10810 4476 11154
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 4540 10690 4568 10950
rect 5072 10908 5368 10928
rect 5128 10906 5152 10908
rect 5208 10906 5232 10908
rect 5288 10906 5312 10908
rect 5150 10854 5152 10906
rect 5214 10854 5226 10906
rect 5288 10854 5290 10906
rect 5128 10852 5152 10854
rect 5208 10852 5232 10854
rect 5288 10852 5312 10854
rect 5072 10832 5368 10852
rect 4448 10662 4568 10690
rect 4448 10606 4476 10662
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 4436 10600 4488 10606
rect 4436 10542 4488 10548
rect 3976 8968 4028 8974
rect 4080 8956 4108 10542
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 4264 10198 4292 10406
rect 4252 10192 4304 10198
rect 4252 10134 4304 10140
rect 4448 9926 4476 10542
rect 4620 10532 4672 10538
rect 4620 10474 4672 10480
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 4028 8928 4108 8956
rect 3976 8910 4028 8916
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 3988 8022 4016 8570
rect 4080 8430 4108 8928
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 3976 8016 4028 8022
rect 3976 7958 4028 7964
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 3884 7948 3936 7954
rect 3884 7890 3936 7896
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 3068 5778 3096 6802
rect 3160 6662 3188 7278
rect 3436 6934 3464 7890
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 3896 7342 3924 7414
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3896 7154 3924 7278
rect 3988 7154 4016 7822
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 3896 7126 4016 7154
rect 3572 7100 3868 7120
rect 3628 7098 3652 7100
rect 3708 7098 3732 7100
rect 3788 7098 3812 7100
rect 3650 7046 3652 7098
rect 3714 7046 3726 7098
rect 3788 7046 3790 7098
rect 3628 7044 3652 7046
rect 3708 7044 3732 7046
rect 3788 7044 3812 7046
rect 3572 7024 3868 7044
rect 3988 7002 4016 7126
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 3424 6928 3476 6934
rect 3424 6870 3476 6876
rect 3884 6928 3936 6934
rect 3884 6870 3936 6876
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3160 6254 3188 6598
rect 3896 6254 3924 6870
rect 4080 6322 4108 7210
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 3068 5574 3096 5714
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 3068 4146 3096 5510
rect 3160 4826 3188 6190
rect 3572 6012 3868 6032
rect 3628 6010 3652 6012
rect 3708 6010 3732 6012
rect 3788 6010 3812 6012
rect 3650 5958 3652 6010
rect 3714 5958 3726 6010
rect 3788 5958 3790 6010
rect 3628 5956 3652 5958
rect 3708 5956 3732 5958
rect 3788 5956 3812 5958
rect 3572 5936 3868 5956
rect 3896 5370 3924 6190
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4080 5846 4108 6054
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 4172 5710 4200 9386
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4356 8634 4384 8978
rect 4436 8900 4488 8906
rect 4436 8842 4488 8848
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4252 8560 4304 8566
rect 4252 8502 4304 8508
rect 4264 8378 4292 8502
rect 4264 8350 4384 8378
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4264 7274 4292 8230
rect 4252 7268 4304 7274
rect 4252 7210 4304 7216
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4264 6254 4292 6938
rect 4356 6730 4384 8350
rect 4448 8090 4476 8842
rect 4540 8362 4568 10066
rect 4528 8356 4580 8362
rect 4528 8298 4580 8304
rect 4436 8084 4488 8090
rect 4436 8026 4488 8032
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 3896 5166 3924 5306
rect 4264 5166 4292 6190
rect 4448 5710 4476 8026
rect 4632 5914 4660 10474
rect 5460 10130 5488 11086
rect 6092 10532 6144 10538
rect 6092 10474 6144 10480
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 5000 9625 5028 9998
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 5072 9820 5368 9840
rect 5128 9818 5152 9820
rect 5208 9818 5232 9820
rect 5288 9818 5312 9820
rect 5150 9766 5152 9818
rect 5214 9766 5226 9818
rect 5288 9766 5290 9818
rect 5128 9764 5152 9766
rect 5208 9764 5232 9766
rect 5288 9764 5312 9766
rect 5072 9744 5368 9764
rect 4986 9616 5042 9625
rect 4986 9551 5042 9560
rect 5460 9042 5488 9862
rect 6104 9722 6132 10474
rect 6380 10266 6408 11154
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6564 10198 6592 10542
rect 6552 10192 6604 10198
rect 6552 10134 6604 10140
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5644 9178 5672 9454
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5736 9110 5764 9658
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6196 9489 6224 9522
rect 5998 9480 6054 9489
rect 5816 9444 5868 9450
rect 5998 9415 6054 9424
rect 6182 9480 6238 9489
rect 6182 9415 6238 9424
rect 5816 9386 5868 9392
rect 5828 9178 5856 9386
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5724 9104 5776 9110
rect 5724 9046 5776 9052
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 5630 8936 5686 8945
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4724 8242 4752 8298
rect 4724 8214 4844 8242
rect 4816 6798 4844 8214
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4448 5234 4476 5646
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 3572 4924 3868 4944
rect 3628 4922 3652 4924
rect 3708 4922 3732 4924
rect 3788 4922 3812 4924
rect 3650 4870 3652 4922
rect 3714 4870 3726 4922
rect 3788 4870 3790 4922
rect 3628 4868 3652 4870
rect 3708 4868 3732 4870
rect 3788 4868 3812 4870
rect 3572 4848 3868 4868
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3516 4752 3568 4758
rect 3516 4694 3568 4700
rect 3528 4282 3556 4694
rect 3896 4486 3924 5102
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 3516 4276 3568 4282
rect 3516 4218 3568 4224
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 2964 4072 3016 4078
rect 3332 4072 3384 4078
rect 2964 4014 3016 4020
rect 3252 4020 3332 4026
rect 3252 4014 3384 4020
rect 3252 3998 3372 4014
rect 2872 3664 2924 3670
rect 2872 3606 2924 3612
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 2072 3292 2368 3312
rect 2128 3290 2152 3292
rect 2208 3290 2232 3292
rect 2288 3290 2312 3292
rect 2150 3238 2152 3290
rect 2214 3238 2226 3290
rect 2288 3238 2290 3290
rect 2128 3236 2152 3238
rect 2208 3236 2232 3238
rect 2288 3236 2312 3238
rect 2072 3216 2368 3236
rect 1676 3120 1728 3126
rect 1676 3062 1728 3068
rect 3252 2990 3280 3998
rect 3572 3836 3868 3856
rect 3628 3834 3652 3836
rect 3708 3834 3732 3836
rect 3788 3834 3812 3836
rect 3650 3782 3652 3834
rect 3714 3782 3726 3834
rect 3788 3782 3790 3834
rect 3628 3780 3652 3782
rect 3708 3780 3732 3782
rect 3788 3780 3812 3782
rect 3572 3760 3868 3780
rect 3424 3664 3476 3670
rect 3424 3606 3476 3612
rect 1584 2984 1636 2990
rect 1584 2926 1636 2932
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 3252 2774 3280 2926
rect 3160 2746 3280 2774
rect 3160 2514 3188 2746
rect 3436 2650 3464 3606
rect 4264 3534 4292 5102
rect 4448 4690 4476 5170
rect 4632 5114 4660 5850
rect 4632 5086 4752 5114
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4436 4684 4488 4690
rect 4436 4626 4488 4632
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4264 2990 4292 3470
rect 4540 2990 4568 4558
rect 4632 4010 4660 4966
rect 4724 4282 4752 5086
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4816 3058 4844 6734
rect 4908 4146 4936 6802
rect 5000 5642 5028 8910
rect 5630 8871 5686 8880
rect 5072 8732 5368 8752
rect 5128 8730 5152 8732
rect 5208 8730 5232 8732
rect 5288 8730 5312 8732
rect 5150 8678 5152 8730
rect 5214 8678 5226 8730
rect 5288 8678 5290 8730
rect 5128 8676 5152 8678
rect 5208 8676 5232 8678
rect 5288 8676 5312 8678
rect 5072 8656 5368 8676
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5072 7644 5368 7664
rect 5128 7642 5152 7644
rect 5208 7642 5232 7644
rect 5288 7642 5312 7644
rect 5150 7590 5152 7642
rect 5214 7590 5226 7642
rect 5288 7590 5290 7642
rect 5128 7588 5152 7590
rect 5208 7588 5232 7590
rect 5288 7588 5312 7590
rect 5072 7568 5368 7588
rect 5072 6556 5368 6576
rect 5128 6554 5152 6556
rect 5208 6554 5232 6556
rect 5288 6554 5312 6556
rect 5150 6502 5152 6554
rect 5214 6502 5226 6554
rect 5288 6502 5290 6554
rect 5128 6500 5152 6502
rect 5208 6500 5232 6502
rect 5288 6500 5312 6502
rect 5072 6480 5368 6500
rect 4988 5636 5040 5642
rect 4988 5578 5040 5584
rect 5072 5468 5368 5488
rect 5128 5466 5152 5468
rect 5208 5466 5232 5468
rect 5288 5466 5312 5468
rect 5150 5414 5152 5466
rect 5214 5414 5226 5466
rect 5288 5414 5290 5466
rect 5128 5412 5152 5414
rect 5208 5412 5232 5414
rect 5288 5412 5312 5414
rect 5072 5392 5368 5412
rect 5460 4826 5488 8230
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5448 4548 5500 4554
rect 5448 4490 5500 4496
rect 5072 4380 5368 4400
rect 5128 4378 5152 4380
rect 5208 4378 5232 4380
rect 5288 4378 5312 4380
rect 5150 4326 5152 4378
rect 5214 4326 5226 4378
rect 5288 4326 5290 4378
rect 5128 4324 5152 4326
rect 5208 4324 5232 4326
rect 5288 4324 5312 4326
rect 5072 4304 5368 4324
rect 5460 4282 5488 4490
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 4252 2984 4304 2990
rect 4252 2926 4304 2932
rect 4528 2984 4580 2990
rect 4528 2926 4580 2932
rect 3572 2748 3868 2768
rect 3628 2746 3652 2748
rect 3708 2746 3732 2748
rect 3788 2746 3812 2748
rect 3650 2694 3652 2746
rect 3714 2694 3726 2746
rect 3788 2694 3790 2746
rect 3628 2692 3652 2694
rect 3708 2692 3732 2694
rect 3788 2692 3812 2694
rect 3572 2672 3868 2692
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 4264 2514 4292 2926
rect 4908 2774 4936 4082
rect 5552 3602 5580 5850
rect 5644 4486 5672 8871
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 6012 4146 6040 9415
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 6184 9376 6236 9382
rect 6288 9364 6316 9590
rect 6236 9336 6316 9364
rect 6184 9318 6236 9324
rect 6104 9178 6132 9318
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6104 8430 6132 8978
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 6104 6254 6132 7890
rect 6196 7342 6224 8774
rect 6288 8090 6316 8978
rect 6276 8084 6328 8090
rect 6276 8026 6328 8032
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6288 6934 6316 7142
rect 6380 7002 6408 10066
rect 6550 9616 6606 9625
rect 6460 9580 6512 9586
rect 6550 9551 6606 9560
rect 6460 9522 6512 9528
rect 6472 9081 6500 9522
rect 6564 9518 6592 9551
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6564 9178 6592 9318
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6458 9072 6514 9081
rect 6458 9007 6514 9016
rect 6656 8362 6684 11086
rect 7194 9480 7250 9489
rect 7194 9415 7196 9424
rect 7248 9415 7250 9424
rect 7196 9386 7248 9392
rect 12452 8498 12480 12446
rect 12544 8974 12572 12718
rect 14094 12608 14150 12617
rect 13740 12566 14094 12594
rect 13740 11218 13768 12566
rect 14094 12543 14150 12552
rect 14200 12510 14228 13087
rect 14188 12504 14240 12510
rect 14188 12446 14240 12452
rect 14094 12064 14150 12073
rect 14094 11999 14150 12008
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 14108 11150 14136 11999
rect 14186 11520 14242 11529
rect 14186 11455 14242 11464
rect 14200 11354 14228 11455
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 14094 10976 14150 10985
rect 14094 10911 14150 10920
rect 14108 10674 14136 10911
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 6276 6928 6328 6934
rect 6276 6870 6328 6876
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 6104 5778 6132 6190
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 6196 5098 6224 5510
rect 6184 5092 6236 5098
rect 6184 5034 6236 5040
rect 6092 4684 6144 4690
rect 6092 4626 6144 4632
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 6012 3942 6040 4082
rect 6104 4010 6132 4626
rect 6184 4548 6236 4554
rect 6184 4490 6236 4496
rect 6196 4078 6224 4490
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 6092 4004 6144 4010
rect 6092 3946 6144 3952
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 6104 3720 6132 3946
rect 6012 3692 6132 3720
rect 6012 3618 6040 3692
rect 5920 3602 6040 3618
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5908 3596 6040 3602
rect 5960 3590 6040 3596
rect 6092 3596 6144 3602
rect 5908 3538 5960 3544
rect 6092 3538 6144 3544
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 4724 2746 4936 2774
rect 4724 2582 4752 2746
rect 5000 2650 5028 3334
rect 5072 3292 5368 3312
rect 5128 3290 5152 3292
rect 5208 3290 5232 3292
rect 5288 3290 5312 3292
rect 5150 3238 5152 3290
rect 5214 3238 5226 3290
rect 5288 3238 5290 3290
rect 5128 3236 5152 3238
rect 5208 3236 5232 3238
rect 5288 3236 5312 3238
rect 5072 3216 5368 3236
rect 5552 2922 5580 3334
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 3148 2508 3200 2514
rect 3148 2450 3200 2456
rect 4252 2508 4304 2514
rect 4252 2450 4304 2456
rect 2072 2204 2368 2224
rect 2128 2202 2152 2204
rect 2208 2202 2232 2204
rect 2288 2202 2312 2204
rect 2150 2150 2152 2202
rect 2214 2150 2226 2202
rect 2288 2150 2290 2202
rect 2128 2148 2152 2150
rect 2208 2148 2232 2150
rect 2288 2148 2312 2150
rect 2072 2128 2368 2148
rect 5072 2204 5368 2224
rect 5128 2202 5152 2204
rect 5208 2202 5232 2204
rect 5288 2202 5312 2204
rect 5150 2150 5152 2202
rect 5214 2150 5226 2202
rect 5288 2150 5290 2202
rect 5128 2148 5152 2150
rect 5208 2148 5232 2150
rect 5288 2148 5312 2150
rect 5072 2128 5368 2148
rect 6104 1562 6132 3538
rect 6288 3058 6316 4014
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 6380 1698 6408 3878
rect 6368 1692 6420 1698
rect 6368 1634 6420 1640
rect 6092 1556 6144 1562
rect 6092 1498 6144 1504
rect 6472 202 6500 6734
rect 6656 5234 6684 8298
rect 13280 6458 13308 10610
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 14096 10532 14148 10538
rect 14096 10474 14148 10480
rect 14108 9897 14136 10474
rect 14200 10441 14228 10542
rect 14186 10432 14242 10441
rect 14186 10367 14242 10376
rect 14094 9888 14150 9897
rect 14094 9823 14150 9832
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14108 8809 14136 9522
rect 14188 9444 14240 9450
rect 14188 9386 14240 9392
rect 14200 9353 14228 9386
rect 14186 9344 14242 9353
rect 14186 9279 14242 9288
rect 14094 8800 14150 8809
rect 14094 8735 14150 8744
rect 14094 8256 14150 8265
rect 14094 8191 14150 8200
rect 14108 7206 14136 8191
rect 14186 7712 14242 7721
rect 14186 7647 14242 7656
rect 14200 7274 14228 7647
rect 14188 7268 14240 7274
rect 14188 7210 14240 7216
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 14186 7168 14242 7177
rect 14186 7103 14242 7112
rect 14200 7002 14228 7103
rect 14188 6996 14240 7002
rect 14188 6938 14240 6944
rect 14094 6624 14150 6633
rect 14094 6559 14150 6568
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 14108 6186 14136 6559
rect 14096 6180 14148 6186
rect 14096 6122 14148 6128
rect 14094 6080 14150 6089
rect 14094 6015 14150 6024
rect 14108 5642 14136 6015
rect 14096 5636 14148 5642
rect 14096 5578 14148 5584
rect 14186 5536 14242 5545
rect 14186 5471 14242 5480
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 14200 5030 14228 5471
rect 14188 5024 14240 5030
rect 14094 4992 14150 5001
rect 14188 4966 14240 4972
rect 14094 4927 14150 4936
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 6552 4548 6604 4554
rect 6552 4490 6604 4496
rect 6564 2582 6592 4490
rect 6552 2576 6604 2582
rect 6552 2518 6604 2524
rect 12452 1358 12480 4558
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 12440 1352 12492 1358
rect 12440 1294 12492 1300
rect 13740 1306 13768 4218
rect 14108 4214 14136 4927
rect 14188 4548 14240 4554
rect 14188 4490 14240 4496
rect 14200 4457 14228 4490
rect 14186 4448 14242 4457
rect 14186 4383 14242 4392
rect 14096 4208 14148 4214
rect 14096 4150 14148 4156
rect 14186 3904 14242 3913
rect 14186 3839 14242 3848
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 14108 2825 14136 3470
rect 14200 2990 14228 3839
rect 14278 3360 14334 3369
rect 14278 3295 14334 3304
rect 14292 3194 14320 3295
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 14094 2816 14150 2825
rect 14094 2751 14150 2760
rect 14094 2272 14150 2281
rect 14094 2207 14150 2216
rect 14108 1562 14136 2207
rect 14186 1728 14242 1737
rect 14186 1663 14188 1672
rect 14240 1663 14242 1672
rect 14188 1634 14240 1640
rect 14096 1556 14148 1562
rect 14096 1498 14148 1504
rect 14188 1352 14240 1358
rect 13740 1278 14136 1306
rect 14188 1294 14240 1300
rect 14108 241 14136 1278
rect 14200 649 14228 1294
rect 14278 1184 14334 1193
rect 14278 1119 14334 1128
rect 14186 640 14242 649
rect 14186 575 14242 584
rect 14094 232 14150 241
rect 6460 196 6512 202
rect 14292 202 14320 1119
rect 14094 167 14150 176
rect 14280 196 14332 202
rect 6460 138 6512 144
rect 14280 138 14332 144
<< via2 >>
rect 14094 13640 14150 13696
rect 14186 13096 14242 13152
rect -1610 11386 -1312 11462
rect 3572 11450 3628 11452
rect 3652 11450 3708 11452
rect 3732 11450 3788 11452
rect 3812 11450 3868 11452
rect 3572 11398 3598 11450
rect 3598 11398 3628 11450
rect 3652 11398 3662 11450
rect 3662 11398 3708 11450
rect 3732 11398 3778 11450
rect 3778 11398 3788 11450
rect 3812 11398 3842 11450
rect 3842 11398 3868 11450
rect 3572 11396 3628 11398
rect 3652 11396 3708 11398
rect 3732 11396 3788 11398
rect 3812 11396 3868 11398
rect -950 10842 -652 10918
rect 2072 10906 2128 10908
rect 2152 10906 2208 10908
rect 2232 10906 2288 10908
rect 2312 10906 2368 10908
rect 2072 10854 2098 10906
rect 2098 10854 2128 10906
rect 2152 10854 2162 10906
rect 2162 10854 2208 10906
rect 2232 10854 2278 10906
rect 2278 10854 2288 10906
rect 2312 10854 2342 10906
rect 2342 10854 2368 10906
rect 2072 10852 2128 10854
rect 2152 10852 2208 10854
rect 2232 10852 2288 10854
rect 2312 10852 2368 10854
rect 2072 9818 2128 9820
rect 2152 9818 2208 9820
rect 2232 9818 2288 9820
rect 2312 9818 2368 9820
rect 2072 9766 2098 9818
rect 2098 9766 2128 9818
rect 2152 9766 2162 9818
rect 2162 9766 2208 9818
rect 2232 9766 2278 9818
rect 2278 9766 2288 9818
rect 2312 9766 2342 9818
rect 2342 9766 2368 9818
rect 2072 9764 2128 9766
rect 2152 9764 2208 9766
rect 2232 9764 2288 9766
rect 2312 9764 2368 9766
rect 2686 9560 2742 9616
rect 3572 10362 3628 10364
rect 3652 10362 3708 10364
rect 3732 10362 3788 10364
rect 3812 10362 3868 10364
rect 3572 10310 3598 10362
rect 3598 10310 3628 10362
rect 3652 10310 3662 10362
rect 3662 10310 3708 10362
rect 3732 10310 3778 10362
rect 3778 10310 3788 10362
rect 3812 10310 3842 10362
rect 3842 10310 3868 10362
rect 3572 10308 3628 10310
rect 3652 10308 3708 10310
rect 3732 10308 3788 10310
rect 3812 10308 3868 10310
rect 2502 8916 2504 8936
rect 2504 8916 2556 8936
rect 2556 8916 2558 8936
rect 2502 8880 2558 8916
rect 2072 8730 2128 8732
rect 2152 8730 2208 8732
rect 2232 8730 2288 8732
rect 2312 8730 2368 8732
rect 2072 8678 2098 8730
rect 2098 8678 2128 8730
rect 2152 8678 2162 8730
rect 2162 8678 2208 8730
rect 2232 8678 2278 8730
rect 2278 8678 2288 8730
rect 2312 8678 2342 8730
rect 2342 8678 2368 8730
rect 2072 8676 2128 8678
rect 2152 8676 2208 8678
rect 2232 8676 2288 8678
rect 2312 8676 2368 8678
rect 2072 7642 2128 7644
rect 2152 7642 2208 7644
rect 2232 7642 2288 7644
rect 2312 7642 2368 7644
rect 2072 7590 2098 7642
rect 2098 7590 2128 7642
rect 2152 7590 2162 7642
rect 2162 7590 2208 7642
rect 2232 7590 2278 7642
rect 2278 7590 2288 7642
rect 2312 7590 2342 7642
rect 2342 7590 2368 7642
rect 2072 7588 2128 7590
rect 2152 7588 2208 7590
rect 2232 7588 2288 7590
rect 2312 7588 2368 7590
rect 2072 6554 2128 6556
rect 2152 6554 2208 6556
rect 2232 6554 2288 6556
rect 2312 6554 2368 6556
rect 2072 6502 2098 6554
rect 2098 6502 2128 6554
rect 2152 6502 2162 6554
rect 2162 6502 2208 6554
rect 2232 6502 2278 6554
rect 2278 6502 2288 6554
rect 2312 6502 2342 6554
rect 2342 6502 2368 6554
rect 2072 6500 2128 6502
rect 2152 6500 2208 6502
rect 2232 6500 2288 6502
rect 2312 6500 2368 6502
rect 2072 5466 2128 5468
rect 2152 5466 2208 5468
rect 2232 5466 2288 5468
rect 2312 5466 2368 5468
rect 2072 5414 2098 5466
rect 2098 5414 2128 5466
rect 2152 5414 2162 5466
rect 2162 5414 2208 5466
rect 2232 5414 2278 5466
rect 2278 5414 2288 5466
rect 2312 5414 2342 5466
rect 2342 5414 2368 5466
rect 2072 5412 2128 5414
rect 2152 5412 2208 5414
rect 2232 5412 2288 5414
rect 2312 5412 2368 5414
rect 2072 4378 2128 4380
rect 2152 4378 2208 4380
rect 2232 4378 2288 4380
rect 2312 4378 2368 4380
rect 2072 4326 2098 4378
rect 2098 4326 2128 4378
rect 2152 4326 2162 4378
rect 2162 4326 2208 4378
rect 2232 4326 2278 4378
rect 2278 4326 2288 4378
rect 2312 4326 2342 4378
rect 2342 4326 2368 4378
rect 2072 4324 2128 4326
rect 2152 4324 2208 4326
rect 2232 4324 2288 4326
rect 2312 4324 2368 4326
rect 2962 9460 2964 9480
rect 2964 9460 3016 9480
rect 3016 9460 3018 9480
rect 2962 9424 3018 9460
rect 3238 9016 3294 9072
rect 3572 9274 3628 9276
rect 3652 9274 3708 9276
rect 3732 9274 3788 9276
rect 3812 9274 3868 9276
rect 3572 9222 3598 9274
rect 3598 9222 3628 9274
rect 3652 9222 3662 9274
rect 3662 9222 3708 9274
rect 3732 9222 3778 9274
rect 3778 9222 3788 9274
rect 3812 9222 3842 9274
rect 3842 9222 3868 9274
rect 3572 9220 3628 9222
rect 3652 9220 3708 9222
rect 3732 9220 3788 9222
rect 3812 9220 3868 9222
rect 3572 8186 3628 8188
rect 3652 8186 3708 8188
rect 3732 8186 3788 8188
rect 3812 8186 3868 8188
rect 3572 8134 3598 8186
rect 3598 8134 3628 8186
rect 3652 8134 3662 8186
rect 3662 8134 3708 8186
rect 3732 8134 3778 8186
rect 3778 8134 3788 8186
rect 3812 8134 3842 8186
rect 3842 8134 3868 8186
rect 3572 8132 3628 8134
rect 3652 8132 3708 8134
rect 3732 8132 3788 8134
rect 3812 8132 3868 8134
rect 5072 10906 5128 10908
rect 5152 10906 5208 10908
rect 5232 10906 5288 10908
rect 5312 10906 5368 10908
rect 5072 10854 5098 10906
rect 5098 10854 5128 10906
rect 5152 10854 5162 10906
rect 5162 10854 5208 10906
rect 5232 10854 5278 10906
rect 5278 10854 5288 10906
rect 5312 10854 5342 10906
rect 5342 10854 5368 10906
rect 5072 10852 5128 10854
rect 5152 10852 5208 10854
rect 5232 10852 5288 10854
rect 5312 10852 5368 10854
rect 3572 7098 3628 7100
rect 3652 7098 3708 7100
rect 3732 7098 3788 7100
rect 3812 7098 3868 7100
rect 3572 7046 3598 7098
rect 3598 7046 3628 7098
rect 3652 7046 3662 7098
rect 3662 7046 3708 7098
rect 3732 7046 3778 7098
rect 3778 7046 3788 7098
rect 3812 7046 3842 7098
rect 3842 7046 3868 7098
rect 3572 7044 3628 7046
rect 3652 7044 3708 7046
rect 3732 7044 3788 7046
rect 3812 7044 3868 7046
rect 3572 6010 3628 6012
rect 3652 6010 3708 6012
rect 3732 6010 3788 6012
rect 3812 6010 3868 6012
rect 3572 5958 3598 6010
rect 3598 5958 3628 6010
rect 3652 5958 3662 6010
rect 3662 5958 3708 6010
rect 3732 5958 3778 6010
rect 3778 5958 3788 6010
rect 3812 5958 3842 6010
rect 3842 5958 3868 6010
rect 3572 5956 3628 5958
rect 3652 5956 3708 5958
rect 3732 5956 3788 5958
rect 3812 5956 3868 5958
rect 5072 9818 5128 9820
rect 5152 9818 5208 9820
rect 5232 9818 5288 9820
rect 5312 9818 5368 9820
rect 5072 9766 5098 9818
rect 5098 9766 5128 9818
rect 5152 9766 5162 9818
rect 5162 9766 5208 9818
rect 5232 9766 5278 9818
rect 5278 9766 5288 9818
rect 5312 9766 5342 9818
rect 5342 9766 5368 9818
rect 5072 9764 5128 9766
rect 5152 9764 5208 9766
rect 5232 9764 5288 9766
rect 5312 9764 5368 9766
rect 4986 9560 5042 9616
rect 5998 9424 6054 9480
rect 6182 9424 6238 9480
rect 3572 4922 3628 4924
rect 3652 4922 3708 4924
rect 3732 4922 3788 4924
rect 3812 4922 3868 4924
rect 3572 4870 3598 4922
rect 3598 4870 3628 4922
rect 3652 4870 3662 4922
rect 3662 4870 3708 4922
rect 3732 4870 3778 4922
rect 3778 4870 3788 4922
rect 3812 4870 3842 4922
rect 3842 4870 3868 4922
rect 3572 4868 3628 4870
rect 3652 4868 3708 4870
rect 3732 4868 3788 4870
rect 3812 4868 3868 4870
rect 2072 3290 2128 3292
rect 2152 3290 2208 3292
rect 2232 3290 2288 3292
rect 2312 3290 2368 3292
rect 2072 3238 2098 3290
rect 2098 3238 2128 3290
rect 2152 3238 2162 3290
rect 2162 3238 2208 3290
rect 2232 3238 2278 3290
rect 2278 3238 2288 3290
rect 2312 3238 2342 3290
rect 2342 3238 2368 3290
rect 2072 3236 2128 3238
rect 2152 3236 2208 3238
rect 2232 3236 2288 3238
rect 2312 3236 2368 3238
rect 3572 3834 3628 3836
rect 3652 3834 3708 3836
rect 3732 3834 3788 3836
rect 3812 3834 3868 3836
rect 3572 3782 3598 3834
rect 3598 3782 3628 3834
rect 3652 3782 3662 3834
rect 3662 3782 3708 3834
rect 3732 3782 3778 3834
rect 3778 3782 3788 3834
rect 3812 3782 3842 3834
rect 3842 3782 3868 3834
rect 3572 3780 3628 3782
rect 3652 3780 3708 3782
rect 3732 3780 3788 3782
rect 3812 3780 3868 3782
rect 5630 8880 5686 8936
rect 5072 8730 5128 8732
rect 5152 8730 5208 8732
rect 5232 8730 5288 8732
rect 5312 8730 5368 8732
rect 5072 8678 5098 8730
rect 5098 8678 5128 8730
rect 5152 8678 5162 8730
rect 5162 8678 5208 8730
rect 5232 8678 5278 8730
rect 5278 8678 5288 8730
rect 5312 8678 5342 8730
rect 5342 8678 5368 8730
rect 5072 8676 5128 8678
rect 5152 8676 5208 8678
rect 5232 8676 5288 8678
rect 5312 8676 5368 8678
rect 5072 7642 5128 7644
rect 5152 7642 5208 7644
rect 5232 7642 5288 7644
rect 5312 7642 5368 7644
rect 5072 7590 5098 7642
rect 5098 7590 5128 7642
rect 5152 7590 5162 7642
rect 5162 7590 5208 7642
rect 5232 7590 5278 7642
rect 5278 7590 5288 7642
rect 5312 7590 5342 7642
rect 5342 7590 5368 7642
rect 5072 7588 5128 7590
rect 5152 7588 5208 7590
rect 5232 7588 5288 7590
rect 5312 7588 5368 7590
rect 5072 6554 5128 6556
rect 5152 6554 5208 6556
rect 5232 6554 5288 6556
rect 5312 6554 5368 6556
rect 5072 6502 5098 6554
rect 5098 6502 5128 6554
rect 5152 6502 5162 6554
rect 5162 6502 5208 6554
rect 5232 6502 5278 6554
rect 5278 6502 5288 6554
rect 5312 6502 5342 6554
rect 5342 6502 5368 6554
rect 5072 6500 5128 6502
rect 5152 6500 5208 6502
rect 5232 6500 5288 6502
rect 5312 6500 5368 6502
rect 5072 5466 5128 5468
rect 5152 5466 5208 5468
rect 5232 5466 5288 5468
rect 5312 5466 5368 5468
rect 5072 5414 5098 5466
rect 5098 5414 5128 5466
rect 5152 5414 5162 5466
rect 5162 5414 5208 5466
rect 5232 5414 5278 5466
rect 5278 5414 5288 5466
rect 5312 5414 5342 5466
rect 5342 5414 5368 5466
rect 5072 5412 5128 5414
rect 5152 5412 5208 5414
rect 5232 5412 5288 5414
rect 5312 5412 5368 5414
rect 5072 4378 5128 4380
rect 5152 4378 5208 4380
rect 5232 4378 5288 4380
rect 5312 4378 5368 4380
rect 5072 4326 5098 4378
rect 5098 4326 5128 4378
rect 5152 4326 5162 4378
rect 5162 4326 5208 4378
rect 5232 4326 5278 4378
rect 5278 4326 5288 4378
rect 5312 4326 5342 4378
rect 5342 4326 5368 4378
rect 5072 4324 5128 4326
rect 5152 4324 5208 4326
rect 5232 4324 5288 4326
rect 5312 4324 5368 4326
rect 3572 2746 3628 2748
rect 3652 2746 3708 2748
rect 3732 2746 3788 2748
rect 3812 2746 3868 2748
rect 3572 2694 3598 2746
rect 3598 2694 3628 2746
rect 3652 2694 3662 2746
rect 3662 2694 3708 2746
rect 3732 2694 3778 2746
rect 3778 2694 3788 2746
rect 3812 2694 3842 2746
rect 3842 2694 3868 2746
rect 3572 2692 3628 2694
rect 3652 2692 3708 2694
rect 3732 2692 3788 2694
rect 3812 2692 3868 2694
rect 6550 9560 6606 9616
rect 6458 9016 6514 9072
rect 7194 9444 7250 9480
rect 7194 9424 7196 9444
rect 7196 9424 7248 9444
rect 7248 9424 7250 9444
rect 14094 12552 14150 12608
rect 14094 12008 14150 12064
rect 14186 11464 14242 11520
rect 14094 10920 14150 10976
rect 5072 3290 5128 3292
rect 5152 3290 5208 3292
rect 5232 3290 5288 3292
rect 5312 3290 5368 3292
rect 5072 3238 5098 3290
rect 5098 3238 5128 3290
rect 5152 3238 5162 3290
rect 5162 3238 5208 3290
rect 5232 3238 5278 3290
rect 5278 3238 5288 3290
rect 5312 3238 5342 3290
rect 5342 3238 5368 3290
rect 5072 3236 5128 3238
rect 5152 3236 5208 3238
rect 5232 3236 5288 3238
rect 5312 3236 5368 3238
rect 2072 2202 2128 2204
rect 2152 2202 2208 2204
rect 2232 2202 2288 2204
rect 2312 2202 2368 2204
rect 2072 2150 2098 2202
rect 2098 2150 2128 2202
rect 2152 2150 2162 2202
rect 2162 2150 2208 2202
rect 2232 2150 2278 2202
rect 2278 2150 2288 2202
rect 2312 2150 2342 2202
rect 2342 2150 2368 2202
rect 2072 2148 2128 2150
rect 2152 2148 2208 2150
rect 2232 2148 2288 2150
rect 2312 2148 2368 2150
rect 5072 2202 5128 2204
rect 5152 2202 5208 2204
rect 5232 2202 5288 2204
rect 5312 2202 5368 2204
rect 5072 2150 5098 2202
rect 5098 2150 5128 2202
rect 5152 2150 5162 2202
rect 5162 2150 5208 2202
rect 5232 2150 5278 2202
rect 5278 2150 5288 2202
rect 5312 2150 5342 2202
rect 5342 2150 5368 2202
rect 5072 2148 5128 2150
rect 5152 2148 5208 2150
rect 5232 2148 5288 2150
rect 5312 2148 5368 2150
rect 14186 10376 14242 10432
rect 14094 9832 14150 9888
rect 14186 9288 14242 9344
rect 14094 8744 14150 8800
rect 14094 8200 14150 8256
rect 14186 7656 14242 7712
rect 14186 7112 14242 7168
rect 14094 6568 14150 6624
rect 14094 6024 14150 6080
rect 14186 5480 14242 5536
rect 14094 4936 14150 4992
rect 14186 4392 14242 4448
rect 14186 3848 14242 3904
rect 14278 3304 14334 3360
rect 14094 2760 14150 2816
rect 14094 2216 14150 2272
rect 14186 1692 14242 1728
rect 14186 1672 14188 1692
rect 14188 1672 14240 1692
rect 14240 1672 14242 1692
rect 14278 1128 14334 1184
rect 14186 584 14242 640
rect 14094 176 14150 232
<< metal3 >>
rect 14000 13696 34000 13728
rect 14000 13640 14094 13696
rect 14150 13640 34000 13696
rect 14000 13608 34000 13640
rect 14000 13152 34000 13184
rect 14000 13096 14186 13152
rect 14242 13096 34000 13152
rect 14000 13064 34000 13096
rect 14000 12608 34000 12640
rect 14000 12552 14094 12608
rect 14150 12552 34000 12608
rect 14000 12520 34000 12552
rect 14000 12064 34000 12096
rect 14000 12008 14094 12064
rect 14150 12008 34000 12064
rect 14000 11976 34000 12008
rect 14000 11520 34000 11552
rect -1620 11462 -1300 11472
rect -1620 11386 -1610 11462
rect -1312 11386 -1300 11462
rect 14000 11464 14186 11520
rect 14242 11464 34000 11520
rect 3560 11456 3880 11457
rect 3560 11392 3568 11456
rect 3632 11392 3648 11456
rect 3712 11392 3728 11456
rect 3792 11392 3808 11456
rect 3872 11392 3880 11456
rect 14000 11432 34000 11464
rect 3560 11391 3880 11392
rect -1620 11376 -1300 11386
rect 14000 10976 34000 11008
rect -960 10918 -640 10928
rect -960 10842 -950 10918
rect -652 10842 -640 10918
rect 14000 10920 14094 10976
rect 14150 10920 34000 10976
rect 2060 10912 2380 10913
rect 2060 10848 2068 10912
rect 2132 10848 2148 10912
rect 2212 10848 2228 10912
rect 2292 10848 2308 10912
rect 2372 10848 2380 10912
rect 2060 10847 2380 10848
rect 5060 10912 5380 10913
rect 5060 10848 5068 10912
rect 5132 10848 5148 10912
rect 5212 10848 5228 10912
rect 5292 10848 5308 10912
rect 5372 10848 5380 10912
rect 14000 10888 34000 10920
rect 5060 10847 5380 10848
rect -960 10832 -640 10842
rect 14000 10432 34000 10464
rect 14000 10376 14186 10432
rect 14242 10376 34000 10432
rect 3560 10368 3880 10369
rect 3560 10304 3568 10368
rect 3632 10304 3648 10368
rect 3712 10304 3728 10368
rect 3792 10304 3808 10368
rect 3872 10304 3880 10368
rect 14000 10344 34000 10376
rect 3560 10303 3880 10304
rect 14000 9888 34000 9920
rect 14000 9832 14094 9888
rect 14150 9832 34000 9888
rect 2060 9824 2380 9825
rect 2060 9760 2068 9824
rect 2132 9760 2148 9824
rect 2212 9760 2228 9824
rect 2292 9760 2308 9824
rect 2372 9760 2380 9824
rect 2060 9759 2380 9760
rect 5060 9824 5380 9825
rect 5060 9760 5068 9824
rect 5132 9760 5148 9824
rect 5212 9760 5228 9824
rect 5292 9760 5308 9824
rect 5372 9760 5380 9824
rect 14000 9800 34000 9832
rect 5060 9759 5380 9760
rect 2681 9618 2747 9621
rect 4981 9618 5047 9621
rect 6545 9618 6611 9621
rect 2681 9616 6611 9618
rect 2681 9560 2686 9616
rect 2742 9560 4986 9616
rect 5042 9560 6550 9616
rect 6606 9560 6611 9616
rect 2681 9558 6611 9560
rect 2681 9555 2747 9558
rect 4981 9555 5047 9558
rect 6545 9555 6611 9558
rect 2957 9482 3023 9485
rect 5993 9482 6059 9485
rect 2957 9480 6059 9482
rect 2957 9424 2962 9480
rect 3018 9424 5998 9480
rect 6054 9424 6059 9480
rect 2957 9422 6059 9424
rect 2957 9419 3023 9422
rect 5993 9419 6059 9422
rect 6177 9482 6243 9485
rect 7189 9482 7255 9485
rect 6177 9480 7255 9482
rect 6177 9424 6182 9480
rect 6238 9424 7194 9480
rect 7250 9424 7255 9480
rect 6177 9422 7255 9424
rect 6177 9419 6243 9422
rect 7189 9419 7255 9422
rect 14000 9344 34000 9376
rect 14000 9288 14186 9344
rect 14242 9288 34000 9344
rect 3560 9280 3880 9281
rect 3560 9216 3568 9280
rect 3632 9216 3648 9280
rect 3712 9216 3728 9280
rect 3792 9216 3808 9280
rect 3872 9216 3880 9280
rect 14000 9256 34000 9288
rect 3560 9215 3880 9216
rect 3233 9074 3299 9077
rect 6453 9074 6519 9077
rect 3233 9072 6519 9074
rect 3233 9016 3238 9072
rect 3294 9016 6458 9072
rect 6514 9016 6519 9072
rect 3233 9014 6519 9016
rect 3233 9011 3299 9014
rect 6453 9011 6519 9014
rect 2497 8938 2563 8941
rect 5625 8938 5691 8941
rect 2497 8936 5691 8938
rect 2497 8880 2502 8936
rect 2558 8880 5630 8936
rect 5686 8880 5691 8936
rect 2497 8878 5691 8880
rect 2497 8875 2563 8878
rect 5625 8875 5691 8878
rect 14000 8800 34000 8832
rect 14000 8744 14094 8800
rect 14150 8744 34000 8800
rect 2060 8736 2380 8737
rect 2060 8672 2068 8736
rect 2132 8672 2148 8736
rect 2212 8672 2228 8736
rect 2292 8672 2308 8736
rect 2372 8672 2380 8736
rect 2060 8671 2380 8672
rect 5060 8736 5380 8737
rect 5060 8672 5068 8736
rect 5132 8672 5148 8736
rect 5212 8672 5228 8736
rect 5292 8672 5308 8736
rect 5372 8672 5380 8736
rect 14000 8712 34000 8744
rect 5060 8671 5380 8672
rect 14000 8256 34000 8288
rect 14000 8200 14094 8256
rect 14150 8200 34000 8256
rect 3560 8192 3880 8193
rect 3560 8128 3568 8192
rect 3632 8128 3648 8192
rect 3712 8128 3728 8192
rect 3792 8128 3808 8192
rect 3872 8128 3880 8192
rect 14000 8168 34000 8200
rect 3560 8127 3880 8128
rect 14000 7712 34000 7744
rect 14000 7656 14186 7712
rect 14242 7656 34000 7712
rect 2060 7648 2380 7649
rect 2060 7584 2068 7648
rect 2132 7584 2148 7648
rect 2212 7584 2228 7648
rect 2292 7584 2308 7648
rect 2372 7584 2380 7648
rect 2060 7583 2380 7584
rect 5060 7648 5380 7649
rect 5060 7584 5068 7648
rect 5132 7584 5148 7648
rect 5212 7584 5228 7648
rect 5292 7584 5308 7648
rect 5372 7584 5380 7648
rect 14000 7624 34000 7656
rect 5060 7583 5380 7584
rect 14000 7168 34000 7200
rect 14000 7112 14186 7168
rect 14242 7112 34000 7168
rect 3560 7104 3880 7105
rect 3560 7040 3568 7104
rect 3632 7040 3648 7104
rect 3712 7040 3728 7104
rect 3792 7040 3808 7104
rect 3872 7040 3880 7104
rect 14000 7080 34000 7112
rect 3560 7039 3880 7040
rect 14000 6624 34000 6656
rect 14000 6568 14094 6624
rect 14150 6568 34000 6624
rect 2060 6560 2380 6561
rect 2060 6496 2068 6560
rect 2132 6496 2148 6560
rect 2212 6496 2228 6560
rect 2292 6496 2308 6560
rect 2372 6496 2380 6560
rect 2060 6495 2380 6496
rect 5060 6560 5380 6561
rect 5060 6496 5068 6560
rect 5132 6496 5148 6560
rect 5212 6496 5228 6560
rect 5292 6496 5308 6560
rect 5372 6496 5380 6560
rect 14000 6536 34000 6568
rect 5060 6495 5380 6496
rect 14000 6080 34000 6112
rect 14000 6024 14094 6080
rect 14150 6024 34000 6080
rect 3560 6016 3880 6017
rect 3560 5952 3568 6016
rect 3632 5952 3648 6016
rect 3712 5952 3728 6016
rect 3792 5952 3808 6016
rect 3872 5952 3880 6016
rect 14000 5992 34000 6024
rect 3560 5951 3880 5952
rect 14000 5536 34000 5568
rect 14000 5480 14186 5536
rect 14242 5480 34000 5536
rect 2060 5472 2380 5473
rect 2060 5408 2068 5472
rect 2132 5408 2148 5472
rect 2212 5408 2228 5472
rect 2292 5408 2308 5472
rect 2372 5408 2380 5472
rect 2060 5407 2380 5408
rect 5060 5472 5380 5473
rect 5060 5408 5068 5472
rect 5132 5408 5148 5472
rect 5212 5408 5228 5472
rect 5292 5408 5308 5472
rect 5372 5408 5380 5472
rect 14000 5448 34000 5480
rect 5060 5407 5380 5408
rect 14000 4992 34000 5024
rect 14000 4936 14094 4992
rect 14150 4936 34000 4992
rect 3560 4928 3880 4929
rect 3560 4864 3568 4928
rect 3632 4864 3648 4928
rect 3712 4864 3728 4928
rect 3792 4864 3808 4928
rect 3872 4864 3880 4928
rect 14000 4904 34000 4936
rect 3560 4863 3880 4864
rect 14000 4448 34000 4480
rect 14000 4392 14186 4448
rect 14242 4392 34000 4448
rect 2060 4384 2380 4385
rect 2060 4320 2068 4384
rect 2132 4320 2148 4384
rect 2212 4320 2228 4384
rect 2292 4320 2308 4384
rect 2372 4320 2380 4384
rect 2060 4319 2380 4320
rect 5060 4384 5380 4385
rect 5060 4320 5068 4384
rect 5132 4320 5148 4384
rect 5212 4320 5228 4384
rect 5292 4320 5308 4384
rect 5372 4320 5380 4384
rect 14000 4360 34000 4392
rect 5060 4319 5380 4320
rect 14000 3904 34000 3936
rect 14000 3848 14186 3904
rect 14242 3848 34000 3904
rect 3560 3840 3880 3841
rect 3560 3776 3568 3840
rect 3632 3776 3648 3840
rect 3712 3776 3728 3840
rect 3792 3776 3808 3840
rect 3872 3776 3880 3840
rect 14000 3816 34000 3848
rect 3560 3775 3880 3776
rect 14000 3360 34000 3392
rect 14000 3304 14278 3360
rect 14334 3304 34000 3360
rect 2060 3296 2380 3297
rect 2060 3232 2068 3296
rect 2132 3232 2148 3296
rect 2212 3232 2228 3296
rect 2292 3232 2308 3296
rect 2372 3232 2380 3296
rect 2060 3231 2380 3232
rect 5060 3296 5380 3297
rect 5060 3232 5068 3296
rect 5132 3232 5148 3296
rect 5212 3232 5228 3296
rect 5292 3232 5308 3296
rect 5372 3232 5380 3296
rect 14000 3272 34000 3304
rect 5060 3231 5380 3232
rect 14000 2816 34000 2848
rect 14000 2760 14094 2816
rect 14150 2760 34000 2816
rect 3560 2752 3880 2753
rect 3560 2688 3568 2752
rect 3632 2688 3648 2752
rect 3712 2688 3728 2752
rect 3792 2688 3808 2752
rect 3872 2688 3880 2752
rect 14000 2728 34000 2760
rect 3560 2687 3880 2688
rect 14000 2272 34000 2304
rect 14000 2216 14094 2272
rect 14150 2216 34000 2272
rect 2060 2208 2380 2209
rect 2060 2144 2068 2208
rect 2132 2144 2148 2208
rect 2212 2144 2228 2208
rect 2292 2144 2308 2208
rect 2372 2144 2380 2208
rect 2060 2143 2380 2144
rect 5060 2208 5380 2209
rect 5060 2144 5068 2208
rect 5132 2144 5148 2208
rect 5212 2144 5228 2208
rect 5292 2144 5308 2208
rect 5372 2144 5380 2208
rect 14000 2184 34000 2216
rect 5060 2143 5380 2144
rect 14000 1728 34000 1760
rect 14000 1672 14186 1728
rect 14242 1672 34000 1728
rect 14000 1640 34000 1672
rect 14000 1184 34000 1216
rect 14000 1128 14278 1184
rect 14334 1128 34000 1184
rect 14000 1096 34000 1128
rect 14000 640 34000 672
rect 14000 584 14186 640
rect 14242 584 34000 640
rect 14000 552 34000 584
rect 14000 232 34000 264
rect 14000 176 14094 232
rect 14150 176 34000 232
rect 14000 144 34000 176
<< via3 >>
rect -1610 11386 -1312 11462
rect 3568 11452 3632 11456
rect 3568 11396 3572 11452
rect 3572 11396 3628 11452
rect 3628 11396 3632 11452
rect 3568 11392 3632 11396
rect 3648 11452 3712 11456
rect 3648 11396 3652 11452
rect 3652 11396 3708 11452
rect 3708 11396 3712 11452
rect 3648 11392 3712 11396
rect 3728 11452 3792 11456
rect 3728 11396 3732 11452
rect 3732 11396 3788 11452
rect 3788 11396 3792 11452
rect 3728 11392 3792 11396
rect 3808 11452 3872 11456
rect 3808 11396 3812 11452
rect 3812 11396 3868 11452
rect 3868 11396 3872 11452
rect 3808 11392 3872 11396
rect -950 10842 -652 10918
rect 2068 10908 2132 10912
rect 2068 10852 2072 10908
rect 2072 10852 2128 10908
rect 2128 10852 2132 10908
rect 2068 10848 2132 10852
rect 2148 10908 2212 10912
rect 2148 10852 2152 10908
rect 2152 10852 2208 10908
rect 2208 10852 2212 10908
rect 2148 10848 2212 10852
rect 2228 10908 2292 10912
rect 2228 10852 2232 10908
rect 2232 10852 2288 10908
rect 2288 10852 2292 10908
rect 2228 10848 2292 10852
rect 2308 10908 2372 10912
rect 2308 10852 2312 10908
rect 2312 10852 2368 10908
rect 2368 10852 2372 10908
rect 2308 10848 2372 10852
rect 5068 10908 5132 10912
rect 5068 10852 5072 10908
rect 5072 10852 5128 10908
rect 5128 10852 5132 10908
rect 5068 10848 5132 10852
rect 5148 10908 5212 10912
rect 5148 10852 5152 10908
rect 5152 10852 5208 10908
rect 5208 10852 5212 10908
rect 5148 10848 5212 10852
rect 5228 10908 5292 10912
rect 5228 10852 5232 10908
rect 5232 10852 5288 10908
rect 5288 10852 5292 10908
rect 5228 10848 5292 10852
rect 5308 10908 5372 10912
rect 5308 10852 5312 10908
rect 5312 10852 5368 10908
rect 5368 10852 5372 10908
rect 5308 10848 5372 10852
rect 3568 10364 3632 10368
rect 3568 10308 3572 10364
rect 3572 10308 3628 10364
rect 3628 10308 3632 10364
rect 3568 10304 3632 10308
rect 3648 10364 3712 10368
rect 3648 10308 3652 10364
rect 3652 10308 3708 10364
rect 3708 10308 3712 10364
rect 3648 10304 3712 10308
rect 3728 10364 3792 10368
rect 3728 10308 3732 10364
rect 3732 10308 3788 10364
rect 3788 10308 3792 10364
rect 3728 10304 3792 10308
rect 3808 10364 3872 10368
rect 3808 10308 3812 10364
rect 3812 10308 3868 10364
rect 3868 10308 3872 10364
rect 3808 10304 3872 10308
rect 2068 9820 2132 9824
rect 2068 9764 2072 9820
rect 2072 9764 2128 9820
rect 2128 9764 2132 9820
rect 2068 9760 2132 9764
rect 2148 9820 2212 9824
rect 2148 9764 2152 9820
rect 2152 9764 2208 9820
rect 2208 9764 2212 9820
rect 2148 9760 2212 9764
rect 2228 9820 2292 9824
rect 2228 9764 2232 9820
rect 2232 9764 2288 9820
rect 2288 9764 2292 9820
rect 2228 9760 2292 9764
rect 2308 9820 2372 9824
rect 2308 9764 2312 9820
rect 2312 9764 2368 9820
rect 2368 9764 2372 9820
rect 2308 9760 2372 9764
rect 5068 9820 5132 9824
rect 5068 9764 5072 9820
rect 5072 9764 5128 9820
rect 5128 9764 5132 9820
rect 5068 9760 5132 9764
rect 5148 9820 5212 9824
rect 5148 9764 5152 9820
rect 5152 9764 5208 9820
rect 5208 9764 5212 9820
rect 5148 9760 5212 9764
rect 5228 9820 5292 9824
rect 5228 9764 5232 9820
rect 5232 9764 5288 9820
rect 5288 9764 5292 9820
rect 5228 9760 5292 9764
rect 5308 9820 5372 9824
rect 5308 9764 5312 9820
rect 5312 9764 5368 9820
rect 5368 9764 5372 9820
rect 5308 9760 5372 9764
rect 3568 9276 3632 9280
rect 3568 9220 3572 9276
rect 3572 9220 3628 9276
rect 3628 9220 3632 9276
rect 3568 9216 3632 9220
rect 3648 9276 3712 9280
rect 3648 9220 3652 9276
rect 3652 9220 3708 9276
rect 3708 9220 3712 9276
rect 3648 9216 3712 9220
rect 3728 9276 3792 9280
rect 3728 9220 3732 9276
rect 3732 9220 3788 9276
rect 3788 9220 3792 9276
rect 3728 9216 3792 9220
rect 3808 9276 3872 9280
rect 3808 9220 3812 9276
rect 3812 9220 3868 9276
rect 3868 9220 3872 9276
rect 3808 9216 3872 9220
rect 2068 8732 2132 8736
rect 2068 8676 2072 8732
rect 2072 8676 2128 8732
rect 2128 8676 2132 8732
rect 2068 8672 2132 8676
rect 2148 8732 2212 8736
rect 2148 8676 2152 8732
rect 2152 8676 2208 8732
rect 2208 8676 2212 8732
rect 2148 8672 2212 8676
rect 2228 8732 2292 8736
rect 2228 8676 2232 8732
rect 2232 8676 2288 8732
rect 2288 8676 2292 8732
rect 2228 8672 2292 8676
rect 2308 8732 2372 8736
rect 2308 8676 2312 8732
rect 2312 8676 2368 8732
rect 2368 8676 2372 8732
rect 2308 8672 2372 8676
rect 5068 8732 5132 8736
rect 5068 8676 5072 8732
rect 5072 8676 5128 8732
rect 5128 8676 5132 8732
rect 5068 8672 5132 8676
rect 5148 8732 5212 8736
rect 5148 8676 5152 8732
rect 5152 8676 5208 8732
rect 5208 8676 5212 8732
rect 5148 8672 5212 8676
rect 5228 8732 5292 8736
rect 5228 8676 5232 8732
rect 5232 8676 5288 8732
rect 5288 8676 5292 8732
rect 5228 8672 5292 8676
rect 5308 8732 5372 8736
rect 5308 8676 5312 8732
rect 5312 8676 5368 8732
rect 5368 8676 5372 8732
rect 5308 8672 5372 8676
rect 3568 8188 3632 8192
rect 3568 8132 3572 8188
rect 3572 8132 3628 8188
rect 3628 8132 3632 8188
rect 3568 8128 3632 8132
rect 3648 8188 3712 8192
rect 3648 8132 3652 8188
rect 3652 8132 3708 8188
rect 3708 8132 3712 8188
rect 3648 8128 3712 8132
rect 3728 8188 3792 8192
rect 3728 8132 3732 8188
rect 3732 8132 3788 8188
rect 3788 8132 3792 8188
rect 3728 8128 3792 8132
rect 3808 8188 3872 8192
rect 3808 8132 3812 8188
rect 3812 8132 3868 8188
rect 3868 8132 3872 8188
rect 3808 8128 3872 8132
rect 2068 7644 2132 7648
rect 2068 7588 2072 7644
rect 2072 7588 2128 7644
rect 2128 7588 2132 7644
rect 2068 7584 2132 7588
rect 2148 7644 2212 7648
rect 2148 7588 2152 7644
rect 2152 7588 2208 7644
rect 2208 7588 2212 7644
rect 2148 7584 2212 7588
rect 2228 7644 2292 7648
rect 2228 7588 2232 7644
rect 2232 7588 2288 7644
rect 2288 7588 2292 7644
rect 2228 7584 2292 7588
rect 2308 7644 2372 7648
rect 2308 7588 2312 7644
rect 2312 7588 2368 7644
rect 2368 7588 2372 7644
rect 2308 7584 2372 7588
rect 5068 7644 5132 7648
rect 5068 7588 5072 7644
rect 5072 7588 5128 7644
rect 5128 7588 5132 7644
rect 5068 7584 5132 7588
rect 5148 7644 5212 7648
rect 5148 7588 5152 7644
rect 5152 7588 5208 7644
rect 5208 7588 5212 7644
rect 5148 7584 5212 7588
rect 5228 7644 5292 7648
rect 5228 7588 5232 7644
rect 5232 7588 5288 7644
rect 5288 7588 5292 7644
rect 5228 7584 5292 7588
rect 5308 7644 5372 7648
rect 5308 7588 5312 7644
rect 5312 7588 5368 7644
rect 5368 7588 5372 7644
rect 5308 7584 5372 7588
rect 3568 7100 3632 7104
rect 3568 7044 3572 7100
rect 3572 7044 3628 7100
rect 3628 7044 3632 7100
rect 3568 7040 3632 7044
rect 3648 7100 3712 7104
rect 3648 7044 3652 7100
rect 3652 7044 3708 7100
rect 3708 7044 3712 7100
rect 3648 7040 3712 7044
rect 3728 7100 3792 7104
rect 3728 7044 3732 7100
rect 3732 7044 3788 7100
rect 3788 7044 3792 7100
rect 3728 7040 3792 7044
rect 3808 7100 3872 7104
rect 3808 7044 3812 7100
rect 3812 7044 3868 7100
rect 3868 7044 3872 7100
rect 3808 7040 3872 7044
rect 2068 6556 2132 6560
rect 2068 6500 2072 6556
rect 2072 6500 2128 6556
rect 2128 6500 2132 6556
rect 2068 6496 2132 6500
rect 2148 6556 2212 6560
rect 2148 6500 2152 6556
rect 2152 6500 2208 6556
rect 2208 6500 2212 6556
rect 2148 6496 2212 6500
rect 2228 6556 2292 6560
rect 2228 6500 2232 6556
rect 2232 6500 2288 6556
rect 2288 6500 2292 6556
rect 2228 6496 2292 6500
rect 2308 6556 2372 6560
rect 2308 6500 2312 6556
rect 2312 6500 2368 6556
rect 2368 6500 2372 6556
rect 2308 6496 2372 6500
rect 5068 6556 5132 6560
rect 5068 6500 5072 6556
rect 5072 6500 5128 6556
rect 5128 6500 5132 6556
rect 5068 6496 5132 6500
rect 5148 6556 5212 6560
rect 5148 6500 5152 6556
rect 5152 6500 5208 6556
rect 5208 6500 5212 6556
rect 5148 6496 5212 6500
rect 5228 6556 5292 6560
rect 5228 6500 5232 6556
rect 5232 6500 5288 6556
rect 5288 6500 5292 6556
rect 5228 6496 5292 6500
rect 5308 6556 5372 6560
rect 5308 6500 5312 6556
rect 5312 6500 5368 6556
rect 5368 6500 5372 6556
rect 5308 6496 5372 6500
rect 3568 6012 3632 6016
rect 3568 5956 3572 6012
rect 3572 5956 3628 6012
rect 3628 5956 3632 6012
rect 3568 5952 3632 5956
rect 3648 6012 3712 6016
rect 3648 5956 3652 6012
rect 3652 5956 3708 6012
rect 3708 5956 3712 6012
rect 3648 5952 3712 5956
rect 3728 6012 3792 6016
rect 3728 5956 3732 6012
rect 3732 5956 3788 6012
rect 3788 5956 3792 6012
rect 3728 5952 3792 5956
rect 3808 6012 3872 6016
rect 3808 5956 3812 6012
rect 3812 5956 3868 6012
rect 3868 5956 3872 6012
rect 3808 5952 3872 5956
rect 2068 5468 2132 5472
rect 2068 5412 2072 5468
rect 2072 5412 2128 5468
rect 2128 5412 2132 5468
rect 2068 5408 2132 5412
rect 2148 5468 2212 5472
rect 2148 5412 2152 5468
rect 2152 5412 2208 5468
rect 2208 5412 2212 5468
rect 2148 5408 2212 5412
rect 2228 5468 2292 5472
rect 2228 5412 2232 5468
rect 2232 5412 2288 5468
rect 2288 5412 2292 5468
rect 2228 5408 2292 5412
rect 2308 5468 2372 5472
rect 2308 5412 2312 5468
rect 2312 5412 2368 5468
rect 2368 5412 2372 5468
rect 2308 5408 2372 5412
rect 5068 5468 5132 5472
rect 5068 5412 5072 5468
rect 5072 5412 5128 5468
rect 5128 5412 5132 5468
rect 5068 5408 5132 5412
rect 5148 5468 5212 5472
rect 5148 5412 5152 5468
rect 5152 5412 5208 5468
rect 5208 5412 5212 5468
rect 5148 5408 5212 5412
rect 5228 5468 5292 5472
rect 5228 5412 5232 5468
rect 5232 5412 5288 5468
rect 5288 5412 5292 5468
rect 5228 5408 5292 5412
rect 5308 5468 5372 5472
rect 5308 5412 5312 5468
rect 5312 5412 5368 5468
rect 5368 5412 5372 5468
rect 5308 5408 5372 5412
rect 3568 4924 3632 4928
rect 3568 4868 3572 4924
rect 3572 4868 3628 4924
rect 3628 4868 3632 4924
rect 3568 4864 3632 4868
rect 3648 4924 3712 4928
rect 3648 4868 3652 4924
rect 3652 4868 3708 4924
rect 3708 4868 3712 4924
rect 3648 4864 3712 4868
rect 3728 4924 3792 4928
rect 3728 4868 3732 4924
rect 3732 4868 3788 4924
rect 3788 4868 3792 4924
rect 3728 4864 3792 4868
rect 3808 4924 3872 4928
rect 3808 4868 3812 4924
rect 3812 4868 3868 4924
rect 3868 4868 3872 4924
rect 3808 4864 3872 4868
rect 2068 4380 2132 4384
rect 2068 4324 2072 4380
rect 2072 4324 2128 4380
rect 2128 4324 2132 4380
rect 2068 4320 2132 4324
rect 2148 4380 2212 4384
rect 2148 4324 2152 4380
rect 2152 4324 2208 4380
rect 2208 4324 2212 4380
rect 2148 4320 2212 4324
rect 2228 4380 2292 4384
rect 2228 4324 2232 4380
rect 2232 4324 2288 4380
rect 2288 4324 2292 4380
rect 2228 4320 2292 4324
rect 2308 4380 2372 4384
rect 2308 4324 2312 4380
rect 2312 4324 2368 4380
rect 2368 4324 2372 4380
rect 2308 4320 2372 4324
rect 5068 4380 5132 4384
rect 5068 4324 5072 4380
rect 5072 4324 5128 4380
rect 5128 4324 5132 4380
rect 5068 4320 5132 4324
rect 5148 4380 5212 4384
rect 5148 4324 5152 4380
rect 5152 4324 5208 4380
rect 5208 4324 5212 4380
rect 5148 4320 5212 4324
rect 5228 4380 5292 4384
rect 5228 4324 5232 4380
rect 5232 4324 5288 4380
rect 5288 4324 5292 4380
rect 5228 4320 5292 4324
rect 5308 4380 5372 4384
rect 5308 4324 5312 4380
rect 5312 4324 5368 4380
rect 5368 4324 5372 4380
rect 5308 4320 5372 4324
rect 3568 3836 3632 3840
rect 3568 3780 3572 3836
rect 3572 3780 3628 3836
rect 3628 3780 3632 3836
rect 3568 3776 3632 3780
rect 3648 3836 3712 3840
rect 3648 3780 3652 3836
rect 3652 3780 3708 3836
rect 3708 3780 3712 3836
rect 3648 3776 3712 3780
rect 3728 3836 3792 3840
rect 3728 3780 3732 3836
rect 3732 3780 3788 3836
rect 3788 3780 3792 3836
rect 3728 3776 3792 3780
rect 3808 3836 3872 3840
rect 3808 3780 3812 3836
rect 3812 3780 3868 3836
rect 3868 3780 3872 3836
rect 3808 3776 3872 3780
rect 2068 3292 2132 3296
rect 2068 3236 2072 3292
rect 2072 3236 2128 3292
rect 2128 3236 2132 3292
rect 2068 3232 2132 3236
rect 2148 3292 2212 3296
rect 2148 3236 2152 3292
rect 2152 3236 2208 3292
rect 2208 3236 2212 3292
rect 2148 3232 2212 3236
rect 2228 3292 2292 3296
rect 2228 3236 2232 3292
rect 2232 3236 2288 3292
rect 2288 3236 2292 3292
rect 2228 3232 2292 3236
rect 2308 3292 2372 3296
rect 2308 3236 2312 3292
rect 2312 3236 2368 3292
rect 2368 3236 2372 3292
rect 2308 3232 2372 3236
rect 5068 3292 5132 3296
rect 5068 3236 5072 3292
rect 5072 3236 5128 3292
rect 5128 3236 5132 3292
rect 5068 3232 5132 3236
rect 5148 3292 5212 3296
rect 5148 3236 5152 3292
rect 5152 3236 5208 3292
rect 5208 3236 5212 3292
rect 5148 3232 5212 3236
rect 5228 3292 5292 3296
rect 5228 3236 5232 3292
rect 5232 3236 5288 3292
rect 5288 3236 5292 3292
rect 5228 3232 5292 3236
rect 5308 3292 5372 3296
rect 5308 3236 5312 3292
rect 5312 3236 5368 3292
rect 5368 3236 5372 3292
rect 5308 3232 5372 3236
rect 3568 2748 3632 2752
rect 3568 2692 3572 2748
rect 3572 2692 3628 2748
rect 3628 2692 3632 2748
rect 3568 2688 3632 2692
rect 3648 2748 3712 2752
rect 3648 2692 3652 2748
rect 3652 2692 3708 2748
rect 3708 2692 3712 2748
rect 3648 2688 3712 2692
rect 3728 2748 3792 2752
rect 3728 2692 3732 2748
rect 3732 2692 3788 2748
rect 3788 2692 3792 2748
rect 3728 2688 3792 2692
rect 3808 2748 3872 2752
rect 3808 2692 3812 2748
rect 3812 2692 3868 2748
rect 3868 2692 3872 2748
rect 3808 2688 3872 2692
rect 2068 2204 2132 2208
rect 2068 2148 2072 2204
rect 2072 2148 2128 2204
rect 2128 2148 2132 2204
rect 2068 2144 2132 2148
rect 2148 2204 2212 2208
rect 2148 2148 2152 2204
rect 2152 2148 2208 2204
rect 2208 2148 2212 2204
rect 2148 2144 2212 2148
rect 2228 2204 2292 2208
rect 2228 2148 2232 2204
rect 2232 2148 2288 2204
rect 2288 2148 2292 2204
rect 2228 2144 2292 2148
rect 2308 2204 2372 2208
rect 2308 2148 2312 2204
rect 2312 2148 2368 2204
rect 2368 2148 2372 2204
rect 2308 2144 2372 2148
rect 5068 2204 5132 2208
rect 5068 2148 5072 2204
rect 5072 2148 5128 2204
rect 5128 2148 5132 2204
rect 5068 2144 5132 2148
rect 5148 2204 5212 2208
rect 5148 2148 5152 2204
rect 5152 2148 5208 2204
rect 5208 2148 5212 2204
rect 5148 2144 5212 2148
rect 5228 2204 5292 2208
rect 5228 2148 5232 2204
rect 5232 2148 5288 2204
rect 5288 2148 5292 2204
rect 5228 2144 5292 2148
rect 5308 2204 5372 2208
rect 5308 2148 5312 2204
rect 5312 2148 5368 2204
rect 5368 2148 5372 2204
rect 5308 2144 5372 2148
<< metal4 >>
rect -1620 13922 -1300 13964
rect -1620 13686 -1578 13922
rect -1342 13686 -1300 13922
rect -1620 11462 -1300 13686
rect -1620 11386 -1610 11462
rect -1312 11386 -1300 11462
rect -1620 9694 -1300 11386
rect -1620 9458 -1578 9694
rect -1342 9458 -1300 9694
rect -1620 6494 -1300 9458
rect -1620 6258 -1578 6494
rect -1342 6258 -1300 6494
rect -1620 -86 -1300 6258
rect -960 13262 -640 13304
rect -960 13026 -918 13262
rect -682 13026 -640 13262
rect -960 10918 -640 13026
rect 2960 13262 3280 13964
rect 2960 13026 3002 13262
rect 3238 13026 3280 13262
rect -960 10842 -950 10918
rect -652 10842 -640 10918
rect -960 8094 -640 10842
rect -960 7858 -918 8094
rect -682 7858 -640 8094
rect -960 4894 -640 7858
rect -960 4658 -918 4894
rect -682 4658 -640 4894
rect -960 574 -640 4658
rect -300 12602 20 12644
rect -300 12366 -258 12602
rect -22 12366 20 12602
rect -300 8794 20 12366
rect -300 8558 -258 8794
rect -22 8558 20 8794
rect -300 5594 20 8558
rect -300 5358 -258 5594
rect -22 5358 20 5594
rect -300 1234 20 5358
rect 360 11942 680 11984
rect 360 11706 402 11942
rect 638 11706 680 11942
rect 360 10394 680 11706
rect 360 10158 402 10394
rect 638 10158 680 10394
rect 360 7194 680 10158
rect 360 6958 402 7194
rect 638 6958 680 7194
rect 360 3994 680 6958
rect 360 3758 402 3994
rect 638 3758 680 3994
rect 360 1894 680 3758
rect 360 1658 402 1894
rect 638 1658 680 1894
rect 360 1616 680 1658
rect 2060 11942 2380 12644
rect 2060 11706 2102 11942
rect 2338 11706 2380 11942
rect 2060 10912 2380 11706
rect 2060 10848 2068 10912
rect 2132 10848 2148 10912
rect 2212 10848 2228 10912
rect 2292 10848 2308 10912
rect 2372 10848 2380 10912
rect 2060 10394 2380 10848
rect 2060 10158 2102 10394
rect 2338 10158 2380 10394
rect 2060 9824 2380 10158
rect 2060 9760 2068 9824
rect 2132 9760 2148 9824
rect 2212 9760 2228 9824
rect 2292 9760 2308 9824
rect 2372 9760 2380 9824
rect 2060 8736 2380 9760
rect 2060 8672 2068 8736
rect 2132 8672 2148 8736
rect 2212 8672 2228 8736
rect 2292 8672 2308 8736
rect 2372 8672 2380 8736
rect 2060 7648 2380 8672
rect 2060 7584 2068 7648
rect 2132 7584 2148 7648
rect 2212 7584 2228 7648
rect 2292 7584 2308 7648
rect 2372 7584 2380 7648
rect 2060 7194 2380 7584
rect 2060 6958 2102 7194
rect 2338 6958 2380 7194
rect 2060 6560 2380 6958
rect 2060 6496 2068 6560
rect 2132 6496 2148 6560
rect 2212 6496 2228 6560
rect 2292 6496 2308 6560
rect 2372 6496 2380 6560
rect 2060 5472 2380 6496
rect 2060 5408 2068 5472
rect 2132 5408 2148 5472
rect 2212 5408 2228 5472
rect 2292 5408 2308 5472
rect 2372 5408 2380 5472
rect 2060 4384 2380 5408
rect 2060 4320 2068 4384
rect 2132 4320 2148 4384
rect 2212 4320 2228 4384
rect 2292 4320 2308 4384
rect 2372 4320 2380 4384
rect 2060 3994 2380 4320
rect 2060 3758 2102 3994
rect 2338 3758 2380 3994
rect 2060 3296 2380 3758
rect 2060 3232 2068 3296
rect 2132 3232 2148 3296
rect 2212 3232 2228 3296
rect 2292 3232 2308 3296
rect 2372 3232 2380 3296
rect 2060 2208 2380 3232
rect 2060 2144 2068 2208
rect 2132 2144 2148 2208
rect 2212 2144 2228 2208
rect 2292 2144 2308 2208
rect 2372 2144 2380 2208
rect 2060 1894 2380 2144
rect 2060 1658 2102 1894
rect 2338 1658 2380 1894
rect -300 998 -258 1234
rect -22 998 20 1234
rect -300 956 20 998
rect 2060 956 2380 1658
rect 2960 8094 3280 13026
rect 4460 13922 4780 13964
rect 4460 13686 4502 13922
rect 4738 13686 4780 13922
rect 2960 7858 3002 8094
rect 3238 7858 3280 8094
rect 2960 4894 3280 7858
rect 2960 4658 3002 4894
rect 3238 4658 3280 4894
rect -960 338 -918 574
rect -682 338 -640 574
rect -960 296 -640 338
rect 2960 574 3280 4658
rect 3560 12602 3880 12644
rect 3560 12366 3602 12602
rect 3838 12366 3880 12602
rect 3560 11456 3880 12366
rect 3560 11392 3568 11456
rect 3632 11392 3648 11456
rect 3712 11392 3728 11456
rect 3792 11392 3808 11456
rect 3872 11392 3880 11456
rect 3560 10368 3880 11392
rect 3560 10304 3568 10368
rect 3632 10304 3648 10368
rect 3712 10304 3728 10368
rect 3792 10304 3808 10368
rect 3872 10304 3880 10368
rect 3560 9280 3880 10304
rect 3560 9216 3568 9280
rect 3632 9216 3648 9280
rect 3712 9216 3728 9280
rect 3792 9216 3808 9280
rect 3872 9216 3880 9280
rect 3560 8794 3880 9216
rect 3560 8558 3602 8794
rect 3838 8558 3880 8794
rect 3560 8192 3880 8558
rect 3560 8128 3568 8192
rect 3632 8128 3648 8192
rect 3712 8128 3728 8192
rect 3792 8128 3808 8192
rect 3872 8128 3880 8192
rect 3560 7104 3880 8128
rect 3560 7040 3568 7104
rect 3632 7040 3648 7104
rect 3712 7040 3728 7104
rect 3792 7040 3808 7104
rect 3872 7040 3880 7104
rect 3560 6016 3880 7040
rect 3560 5952 3568 6016
rect 3632 5952 3648 6016
rect 3712 5952 3728 6016
rect 3792 5952 3808 6016
rect 3872 5952 3880 6016
rect 3560 5594 3880 5952
rect 3560 5358 3602 5594
rect 3838 5358 3880 5594
rect 3560 4928 3880 5358
rect 3560 4864 3568 4928
rect 3632 4864 3648 4928
rect 3712 4864 3728 4928
rect 3792 4864 3808 4928
rect 3872 4864 3880 4928
rect 3560 3840 3880 4864
rect 3560 3776 3568 3840
rect 3632 3776 3648 3840
rect 3712 3776 3728 3840
rect 3792 3776 3808 3840
rect 3872 3776 3880 3840
rect 3560 2752 3880 3776
rect 3560 2688 3568 2752
rect 3632 2688 3648 2752
rect 3712 2688 3728 2752
rect 3792 2688 3808 2752
rect 3872 2688 3880 2752
rect 3560 1234 3880 2688
rect 3560 998 3602 1234
rect 3838 998 3880 1234
rect 3560 956 3880 998
rect 4460 9694 4780 13686
rect 5960 13262 6280 13964
rect 9304 13922 9624 13964
rect 9304 13686 9346 13922
rect 9582 13686 9624 13922
rect 5960 13026 6002 13262
rect 6238 13026 6280 13262
rect 4460 9458 4502 9694
rect 4738 9458 4780 9694
rect 4460 6494 4780 9458
rect 4460 6258 4502 6494
rect 4738 6258 4780 6494
rect 2960 338 3002 574
rect 3238 338 3280 574
rect -1620 -322 -1578 -86
rect -1342 -322 -1300 -86
rect -1620 -364 -1300 -322
rect 2960 -364 3280 338
rect 4460 -86 4780 6258
rect 5060 11942 5380 12644
rect 5060 11706 5102 11942
rect 5338 11706 5380 11942
rect 5060 10912 5380 11706
rect 5060 10848 5068 10912
rect 5132 10848 5148 10912
rect 5212 10848 5228 10912
rect 5292 10848 5308 10912
rect 5372 10848 5380 10912
rect 5060 10394 5380 10848
rect 5060 10158 5102 10394
rect 5338 10158 5380 10394
rect 5060 9824 5380 10158
rect 5060 9760 5068 9824
rect 5132 9760 5148 9824
rect 5212 9760 5228 9824
rect 5292 9760 5308 9824
rect 5372 9760 5380 9824
rect 5060 8736 5380 9760
rect 5060 8672 5068 8736
rect 5132 8672 5148 8736
rect 5212 8672 5228 8736
rect 5292 8672 5308 8736
rect 5372 8672 5380 8736
rect 5060 7648 5380 8672
rect 5060 7584 5068 7648
rect 5132 7584 5148 7648
rect 5212 7584 5228 7648
rect 5292 7584 5308 7648
rect 5372 7584 5380 7648
rect 5060 7194 5380 7584
rect 5060 6958 5102 7194
rect 5338 6958 5380 7194
rect 5060 6560 5380 6958
rect 5060 6496 5068 6560
rect 5132 6496 5148 6560
rect 5212 6496 5228 6560
rect 5292 6496 5308 6560
rect 5372 6496 5380 6560
rect 5060 5472 5380 6496
rect 5060 5408 5068 5472
rect 5132 5408 5148 5472
rect 5212 5408 5228 5472
rect 5292 5408 5308 5472
rect 5372 5408 5380 5472
rect 5060 4384 5380 5408
rect 5060 4320 5068 4384
rect 5132 4320 5148 4384
rect 5212 4320 5228 4384
rect 5292 4320 5308 4384
rect 5372 4320 5380 4384
rect 5060 3994 5380 4320
rect 5060 3758 5102 3994
rect 5338 3758 5380 3994
rect 5060 3296 5380 3758
rect 5060 3232 5068 3296
rect 5132 3232 5148 3296
rect 5212 3232 5228 3296
rect 5292 3232 5308 3296
rect 5372 3232 5380 3296
rect 5060 2208 5380 3232
rect 5060 2144 5068 2208
rect 5132 2144 5148 2208
rect 5212 2144 5228 2208
rect 5292 2144 5308 2208
rect 5372 2144 5380 2208
rect 5060 1894 5380 2144
rect 5060 1658 5102 1894
rect 5338 1658 5380 1894
rect 5060 956 5380 1658
rect 5960 8094 6280 13026
rect 8644 13262 8964 13304
rect 8644 13026 8686 13262
rect 8922 13026 8964 13262
rect 7984 12602 8304 12644
rect 7984 12366 8026 12602
rect 8262 12366 8304 12602
rect 5960 7858 6002 8094
rect 6238 7858 6280 8094
rect 5960 4894 6280 7858
rect 5960 4658 6002 4894
rect 6238 4658 6280 4894
rect 4460 -322 4502 -86
rect 4738 -322 4780 -86
rect 4460 -364 4780 -322
rect 5960 574 6280 4658
rect 7324 11942 7644 11984
rect 7324 11706 7366 11942
rect 7602 11706 7644 11942
rect 7324 10394 7644 11706
rect 7324 10158 7366 10394
rect 7602 10158 7644 10394
rect 7324 7194 7644 10158
rect 7324 6958 7366 7194
rect 7602 6958 7644 7194
rect 7324 3994 7644 6958
rect 7324 3758 7366 3994
rect 7602 3758 7644 3994
rect 7324 1894 7644 3758
rect 7324 1658 7366 1894
rect 7602 1658 7644 1894
rect 7324 1616 7644 1658
rect 7984 8794 8304 12366
rect 7984 8558 8026 8794
rect 8262 8558 8304 8794
rect 7984 5594 8304 8558
rect 7984 5358 8026 5594
rect 8262 5358 8304 5594
rect 7984 1234 8304 5358
rect 7984 998 8026 1234
rect 8262 998 8304 1234
rect 7984 956 8304 998
rect 8644 8094 8964 13026
rect 8644 7858 8686 8094
rect 8922 7858 8964 8094
rect 8644 4894 8964 7858
rect 8644 4658 8686 4894
rect 8922 4658 8964 4894
rect 5960 338 6002 574
rect 6238 338 6280 574
rect 5960 -364 6280 338
rect 8644 574 8964 4658
rect 8644 338 8686 574
rect 8922 338 8964 574
rect 8644 296 8964 338
rect 9304 9694 9624 13686
rect 9304 9458 9346 9694
rect 9582 9458 9624 9694
rect 9304 6494 9624 9458
rect 9304 6258 9346 6494
rect 9582 6258 9624 6494
rect 9304 -86 9624 6258
rect 9304 -322 9346 -86
rect 9582 -322 9624 -86
rect 9304 -364 9624 -322
<< via4 >>
rect -1578 13686 -1342 13922
rect -1578 9458 -1342 9694
rect -1578 6258 -1342 6494
rect -918 13026 -682 13262
rect 3002 13026 3238 13262
rect -918 7858 -682 8094
rect -918 4658 -682 4894
rect -258 12366 -22 12602
rect -258 8558 -22 8794
rect -258 5358 -22 5594
rect 402 11706 638 11942
rect 402 10158 638 10394
rect 402 6958 638 7194
rect 402 3758 638 3994
rect 402 1658 638 1894
rect 2102 11706 2338 11942
rect 2102 10158 2338 10394
rect 2102 6958 2338 7194
rect 2102 3758 2338 3994
rect 2102 1658 2338 1894
rect -258 998 -22 1234
rect 4502 13686 4738 13922
rect 3002 7858 3238 8094
rect 3002 4658 3238 4894
rect -918 338 -682 574
rect 3602 12366 3838 12602
rect 3602 8558 3838 8794
rect 3602 5358 3838 5594
rect 3602 998 3838 1234
rect 9346 13686 9582 13922
rect 6002 13026 6238 13262
rect 4502 9458 4738 9694
rect 4502 6258 4738 6494
rect 3002 338 3238 574
rect -1578 -322 -1342 -86
rect 5102 11706 5338 11942
rect 5102 10158 5338 10394
rect 5102 6958 5338 7194
rect 5102 3758 5338 3994
rect 5102 1658 5338 1894
rect 8686 13026 8922 13262
rect 8026 12366 8262 12602
rect 6002 7858 6238 8094
rect 6002 4658 6238 4894
rect 4502 -322 4738 -86
rect 7366 11706 7602 11942
rect 7366 10158 7602 10394
rect 7366 6958 7602 7194
rect 7366 3758 7602 3994
rect 7366 1658 7602 1894
rect 8026 8558 8262 8794
rect 8026 5358 8262 5594
rect 8026 998 8262 1234
rect 8686 7858 8922 8094
rect 8686 4658 8922 4894
rect 6002 338 6238 574
rect 8686 338 8922 574
rect 9346 9458 9582 9694
rect 9346 6258 9582 6494
rect 9346 -322 9582 -86
<< metal5 >>
rect -1620 13922 9624 13964
rect -1620 13686 -1578 13922
rect -1342 13686 4502 13922
rect 4738 13686 9346 13922
rect 9582 13686 9624 13922
rect -1620 13644 9624 13686
rect -960 13262 8964 13304
rect -960 13026 -918 13262
rect -682 13026 3002 13262
rect 3238 13026 6002 13262
rect 6238 13026 8686 13262
rect 8922 13026 8964 13262
rect -960 12984 8964 13026
rect -300 12602 8304 12644
rect -300 12366 -258 12602
rect -22 12366 3602 12602
rect 3838 12366 8026 12602
rect 8262 12366 8304 12602
rect -300 12324 8304 12366
rect 360 11942 7644 11984
rect 360 11706 402 11942
rect 638 11706 2102 11942
rect 2338 11706 5102 11942
rect 5338 11706 7366 11942
rect 7602 11706 7644 11942
rect 360 11664 7644 11706
rect -300 10394 8304 10436
rect -300 10158 402 10394
rect 638 10158 2102 10394
rect 2338 10158 5102 10394
rect 5338 10158 7366 10394
rect 7602 10158 8304 10394
rect -300 10116 8304 10158
rect -1620 9694 9624 9736
rect -1620 9458 -1578 9694
rect -1342 9458 4502 9694
rect 4738 9458 9346 9694
rect 9582 9458 9624 9694
rect -1620 9416 9624 9458
rect -300 8794 8304 8836
rect -300 8558 -258 8794
rect -22 8558 3602 8794
rect 3838 8558 8026 8794
rect 8262 8558 8304 8794
rect -300 8516 8304 8558
rect -1620 8094 9624 8136
rect -1620 7858 -918 8094
rect -682 7858 3002 8094
rect 3238 7858 6002 8094
rect 6238 7858 8686 8094
rect 8922 7858 9624 8094
rect -1620 7816 9624 7858
rect -300 7194 8304 7236
rect -300 6958 402 7194
rect 638 6958 2102 7194
rect 2338 6958 5102 7194
rect 5338 6958 7366 7194
rect 7602 6958 8304 7194
rect -300 6916 8304 6958
rect -1620 6494 9624 6536
rect -1620 6258 -1578 6494
rect -1342 6258 4502 6494
rect 4738 6258 9346 6494
rect 9582 6258 9624 6494
rect -1620 6216 9624 6258
rect -300 5594 8304 5636
rect -300 5358 -258 5594
rect -22 5358 3602 5594
rect 3838 5358 8026 5594
rect 8262 5358 8304 5594
rect -300 5316 8304 5358
rect -1620 4894 9624 4936
rect -1620 4658 -918 4894
rect -682 4658 3002 4894
rect 3238 4658 6002 4894
rect 6238 4658 8686 4894
rect 8922 4658 9624 4894
rect -1620 4616 9624 4658
rect -300 3994 8304 4036
rect -300 3758 402 3994
rect 638 3758 2102 3994
rect 2338 3758 5102 3994
rect 5338 3758 7366 3994
rect 7602 3758 8304 3994
rect -300 3716 8304 3758
rect 360 1894 7644 1936
rect 360 1658 402 1894
rect 638 1658 2102 1894
rect 2338 1658 5102 1894
rect 5338 1658 7366 1894
rect 7602 1658 7644 1894
rect 360 1616 7644 1658
rect -300 1234 8304 1276
rect -300 998 -258 1234
rect -22 998 3602 1234
rect 3838 998 8026 1234
rect 8262 998 8304 1234
rect -300 956 8304 998
rect -960 574 8964 616
rect -960 338 -918 574
rect -682 338 3002 574
rect 3238 338 6002 574
rect 6238 338 8686 574
rect 8922 338 8964 574
rect -960 296 8964 338
rect -1620 -86 9624 -44
rect -1620 -322 -1578 -86
rect -1342 -322 4502 -86
rect 4738 -322 9346 -86
rect 9582 -322 9624 -86
rect -1620 -364 9624 -322
use sky130_fd_sc_hd__dfrtp_4  _098_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 1656 0 1 2720
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 920 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1611581575
transform 1 0 920 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 1196 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 2300 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 3036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 1196 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 1564 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _057_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 3864 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1611581575
transform 1 0 3220 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_36
timestamp 1611581575
transform 1 0 3772 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1611581575
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 3864 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_36
timestamp 1611581575
transform 1 0 4232 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38
timestamp 1611581575
transform 1 0 4416 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _093_
timestamp 1611581575
transform 1 0 4508 0 -1 2720
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_4  _094_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 4416 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1611581575
transform -1 0 7084 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1611581575
transform -1 0 7084 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_35
timestamp 1611581575
transform 1 0 6624 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63
timestamp 1611581575
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_62
timestamp 1611581575
transform 1 0 6624 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _096_
timestamp 1611581575
transform 1 0 2576 0 -1 3808
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1611581575
transform 1 0 920 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1611581575
transform 1 0 1196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_15
timestamp 1611581575
transform 1 0 2300 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1611581575
transform 1 0 5152 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1611581575
transform 1 0 4784 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_41
timestamp 1611581575
transform 1 0 4692 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _078_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 5888 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1611581575
transform -1 0 7084 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_37
timestamp 1611581575
transform 1 0 6532 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 5704 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_50
timestamp 1611581575
transform 1 0 5520 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_62
timestamp 1611581575
transform 1 0 6624 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _106_
timestamp 1611581575
transform 1 0 1196 0 1 3808
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1611581575
transform 1 0 920 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1611581575
transform 1 0 3312 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _109_
timestamp 1611581575
transform 1 0 3864 0 1 3808
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_38
timestamp 1611581575
transform 1 0 3772 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_30
timestamp 1611581575
transform 1 0 3680 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _077_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 5980 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1611581575
transform -1 0 7084 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _046_
timestamp 1611581575
transform 1 0 2116 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _047_
timestamp 1611581575
transform 1 0 1748 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _049_
timestamp 1611581575
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _097_
timestamp 1611581575
transform 1 0 2484 0 -1 4896
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1611581575
transform 1 0 920 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1611581575
transform 1 0 1196 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _076_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 5428 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1611581575
transform 1 0 5060 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 4784 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_40
timestamp 1611581575
transform 1 0 4600 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _079_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 5704 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1611581575
transform -1 0 7084 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_39
timestamp 1611581575
transform 1 0 6532 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_62
timestamp 1611581575
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _105_
timestamp 1611581575
transform 1 0 1196 0 1 4896
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1611581575
transform 1 0 920 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _043_
timestamp 1611581575
transform 1 0 3312 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _044_
timestamp 1611581575
transform 1 0 3956 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_4  _095_
timestamp 1611581575
transform 1 0 4600 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_40
timestamp 1611581575
transform 1 0 3772 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_30
timestamp 1611581575
transform 1 0 3680 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_32
timestamp 1611581575
transform 1 0 3864 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_37
timestamp 1611581575
transform 1 0 4324 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1611581575
transform -1 0 7084 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _104_
timestamp 1611581575
transform 1 0 1196 0 1 5984
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _107_
timestamp 1611581575
transform 1 0 1380 0 -1 5984
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1611581575
transform 1 0 920 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1611581575
transform 1 0 920 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1611581575
transform 1 0 1196 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _045_
timestamp 1611581575
transform 1 0 3864 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _050_
timestamp 1611581575
transform 1 0 3312 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _091_
timestamp 1611581575
transform 1 0 4324 0 1 5984
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _108_
timestamp 1611581575
transform 1 0 3496 0 -1 5984
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_42
timestamp 1611581575
transform 1 0 3772 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_30
timestamp 1611581575
transform 1 0 3680 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_36
timestamp 1611581575
transform 1 0 4232 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1611581575
transform 1 0 5612 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1611581575
transform 1 0 5980 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1611581575
transform 1 0 6440 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1611581575
transform -1 0 7084 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1611581575
transform -1 0 7084 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_41
timestamp 1611581575
transform 1 0 6532 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_59
timestamp 1611581575
transform 1 0 6348 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_62
timestamp 1611581575
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _110_
timestamp 1611581575
transform 1 0 3036 0 -1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1611581575
transform 1 0 920 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 1196 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  _053_
timestamp 1611581575
transform 1 0 5152 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_2  _085_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 5704 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1611581575
transform -1 0 7084 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_43
timestamp 1611581575
transform 1 0 6532 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_50
timestamp 1611581575
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_62
timestamp 1611581575
transform 1 0 6624 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _103_
timestamp 1611581575
transform 1 0 1288 0 1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1611581575
transform 1 0 920 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1611581575
transform 1 0 1196 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _051_
timestamp 1611581575
transform 1 0 3404 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _090_
timestamp 1611581575
transform 1 0 3864 0 1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_44
timestamp 1611581575
transform 1 0 3772 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _073_
timestamp 1611581575
transform 1 0 5980 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1611581575
transform -1 0 7084 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_62
timestamp 1611581575
transform 1 0 6624 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _102_
timestamp 1611581575
transform 1 0 1196 0 -1 8160
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1611581575
transform 1 0 920 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _048_
timestamp 1611581575
transform 1 0 3312 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_4  _092_
timestamp 1611581575
transform 1 0 3956 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 3680 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1611581575
transform 1 0 6164 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1611581575
transform -1 0 7084 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_45
timestamp 1611581575
transform 1 0 6532 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_62
timestamp 1611581575
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _101_
timestamp 1611581575
transform 1 0 1196 0 1 8160
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1611581575
transform 1 0 920 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _052_
timestamp 1611581575
transform 1 0 3312 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1611581575
transform 1 0 3956 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _111_
timestamp 1611581575
transform 1 0 4324 0 1 8160
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46
timestamp 1611581575
transform 1 0 3772 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_30
timestamp 1611581575
transform 1 0 3680 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_32
timestamp 1611581575
transform 1 0 3864 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1611581575
transform 1 0 6440 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1611581575
transform -1 0 7084 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_4  _080_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 1380 0 -1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_4  _087_
timestamp 1611581575
transform 1 0 2944 0 -1 9248
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1611581575
transform 1 0 920 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1611581575
transform 1 0 1196 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _042_
timestamp 1611581575
transform 1 0 5060 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1611581575
transform 1 0 5428 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1611581575
transform 1 0 5796 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _072_
timestamp 1611581575
transform 1 0 6256 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1611581575
transform -1 0 7084 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1611581575
transform 1 0 6532 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_57
timestamp 1611581575
transform 1 0 6164 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_62
timestamp 1611581575
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _054_
timestamp 1611581575
transform 1 0 1840 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_4  _075_
timestamp 1611581575
transform 1 0 2208 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_4  _100_
timestamp 1611581575
transform 1 0 1196 0 -1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1611581575
transform 1 0 920 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1611581575
transform 1 0 920 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1611581575
transform 1 0 1196 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_9
timestamp 1611581575
transform 1 0 1748 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_4  _086_
timestamp 1611581575
transform 1 0 3312 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrtp_4  _088_
timestamp 1611581575
transform 1 0 3864 0 1 9248
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1611581575
transform 1 0 3772 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _041_
timestamp 1611581575
transform 1 0 5520 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1611581575
transform 1 0 5980 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_57
timestamp 1611581575
transform 1 0 6164 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _074_
timestamp 1611581575
transform 1 0 6348 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _081_
timestamp 1611581575
transform 1 0 6256 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1611581575
transform -1 0 7084 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1611581575
transform -1 0 7084 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1611581575
transform 1 0 6532 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1611581575
transform 1 0 6624 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_62
timestamp 1611581575
transform 1 0 6624 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _099_
timestamp 1611581575
transform 1 0 1656 0 1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1611581575
transform 1 0 920 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1611581575
transform 1 0 1472 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1611581575
transform 1 0 1196 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1611581575
transform 1 0 4048 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _089_
timestamp 1611581575
transform 1 0 4416 0 1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1611581575
transform 1 0 3772 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_32
timestamp 1611581575
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _082_
timestamp 1611581575
transform 1 0 6532 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1611581575
transform -1 0 7084 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1611581575
transform 1 0 1196 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _055_
timestamp 1611581575
transform 1 0 2760 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1611581575
transform 1 0 3128 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_6
timestamp 1611581575
transform 1 0 1472 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_18
timestamp 1611581575
transform 1 0 2576 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _083_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 4324 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_8  gpio_in_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611581575
transform 1 0 4968 0 -1 11424
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1611581575
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_serial_clock
timestamp 1611581575
transform 1 0 3496 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_32
timestamp 1611581575
transform 1 0 3864 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_36
timestamp 1611581575
transform 1 0 4232 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1611581575
transform -1 0 7084 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1611581575
transform 1 0 6624 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_63
timestamp 1611581575
transform 1 0 6716 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1611581575
transform -1 0 460 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  gpio_logic_high
timestamp 1611581575
transform 1 0 92 0 -1 11424
box -38 -48 314 592
<< labels >>
rlabel metal3 s 14000 1096 34000 1216 6 mgmt_gpio_in
port 0 nsew signal tristate
rlabel metal3 s 14000 1640 34000 1760 6 mgmt_gpio_oeb
port 1 nsew signal input
rlabel metal3 s 14000 2184 34000 2304 6 mgmt_gpio_out
port 2 nsew signal input
rlabel metal3 s 14000 552 34000 672 6 one
port 3 nsew signal tristate
rlabel metal3 s 14000 2728 34000 2848 6 pad_gpio_ana_en
port 4 nsew signal tristate
rlabel metal3 s 14000 3272 34000 3392 6 pad_gpio_ana_pol
port 5 nsew signal tristate
rlabel metal3 s 14000 3816 34000 3936 6 pad_gpio_ana_sel
port 6 nsew signal tristate
rlabel metal3 s 14000 4360 34000 4480 6 pad_gpio_dm[0]
port 7 nsew signal tristate
rlabel metal3 s 14000 4904 34000 5024 6 pad_gpio_dm[1]
port 8 nsew signal tristate
rlabel metal3 s 14000 5448 34000 5568 6 pad_gpio_dm[2]
port 9 nsew signal tristate
rlabel metal3 s 14000 5992 34000 6112 6 pad_gpio_holdover
port 10 nsew signal tristate
rlabel metal3 s 14000 6536 34000 6656 6 pad_gpio_ib_mode_sel
port 11 nsew signal tristate
rlabel metal3 s 14000 7080 34000 7200 6 pad_gpio_in
port 12 nsew signal input
rlabel metal3 s 14000 7624 34000 7744 6 pad_gpio_inenb
port 13 nsew signal tristate
rlabel metal3 s 14000 8168 34000 8288 6 pad_gpio_out
port 14 nsew signal tristate
rlabel metal3 s 14000 8712 34000 8832 6 pad_gpio_outenb
port 15 nsew signal tristate
rlabel metal3 s 14000 9256 34000 9376 6 pad_gpio_slow_sel
port 16 nsew signal tristate
rlabel metal3 s 14000 9800 34000 9920 6 pad_gpio_vtrip_sel
port 17 nsew signal tristate
rlabel metal3 s 14000 10344 34000 10464 6 resetn
port 18 nsew signal input
rlabel metal3 s 14000 10888 34000 11008 6 serial_clock
port 19 nsew signal input
rlabel metal3 s 14000 11432 34000 11552 6 serial_data_in
port 20 nsew signal input
rlabel metal3 s 14000 11976 34000 12096 6 serial_data_out
port 21 nsew signal tristate
rlabel metal3 s 14000 12520 34000 12640 6 user_gpio_in
port 22 nsew signal tristate
rlabel metal3 s 14000 13064 34000 13184 6 user_gpio_oeb
port 23 nsew signal input
rlabel metal3 s 14000 13608 34000 13728 6 user_gpio_out
port 24 nsew signal input
rlabel metal3 s 14000 144 34000 264 6 zero
port 25 nsew signal tristate
rlabel metal4 s 5060 956 5380 12644 6 vccd
port 26 nsew power bidirectional
rlabel metal4 s 2060 956 2380 12644 6 vccd
port 27 nsew power bidirectional
rlabel metal4 s 7324 1616 7644 11984 6 vccd
port 28 nsew power bidirectional
rlabel metal4 s 360 1616 680 11984 6 vccd
port 29 nsew power bidirectional
rlabel metal5 s 360 11664 7644 11984 6 vccd
port 30 nsew power bidirectional
rlabel metal5 s -300 10116 8304 10436 6 vccd
port 31 nsew power bidirectional
rlabel metal5 s -300 6916 8304 7236 6 vccd
port 32 nsew power bidirectional
rlabel metal5 s -300 3716 8304 4036 6 vccd
port 33 nsew power bidirectional
rlabel metal5 s 360 1616 7644 1936 6 vccd
port 34 nsew power bidirectional
rlabel metal4 s 7984 956 8304 12644 6 vssd
port 35 nsew ground bidirectional
rlabel metal4 s 3560 956 3880 12644 6 vssd
port 36 nsew ground bidirectional
rlabel metal4 s -300 956 20 12644 4 vssd
port 37 nsew ground bidirectional
rlabel metal5 s -300 12324 8304 12644 6 vssd
port 38 nsew ground bidirectional
rlabel metal5 s -300 8516 8304 8836 6 vssd
port 39 nsew ground bidirectional
rlabel metal5 s -300 5316 8304 5636 6 vssd
port 40 nsew ground bidirectional
rlabel metal5 s -300 956 8304 1276 6 vssd
port 41 nsew ground bidirectional
rlabel metal4 s 5960 -364 6280 13964 6 vccd1
port 42 nsew power bidirectional
rlabel metal4 s 2960 -364 3280 13964 6 vccd1
port 43 nsew power bidirectional
rlabel metal4 s 8644 296 8964 13304 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s -960 296 -640 13304 4 vccd1
port 45 nsew power bidirectional
rlabel metal5 s -960 12984 8964 13304 6 vccd1
port 46 nsew power bidirectional
rlabel metal5 s -1620 7816 9624 8136 6 vccd1
port 47 nsew power bidirectional
rlabel metal5 s -1620 4616 9624 4936 6 vccd1
port 48 nsew power bidirectional
rlabel metal5 s -960 296 8964 616 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 9304 -364 9624 13964 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 4460 -364 4780 13964 6 vssd1
port 51 nsew ground bidirectional
rlabel metal4 s -1620 -364 -1300 13964 4 vssd1
port 52 nsew ground bidirectional
rlabel metal5 s -1620 13644 9624 13964 6 vssd1
port 53 nsew ground bidirectional
rlabel metal5 s -1620 9416 9624 9736 6 vssd1
port 54 nsew ground bidirectional
rlabel metal5 s -1620 6216 9624 6536 6 vssd1
port 55 nsew ground bidirectional
rlabel metal5 s -1620 -364 9624 -44 8 vssd1
port 56 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 34000 14000
<< end >>
