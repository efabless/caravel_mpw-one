* SPICE NETLIST
***************************************

.SUBCKT MN g s d b
.ENDS
***************************************
.SUBCKT MP g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT condiodeHvPsub pin0 pin1
.ENDS
***************************************
.SUBCKT nvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20nativevhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT n20nativevhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT pvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT p20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcnwvc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcnwvc2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xchvnwc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT xcmvpp pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_nhvnative10x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_phv5x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap2_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l40 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l20 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l10 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvppx4_2xnhvnative10x4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym50p4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_lim4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp3 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT ind4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_55959141808692 2 3
** N=7 EP=2 IP=0 FDC=1
R0 3 2 L=900 W=0.33 m=1 mult=1 model="mrp1" $[mrp1] $X=-250 $Y=-3240 $D=257
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd2__example_55959141808666
** N=23 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808687 2 3 4
** N=55 EP=3 IP=33 FDC=10
*.SEEDPROM
M0 4 3 2 2 pshort L=0.18 W=7 AD=0.98 AS=1.96 PD=7.28 PS=14.56 NRD=0 NRS=0 m=1 r=38.8889 sa=90000.2 sb=90004.3 a=1.26 p=14.36 mult=1 $X=0 $Y=0 $D=79
M1 2 3 4 2 pshort L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=38.8889 sa=90000.7 sb=90003.9 a=1.26 p=14.36 mult=1 $X=460 $Y=0 $D=79
M2 4 3 2 2 pshort L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=38.8889 sa=90001.1 sb=90003.4 a=1.26 p=14.36 mult=1 $X=920 $Y=0 $D=79
M3 2 3 4 2 pshort L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=38.8889 sa=90001.6 sb=90002.9 a=1.26 p=14.36 mult=1 $X=1380 $Y=0 $D=79
M4 4 3 2 2 pshort L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=38.8889 sa=90002 sb=90002.5 a=1.26 p=14.36 mult=1 $X=1840 $Y=0 $D=79
M5 2 3 4 2 pshort L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=38.8889 sa=90002.5 sb=90002 a=1.26 p=14.36 mult=1 $X=2300 $Y=0 $D=79
M6 4 3 2 2 pshort L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=38.8889 sa=90002.9 sb=90001.6 a=1.26 p=14.36 mult=1 $X=2760 $Y=0 $D=79
M7 2 3 4 2 pshort L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=38.8889 sa=90003.4 sb=90001.1 a=1.26 p=14.36 mult=1 $X=3220 $Y=0 $D=79
M8 4 3 2 2 pshort L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=38.8889 sa=90003.9 sb=90000.7 a=1.26 p=14.36 mult=1 $X=3680 $Y=0 $D=79
M9 2 3 4 2 pshort L=0.18 W=7 AD=1.96 AS=0.98 PD=14.56 PS=7.28 NRD=0 NRS=0 m=1 r=38.8889 sa=90004.3 sb=90000.2 a=1.26 p=14.36 mult=1 $X=4140 $Y=0 $D=79
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1__example_55959141808682
** N=24 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_4
** N=4 EP=0 IP=8 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1__example_55959141808681
** N=18 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_5
** N=4 EP=0 IP=8 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_55959141808691 2 3
** N=7 EP=2 IP=0 FDC=1
R0 3 2 L=200 W=0.33 m=1 mult=1 model="mrp1" $[mrp1] $X=-250 $Y=-9720 $D=257
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd__example_55959141808700
** N=21 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd2__example_55959141808559
** N=21 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808699
** N=68 EP=0 IP=46 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dftpl1s2__example_55959141808702
** N=63 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808704 2
** N=25 EP=1 IP=33 FDC=2
*.SEEDPROM
X0 2 2 Dpar a=2.1 p=14.6 m=1 $[ndiode] $X=-1825 $Y=0 $D=181
X1 2 2 Dpar a=2.1 p=14.6 m=1 $[ndiode] $X=40675 $Y=0 $D=181
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dftpl1s2__example_55959141808694
** N=45 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808695 2
** N=25 EP=1 IP=33 FDC=2
*.SEEDPROM
X0 2 2 Dpar a=1.5 p=10.6 m=1 $[ndiode] $X=-1825 $Y=0 $D=181
X1 2 2 Dpar a=1.5 p=10.6 m=1 $[ndiode] $X=40675 $Y=0 $D=181
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd2__example_55959141808679
** N=24 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808696
** N=46 EP=0 IP=48 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd__example_5595914180851
** N=17 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd2__example_55959141808378
** N=18 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808698
** N=61 EP=0 IP=54 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__tpl1__example_55959141808685
** N=48 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__tpl1__example_55959141808686
** N=57 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_io__gnd2gnd_tap
** N=174 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_io__gnd2gnd_diff
** N=174 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_io__gnd2gnd_sub_dnwl 1 2
** N=3 EP=2 IP=22 FDC=1
X0 1 2 Dpar a=283.052 p=67.56 m=1 $[nwdiode] $X=900 $Y=900 $D=191
.ENDS
***************************************
.SUBCKT sky130_fd_io__gnd2gnd_120x2_lv_isosub VSUB VSSI VSS_N
** N=3 EP=3 IP=6 FDC=10
D0 VSS_N VSSI pdiode AREA=22.5 PJ=33 m=1 ahftempperim=33 $X=3160 $Y=1100 $D=172
D1 VSS_N VSSI pdiode AREA=22.5 PJ=33 m=1 ahftempperim=33 $X=7280 $Y=1100 $D=172
D2 VSS_N VSSI pdiode AREA=22.5 PJ=33 m=1 ahftempperim=33 $X=11400 $Y=1100 $D=172
D3 VSS_N VSSI pdiode AREA=22.5 PJ=33 m=1 ahftempperim=33 $X=15520 $Y=1100 $D=172
D4 VSSI VSS_N pdiode AREA=22.5 PJ=33 m=1 ahftempperim=33 $X=23150 $Y=1100 $D=172
D5 VSSI VSS_N pdiode AREA=22.5 PJ=33 m=1 ahftempperim=33 $X=27270 $Y=1100 $D=172
D6 VSSI VSS_N pdiode AREA=22.5 PJ=33 m=1 ahftempperim=33 $X=31390 $Y=1100 $D=172
D7 VSSI VSS_N pdiode AREA=22.5 PJ=33 m=1 ahftempperim=33 $X=35510 $Y=1100 $D=172
X8 VSUB VSSI sky130_fd_io__gnd2gnd_sub_dnwl $T=0 0 0 0 $X=0 $Y=0
X9 VSUB VSS_N sky130_fd_io__gnd2gnd_sub_dnwl $T=40170 0 1 180 $X=19990 $Y=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808701 2
** N=41 EP=1 IP=57 FDC=2
*.SEEDPROM
X0 2 2 Dpar a=2.1 p=14.6 m=1 $[ndiode] $X=-1200 $Y=0 $D=181
X1 2 2 Dpar a=2.1 p=14.6 m=1 $[ndiode] $X=49360 $Y=0 $D=181
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808703 2
** N=29 EP=1 IP=39 FDC=2
*.SEEDPROM
X0 2 2 Dpar a=2.1 p=14.6 m=1 $[ndiode] $X=-1825 $Y=0 $D=181
X1 2 2 Dpar a=2.1 p=14.6 m=1 $[ndiode] $X=49035 $Y=0 $D=181
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808705 2
** N=43 EP=1 IP=60 FDC=2
*.SEEDPROM
X0 2 2 Dpar a=2.1 p=14.6 m=1 $[ndiode] $X=-1200 $Y=0 $D=181
X1 2 2 Dpar a=2.1 p=14.6 m=1 $[ndiode] $X=52130 $Y=0 $D=181
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808693 2
** N=43 EP=1 IP=60 FDC=2
*.SEEDPROM
X0 2 2 Dpar a=1.5 p=10.6 m=1 $[ndiode] $X=-1200 $Y=0 $D=181
X1 2 2 Dpar a=1.5 p=10.6 m=1 $[ndiode] $X=52130 $Y=0 $D=181
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808697
** N=37 EP=0 IP=34 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_55959141808688 3 4
** N=8 EP=2 IP=0 FDC=1
*.SEEDPROM
R0 3 4 L=720 W=0.33 m=1 mult=1 model="mrp1" $[mrp1] $X=-250 $Y=-8100 $D=257
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_55959141808690 2 3
** N=6 EP=2 IP=0 FDC=1
R0 3 2 L=300 W=0.33 m=1 mult=1 model="mrp1" $[mrp1] $X=-250 $Y=-3240 $D=257
.ENDS
***************************************
.SUBCKT sky130_fd_io__top_power_lvc_wpad VSSD SRC_BDY_LVC2 SRC_BDY_LVC1 DRN_LVC1 VDDIO DRN_LVC2 BDY2_B2B P_CORE P_PAD
** N=12422 EP=9 IP=1228 FDC=501
*.CALIBRE ISOLATED NETS: OGC_LVC VCCHIB VCCD VDDA VSSIO VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
M0 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90001.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=14360 $Y=26860 $D=9
M1 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90001.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=14360 $Y=36860 $D=9
M2 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90001.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=14360 $Y=46860 $D=9
M3 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90001.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=14360 $Y=56860 $D=9
M4 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90001.1 sb=90019.9 a=0.9 p=10.36 mult=1 $X=14360 $Y=66860 $D=9
M5 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90001.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=14360 $Y=186860 $D=9
M6 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90002.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=15550 $Y=26860 $D=9
M7 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90002.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=15550 $Y=36860 $D=9
M8 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90002.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=15550 $Y=46860 $D=9
M9 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90002.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=15550 $Y=56860 $D=9
M10 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90002.3 sb=90019.9 a=0.9 p=10.36 mult=1 $X=15550 $Y=66860 $D=9
M11 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90002.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=15550 $Y=186860 $D=9
M12 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=4 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 r=1.25 sa=2e+06 sb=2.00002e+06 a=20 p=18 mult=1 $X=12975 $Y=75805 $D=9
M13 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90003.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=17130 $Y=26860 $D=9
M14 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90003.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=17130 $Y=36860 $D=9
M15 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90003.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=17130 $Y=46860 $D=9
M16 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90003.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=17130 $Y=56860 $D=9
M17 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90003.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=17130 $Y=66860 $D=9
M18 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90001.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=17130 $Y=176860 $D=9
M19 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90003.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=17130 $Y=186860 $D=9
M20 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90001.7 sb=90019.9 a=1.26 p=14.36 mult=1 $X=17455 $Y=146860 $D=9
M21 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90001.7 sb=90019.9 a=1.26 p=14.36 mult=1 $X=17455 $Y=156860 $D=9
M22 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90001.7 sb=90019.9 a=1.26 p=14.36 mult=1 $X=17455 $Y=166860 $D=9
M23 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90005.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=18320 $Y=26860 $D=9
M24 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90005.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=18320 $Y=36860 $D=9
M25 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90005.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=18320 $Y=46860 $D=9
M26 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90005.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=18320 $Y=56860 $D=9
M27 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90005.1 sb=90019.9 a=0.9 p=10.36 mult=1 $X=18320 $Y=66860 $D=9
M28 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90002.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=18320 $Y=176860 $D=9
M29 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90005.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=18320 $Y=186860 $D=9
M30 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90003.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=18805 $Y=146860 $D=9
M31 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90003.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=18805 $Y=156860 $D=9
M32 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90003.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=18805 $Y=166860 $D=9
M33 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90006.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=19900 $Y=26860 $D=9
M34 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90006.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=19900 $Y=36860 $D=9
M35 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90006.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=19900 $Y=46860 $D=9
M36 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90006.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=19900 $Y=56860 $D=9
M37 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90006.6 sb=90019.9 a=0.9 p=10.36 mult=1 $X=19900 $Y=66860 $D=9
M38 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90003.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=19900 $Y=176860 $D=9
M39 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90006.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=19900 $Y=186860 $D=9
M40 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90007.8 sb=90019.9 a=1.26 p=14.36 mult=1 $X=21090 $Y=26860 $D=9
M41 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90007.8 sb=90019.9 a=1.26 p=14.36 mult=1 $X=21090 $Y=36860 $D=9
M42 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90007.8 sb=90019.9 a=1.26 p=14.36 mult=1 $X=21090 $Y=46860 $D=9
M43 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90007.8 sb=90019.9 a=1.26 p=14.36 mult=1 $X=21090 $Y=56860 $D=9
M44 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90007.8 sb=90019.9 a=0.9 p=10.36 mult=1 $X=21090 $Y=66860 $D=9
M45 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90005.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=21090 $Y=176860 $D=9
M46 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90007.8 sb=90019.9 a=1.26 p=14.36 mult=1 $X=21090 $Y=186860 $D=9
M47 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90005.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=21635 $Y=146860 $D=9
M48 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90005.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=21635 $Y=156860 $D=9
M49 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90005.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=21635 $Y=166860 $D=9
M50 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90009.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=22670 $Y=26860 $D=9
M51 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90009.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=22670 $Y=36860 $D=9
M52 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90009.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=22670 $Y=46860 $D=9
M53 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90009.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=22670 $Y=56860 $D=9
M54 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90009.4 sb=90019.9 a=0.9 p=10.36 mult=1 $X=22670 $Y=66860 $D=9
M55 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90006.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=22670 $Y=176860 $D=9
M56 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90009.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=22670 $Y=186860 $D=9
M57 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90007.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=22985 $Y=146860 $D=9
M58 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90007.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=22985 $Y=156860 $D=9
M59 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90007.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=22985 $Y=166860 $D=9
M60 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90010.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=23860 $Y=26860 $D=9
M61 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90010.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=23860 $Y=36860 $D=9
M62 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90010.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=23860 $Y=46860 $D=9
M63 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90010.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=23860 $Y=56860 $D=9
M64 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90010.6 sb=90019.9 a=0.9 p=10.36 mult=1 $X=23860 $Y=66860 $D=9
M65 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90007.8 sb=90019.9 a=1.26 p=14.36 mult=1 $X=23860 $Y=176860 $D=9
M66 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90010.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=23860 $Y=186860 $D=9
M67 SRC_BDY_LVC2 23 25 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 r=38.8889 sa=90000.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=24670 $Y=82805 $D=9
M68 SRC_BDY_LVC2 23 25 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 r=38.8889 sa=90000.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=24670 $Y=91300 $D=9
M69 SRC_BDY_LVC1 21 24 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 r=38.8889 sa=90000.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=24670 $Y=101405 $D=9
M70 SRC_BDY_LVC1 21 24 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 r=38.8889 sa=90000.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=24670 $Y=109900 $D=9
M71 SRC_BDY_LVC1 21 24 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 r=38.8889 sa=90000.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=24670 $Y=118725 $D=9
M72 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=0.625 sa=4e+06 sb=4.00002e+06 a=40 p=26 mult=1 $X=17255 $Y=75805 $D=9
M73 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90012.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=25440 $Y=26860 $D=9
M74 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90012.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=25440 $Y=36860 $D=9
M75 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90012.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=25440 $Y=46860 $D=9
M76 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90012.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=25440 $Y=56860 $D=9
M77 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90012.2 sb=90019.9 a=0.9 p=10.36 mult=1 $X=25440 $Y=66860 $D=9
M78 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90009.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=25440 $Y=176860 $D=9
M79 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90012.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=25440 $Y=186860 $D=9
M80 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 r=27.7778 sa=90001.7 sb=90019.9 a=0.9 p=10.36 mult=1 $X=25815 $Y=128755 $D=9
M81 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90001.7 sb=90019.9 a=1.26 p=14.36 mult=1 $X=25815 $Y=136860 $D=9
M82 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90010.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=25815 $Y=146860 $D=9
M83 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90010.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=25815 $Y=156860 $D=9
M84 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90010.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=25815 $Y=166860 $D=9
M85 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90013.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=26630 $Y=26860 $D=9
M86 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90013.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=26630 $Y=36860 $D=9
M87 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90013.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=26630 $Y=46860 $D=9
M88 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90013.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=26630 $Y=56860 $D=9
M89 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90013.4 sb=90019.9 a=0.9 p=10.36 mult=1 $X=26630 $Y=66860 $D=9
M90 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90010.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=26630 $Y=176860 $D=9
M91 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90013.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=26630 $Y=186860 $D=9
M92 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 r=27.7778 sa=90003.1 sb=90019.9 a=0.9 p=10.36 mult=1 $X=27165 $Y=128755 $D=9
M93 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90003.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=27165 $Y=136860 $D=9
M94 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90011.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=27165 $Y=146860 $D=9
M95 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90011.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=27165 $Y=156860 $D=9
M96 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90011.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=27165 $Y=166860 $D=9
M97 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90015 sb=90019.9 a=1.26 p=14.36 mult=1 $X=28210 $Y=26860 $D=9
M98 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90015 sb=90019.9 a=1.26 p=14.36 mult=1 $X=28210 $Y=36860 $D=9
M99 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90015 sb=90019.9 a=1.26 p=14.36 mult=1 $X=28210 $Y=46860 $D=9
M100 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90015 sb=90019.9 a=1.26 p=14.36 mult=1 $X=28210 $Y=56860 $D=9
M101 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90015 sb=90019.9 a=0.9 p=10.36 mult=1 $X=28210 $Y=66860 $D=9
M102 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90012.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=28210 $Y=176860 $D=9
M103 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90015 sb=90019.9 a=1.26 p=14.36 mult=1 $X=28210 $Y=186860 $D=9
M104 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90016.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=29400 $Y=26860 $D=9
M105 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90016.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=29400 $Y=36860 $D=9
M106 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90016.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=29400 $Y=46860 $D=9
M107 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90016.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=29400 $Y=56860 $D=9
M108 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90016.1 sb=90019.9 a=0.9 p=10.36 mult=1 $X=29400 $Y=66860 $D=9
M109 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90013.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=29400 $Y=176860 $D=9
M110 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90016.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=29400 $Y=186860 $D=9
M111 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 r=27.7778 sa=90005.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=29995 $Y=128755 $D=9
M112 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90005.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=29995 $Y=136860 $D=9
M113 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90014.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=29995 $Y=146860 $D=9
M114 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90014.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=29995 $Y=156860 $D=9
M115 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90014.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=29995 $Y=166860 $D=9
M116 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90017.7 sb=90019.9 a=1.26 p=14.36 mult=1 $X=30980 $Y=26860 $D=9
M117 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90017.7 sb=90019.9 a=1.26 p=14.36 mult=1 $X=30980 $Y=36860 $D=9
M118 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90017.7 sb=90019.9 a=1.26 p=14.36 mult=1 $X=30980 $Y=46860 $D=9
M119 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90017.7 sb=90019.9 a=1.26 p=14.36 mult=1 $X=30980 $Y=56860 $D=9
M120 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90017.7 sb=90019.9 a=0.9 p=10.36 mult=1 $X=30980 $Y=66860 $D=9
M121 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90015 sb=90019.9 a=1.26 p=14.36 mult=1 $X=30980 $Y=176860 $D=9
M122 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90017.7 sb=90019.9 a=1.26 p=14.36 mult=1 $X=30980 $Y=186860 $D=9
M123 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 r=27.7778 sa=90007.3 sb=90019.9 a=0.9 p=10.36 mult=1 $X=31345 $Y=128755 $D=9
M124 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90007.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=31345 $Y=136860 $D=9
M125 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90015.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=31345 $Y=146860 $D=9
M126 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90015.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=31345 $Y=156860 $D=9
M127 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90015.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=31345 $Y=166860 $D=9
M128 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90018.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=32170 $Y=26860 $D=9
M129 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90018.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=32170 $Y=36860 $D=9
M130 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90018.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=32170 $Y=46860 $D=9
M131 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90018.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=32170 $Y=56860 $D=9
M132 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90018.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=32170 $Y=66860 $D=9
M133 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90016.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=32170 $Y=176860 $D=9
M134 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90018.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=32170 $Y=186860 $D=9
M135 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=0.625 sa=4.00001e+06 sb=4.00002e+06 a=40 p=26 mult=1 $X=25535 $Y=75805 $D=9
M136 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 r=0.875 sa=4e+06 sb=4.00002e+06 a=56 p=30 mult=1 $X=25535 $Y=82805 $D=9
M137 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 r=0.875 sa=4e+06 sb=4.00002e+06 a=56 p=30 mult=1 $X=25535 $Y=91300 $D=9
M138 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 r=0.875 sa=4e+06 sb=4.00002e+06 a=56 p=30 mult=1 $X=25535 $Y=101405 $D=9
M139 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 r=0.875 sa=4e+06 sb=4.00002e+06 a=56 p=30 mult=1 $X=25535 $Y=109900 $D=9
M140 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 r=0.875 sa=4e+06 sb=4.00002e+06 a=56 p=30 mult=1 $X=25535 $Y=118725 $D=9
M141 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=33750 $Y=26860 $D=9
M142 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=33750 $Y=36860 $D=9
M143 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=33750 $Y=46860 $D=9
M144 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=33750 $Y=56860 $D=9
M145 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=33750 $Y=66860 $D=9
M146 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90017.7 sb=90019.9 a=1.26 p=14.36 mult=1 $X=33750 $Y=176860 $D=9
M147 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=33750 $Y=186860 $D=9
M148 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 r=27.7778 sa=90010.1 sb=90019.9 a=0.9 p=10.36 mult=1 $X=34175 $Y=128755 $D=9
M149 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90010.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=34175 $Y=136860 $D=9
M150 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90018.5 sb=90019.9 a=1.26 p=14.36 mult=1 $X=34175 $Y=146860 $D=9
M151 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90018.5 sb=90019.9 a=1.26 p=14.36 mult=1 $X=34175 $Y=156860 $D=9
M152 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90018.5 sb=90019.9 a=1.26 p=14.36 mult=1 $X=34175 $Y=166860 $D=9
M153 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=34940 $Y=26860 $D=9
M154 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=34940 $Y=36860 $D=9
M155 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=34940 $Y=46860 $D=9
M156 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=34940 $Y=56860 $D=9
M157 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=34940 $Y=66860 $D=9
M158 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90018.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=34940 $Y=176860 $D=9
M159 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=34940 $Y=186860 $D=9
M160 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 r=27.7778 sa=90011.4 sb=90019.9 a=0.9 p=10.36 mult=1 $X=35525 $Y=128755 $D=9
M161 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90011.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=35525 $Y=136860 $D=9
M162 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.8 sb=90019.9 a=1.26 p=14.36 mult=1 $X=35525 $Y=146860 $D=9
M163 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.8 sb=90019.9 a=1.26 p=14.36 mult=1 $X=35525 $Y=156860 $D=9
M164 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.8 sb=90019.9 a=1.26 p=14.36 mult=1 $X=35525 $Y=166860 $D=9
M165 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=36520 $Y=26860 $D=9
M166 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=36520 $Y=36860 $D=9
M167 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=36520 $Y=46860 $D=9
M168 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=36520 $Y=56860 $D=9
M169 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=36520 $Y=66860 $D=9
M170 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=36520 $Y=176860 $D=9
M171 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=36520 $Y=186860 $D=9
M172 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=37710 $Y=26860 $D=9
M173 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=37710 $Y=36860 $D=9
M174 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=37710 $Y=46860 $D=9
M175 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=37710 $Y=56860 $D=9
M176 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=37710 $Y=66860 $D=9
M177 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=37710 $Y=176860 $D=9
M178 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=37710 $Y=186860 $D=9
M179 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 r=27.7778 sa=90014.3 sb=90019.9 a=0.9 p=10.36 mult=1 $X=38355 $Y=128755 $D=9
M180 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90014.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=38355 $Y=136860 $D=9
M181 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=38355 $Y=146860 $D=9
M182 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=38355 $Y=156860 $D=9
M183 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=38355 $Y=166860 $D=9
M184 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=39290 $Y=26860 $D=9
M185 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=39290 $Y=36860 $D=9
M186 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=39290 $Y=46860 $D=9
M187 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=39290 $Y=56860 $D=9
M188 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=39290 $Y=66860 $D=9
M189 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=39290 $Y=176860 $D=9
M190 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=39290 $Y=186860 $D=9
M191 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 r=27.7778 sa=90015.6 sb=90019.9 a=0.9 p=10.36 mult=1 $X=39705 $Y=128755 $D=9
M192 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90015.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=39705 $Y=136860 $D=9
M193 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=39705 $Y=146860 $D=9
M194 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=39705 $Y=156860 $D=9
M195 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=39705 $Y=166860 $D=9
M196 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=40480 $Y=26860 $D=9
M197 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=40480 $Y=36860 $D=9
M198 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=40480 $Y=46860 $D=9
M199 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=40480 $Y=56860 $D=9
M200 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=40480 $Y=66860 $D=9
M201 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=40480 $Y=176860 $D=9
M202 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=40480 $Y=186860 $D=9
M203 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=0.625 sa=4.00002e+06 sb=4.00002e+06 a=40 p=26 mult=1 $X=33815 $Y=75805 $D=9
M204 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30 mult=1 $X=33815 $Y=82805 $D=9
M205 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30 mult=1 $X=33815 $Y=91300 $D=9
M206 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30 mult=1 $X=33815 $Y=101405 $D=9
M207 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30 mult=1 $X=33815 $Y=109900 $D=9
M208 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30 mult=1 $X=33815 $Y=118725 $D=9
M209 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=42060 $Y=26860 $D=9
M210 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=42060 $Y=36860 $D=9
M211 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=42060 $Y=46860 $D=9
M212 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=42060 $Y=56860 $D=9
M213 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=42060 $Y=66860 $D=9
M214 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=42060 $Y=176860 $D=9
M215 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=42060 $Y=186860 $D=9
M216 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 r=27.7778 sa=90018.5 sb=90019.9 a=0.9 p=10.36 mult=1 $X=42535 $Y=128755 $D=9
M217 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90018.5 sb=90019.9 a=1.26 p=14.36 mult=1 $X=42535 $Y=136860 $D=9
M218 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=42535 $Y=146860 $D=9
M219 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=42535 $Y=156860 $D=9
M220 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=42535 $Y=166860 $D=9
M221 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=43250 $Y=26860 $D=9
M222 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=43250 $Y=36860 $D=9
M223 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=43250 $Y=46860 $D=9
M224 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=43250 $Y=56860 $D=9
M225 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=43250 $Y=66860 $D=9
M226 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=43250 $Y=176860 $D=9
M227 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=43250 $Y=186860 $D=9
M228 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 r=27.7778 sa=90019.8 sb=90019.9 a=0.9 p=10.36 mult=1 $X=43885 $Y=128755 $D=9
M229 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.8 sb=90019.9 a=1.26 p=14.36 mult=1 $X=43885 $Y=136860 $D=9
M230 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=43885 $Y=146860 $D=9
M231 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=43885 $Y=156860 $D=9
M232 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=43885 $Y=166860 $D=9
M233 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=44830 $Y=26860 $D=9
M234 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=44830 $Y=36860 $D=9
M235 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=44830 $Y=46860 $D=9
M236 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=44830 $Y=56860 $D=9
M237 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=44830 $Y=66860 $D=9
M238 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=44830 $Y=176860 $D=9
M239 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=44830 $Y=186860 $D=9
M240 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=46020 $Y=26860 $D=9
M241 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=46020 $Y=36860 $D=9
M242 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=46020 $Y=46860 $D=9
M243 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=46020 $Y=56860 $D=9
M244 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=46020 $Y=66860 $D=9
M245 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=46020 $Y=176860 $D=9
M246 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=46020 $Y=186860 $D=9
M247 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 r=27.7778 sa=90019.9 sb=90019.8 a=0.9 p=10.36 mult=1 $X=46715 $Y=128755 $D=9
M248 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90019.8 a=1.26 p=14.36 mult=1 $X=46715 $Y=136860 $D=9
M249 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90019.8 a=1.26 p=14.36 mult=1 $X=46715 $Y=146860 $D=9
M250 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90019.8 a=1.26 p=14.36 mult=1 $X=46715 $Y=156860 $D=9
M251 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90019.8 a=1.26 p=14.36 mult=1 $X=46715 $Y=166860 $D=9
M252 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90018.9 a=1.26 p=14.36 mult=1 $X=47600 $Y=26860 $D=9
M253 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90018.9 a=1.26 p=14.36 mult=1 $X=47600 $Y=36860 $D=9
M254 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90018.9 a=1.26 p=14.36 mult=1 $X=47600 $Y=46860 $D=9
M255 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90018.9 a=1.26 p=14.36 mult=1 $X=47600 $Y=56860 $D=9
M256 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90018.9 a=0.9 p=10.36 mult=1 $X=47600 $Y=66860 $D=9
M257 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90018.9 a=1.26 p=14.36 mult=1 $X=47600 $Y=176860 $D=9
M258 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90018.9 a=1.26 p=14.36 mult=1 $X=47600 $Y=186860 $D=9
M259 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 r=27.7778 sa=90019.9 sb=90018.5 a=0.9 p=10.36 mult=1 $X=48065 $Y=128755 $D=9
M260 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90018.5 a=1.26 p=14.36 mult=1 $X=48065 $Y=136860 $D=9
M261 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90018.5 a=1.26 p=14.36 mult=1 $X=48065 $Y=146860 $D=9
M262 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90018.5 a=1.26 p=14.36 mult=1 $X=48065 $Y=156860 $D=9
M263 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90018.5 a=1.26 p=14.36 mult=1 $X=48065 $Y=166860 $D=9
M264 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90017.7 a=1.26 p=14.36 mult=1 $X=48790 $Y=26860 $D=9
M265 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90017.7 a=1.26 p=14.36 mult=1 $X=48790 $Y=36860 $D=9
M266 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90017.7 a=1.26 p=14.36 mult=1 $X=48790 $Y=46860 $D=9
M267 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90017.7 a=1.26 p=14.36 mult=1 $X=48790 $Y=56860 $D=9
M268 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90017.7 a=0.9 p=10.36 mult=1 $X=48790 $Y=66860 $D=9
M269 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90017.7 a=1.26 p=14.36 mult=1 $X=48790 $Y=176860 $D=9
M270 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90017.7 a=1.26 p=14.36 mult=1 $X=48790 $Y=186860 $D=9
M271 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=0.625 sa=4.00002e+06 sb=4.00001e+06 a=40 p=26 mult=1 $X=42095 $Y=75805 $D=9
M272 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30 mult=1 $X=42095 $Y=82805 $D=9
M273 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30 mult=1 $X=42095 $Y=91300 $D=9
M274 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30 mult=1 $X=42095 $Y=101405 $D=9
M275 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30 mult=1 $X=42095 $Y=109900 $D=9
M276 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30 mult=1 $X=42095 $Y=118725 $D=9
M277 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90016.2 a=1.26 p=14.36 mult=1 $X=50370 $Y=26860 $D=9
M278 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90016.2 a=1.26 p=14.36 mult=1 $X=50370 $Y=36860 $D=9
M279 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90016.2 a=1.26 p=14.36 mult=1 $X=50370 $Y=46860 $D=9
M280 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90016.2 a=1.26 p=14.36 mult=1 $X=50370 $Y=56860 $D=9
M281 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90016.1 a=0.9 p=10.36 mult=1 $X=50370 $Y=66860 $D=9
M282 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90016.2 a=1.26 p=14.36 mult=1 $X=50370 $Y=176860 $D=9
M283 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90016.2 a=1.26 p=14.36 mult=1 $X=50370 $Y=186860 $D=9
M284 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 r=27.7778 sa=90019.9 sb=90015.6 a=0.9 p=10.36 mult=1 $X=50895 $Y=128755 $D=9
M285 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90015.6 a=1.26 p=14.36 mult=1 $X=50895 $Y=136860 $D=9
M286 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90015.6 a=1.26 p=14.36 mult=1 $X=50895 $Y=146860 $D=9
M287 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90015.6 a=1.26 p=14.36 mult=1 $X=50895 $Y=156860 $D=9
M288 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90015.6 a=1.26 p=14.36 mult=1 $X=50895 $Y=166860 $D=9
M289 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90015 a=1.26 p=14.36 mult=1 $X=51560 $Y=26860 $D=9
M290 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90015 a=1.26 p=14.36 mult=1 $X=51560 $Y=36860 $D=9
M291 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90015 a=1.26 p=14.36 mult=1 $X=51560 $Y=46860 $D=9
M292 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90015 a=1.26 p=14.36 mult=1 $X=51560 $Y=56860 $D=9
M293 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90015 a=0.9 p=10.36 mult=1 $X=51560 $Y=66860 $D=9
M294 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90015 a=1.26 p=14.36 mult=1 $X=51560 $Y=176860 $D=9
M295 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90015 a=1.26 p=14.36 mult=1 $X=51560 $Y=186860 $D=9
M296 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 r=27.7778 sa=90019.9 sb=90014.3 a=0.9 p=10.36 mult=1 $X=52245 $Y=128755 $D=9
M297 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90014.3 a=1.26 p=14.36 mult=1 $X=52245 $Y=136860 $D=9
M298 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90014.3 a=1.26 p=14.36 mult=1 $X=52245 $Y=146860 $D=9
M299 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90014.3 a=1.26 p=14.36 mult=1 $X=52245 $Y=156860 $D=9
M300 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90014.3 a=1.26 p=14.36 mult=1 $X=52245 $Y=166860 $D=9
M301 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90013.4 a=1.26 p=14.36 mult=1 $X=53140 $Y=26860 $D=9
M302 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90013.4 a=1.26 p=14.36 mult=1 $X=53140 $Y=36860 $D=9
M303 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90013.4 a=1.26 p=14.36 mult=1 $X=53140 $Y=46860 $D=9
M304 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90013.4 a=1.26 p=14.36 mult=1 $X=53140 $Y=56860 $D=9
M305 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90013.4 a=0.9 p=10.36 mult=1 $X=53140 $Y=66860 $D=9
M306 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90013.4 a=1.26 p=14.36 mult=1 $X=53140 $Y=176860 $D=9
M307 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90013.4 a=1.26 p=14.36 mult=1 $X=53140 $Y=186860 $D=9
M308 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90012.2 a=1.26 p=14.36 mult=1 $X=54330 $Y=26860 $D=9
M309 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90012.2 a=1.26 p=14.36 mult=1 $X=54330 $Y=36860 $D=9
M310 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90012.2 a=1.26 p=14.36 mult=1 $X=54330 $Y=46860 $D=9
M311 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90012.2 a=1.26 p=14.36 mult=1 $X=54330 $Y=56860 $D=9
M312 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90012.2 a=0.9 p=10.36 mult=1 $X=54330 $Y=66860 $D=9
M313 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90012.2 a=1.26 p=14.36 mult=1 $X=54330 $Y=176860 $D=9
M314 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90012.2 a=1.26 p=14.36 mult=1 $X=54330 $Y=186860 $D=9
M315 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 r=27.7778 sa=90019.9 sb=90011.4 a=0.9 p=10.36 mult=1 $X=55075 $Y=128755 $D=9
M316 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90011.4 a=1.26 p=14.36 mult=1 $X=55075 $Y=136860 $D=9
M317 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90011.4 a=1.26 p=14.36 mult=1 $X=55075 $Y=146860 $D=9
M318 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90011.4 a=1.26 p=14.36 mult=1 $X=55075 $Y=156860 $D=9
M319 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90011.4 a=1.26 p=14.36 mult=1 $X=55075 $Y=166860 $D=9
M320 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90010.6 a=1.26 p=14.36 mult=1 $X=55910 $Y=26860 $D=9
M321 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90010.6 a=1.26 p=14.36 mult=1 $X=55910 $Y=36860 $D=9
M322 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90010.6 a=1.26 p=14.36 mult=1 $X=55910 $Y=46860 $D=9
M323 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90010.6 a=1.26 p=14.36 mult=1 $X=55910 $Y=56860 $D=9
M324 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90010.6 a=0.9 p=10.36 mult=1 $X=55910 $Y=66860 $D=9
M325 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90010.6 a=1.26 p=14.36 mult=1 $X=55910 $Y=176860 $D=9
M326 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90010.6 a=1.26 p=14.36 mult=1 $X=55910 $Y=186860 $D=9
M327 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 r=27.7778 sa=90019.9 sb=90010.1 a=0.9 p=10.36 mult=1 $X=56425 $Y=128755 $D=9
M328 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90010.1 a=1.26 p=14.36 mult=1 $X=56425 $Y=136860 $D=9
M329 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90010.1 a=1.26 p=14.36 mult=1 $X=56425 $Y=146860 $D=9
M330 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90010.1 a=1.26 p=14.36 mult=1 $X=56425 $Y=156860 $D=9
M331 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90010.1 a=1.26 p=14.36 mult=1 $X=56425 $Y=166860 $D=9
M332 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90009.4 a=1.26 p=14.36 mult=1 $X=57100 $Y=26860 $D=9
M333 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90009.4 a=1.26 p=14.36 mult=1 $X=57100 $Y=36860 $D=9
M334 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90009.4 a=1.26 p=14.36 mult=1 $X=57100 $Y=46860 $D=9
M335 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90009.4 a=1.26 p=14.36 mult=1 $X=57100 $Y=56860 $D=9
M336 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90009.4 a=0.9 p=10.36 mult=1 $X=57100 $Y=66860 $D=9
M337 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90009.4 a=1.26 p=14.36 mult=1 $X=57100 $Y=176860 $D=9
M338 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90009.4 a=1.26 p=14.36 mult=1 $X=57100 $Y=186860 $D=9
M339 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=0.625 sa=4.00002e+06 sb=4e+06 a=40 p=26 mult=1 $X=50375 $Y=75805 $D=9
M340 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00002e+06 sb=4e+06 a=56 p=30 mult=1 $X=50375 $Y=82805 $D=9
M341 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00002e+06 sb=4e+06 a=56 p=30 mult=1 $X=50375 $Y=91300 $D=9
M342 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00002e+06 sb=4e+06 a=56 p=30 mult=1 $X=50375 $Y=101405 $D=9
M343 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00002e+06 sb=4e+06 a=56 p=30 mult=1 $X=50375 $Y=109900 $D=9
M344 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00002e+06 sb=4e+06 a=56 p=30 mult=1 $X=50375 $Y=118725 $D=9
M345 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90007.8 a=1.26 p=14.36 mult=1 $X=58680 $Y=26860 $D=9
M346 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90007.8 a=1.26 p=14.36 mult=1 $X=58680 $Y=36860 $D=9
M347 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90007.8 a=1.26 p=14.36 mult=1 $X=58680 $Y=46860 $D=9
M348 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90007.8 a=1.26 p=14.36 mult=1 $X=58680 $Y=56860 $D=9
M349 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90007.8 a=0.9 p=10.36 mult=1 $X=58680 $Y=66860 $D=9
M350 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90007.8 a=1.26 p=14.36 mult=1 $X=58680 $Y=176860 $D=9
M351 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90007.8 a=1.26 p=14.36 mult=1 $X=58680 $Y=186860 $D=9
M352 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 r=27.7778 sa=90019.9 sb=90007.3 a=0.9 p=10.36 mult=1 $X=59255 $Y=128755 $D=9
M353 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90007.3 a=1.26 p=14.36 mult=1 $X=59255 $Y=136860 $D=9
M354 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90007.3 a=1.26 p=14.36 mult=1 $X=59255 $Y=146860 $D=9
M355 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90007.3 a=1.26 p=14.36 mult=1 $X=59255 $Y=156860 $D=9
M356 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90007.3 a=1.26 p=14.36 mult=1 $X=59255 $Y=166860 $D=9
M357 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90006.6 a=1.26 p=14.36 mult=1 $X=59870 $Y=26860 $D=9
M358 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90006.6 a=1.26 p=14.36 mult=1 $X=59870 $Y=36860 $D=9
M359 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90006.6 a=1.26 p=14.36 mult=1 $X=59870 $Y=46860 $D=9
M360 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90006.6 a=1.26 p=14.36 mult=1 $X=59870 $Y=56860 $D=9
M361 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90006.6 a=0.9 p=10.36 mult=1 $X=59870 $Y=66860 $D=9
M362 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90006.6 a=1.26 p=14.36 mult=1 $X=59870 $Y=176860 $D=9
M363 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90006.6 a=1.26 p=14.36 mult=1 $X=59870 $Y=186860 $D=9
M364 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 r=27.7778 sa=90019.9 sb=90005.9 a=0.9 p=10.36 mult=1 $X=60605 $Y=128755 $D=9
M365 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90005.9 a=1.26 p=14.36 mult=1 $X=60605 $Y=136860 $D=9
M366 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90005.9 a=1.26 p=14.36 mult=1 $X=60605 $Y=146860 $D=9
M367 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90005.9 a=1.26 p=14.36 mult=1 $X=60605 $Y=156860 $D=9
M368 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90005.9 a=1.26 p=14.36 mult=1 $X=60605 $Y=166860 $D=9
M369 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90005.1 a=1.26 p=14.36 mult=1 $X=61450 $Y=26860 $D=9
M370 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90005.1 a=1.26 p=14.36 mult=1 $X=61450 $Y=36860 $D=9
M371 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90005.1 a=1.26 p=14.36 mult=1 $X=61450 $Y=46860 $D=9
M372 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90005.1 a=1.26 p=14.36 mult=1 $X=61450 $Y=56860 $D=9
M373 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90005.1 a=0.9 p=10.36 mult=1 $X=61450 $Y=66860 $D=9
M374 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90005.1 a=1.26 p=14.36 mult=1 $X=61450 $Y=176860 $D=9
M375 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90005.1 a=1.26 p=14.36 mult=1 $X=61450 $Y=186860 $D=9
M376 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90003.9 a=1.26 p=14.36 mult=1 $X=62640 $Y=26860 $D=9
M377 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90003.9 a=1.26 p=14.36 mult=1 $X=62640 $Y=36860 $D=9
M378 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90003.9 a=1.26 p=14.36 mult=1 $X=62640 $Y=46860 $D=9
M379 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90003.9 a=1.26 p=14.36 mult=1 $X=62640 $Y=56860 $D=9
M380 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90003.9 a=0.9 p=10.36 mult=1 $X=62640 $Y=66860 $D=9
M381 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90003.9 a=1.26 p=14.36 mult=1 $X=62640 $Y=176860 $D=9
M382 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90003.9 a=1.26 p=14.36 mult=1 $X=62640 $Y=186860 $D=9
M383 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 r=27.7778 sa=90019.9 sb=90003.1 a=0.9 p=10.36 mult=1 $X=63435 $Y=128755 $D=9
M384 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90003.1 a=1.26 p=14.36 mult=1 $X=63435 $Y=136860 $D=9
M385 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90003.1 a=1.26 p=14.36 mult=1 $X=63435 $Y=146860 $D=9
M386 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90003.1 a=1.26 p=14.36 mult=1 $X=63435 $Y=156860 $D=9
M387 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90003.1 a=1.26 p=14.36 mult=1 $X=63435 $Y=166860 $D=9
M388 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90002.3 a=1.26 p=14.36 mult=1 $X=64220 $Y=26860 $D=9
M389 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90002.3 a=1.26 p=14.36 mult=1 $X=64220 $Y=36860 $D=9
M390 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90002.3 a=1.26 p=14.36 mult=1 $X=64220 $Y=46860 $D=9
M391 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90002.3 a=1.26 p=14.36 mult=1 $X=64220 $Y=56860 $D=9
M392 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90002.3 a=0.9 p=10.36 mult=1 $X=64220 $Y=66860 $D=9
M393 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90002.3 a=1.26 p=14.36 mult=1 $X=64220 $Y=176860 $D=9
M394 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90002.3 a=1.26 p=14.36 mult=1 $X=64220 $Y=186860 $D=9
M395 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 r=27.7778 sa=90019.9 sb=90001.7 a=0.9 p=10.36 mult=1 $X=64785 $Y=128755 $D=9
M396 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90001.7 a=1.26 p=14.36 mult=1 $X=64785 $Y=136860 $D=9
M397 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90001.7 a=1.26 p=14.36 mult=1 $X=64785 $Y=146860 $D=9
M398 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90001.7 a=1.26 p=14.36 mult=1 $X=64785 $Y=156860 $D=9
M399 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90001.7 a=1.26 p=14.36 mult=1 $X=64785 $Y=166860 $D=9
M400 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90001.1 a=1.26 p=14.36 mult=1 $X=65410 $Y=26860 $D=9
M401 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90001.1 a=1.26 p=14.36 mult=1 $X=65410 $Y=36860 $D=9
M402 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90001.1 a=1.26 p=14.36 mult=1 $X=65410 $Y=46860 $D=9
M403 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90001.1 a=1.26 p=14.36 mult=1 $X=65410 $Y=56860 $D=9
M404 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90001.1 a=0.9 p=10.36 mult=1 $X=65410 $Y=66860 $D=9
M405 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90001.1 a=1.26 p=14.36 mult=1 $X=65410 $Y=176860 $D=9
M406 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90001.1 a=1.26 p=14.36 mult=1 $X=65410 $Y=186860 $D=9
M407 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 r=0.625 sa=4.00002e+06 sb=4e+06 a=40 p=26 mult=1 $X=58655 $Y=75805 $D=9
M408 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00002e+06 sb=4e+06 a=56 p=30 mult=1 $X=58655 $Y=82805 $D=9
M409 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00002e+06 sb=4e+06 a=56 p=30 mult=1 $X=58655 $Y=91300 $D=9
M410 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00002e+06 sb=4e+06 a=56 p=30 mult=1 $X=58655 $Y=101405 $D=9
M411 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00002e+06 sb=4e+06 a=56 p=30 mult=1 $X=58655 $Y=109900 $D=9
M412 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00002e+06 sb=4e+06 a=56 p=30 mult=1 $X=58655 $Y=118725 $D=9
X413 SRC_BDY_LVC1 VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=40185 $Y=114790 $D=150
X414 SRC_BDY_LVC2 VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=40605 $Y=34930 $D=150
X415 SRC_BDY_LVC1 VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=40640 $Y=196080 $D=150
X416 VSSD DRN_LVC1 Dpar a=108.41 p=46.58 m=1 $[nwdiode] $X=1015 $Y=685 $D=191
X417 VSSD DRN_LVC2 Dpar a=108.41 p=46.58 m=1 $[nwdiode] $X=67280 $Y=745 $D=191
X418 VSSD VDDIO Dpar a=10516.3 p=468.87 m=1 $[dnwdiode_psub] $X=9500 $Y=23605 $D=193
X419 SRC_BDY_LVC2 VDDIO Dpar a=4115.42 p=264.63 m=1 $[dnwdiode_pw] $X=10870 $Y=24975 $D=194
X420 SRC_BDY_LVC1 VDDIO Dpar a=5703.29 p=340.89 m=1 $[dnwdiode_pw] $X=10870 $Y=83485 $D=194
R421 DRN_LVC1 21 L=1950 W=0.33 m=1 mult=1 model="mrp1" $[mrp1] $X=240 $Y=19200 $D=257
R422 P_CORE P_PAD 0.01 m=1 $[short] $X=6670 $Y=103345 $D=286
X423 27 DRN_LVC2 sky130_fd_pr__res_bent_po__example_55959141808692 $T=70965 18130 0 90 $X=70615 $Y=17860
X424 DRN_LVC1 21 24 sky130_fd_pr__pfet_01v8__example_55959141808687 $T=2070 2020 0 0 $X=1610 $Y=1840
X425 DRN_LVC1 21 24 sky130_fd_pr__pfet_01v8__example_55959141808687 $T=2070 9670 0 0 $X=1610 $Y=9490
X426 DRN_LVC2 23 25 sky130_fd_pr__pfet_01v8__example_55959141808687 $T=68335 2080 0 0 $X=67875 $Y=1900
X427 DRN_LVC2 23 25 sky130_fd_pr__pfet_01v8__example_55959141808687 $T=68335 9730 0 0 $X=67875 $Y=9550
X616 23 26 sky130_fd_pr__res_bent_po__example_55959141808691 $T=66785 1745 1 90 $X=57045 $Y=1475
X622 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808704 $T=25815 136860 0 0 $X=23860 $Y=136700
X623 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808695 $T=25815 128755 0 0 $X=23860 $Y=128595
X630 VSSD BDY2_B2B SRC_BDY_LVC1 sky130_fd_io__gnd2gnd_120x2_lv_isosub $T=16525 18480 1 0 $X=16525 $Y=320
X631 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808701 $T=17130 176860 0 0 $X=15800 $Y=176700
X632 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808703 $T=17455 146860 0 0 $X=15500 $Y=146700
X633 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808703 $T=17455 156860 0 0 $X=15500 $Y=156700
X634 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808703 $T=17455 166860 0 0 $X=15500 $Y=166700
X635 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705 $T=14360 26860 0 0 $X=13030 $Y=26700
X636 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705 $T=14360 36860 0 0 $X=13030 $Y=36700
X637 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705 $T=14360 46860 0 0 $X=13030 $Y=46700
X638 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705 $T=14360 56860 0 0 $X=13030 $Y=56700
X639 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808705 $T=14360 186860 0 0 $X=13030 $Y=186700
X640 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808693 $T=14360 66860 0 0 $X=13030 $Y=66700
X642 22 26 sky130_fd_pr__res_bent_po__example_55959141808688 $T=11245 84330 0 90 $X=10895 $Y=84060
X643 27 22 sky130_fd_pr__res_bent_po__example_55959141808690 $T=69775 19510 0 180 $X=10025 $Y=19160
.ENDS
***************************************
.SUBCKT sky130_ef_io__vccd_lvc_clamped2_pad VSSD VSSA VSSIO VCCD VDDIO VCCD_PAD
** N=13 EP=6 IP=20 FDC=501
*.CALIBRE ISOLATED NETS: VCCHIB VDDA VSWITCH AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
X0 VSSD VSSD VSSIO VCCD VDDIO VCCD VSSA VCCD VCCD_PAD sky130_fd_io__top_power_lvc_wpad $T=0 -35 0 0 $X=0 $Y=-35
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_55959141808669 2 3
** N=6 EP=2 IP=0 FDC=1
R0 2 3 L=470 W=0.33 m=1 mult=1 model="mrp1" $[mrp1] $X=-250 $Y=-1620 $D=257
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1__example_55959141808662
** N=60 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1__example_55959141808663
** N=120 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__model__nfet_highvoltage__example_55959141808664 2 3
** N=38 EP=2 IP=34 FDC=1
*.SEEDPROM
M0 2 3 2 2 nhv L=4 W=5 AD=1.325 AS=1.325 PD=10.53 PS=10.53 NRD=0 NRS=0 m=1 r=1.25 sa=2e+06 sb=2e+06 a=20 p=18 mult=1 $X=0 $Y=0 $D=49
.ENDS
***************************************
.SUBCKT sky130_fd_io__sio_clamp_pcap_4x5 2 3
** N=84 EP=2 IP=7 FDC=1
*.SEEDPROM
X0 2 3 sky130_fd_pr__model__nfet_highvoltage__example_55959141808664 $T=1145 720 0 0 $X=700 $Y=540
.ENDS
***************************************
.SUBCKT sky130_fd_io__esd_rcclamp_nfetcap 2 3
** N=150 EP=2 IP=34 FDC=1
*.SEEDPROM
M0 2 3 2 2 nhv L=8 W=5 AD=1.325 AS=1.325 PD=10.53 PS=10.53 NRD=0 NRS=0 m=1 r=0.625 sa=4e+06 sb=4e+06 a=40 p=26 mult=1 $X=895 $Y=630 $D=49
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd__example_55959141808678
** N=23 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_6
** N=45 EP=0 IP=48 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_7
** N=5 EP=0 IP=10 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808677 2 3 4
** N=81 EP=3 IP=26 FDC=15
*.SEEDPROM
M0 4 3 2 2 nhv L=0.5 W=7 AD=0.98 AS=1.855 PD=7.28 PS=14.53 NRD=0 NRS=0 m=1 r=14 sa=250000 sb=250011 a=3.5 p=15 mult=1 $X=0 $Y=0 $D=49
M1 2 3 4 2 nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250001 sb=250010 a=3.5 p=15 mult=1 $X=780 $Y=0 $D=49
M2 4 3 2 2 nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250002 sb=250009 a=3.5 p=15 mult=1 $X=1560 $Y=0 $D=49
M3 2 3 4 2 nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250002 sb=250009 a=3.5 p=15 mult=1 $X=2340 $Y=0 $D=49
M4 4 3 2 2 nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250003 sb=250008 a=3.5 p=15 mult=1 $X=3120 $Y=0 $D=49
M5 2 3 4 2 nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250004 sb=250007 a=3.5 p=15 mult=1 $X=3900 $Y=0 $D=49
M6 4 3 2 2 nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250005 sb=250006 a=3.5 p=15 mult=1 $X=4680 $Y=0 $D=49
M7 2 3 4 2 nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250005 sb=250005 a=3.5 p=15 mult=1 $X=5460 $Y=0 $D=49
M8 4 3 2 2 nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250006 sb=250005 a=3.5 p=15 mult=1 $X=6240 $Y=0 $D=49
M9 2 3 4 2 nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250007 sb=250004 a=3.5 p=15 mult=1 $X=7020 $Y=0 $D=49
M10 4 3 2 2 nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250008 sb=250003 a=3.5 p=15 mult=1 $X=7800 $Y=0 $D=49
M11 2 3 4 2 nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250009 sb=250002 a=3.5 p=15 mult=1 $X=8580 $Y=0 $D=49
M12 4 3 2 2 nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250009 sb=250002 a=3.5 p=15 mult=1 $X=9360 $Y=0 $D=49
M13 2 3 4 2 nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250010 sb=250001 a=3.5 p=15 mult=1 $X=10140 $Y=0 $D=49
M14 4 3 2 2 nhv L=0.5 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250011 sb=250000 a=3.5 p=15 mult=1 $X=10920 $Y=0 $D=49
.ENDS
***************************************
.SUBCKT ICV_8 2 3
** N=167 EP=2 IP=188 FDC=2
*.SEEDPROM
X0 2 3 sky130_fd_io__esd_rcclamp_nfetcap $T=-9760 0 0 0 $X=-10010 $Y=-90
X1 2 3 sky130_fd_io__esd_rcclamp_nfetcap $T=0 0 0 0 $X=-250 $Y=-90
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s__example_55959141808671
** N=119 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s2__example_55959141808672
** N=177 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808670
** N=23 EP=0 IP=30 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s__example_55959141808675
** N=61 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s2__example_55959141808676
** N=90 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808674
** N=27 EP=0 IP=36 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808673
** N=27 EP=0 IP=36 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_55959141808668 2 3
** N=6 EP=2 IP=0 FDC=1
R0 2 3 L=700 W=0.33 m=1 mult=1 model="mrp1" $[mrp1] $X=-250 $Y=-8100 $D=257
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd__example_55959141808336
** N=22 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_9
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_10
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_11
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_12
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808665 2 3 4
** N=254 EP=3 IP=16 FDC=50
*.SEEDPROM
M0 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=1.855 PD=7.28 PS=14.53 NRD=0 NRS=0 m=1 r=14 sa=250000 sb=250020 a=3.5 p=15 mult=1 $X=0 $Y=0 $D=109
M1 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250001 sb=250020 a=3.5 p=15 mult=1 $X=780 $Y=0 $D=109
M2 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250002 sb=250020 a=3.5 p=15 mult=1 $X=1560 $Y=0 $D=109
M3 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250002 sb=250020 a=3.5 p=15 mult=1 $X=2340 $Y=0 $D=109
M4 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250003 sb=250020 a=3.5 p=15 mult=1 $X=3120 $Y=0 $D=109
M5 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250004 sb=250020 a=3.5 p=15 mult=1 $X=3900 $Y=0 $D=109
M6 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250005 sb=250020 a=3.5 p=15 mult=1 $X=4680 $Y=0 $D=109
M7 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250005 sb=250020 a=3.5 p=15 mult=1 $X=5460 $Y=0 $D=109
M8 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250006 sb=250020 a=3.5 p=15 mult=1 $X=6240 $Y=0 $D=109
M9 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250007 sb=250020 a=3.5 p=15 mult=1 $X=7020 $Y=0 $D=109
M10 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250008 sb=250020 a=3.5 p=15 mult=1 $X=7800 $Y=0 $D=109
M11 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250009 sb=250020 a=3.5 p=15 mult=1 $X=8580 $Y=0 $D=109
M12 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250009 sb=250020 a=3.5 p=15 mult=1 $X=9360 $Y=0 $D=109
M13 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250010 sb=250020 a=3.5 p=15 mult=1 $X=10140 $Y=0 $D=109
M14 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250011 sb=250020 a=3.5 p=15 mult=1 $X=10920 $Y=0 $D=109
M15 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250012 sb=250020 a=3.5 p=15 mult=1 $X=11700 $Y=0 $D=109
M16 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250012 sb=250020 a=3.5 p=15 mult=1 $X=12480 $Y=0 $D=109
M17 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250013 sb=250020 a=3.5 p=15 mult=1 $X=13260 $Y=0 $D=109
M18 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250014 sb=250020 a=3.5 p=15 mult=1 $X=14040 $Y=0 $D=109
M19 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250015 sb=250020 a=3.5 p=15 mult=1 $X=14820 $Y=0 $D=109
M20 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250016 sb=250020 a=3.5 p=15 mult=1 $X=15600 $Y=0 $D=109
M21 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250016 sb=250020 a=3.5 p=15 mult=1 $X=16380 $Y=0 $D=109
M22 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250017 sb=250020 a=3.5 p=15 mult=1 $X=17160 $Y=0 $D=109
M23 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250018 sb=250020 a=3.5 p=15 mult=1 $X=17940 $Y=0 $D=109
M24 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250019 sb=250020 a=3.5 p=15 mult=1 $X=18720 $Y=0 $D=109
M25 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250019 a=3.5 p=15 mult=1 $X=19500 $Y=0 $D=109
M26 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250018 a=3.5 p=15 mult=1 $X=20280 $Y=0 $D=109
M27 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250017 a=3.5 p=15 mult=1 $X=21060 $Y=0 $D=109
M28 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250016 a=3.5 p=15 mult=1 $X=21840 $Y=0 $D=109
M29 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250016 a=3.5 p=15 mult=1 $X=22620 $Y=0 $D=109
M30 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250015 a=3.5 p=15 mult=1 $X=23400 $Y=0 $D=109
M31 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250014 a=3.5 p=15 mult=1 $X=24180 $Y=0 $D=109
M32 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250013 a=3.5 p=15 mult=1 $X=24960 $Y=0 $D=109
M33 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250012 a=3.5 p=15 mult=1 $X=25740 $Y=0 $D=109
M34 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250012 a=3.5 p=15 mult=1 $X=26520 $Y=0 $D=109
M35 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250011 a=3.5 p=15 mult=1 $X=27300 $Y=0 $D=109
M36 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250010 a=3.5 p=15 mult=1 $X=28080 $Y=0 $D=109
M37 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250009 a=3.5 p=15 mult=1 $X=28860 $Y=0 $D=109
M38 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250009 a=3.5 p=15 mult=1 $X=29640 $Y=0 $D=109
M39 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250008 a=3.5 p=15 mult=1 $X=30420 $Y=0 $D=109
M40 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250007 a=3.5 p=15 mult=1 $X=31200 $Y=0 $D=109
M41 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250006 a=3.5 p=15 mult=1 $X=31980 $Y=0 $D=109
M42 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250005 a=3.5 p=15 mult=1 $X=32760 $Y=0 $D=109
M43 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250005 a=3.5 p=15 mult=1 $X=33540 $Y=0 $D=109
M44 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250004 a=3.5 p=15 mult=1 $X=34320 $Y=0 $D=109
M45 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250003 a=3.5 p=15 mult=1 $X=35100 $Y=0 $D=109
M46 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250002 a=3.5 p=15 mult=1 $X=35880 $Y=0 $D=109
M47 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250002 a=3.5 p=15 mult=1 $X=36660 $Y=0 $D=109
M48 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250001 a=3.5 p=15 mult=1 $X=37440 $Y=0 $D=109
M49 2 3 4 2 phv L=0.5 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250000 a=3.5 p=15 mult=1 $X=38220 $Y=0 $D=109
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_55959141808667 2 3
** N=6 EP=2 IP=0 FDC=1
R0 2 3 L=1550 W=0.33 m=1 mult=1 model="mrp1" $[mrp1] $X=-250 $Y=-6480 $D=257
.ENDS
***************************************
.SUBCKT sky130_fd_io__top_ground_hvc_wpad VSSD SRC_BDY_HVC DRN_HVC VDDIO G_CORE G_PAD
** N=14148 EP=6 IP=1976 FDC=241
*.CALIBRE ISOLATED NETS: OGC_HVC VCCHIB VCCD VDDA VSSIO VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
M0 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=15885 $Y=47180 $D=49
M1 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=15885 $Y=139180 $D=49
M2 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=15885 $Y=162180 $D=49
M3 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250001 sb=250020 a=5 p=21 mult=1 $X=15885 $Y=185180 $D=49
M4 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=17895 $Y=47180 $D=49
M5 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=17895 $Y=139180 $D=49
M6 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=17895 $Y=162180 $D=49
M7 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250003 sb=250020 a=5 p=21 mult=1 $X=17895 $Y=185180 $D=49
M8 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=20485 $Y=47180 $D=49
M9 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=20485 $Y=139180 $D=49
M10 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=20485 $Y=162180 $D=49
M11 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250006 sb=250020 a=5 p=21 mult=1 $X=20485 $Y=185180 $D=49
M12 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=22495 $Y=47180 $D=49
M13 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=22495 $Y=139180 $D=49
M14 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=22495 $Y=162180 $D=49
M15 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250008 sb=250020 a=5 p=21 mult=1 $X=22495 $Y=185180 $D=49
M16 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=25085 $Y=47180 $D=49
M17 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=25085 $Y=70180 $D=49
M18 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=25085 $Y=93180 $D=49
M19 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=25085 $Y=116180 $D=49
M20 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=25085 $Y=139180 $D=49
M21 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=25085 $Y=162180 $D=49
M22 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250010 sb=250020 a=5 p=21 mult=1 $X=25085 $Y=185180 $D=49
M23 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=27095 $Y=47180 $D=49
M24 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=27095 $Y=70180 $D=49
M25 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=27095 $Y=93180 $D=49
M26 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=27095 $Y=116180 $D=49
M27 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=27095 $Y=139180 $D=49
M28 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=27095 $Y=162180 $D=49
M29 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250012 sb=250020 a=5 p=21 mult=1 $X=27095 $Y=185180 $D=49
M30 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=29685 $Y=47180 $D=49
M31 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=29685 $Y=70180 $D=49
M32 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=29685 $Y=93180 $D=49
M33 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=29685 $Y=116180 $D=49
M34 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=29685 $Y=139180 $D=49
M35 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=29685 $Y=162180 $D=49
M36 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250015 sb=250020 a=5 p=21 mult=1 $X=29685 $Y=185180 $D=49
M37 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=31695 $Y=47180 $D=49
M38 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=31695 $Y=70180 $D=49
M39 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=31695 $Y=93180 $D=49
M40 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=31695 $Y=116180 $D=49
M41 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=31695 $Y=139180 $D=49
M42 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=31695 $Y=162180 $D=49
M43 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250017 sb=250020 a=5 p=21 mult=1 $X=31695 $Y=185180 $D=49
M44 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=34285 $Y=47180 $D=49
M45 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=34285 $Y=70180 $D=49
M46 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=34285 $Y=93180 $D=49
M47 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=34285 $Y=116180 $D=49
M48 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=34285 $Y=139180 $D=49
M49 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=34285 $Y=162180 $D=49
M50 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=34285 $Y=185180 $D=49
M51 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=36295 $Y=47180 $D=49
M52 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=36295 $Y=70180 $D=49
M53 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=36295 $Y=93180 $D=49
M54 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=36295 $Y=116180 $D=49
M55 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=36295 $Y=139180 $D=49
M56 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=36295 $Y=162180 $D=49
M57 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=36295 $Y=185180 $D=49
M58 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=38885 $Y=47180 $D=49
M59 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=38885 $Y=70180 $D=49
M60 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=38885 $Y=93180 $D=49
M61 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=38885 $Y=116180 $D=49
M62 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=38885 $Y=139180 $D=49
M63 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=38885 $Y=162180 $D=49
M64 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=38885 $Y=185180 $D=49
M65 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=40895 $Y=47180 $D=49
M66 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=40895 $Y=70180 $D=49
M67 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=40895 $Y=93180 $D=49
M68 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=40895 $Y=116180 $D=49
M69 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=40895 $Y=139180 $D=49
M70 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=40895 $Y=162180 $D=49
M71 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=40895 $Y=185180 $D=49
M72 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=43485 $Y=47180 $D=49
M73 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=43485 $Y=70180 $D=49
M74 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=43485 $Y=93180 $D=49
M75 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=43485 $Y=116180 $D=49
M76 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=43485 $Y=139180 $D=49
M77 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=43485 $Y=162180 $D=49
M78 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=43485 $Y=185180 $D=49
M79 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=45495 $Y=47180 $D=49
M80 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=45495 $Y=70180 $D=49
M81 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=45495 $Y=93180 $D=49
M82 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=45495 $Y=116180 $D=49
M83 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=45495 $Y=139180 $D=49
M84 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=45495 $Y=162180 $D=49
M85 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=45495 $Y=185180 $D=49
M86 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=48085 $Y=47180 $D=49
M87 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=48085 $Y=70180 $D=49
M88 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=48085 $Y=93180 $D=49
M89 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=48085 $Y=116180 $D=49
M90 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=48085 $Y=139180 $D=49
M91 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=48085 $Y=162180 $D=49
M92 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250017 a=5 p=21 mult=1 $X=48085 $Y=185180 $D=49
M93 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=50095 $Y=47180 $D=49
M94 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=50095 $Y=70180 $D=49
M95 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=50095 $Y=93180 $D=49
M96 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=50095 $Y=116180 $D=49
M97 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=50095 $Y=139180 $D=49
M98 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=50095 $Y=162180 $D=49
M99 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250015 a=5 p=21 mult=1 $X=50095 $Y=185180 $D=49
M100 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=52685 $Y=47180 $D=49
M101 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=52685 $Y=70180 $D=49
M102 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=52685 $Y=93180 $D=49
M103 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=52685 $Y=116180 $D=49
M104 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=52685 $Y=139180 $D=49
M105 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=52685 $Y=162180 $D=49
M106 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250012 a=5 p=21 mult=1 $X=52685 $Y=185180 $D=49
M107 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=54695 $Y=47180 $D=49
M108 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=54695 $Y=70180 $D=49
M109 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=54695 $Y=93180 $D=49
M110 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=54695 $Y=116180 $D=49
M111 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=54695 $Y=139180 $D=49
M112 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=54695 $Y=162180 $D=49
M113 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250010 a=5 p=21 mult=1 $X=54695 $Y=185180 $D=49
M114 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=57285 $Y=47180 $D=49
M115 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=57285 $Y=70180 $D=49
M116 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=57285 $Y=93180 $D=49
M117 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=57285 $Y=116180 $D=49
M118 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=57285 $Y=139180 $D=49
M119 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=57285 $Y=162180 $D=49
M120 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250008 a=5 p=21 mult=1 $X=57285 $Y=185180 $D=49
M121 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=59295 $Y=47180 $D=49
M122 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=59295 $Y=70180 $D=49
M123 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=59295 $Y=93180 $D=49
M124 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=59295 $Y=116180 $D=49
M125 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=59295 $Y=139180 $D=49
M126 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=59295 $Y=162180 $D=49
M127 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250006 a=5 p=21 mult=1 $X=59295 $Y=185180 $D=49
M128 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=61885 $Y=47180 $D=49
M129 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=61885 $Y=70180 $D=49
M130 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=61885 $Y=93180 $D=49
M131 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=61885 $Y=116180 $D=49
M132 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=61885 $Y=139180 $D=49
M133 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=61885 $Y=162180 $D=49
M134 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250003 a=5 p=21 mult=1 $X=61885 $Y=185180 $D=49
M135 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=63895 $Y=47180 $D=49
M136 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=63895 $Y=70180 $D=49
M137 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=63895 $Y=93180 $D=49
M138 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=63895 $Y=116180 $D=49
M139 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=63895 $Y=139180 $D=49
M140 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=63895 $Y=162180 $D=49
M141 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250001 a=5 p=21 mult=1 $X=63895 $Y=185180 $D=49
X142 SRC_BDY_HVC VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=51225 $Y=21735 $D=150
X143 SRC_BDY_HVC VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=51225 $Y=45310 $D=150
X144 SRC_BDY_HVC VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=64770 $Y=40835 $D=150
X145 SRC_BDY_HVC VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=68375 $Y=197675 $D=150
X146 VSSD VDDIO Dpar a=126.883 p=0 m=1 $[nwdiode] $X=8835 $Y=43175 $D=189
X147 VSSD DRN_HVC Dpar a=376.949 p=101.73 m=1 $[nwdiode] $X=4400 $Y=28925 $D=191
X148 VSSD VDDIO Dpar a=10358.7 p=619.08 m=1 $[dnwdiode_psub] $X=9500 $Y=133835 $D=193
X149 SRC_BDY_HVC VDDIO Dpar a=137.463 p=47.72 m=1 $[dnwdiode_pw] $X=53530 $Y=31395 $D=194
X150 SRC_BDY_HVC VDDIO Dpar a=8184.99 p=443.22 m=1 $[dnwdiode_pw] $X=10695 $Y=45035 $D=194
X151 SRC_BDY_HVC VDDIO Dpar a=1172.63 p=163 m=1 $[dnwdiode_pw] $X=13380 $Y=2205 $D=194
R152 G_CORE G_PAD 0.01 m=1 $[short] $X=6670 $Y=105345 $D=286
X153 18 20 sky130_fd_pr__res_bent_po__example_55959141808669 $T=71055 43015 0 90 $X=70705 $Y=42745
X225 SRC_BDY_HVC 18 sky130_fd_pr__model__nfet_highvoltage__example_55959141808664 $T=61815 27145 0 180 $X=57370 $Y=21965
X226 SRC_BDY_HVC 18 sky130_fd_io__sio_clamp_pcap_4x5 $T=19920 9205 0 180 $X=13630 $Y=2455
X227 SRC_BDY_HVC 18 sky130_fd_io__sio_clamp_pcap_4x5 $T=19920 15425 0 180 $X=13630 $Y=8675
X228 SRC_BDY_HVC 18 sky130_fd_io__sio_clamp_pcap_4x5 $T=19920 21645 0 180 $X=13630 $Y=14895
X229 SRC_BDY_HVC 18 sky130_fd_io__sio_clamp_pcap_4x5 $T=68720 27865 0 180 $X=62430 $Y=21115
X230 SRC_BDY_HVC 18 sky130_fd_io__esd_rcclamp_nfetcap $T=68470 9115 0 180 $X=58430 $Y=2455
X231 SRC_BDY_HVC 18 sky130_fd_io__esd_rcclamp_nfetcap $T=68470 15335 0 180 $X=58430 $Y=8675
X232 SRC_BDY_HVC 18 sky130_fd_io__esd_rcclamp_nfetcap $T=68470 21555 0 180 $X=58430 $Y=14895
X233 SRC_BDY_HVC 18 19 sky130_fd_pr__nfet_01v8__example_55959141808677 $T=54915 32580 0 0 $X=54470 $Y=32400
X234 SRC_BDY_HVC 18 ICV_8 $T=29430 9115 0 180 $X=19390 $Y=2455
X235 SRC_BDY_HVC 18 ICV_8 $T=29430 15335 0 180 $X=19390 $Y=8675
X236 SRC_BDY_HVC 18 ICV_8 $T=29430 21555 0 180 $X=19390 $Y=14895
X237 SRC_BDY_HVC 18 ICV_8 $T=48950 9115 0 180 $X=38910 $Y=2455
X238 SRC_BDY_HVC 18 ICV_8 $T=48950 15335 0 180 $X=38910 $Y=8675
X239 SRC_BDY_HVC 18 ICV_8 $T=48950 21555 0 180 $X=38910 $Y=14895
X247 DRN_HVC 21 sky130_fd_pr__res_bent_po__example_55959141808668 $T=9830 74355 0 90 $X=9480 $Y=74085
X248 DRN_HVC 18 19 sky130_fd_pr__pfet_01v8__example_55959141808665 $T=6340 29800 0 0 $X=5745 $Y=29470
X249 21 20 sky130_fd_pr__res_bent_po__example_55959141808667 $T=8360 43440 1 90 $X=1050 $Y=43170
.ENDS
***************************************
.SUBCKT sky130_ef_io__vssio_hvc_clamped_pad VSSD VDDIO VSSIO VSSIO_PAD
** N=12 EP=4 IP=17 FDC=241
*.CALIBRE ISOLATED NETS: VCCHIB VCCD VDDA VSWITCH VSSA AMUXBUS_B AMUXBUS_A VDDIO_Q
X0 VSSD VSSIO VDDIO VDDIO VSSIO VSSIO_PAD sky130_fd_io__top_ground_hvc_wpad $T=0 -2035 0 0 $X=0 $Y=-2035
*.CALIBRE WARNING SHORT Short circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT sky130_ef_io__vssa_hvc_clamped_pad VSSD VDDIO VSSA VDDA VSSA_PAD
** N=13 EP=5 IP=17 FDC=241
*.CALIBRE ISOLATED NETS: VCCHIB VCCD VSSIO VSWITCH AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
X0 VSSD VSSA VDDA VDDIO VSSA VSSA_PAD sky130_fd_io__top_ground_hvc_wpad $T=0 -2035 0 0 $X=0 $Y=-2035
.ENDS
***************************************
.SUBCKT ICV_13 1 16 115 193 195 199 206 207 212 213 214 215
** N=281 EP=12 IP=51 FDC=1484
X0 1 193 16 199 195 212 sky130_ef_io__vccd_lvc_clamped2_pad $T=197965 4560000 0 90 $X=0 $Y=4560000
X1 1 115 16 207 195 215 sky130_ef_io__vccd_lvc_clamped2_pad $T=3390035 4613000 0 270 $X=3379500 $Y=4526805
X2 1 195 16 213 sky130_ef_io__vssio_hvc_clamped_pad $T=1667000 4990035 0 0 $X=1667000 $Y=4988000
X3 1 195 115 206 214 sky130_ef_io__vssa_hvc_clamped_pad $T=2878000 4990035 0 0 $X=2878000 $Y=4988000
.ENDS
***************************************
.SUBCKT sky130_fd_io__top_power_hvc_wpadv2 VSSD SRC_BDY_HVC DRN_HVC VDDIO P_CORE P_PAD
** N=18956 EP=6 IP=1976 FDC=241
*.CALIBRE ISOLATED NETS: OGC_HVC VCCHIB VCCD VDDA VSSIO VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
M0 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=15885 $Y=47180 $D=49
M1 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=15885 $Y=139180 $D=49
M2 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=15885 $Y=162180 $D=49
M3 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250001 sb=250020 a=5 p=21 mult=1 $X=15885 $Y=185180 $D=49
M4 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=17895 $Y=47180 $D=49
M5 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=17895 $Y=139180 $D=49
M6 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=17895 $Y=162180 $D=49
M7 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250003 sb=250020 a=5 p=21 mult=1 $X=17895 $Y=185180 $D=49
M8 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=20485 $Y=47180 $D=49
M9 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=20485 $Y=139180 $D=49
M10 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=20485 $Y=162180 $D=49
M11 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250006 sb=250020 a=5 p=21 mult=1 $X=20485 $Y=185180 $D=49
M12 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=22495 $Y=47180 $D=49
M13 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=22495 $Y=139180 $D=49
M14 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=22495 $Y=162180 $D=49
M15 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250008 sb=250020 a=5 p=21 mult=1 $X=22495 $Y=185180 $D=49
M16 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=25085 $Y=47180 $D=49
M17 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=25085 $Y=70180 $D=49
M18 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=25085 $Y=93180 $D=49
M19 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=25085 $Y=116180 $D=49
M20 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=25085 $Y=139180 $D=49
M21 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=25085 $Y=162180 $D=49
M22 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250010 sb=250020 a=5 p=21 mult=1 $X=25085 $Y=185180 $D=49
M23 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=27095 $Y=47180 $D=49
M24 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=27095 $Y=70180 $D=49
M25 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=27095 $Y=93180 $D=49
M26 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=27095 $Y=116180 $D=49
M27 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=27095 $Y=139180 $D=49
M28 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=27095 $Y=162180 $D=49
M29 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250012 sb=250020 a=5 p=21 mult=1 $X=27095 $Y=185180 $D=49
M30 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=29685 $Y=47180 $D=49
M31 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=29685 $Y=70180 $D=49
M32 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=29685 $Y=93180 $D=49
M33 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=29685 $Y=116180 $D=49
M34 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=29685 $Y=139180 $D=49
M35 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=29685 $Y=162180 $D=49
M36 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250015 sb=250020 a=5 p=21 mult=1 $X=29685 $Y=185180 $D=49
M37 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=31695 $Y=47180 $D=49
M38 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=31695 $Y=70180 $D=49
M39 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=31695 $Y=93180 $D=49
M40 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=31695 $Y=116180 $D=49
M41 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=31695 $Y=139180 $D=49
M42 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=31695 $Y=162180 $D=49
M43 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250017 sb=250020 a=5 p=21 mult=1 $X=31695 $Y=185180 $D=49
M44 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=34285 $Y=47180 $D=49
M45 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=34285 $Y=70180 $D=49
M46 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=34285 $Y=93180 $D=49
M47 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=34285 $Y=116180 $D=49
M48 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=34285 $Y=139180 $D=49
M49 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=34285 $Y=162180 $D=49
M50 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=34285 $Y=185180 $D=49
M51 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=36295 $Y=47180 $D=49
M52 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=36295 $Y=70180 $D=49
M53 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=36295 $Y=93180 $D=49
M54 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=36295 $Y=116180 $D=49
M55 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=36295 $Y=139180 $D=49
M56 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=36295 $Y=162180 $D=49
M57 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=36295 $Y=185180 $D=49
M58 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=38885 $Y=47180 $D=49
M59 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=38885 $Y=70180 $D=49
M60 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=38885 $Y=93180 $D=49
M61 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=38885 $Y=116180 $D=49
M62 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=38885 $Y=139180 $D=49
M63 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=38885 $Y=162180 $D=49
M64 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=38885 $Y=185180 $D=49
M65 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=40895 $Y=47180 $D=49
M66 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=40895 $Y=70180 $D=49
M67 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=40895 $Y=93180 $D=49
M68 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=40895 $Y=116180 $D=49
M69 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=40895 $Y=139180 $D=49
M70 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=40895 $Y=162180 $D=49
M71 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=40895 $Y=185180 $D=49
M72 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=43485 $Y=47180 $D=49
M73 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=43485 $Y=70180 $D=49
M74 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=43485 $Y=93180 $D=49
M75 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=43485 $Y=116180 $D=49
M76 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=43485 $Y=139180 $D=49
M77 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=43485 $Y=162180 $D=49
M78 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=43485 $Y=185180 $D=49
M79 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=45495 $Y=47180 $D=49
M80 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=45495 $Y=70180 $D=49
M81 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=45495 $Y=93180 $D=49
M82 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=45495 $Y=116180 $D=49
M83 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=45495 $Y=139180 $D=49
M84 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=45495 $Y=162180 $D=49
M85 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=45495 $Y=185180 $D=49
M86 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=48085 $Y=47180 $D=49
M87 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=48085 $Y=70180 $D=49
M88 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=48085 $Y=93180 $D=49
M89 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=48085 $Y=116180 $D=49
M90 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=48085 $Y=139180 $D=49
M91 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=48085 $Y=162180 $D=49
M92 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250017 a=5 p=21 mult=1 $X=48085 $Y=185180 $D=49
M93 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=50095 $Y=47180 $D=49
M94 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=50095 $Y=70180 $D=49
M95 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=50095 $Y=93180 $D=49
M96 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=50095 $Y=116180 $D=49
M97 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=50095 $Y=139180 $D=49
M98 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=50095 $Y=162180 $D=49
M99 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250015 a=5 p=21 mult=1 $X=50095 $Y=185180 $D=49
M100 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=52685 $Y=47180 $D=49
M101 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=52685 $Y=70180 $D=49
M102 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=52685 $Y=93180 $D=49
M103 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=52685 $Y=116180 $D=49
M104 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=52685 $Y=139180 $D=49
M105 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=52685 $Y=162180 $D=49
M106 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250012 a=5 p=21 mult=1 $X=52685 $Y=185180 $D=49
M107 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=54695 $Y=47180 $D=49
M108 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=54695 $Y=70180 $D=49
M109 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=54695 $Y=93180 $D=49
M110 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=54695 $Y=116180 $D=49
M111 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=54695 $Y=139180 $D=49
M112 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=54695 $Y=162180 $D=49
M113 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250010 a=5 p=21 mult=1 $X=54695 $Y=185180 $D=49
M114 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=57285 $Y=47180 $D=49
M115 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=57285 $Y=70180 $D=49
M116 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=57285 $Y=93180 $D=49
M117 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=57285 $Y=116180 $D=49
M118 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=57285 $Y=139180 $D=49
M119 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=57285 $Y=162180 $D=49
M120 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250008 a=5 p=21 mult=1 $X=57285 $Y=185180 $D=49
M121 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=59295 $Y=47180 $D=49
M122 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=59295 $Y=70180 $D=49
M123 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=59295 $Y=93180 $D=49
M124 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=59295 $Y=116180 $D=49
M125 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=59295 $Y=139180 $D=49
M126 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=59295 $Y=162180 $D=49
M127 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250006 a=5 p=21 mult=1 $X=59295 $Y=185180 $D=49
M128 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=61885 $Y=47180 $D=49
M129 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=61885 $Y=70180 $D=49
M130 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=61885 $Y=93180 $D=49
M131 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=61885 $Y=116180 $D=49
M132 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=61885 $Y=139180 $D=49
M133 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=61885 $Y=162180 $D=49
M134 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250003 a=5 p=21 mult=1 $X=61885 $Y=185180 $D=49
M135 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=63895 $Y=47180 $D=49
M136 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=63895 $Y=70180 $D=49
M137 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=63895 $Y=93180 $D=49
M138 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=63895 $Y=116180 $D=49
M139 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=63895 $Y=139180 $D=49
M140 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=63895 $Y=162180 $D=49
M141 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250001 a=5 p=21 mult=1 $X=63895 $Y=185180 $D=49
X142 SRC_BDY_HVC VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=51225 $Y=21735 $D=150
X143 SRC_BDY_HVC VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=51225 $Y=45310 $D=150
X144 SRC_BDY_HVC VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=64770 $Y=40835 $D=150
X145 SRC_BDY_HVC VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=68375 $Y=197675 $D=150
X146 VSSD VDDIO Dpar a=126.766 p=0 m=1 $[nwdiode] $X=8835 $Y=43175 $D=189
X147 VSSD DRN_HVC Dpar a=369.745 p=100.13 m=1 $[nwdiode] $X=5200 $Y=28925 $D=191
X148 VSSD VDDIO Dpar a=10358.7 p=619.08 m=1 $[dnwdiode_psub] $X=9500 $Y=133835 $D=193
X149 SRC_BDY_HVC VDDIO Dpar a=137.463 p=47.72 m=1 $[dnwdiode_pw] $X=53530 $Y=31395 $D=194
X150 SRC_BDY_HVC VDDIO Dpar a=8184.99 p=443.22 m=1 $[dnwdiode_pw] $X=10695 $Y=45035 $D=194
X151 SRC_BDY_HVC VDDIO Dpar a=1172.63 p=163 m=1 $[dnwdiode_pw] $X=13380 $Y=2205 $D=194
R152 P_CORE P_PAD 0.01 m=1 $[short] $X=6670 $Y=105345 $D=286
X153 19 20 sky130_fd_pr__res_bent_po__example_55959141808669 $T=71055 42015 0 90 $X=70705 $Y=41745
X225 SRC_BDY_HVC 19 sky130_fd_pr__model__nfet_highvoltage__example_55959141808664 $T=61815 27145 0 180 $X=57370 $Y=21965
X226 SRC_BDY_HVC 19 sky130_fd_io__sio_clamp_pcap_4x5 $T=19920 9205 0 180 $X=13630 $Y=2455
X227 SRC_BDY_HVC 19 sky130_fd_io__sio_clamp_pcap_4x5 $T=19920 15425 0 180 $X=13630 $Y=8675
X228 SRC_BDY_HVC 19 sky130_fd_io__sio_clamp_pcap_4x5 $T=19920 21645 0 180 $X=13630 $Y=14895
X229 SRC_BDY_HVC 19 sky130_fd_io__sio_clamp_pcap_4x5 $T=68720 27865 0 180 $X=62430 $Y=21115
X230 SRC_BDY_HVC 19 sky130_fd_io__esd_rcclamp_nfetcap $T=68470 9115 0 180 $X=58430 $Y=2455
X231 SRC_BDY_HVC 19 sky130_fd_io__esd_rcclamp_nfetcap $T=68470 15335 0 180 $X=58430 $Y=8675
X232 SRC_BDY_HVC 19 sky130_fd_io__esd_rcclamp_nfetcap $T=68470 21555 0 180 $X=58430 $Y=14895
X233 SRC_BDY_HVC 19 21 sky130_fd_pr__nfet_01v8__example_55959141808677 $T=54915 32580 0 0 $X=54470 $Y=32400
X234 SRC_BDY_HVC 19 ICV_8 $T=29430 9115 0 180 $X=19390 $Y=2455
X235 SRC_BDY_HVC 19 ICV_8 $T=29430 15335 0 180 $X=19390 $Y=8675
X236 SRC_BDY_HVC 19 ICV_8 $T=29430 21555 0 180 $X=19390 $Y=14895
X237 SRC_BDY_HVC 19 ICV_8 $T=48950 9115 0 180 $X=38910 $Y=2455
X238 SRC_BDY_HVC 19 ICV_8 $T=48950 15335 0 180 $X=38910 $Y=8675
X239 SRC_BDY_HVC 19 ICV_8 $T=48950 21555 0 180 $X=38910 $Y=14895
X247 DRN_HVC 18 sky130_fd_pr__res_bent_po__example_55959141808668 $T=9830 74355 0 90 $X=9480 $Y=74085
X248 DRN_HVC 19 21 sky130_fd_pr__pfet_01v8__example_55959141808665 $T=6340 29800 0 0 $X=5745 $Y=29470
X249 18 20 sky130_fd_pr__res_bent_po__example_55959141808667 $T=8360 43440 1 90 $X=1050 $Y=43170
.ENDS
***************************************
.SUBCKT sky130_ef_io__vddio_hvc_clamped_pad VSSD VSSIO VDDIO VDDIO_PAD
** N=12 EP=4 IP=17 FDC=241
*.CALIBRE ISOLATED NETS: VCCHIB VCCD VDDA VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q
X0 VSSD VSSIO VDDIO VDDIO VDDIO VDDIO_PAD sky130_fd_io__top_power_hvc_wpadv2 $T=0 -2035 0 0 $X=0 $Y=-2035
*.CALIBRE WARNING SHORT Short circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT ICV_14 1 3 16
** N=38 EP=3 IP=12 FDC=241
X0 1 3 16 38 sky130_ef_io__vddio_hvc_clamped_pad $T=197965 4349000 0 90 $X=0 $Y=4349000
.ENDS
***************************************
.SUBCKT sky130_ef_io__vdda_hvc_clamped_pad VSSD VSSA VDDIO VDDA VDDA_PAD
** N=13 EP=5 IP=17 FDC=241
*.CALIBRE ISOLATED NETS: VCCHIB VCCD VSSIO VSWITCH AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
X0 VSSD VSSA VDDA VDDIO VDDA VDDA_PAD sky130_fd_io__top_power_hvc_wpadv2 $T=0 -2035 0 0 $X=0 $Y=-2035
.ENDS
***************************************
.SUBCKT ICV_15 1 142 191 192 229 239 248 249
** N=327 EP=8 IP=26 FDC=482
X0 1 191 229 239 248 sky130_ef_io__vssa_hvc_clamped_pad $T=197965 4138000 0 90 $X=0 $Y=4138000
X1 1 192 191 142 249 sky130_ef_io__vdda_hvc_clamped_pad $T=3390035 4167000 0 270 $X=3388000 $Y=4092000
.ENDS
***************************************
.SUBCKT sky130_fd_io__top_ground_lvc_wpad VSSD SRC_BDY_LVC2 SRC_BDY_LVC1 DRN_LVC1 VDDIO DRN_LVC2 BDY2_B2B G_CORE G_PAD
** N=12725 EP=9 IP=1228 FDC=501
*.CALIBRE ISOLATED NETS: OGC_LVC VCCHIB VCCD VDDA VSSIO VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
M0 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90001.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=14360 $Y=26860 $D=9
M1 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90001.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=14360 $Y=36860 $D=9
M2 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90001.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=14360 $Y=46860 $D=9
M3 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90001.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=14360 $Y=56860 $D=9
M4 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90001.1 sb=90019.9 a=0.9 p=10.36 mult=1 $X=14360 $Y=66860 $D=9
M5 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90001.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=14360 $Y=186860 $D=9
M6 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90002.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=15550 $Y=26860 $D=9
M7 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90002.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=15550 $Y=36860 $D=9
M8 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90002.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=15550 $Y=46860 $D=9
M9 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90002.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=15550 $Y=56860 $D=9
M10 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90002.3 sb=90019.9 a=0.9 p=10.36 mult=1 $X=15550 $Y=66860 $D=9
M11 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90002.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=15550 $Y=186860 $D=9
M12 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=4 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 r=1.25 sa=2e+06 sb=2.00002e+06 a=20 p=18 mult=1 $X=12975 $Y=75805 $D=9
M13 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90003.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=17130 $Y=26860 $D=9
M14 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90003.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=17130 $Y=36860 $D=9
M15 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90003.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=17130 $Y=46860 $D=9
M16 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90003.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=17130 $Y=56860 $D=9
M17 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90003.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=17130 $Y=66860 $D=9
M18 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90001.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=17130 $Y=176860 $D=9
M19 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90003.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=17130 $Y=186860 $D=9
M20 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90001.7 sb=90019.9 a=1.26 p=14.36 mult=1 $X=17455 $Y=146860 $D=9
M21 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90001.7 sb=90019.9 a=1.26 p=14.36 mult=1 $X=17455 $Y=156860 $D=9
M22 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90001.7 sb=90019.9 a=1.26 p=14.36 mult=1 $X=17455 $Y=166860 $D=9
M23 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90005.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=18320 $Y=26860 $D=9
M24 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90005.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=18320 $Y=36860 $D=9
M25 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90005.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=18320 $Y=46860 $D=9
M26 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90005.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=18320 $Y=56860 $D=9
M27 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90005.1 sb=90019.9 a=0.9 p=10.36 mult=1 $X=18320 $Y=66860 $D=9
M28 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90002.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=18320 $Y=176860 $D=9
M29 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90005.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=18320 $Y=186860 $D=9
M30 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90003.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=18805 $Y=146860 $D=9
M31 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90003.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=18805 $Y=156860 $D=9
M32 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90003.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=18805 $Y=166860 $D=9
M33 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90006.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=19900 $Y=26860 $D=9
M34 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90006.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=19900 $Y=36860 $D=9
M35 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90006.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=19900 $Y=46860 $D=9
M36 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90006.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=19900 $Y=56860 $D=9
M37 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90006.6 sb=90019.9 a=0.9 p=10.36 mult=1 $X=19900 $Y=66860 $D=9
M38 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90003.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=19900 $Y=176860 $D=9
M39 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90006.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=19900 $Y=186860 $D=9
M40 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90007.8 sb=90019.9 a=1.26 p=14.36 mult=1 $X=21090 $Y=26860 $D=9
M41 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90007.8 sb=90019.9 a=1.26 p=14.36 mult=1 $X=21090 $Y=36860 $D=9
M42 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90007.8 sb=90019.9 a=1.26 p=14.36 mult=1 $X=21090 $Y=46860 $D=9
M43 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90007.8 sb=90019.9 a=1.26 p=14.36 mult=1 $X=21090 $Y=56860 $D=9
M44 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90007.8 sb=90019.9 a=0.9 p=10.36 mult=1 $X=21090 $Y=66860 $D=9
M45 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90005.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=21090 $Y=176860 $D=9
M46 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90007.8 sb=90019.9 a=1.26 p=14.36 mult=1 $X=21090 $Y=186860 $D=9
M47 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90005.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=21635 $Y=146860 $D=9
M48 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90005.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=21635 $Y=156860 $D=9
M49 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90005.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=21635 $Y=166860 $D=9
M50 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90009.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=22670 $Y=26860 $D=9
M51 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90009.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=22670 $Y=36860 $D=9
M52 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90009.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=22670 $Y=46860 $D=9
M53 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90009.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=22670 $Y=56860 $D=9
M54 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90009.4 sb=90019.9 a=0.9 p=10.36 mult=1 $X=22670 $Y=66860 $D=9
M55 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90006.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=22670 $Y=176860 $D=9
M56 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90009.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=22670 $Y=186860 $D=9
M57 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90007.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=22985 $Y=146860 $D=9
M58 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90007.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=22985 $Y=156860 $D=9
M59 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90007.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=22985 $Y=166860 $D=9
M60 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90010.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=23860 $Y=26860 $D=9
M61 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90010.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=23860 $Y=36860 $D=9
M62 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90010.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=23860 $Y=46860 $D=9
M63 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90010.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=23860 $Y=56860 $D=9
M64 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90010.6 sb=90019.9 a=0.9 p=10.36 mult=1 $X=23860 $Y=66860 $D=9
M65 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90007.8 sb=90019.9 a=1.26 p=14.36 mult=1 $X=23860 $Y=176860 $D=9
M66 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90010.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=23860 $Y=186860 $D=9
M67 SRC_BDY_LVC2 23 25 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 r=38.8889 sa=90000.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=24670 $Y=82805 $D=9
M68 SRC_BDY_LVC2 23 25 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 r=38.8889 sa=90000.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=24670 $Y=91300 $D=9
M69 SRC_BDY_LVC1 21 24 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 r=38.8889 sa=90000.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=24670 $Y=101405 $D=9
M70 SRC_BDY_LVC1 21 24 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 r=38.8889 sa=90000.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=24670 $Y=109900 $D=9
M71 SRC_BDY_LVC1 21 24 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 r=38.8889 sa=90000.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=24670 $Y=118725 $D=9
M72 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=0.625 sa=4e+06 sb=4.00002e+06 a=40 p=26 mult=1 $X=17255 $Y=75805 $D=9
M73 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90012.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=25440 $Y=26860 $D=9
M74 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90012.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=25440 $Y=36860 $D=9
M75 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90012.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=25440 $Y=46860 $D=9
M76 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90012.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=25440 $Y=56860 $D=9
M77 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90012.2 sb=90019.9 a=0.9 p=10.36 mult=1 $X=25440 $Y=66860 $D=9
M78 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90009.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=25440 $Y=176860 $D=9
M79 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90012.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=25440 $Y=186860 $D=9
M80 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 r=27.7778 sa=90001.7 sb=90019.9 a=0.9 p=10.36 mult=1 $X=25815 $Y=128755 $D=9
M81 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90001.7 sb=90019.9 a=1.26 p=14.36 mult=1 $X=25815 $Y=136860 $D=9
M82 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90010.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=25815 $Y=146860 $D=9
M83 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90010.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=25815 $Y=156860 $D=9
M84 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90010.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=25815 $Y=166860 $D=9
M85 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90013.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=26630 $Y=26860 $D=9
M86 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90013.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=26630 $Y=36860 $D=9
M87 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90013.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=26630 $Y=46860 $D=9
M88 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90013.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=26630 $Y=56860 $D=9
M89 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90013.4 sb=90019.9 a=0.9 p=10.36 mult=1 $X=26630 $Y=66860 $D=9
M90 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90010.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=26630 $Y=176860 $D=9
M91 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90013.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=26630 $Y=186860 $D=9
M92 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 r=27.7778 sa=90003.1 sb=90019.9 a=0.9 p=10.36 mult=1 $X=27165 $Y=128755 $D=9
M93 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90003.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=27165 $Y=136860 $D=9
M94 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90011.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=27165 $Y=146860 $D=9
M95 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90011.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=27165 $Y=156860 $D=9
M96 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90011.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=27165 $Y=166860 $D=9
M97 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90015 sb=90019.9 a=1.26 p=14.36 mult=1 $X=28210 $Y=26860 $D=9
M98 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90015 sb=90019.9 a=1.26 p=14.36 mult=1 $X=28210 $Y=36860 $D=9
M99 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90015 sb=90019.9 a=1.26 p=14.36 mult=1 $X=28210 $Y=46860 $D=9
M100 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90015 sb=90019.9 a=1.26 p=14.36 mult=1 $X=28210 $Y=56860 $D=9
M101 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90015 sb=90019.9 a=0.9 p=10.36 mult=1 $X=28210 $Y=66860 $D=9
M102 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90012.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=28210 $Y=176860 $D=9
M103 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90015 sb=90019.9 a=1.26 p=14.36 mult=1 $X=28210 $Y=186860 $D=9
M104 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90016.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=29400 $Y=26860 $D=9
M105 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90016.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=29400 $Y=36860 $D=9
M106 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90016.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=29400 $Y=46860 $D=9
M107 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90016.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=29400 $Y=56860 $D=9
M108 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90016.1 sb=90019.9 a=0.9 p=10.36 mult=1 $X=29400 $Y=66860 $D=9
M109 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90013.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=29400 $Y=176860 $D=9
M110 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90016.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=29400 $Y=186860 $D=9
M111 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 r=27.7778 sa=90005.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=29995 $Y=128755 $D=9
M112 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90005.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=29995 $Y=136860 $D=9
M113 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90014.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=29995 $Y=146860 $D=9
M114 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90014.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=29995 $Y=156860 $D=9
M115 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90014.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=29995 $Y=166860 $D=9
M116 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90017.7 sb=90019.9 a=1.26 p=14.36 mult=1 $X=30980 $Y=26860 $D=9
M117 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90017.7 sb=90019.9 a=1.26 p=14.36 mult=1 $X=30980 $Y=36860 $D=9
M118 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90017.7 sb=90019.9 a=1.26 p=14.36 mult=1 $X=30980 $Y=46860 $D=9
M119 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90017.7 sb=90019.9 a=1.26 p=14.36 mult=1 $X=30980 $Y=56860 $D=9
M120 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90017.7 sb=90019.9 a=0.9 p=10.36 mult=1 $X=30980 $Y=66860 $D=9
M121 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90015 sb=90019.9 a=1.26 p=14.36 mult=1 $X=30980 $Y=176860 $D=9
M122 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90017.7 sb=90019.9 a=1.26 p=14.36 mult=1 $X=30980 $Y=186860 $D=9
M123 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 r=27.7778 sa=90007.3 sb=90019.9 a=0.9 p=10.36 mult=1 $X=31345 $Y=128755 $D=9
M124 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90007.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=31345 $Y=136860 $D=9
M125 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90015.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=31345 $Y=146860 $D=9
M126 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90015.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=31345 $Y=156860 $D=9
M127 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90015.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=31345 $Y=166860 $D=9
M128 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90018.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=32170 $Y=26860 $D=9
M129 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90018.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=32170 $Y=36860 $D=9
M130 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90018.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=32170 $Y=46860 $D=9
M131 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90018.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=32170 $Y=56860 $D=9
M132 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90018.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=32170 $Y=66860 $D=9
M133 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90016.2 sb=90019.9 a=1.26 p=14.36 mult=1 $X=32170 $Y=176860 $D=9
M134 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90018.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=32170 $Y=186860 $D=9
M135 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=0.625 sa=4.00001e+06 sb=4.00002e+06 a=40 p=26 mult=1 $X=25535 $Y=75805 $D=9
M136 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 r=0.875 sa=4e+06 sb=4.00002e+06 a=56 p=30 mult=1 $X=25535 $Y=82805 $D=9
M137 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 r=0.875 sa=4e+06 sb=4.00002e+06 a=56 p=30 mult=1 $X=25535 $Y=91300 $D=9
M138 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 r=0.875 sa=4e+06 sb=4.00002e+06 a=56 p=30 mult=1 $X=25535 $Y=101405 $D=9
M139 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 r=0.875 sa=4e+06 sb=4.00002e+06 a=56 p=30 mult=1 $X=25535 $Y=109900 $D=9
M140 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 r=0.875 sa=4e+06 sb=4.00002e+06 a=56 p=30 mult=1 $X=25535 $Y=118725 $D=9
M141 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=33750 $Y=26860 $D=9
M142 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=33750 $Y=36860 $D=9
M143 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=33750 $Y=46860 $D=9
M144 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=33750 $Y=56860 $D=9
M145 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=33750 $Y=66860 $D=9
M146 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90017.7 sb=90019.9 a=1.26 p=14.36 mult=1 $X=33750 $Y=176860 $D=9
M147 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=33750 $Y=186860 $D=9
M148 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 r=27.7778 sa=90010.1 sb=90019.9 a=0.9 p=10.36 mult=1 $X=34175 $Y=128755 $D=9
M149 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90010.1 sb=90019.9 a=1.26 p=14.36 mult=1 $X=34175 $Y=136860 $D=9
M150 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90018.5 sb=90019.9 a=1.26 p=14.36 mult=1 $X=34175 $Y=146860 $D=9
M151 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90018.5 sb=90019.9 a=1.26 p=14.36 mult=1 $X=34175 $Y=156860 $D=9
M152 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90018.5 sb=90019.9 a=1.26 p=14.36 mult=1 $X=34175 $Y=166860 $D=9
M153 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=34940 $Y=26860 $D=9
M154 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=34940 $Y=36860 $D=9
M155 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=34940 $Y=46860 $D=9
M156 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=34940 $Y=56860 $D=9
M157 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=34940 $Y=66860 $D=9
M158 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90018.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=34940 $Y=176860 $D=9
M159 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=34940 $Y=186860 $D=9
M160 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 r=27.7778 sa=90011.4 sb=90019.9 a=0.9 p=10.36 mult=1 $X=35525 $Y=128755 $D=9
M161 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90011.4 sb=90019.9 a=1.26 p=14.36 mult=1 $X=35525 $Y=136860 $D=9
M162 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.8 sb=90019.9 a=1.26 p=14.36 mult=1 $X=35525 $Y=146860 $D=9
M163 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.8 sb=90019.9 a=1.26 p=14.36 mult=1 $X=35525 $Y=156860 $D=9
M164 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.8 sb=90019.9 a=1.26 p=14.36 mult=1 $X=35525 $Y=166860 $D=9
M165 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=36520 $Y=26860 $D=9
M166 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=36520 $Y=36860 $D=9
M167 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=36520 $Y=46860 $D=9
M168 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=36520 $Y=56860 $D=9
M169 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=36520 $Y=66860 $D=9
M170 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=36520 $Y=176860 $D=9
M171 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=36520 $Y=186860 $D=9
M172 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=37710 $Y=26860 $D=9
M173 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=37710 $Y=36860 $D=9
M174 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=37710 $Y=46860 $D=9
M175 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=37710 $Y=56860 $D=9
M176 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=37710 $Y=66860 $D=9
M177 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=37710 $Y=176860 $D=9
M178 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=37710 $Y=186860 $D=9
M179 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 r=27.7778 sa=90014.3 sb=90019.9 a=0.9 p=10.36 mult=1 $X=38355 $Y=128755 $D=9
M180 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90014.3 sb=90019.9 a=1.26 p=14.36 mult=1 $X=38355 $Y=136860 $D=9
M181 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=38355 $Y=146860 $D=9
M182 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=38355 $Y=156860 $D=9
M183 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=38355 $Y=166860 $D=9
M184 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=39290 $Y=26860 $D=9
M185 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=39290 $Y=36860 $D=9
M186 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=39290 $Y=46860 $D=9
M187 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=39290 $Y=56860 $D=9
M188 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=39290 $Y=66860 $D=9
M189 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=39290 $Y=176860 $D=9
M190 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=39290 $Y=186860 $D=9
M191 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 r=27.7778 sa=90015.6 sb=90019.9 a=0.9 p=10.36 mult=1 $X=39705 $Y=128755 $D=9
M192 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90015.6 sb=90019.9 a=1.26 p=14.36 mult=1 $X=39705 $Y=136860 $D=9
M193 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=39705 $Y=146860 $D=9
M194 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=39705 $Y=156860 $D=9
M195 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=39705 $Y=166860 $D=9
M196 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=40480 $Y=26860 $D=9
M197 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=40480 $Y=36860 $D=9
M198 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=40480 $Y=46860 $D=9
M199 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=40480 $Y=56860 $D=9
M200 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=40480 $Y=66860 $D=9
M201 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=40480 $Y=176860 $D=9
M202 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=40480 $Y=186860 $D=9
M203 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=0.625 sa=4.00002e+06 sb=4.00002e+06 a=40 p=26 mult=1 $X=33815 $Y=75805 $D=9
M204 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30 mult=1 $X=33815 $Y=82805 $D=9
M205 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30 mult=1 $X=33815 $Y=91300 $D=9
M206 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30 mult=1 $X=33815 $Y=101405 $D=9
M207 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30 mult=1 $X=33815 $Y=109900 $D=9
M208 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30 mult=1 $X=33815 $Y=118725 $D=9
M209 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=42060 $Y=26860 $D=9
M210 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=42060 $Y=36860 $D=9
M211 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=42060 $Y=46860 $D=9
M212 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=42060 $Y=56860 $D=9
M213 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=42060 $Y=66860 $D=9
M214 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=42060 $Y=176860 $D=9
M215 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=42060 $Y=186860 $D=9
M216 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 r=27.7778 sa=90018.5 sb=90019.9 a=0.9 p=10.36 mult=1 $X=42535 $Y=128755 $D=9
M217 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90018.5 sb=90019.9 a=1.26 p=14.36 mult=1 $X=42535 $Y=136860 $D=9
M218 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=42535 $Y=146860 $D=9
M219 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=42535 $Y=156860 $D=9
M220 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=42535 $Y=166860 $D=9
M221 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=43250 $Y=26860 $D=9
M222 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=43250 $Y=36860 $D=9
M223 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=43250 $Y=46860 $D=9
M224 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=43250 $Y=56860 $D=9
M225 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=43250 $Y=66860 $D=9
M226 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=43250 $Y=176860 $D=9
M227 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=43250 $Y=186860 $D=9
M228 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 r=27.7778 sa=90019.8 sb=90019.9 a=0.9 p=10.36 mult=1 $X=43885 $Y=128755 $D=9
M229 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.8 sb=90019.9 a=1.26 p=14.36 mult=1 $X=43885 $Y=136860 $D=9
M230 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=43885 $Y=146860 $D=9
M231 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=43885 $Y=156860 $D=9
M232 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=43885 $Y=166860 $D=9
M233 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=44830 $Y=26860 $D=9
M234 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=44830 $Y=36860 $D=9
M235 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=44830 $Y=46860 $D=9
M236 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=44830 $Y=56860 $D=9
M237 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=44830 $Y=66860 $D=9
M238 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=44830 $Y=176860 $D=9
M239 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=44830 $Y=186860 $D=9
M240 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=46020 $Y=26860 $D=9
M241 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=46020 $Y=36860 $D=9
M242 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=46020 $Y=46860 $D=9
M243 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=46020 $Y=56860 $D=9
M244 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90019.9 a=0.9 p=10.36 mult=1 $X=46020 $Y=66860 $D=9
M245 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=46020 $Y=176860 $D=9
M246 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90019.9 a=1.26 p=14.36 mult=1 $X=46020 $Y=186860 $D=9
M247 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 r=27.7778 sa=90019.9 sb=90019.8 a=0.9 p=10.36 mult=1 $X=46715 $Y=128755 $D=9
M248 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90019.8 a=1.26 p=14.36 mult=1 $X=46715 $Y=136860 $D=9
M249 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90019.8 a=1.26 p=14.36 mult=1 $X=46715 $Y=146860 $D=9
M250 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90019.8 a=1.26 p=14.36 mult=1 $X=46715 $Y=156860 $D=9
M251 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90019.8 a=1.26 p=14.36 mult=1 $X=46715 $Y=166860 $D=9
M252 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90018.9 a=1.26 p=14.36 mult=1 $X=47600 $Y=26860 $D=9
M253 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90018.9 a=1.26 p=14.36 mult=1 $X=47600 $Y=36860 $D=9
M254 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90018.9 a=1.26 p=14.36 mult=1 $X=47600 $Y=46860 $D=9
M255 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90018.9 a=1.26 p=14.36 mult=1 $X=47600 $Y=56860 $D=9
M256 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90018.9 a=0.9 p=10.36 mult=1 $X=47600 $Y=66860 $D=9
M257 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90018.9 a=1.26 p=14.36 mult=1 $X=47600 $Y=176860 $D=9
M258 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90018.9 a=1.26 p=14.36 mult=1 $X=47600 $Y=186860 $D=9
M259 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 r=27.7778 sa=90019.9 sb=90018.5 a=0.9 p=10.36 mult=1 $X=48065 $Y=128755 $D=9
M260 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90018.5 a=1.26 p=14.36 mult=1 $X=48065 $Y=136860 $D=9
M261 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90018.5 a=1.26 p=14.36 mult=1 $X=48065 $Y=146860 $D=9
M262 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90018.5 a=1.26 p=14.36 mult=1 $X=48065 $Y=156860 $D=9
M263 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90018.5 a=1.26 p=14.36 mult=1 $X=48065 $Y=166860 $D=9
M264 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90017.7 a=1.26 p=14.36 mult=1 $X=48790 $Y=26860 $D=9
M265 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90017.7 a=1.26 p=14.36 mult=1 $X=48790 $Y=36860 $D=9
M266 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90017.7 a=1.26 p=14.36 mult=1 $X=48790 $Y=46860 $D=9
M267 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90017.7 a=1.26 p=14.36 mult=1 $X=48790 $Y=56860 $D=9
M268 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90017.7 a=0.9 p=10.36 mult=1 $X=48790 $Y=66860 $D=9
M269 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90017.7 a=1.26 p=14.36 mult=1 $X=48790 $Y=176860 $D=9
M270 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90017.7 a=1.26 p=14.36 mult=1 $X=48790 $Y=186860 $D=9
M271 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=0.625 sa=4.00002e+06 sb=4.00001e+06 a=40 p=26 mult=1 $X=42095 $Y=75805 $D=9
M272 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30 mult=1 $X=42095 $Y=82805 $D=9
M273 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30 mult=1 $X=42095 $Y=91300 $D=9
M274 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30 mult=1 $X=42095 $Y=101405 $D=9
M275 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30 mult=1 $X=42095 $Y=109900 $D=9
M276 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30 mult=1 $X=42095 $Y=118725 $D=9
M277 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90016.2 a=1.26 p=14.36 mult=1 $X=50370 $Y=26860 $D=9
M278 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90016.2 a=1.26 p=14.36 mult=1 $X=50370 $Y=36860 $D=9
M279 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90016.2 a=1.26 p=14.36 mult=1 $X=50370 $Y=46860 $D=9
M280 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90016.2 a=1.26 p=14.36 mult=1 $X=50370 $Y=56860 $D=9
M281 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90016.1 a=0.9 p=10.36 mult=1 $X=50370 $Y=66860 $D=9
M282 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90016.2 a=1.26 p=14.36 mult=1 $X=50370 $Y=176860 $D=9
M283 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90016.2 a=1.26 p=14.36 mult=1 $X=50370 $Y=186860 $D=9
M284 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 r=27.7778 sa=90019.9 sb=90015.6 a=0.9 p=10.36 mult=1 $X=50895 $Y=128755 $D=9
M285 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90015.6 a=1.26 p=14.36 mult=1 $X=50895 $Y=136860 $D=9
M286 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90015.6 a=1.26 p=14.36 mult=1 $X=50895 $Y=146860 $D=9
M287 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90015.6 a=1.26 p=14.36 mult=1 $X=50895 $Y=156860 $D=9
M288 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90015.6 a=1.26 p=14.36 mult=1 $X=50895 $Y=166860 $D=9
M289 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90015 a=1.26 p=14.36 mult=1 $X=51560 $Y=26860 $D=9
M290 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90015 a=1.26 p=14.36 mult=1 $X=51560 $Y=36860 $D=9
M291 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90015 a=1.26 p=14.36 mult=1 $X=51560 $Y=46860 $D=9
M292 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90015 a=1.26 p=14.36 mult=1 $X=51560 $Y=56860 $D=9
M293 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90015 a=0.9 p=10.36 mult=1 $X=51560 $Y=66860 $D=9
M294 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90015 a=1.26 p=14.36 mult=1 $X=51560 $Y=176860 $D=9
M295 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90015 a=1.26 p=14.36 mult=1 $X=51560 $Y=186860 $D=9
M296 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 r=27.7778 sa=90019.9 sb=90014.3 a=0.9 p=10.36 mult=1 $X=52245 $Y=128755 $D=9
M297 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90014.3 a=1.26 p=14.36 mult=1 $X=52245 $Y=136860 $D=9
M298 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90014.3 a=1.26 p=14.36 mult=1 $X=52245 $Y=146860 $D=9
M299 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90014.3 a=1.26 p=14.36 mult=1 $X=52245 $Y=156860 $D=9
M300 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90014.3 a=1.26 p=14.36 mult=1 $X=52245 $Y=166860 $D=9
M301 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90013.4 a=1.26 p=14.36 mult=1 $X=53140 $Y=26860 $D=9
M302 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90013.4 a=1.26 p=14.36 mult=1 $X=53140 $Y=36860 $D=9
M303 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90013.4 a=1.26 p=14.36 mult=1 $X=53140 $Y=46860 $D=9
M304 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90013.4 a=1.26 p=14.36 mult=1 $X=53140 $Y=56860 $D=9
M305 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90013.4 a=0.9 p=10.36 mult=1 $X=53140 $Y=66860 $D=9
M306 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90013.4 a=1.26 p=14.36 mult=1 $X=53140 $Y=176860 $D=9
M307 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90013.4 a=1.26 p=14.36 mult=1 $X=53140 $Y=186860 $D=9
M308 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90012.2 a=1.26 p=14.36 mult=1 $X=54330 $Y=26860 $D=9
M309 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90012.2 a=1.26 p=14.36 mult=1 $X=54330 $Y=36860 $D=9
M310 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90012.2 a=1.26 p=14.36 mult=1 $X=54330 $Y=46860 $D=9
M311 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90012.2 a=1.26 p=14.36 mult=1 $X=54330 $Y=56860 $D=9
M312 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90012.2 a=0.9 p=10.36 mult=1 $X=54330 $Y=66860 $D=9
M313 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90012.2 a=1.26 p=14.36 mult=1 $X=54330 $Y=176860 $D=9
M314 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90012.2 a=1.26 p=14.36 mult=1 $X=54330 $Y=186860 $D=9
M315 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 r=27.7778 sa=90019.9 sb=90011.4 a=0.9 p=10.36 mult=1 $X=55075 $Y=128755 $D=9
M316 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90011.4 a=1.26 p=14.36 mult=1 $X=55075 $Y=136860 $D=9
M317 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90011.4 a=1.26 p=14.36 mult=1 $X=55075 $Y=146860 $D=9
M318 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90011.4 a=1.26 p=14.36 mult=1 $X=55075 $Y=156860 $D=9
M319 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90011.4 a=1.26 p=14.36 mult=1 $X=55075 $Y=166860 $D=9
M320 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90010.6 a=1.26 p=14.36 mult=1 $X=55910 $Y=26860 $D=9
M321 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90010.6 a=1.26 p=14.36 mult=1 $X=55910 $Y=36860 $D=9
M322 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90010.6 a=1.26 p=14.36 mult=1 $X=55910 $Y=46860 $D=9
M323 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90010.6 a=1.26 p=14.36 mult=1 $X=55910 $Y=56860 $D=9
M324 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90010.6 a=0.9 p=10.36 mult=1 $X=55910 $Y=66860 $D=9
M325 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90010.6 a=1.26 p=14.36 mult=1 $X=55910 $Y=176860 $D=9
M326 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90010.6 a=1.26 p=14.36 mult=1 $X=55910 $Y=186860 $D=9
M327 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 r=27.7778 sa=90019.9 sb=90010.1 a=0.9 p=10.36 mult=1 $X=56425 $Y=128755 $D=9
M328 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90010.1 a=1.26 p=14.36 mult=1 $X=56425 $Y=136860 $D=9
M329 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90010.1 a=1.26 p=14.36 mult=1 $X=56425 $Y=146860 $D=9
M330 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90010.1 a=1.26 p=14.36 mult=1 $X=56425 $Y=156860 $D=9
M331 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90010.1 a=1.26 p=14.36 mult=1 $X=56425 $Y=166860 $D=9
M332 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90009.4 a=1.26 p=14.36 mult=1 $X=57100 $Y=26860 $D=9
M333 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90009.4 a=1.26 p=14.36 mult=1 $X=57100 $Y=36860 $D=9
M334 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90009.4 a=1.26 p=14.36 mult=1 $X=57100 $Y=46860 $D=9
M335 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90009.4 a=1.26 p=14.36 mult=1 $X=57100 $Y=56860 $D=9
M336 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90009.4 a=0.9 p=10.36 mult=1 $X=57100 $Y=66860 $D=9
M337 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90009.4 a=1.26 p=14.36 mult=1 $X=57100 $Y=176860 $D=9
M338 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90009.4 a=1.26 p=14.36 mult=1 $X=57100 $Y=186860 $D=9
M339 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=0.625 sa=4.00002e+06 sb=4e+06 a=40 p=26 mult=1 $X=50375 $Y=75805 $D=9
M340 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00002e+06 sb=4e+06 a=56 p=30 mult=1 $X=50375 $Y=82805 $D=9
M341 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00002e+06 sb=4e+06 a=56 p=30 mult=1 $X=50375 $Y=91300 $D=9
M342 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00002e+06 sb=4e+06 a=56 p=30 mult=1 $X=50375 $Y=101405 $D=9
M343 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00002e+06 sb=4e+06 a=56 p=30 mult=1 $X=50375 $Y=109900 $D=9
M344 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00002e+06 sb=4e+06 a=56 p=30 mult=1 $X=50375 $Y=118725 $D=9
M345 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90007.8 a=1.26 p=14.36 mult=1 $X=58680 $Y=26860 $D=9
M346 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90007.8 a=1.26 p=14.36 mult=1 $X=58680 $Y=36860 $D=9
M347 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90007.8 a=1.26 p=14.36 mult=1 $X=58680 $Y=46860 $D=9
M348 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90007.8 a=1.26 p=14.36 mult=1 $X=58680 $Y=56860 $D=9
M349 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90007.8 a=0.9 p=10.36 mult=1 $X=58680 $Y=66860 $D=9
M350 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90007.8 a=1.26 p=14.36 mult=1 $X=58680 $Y=176860 $D=9
M351 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90007.8 a=1.26 p=14.36 mult=1 $X=58680 $Y=186860 $D=9
M352 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 r=27.7778 sa=90019.9 sb=90007.3 a=0.9 p=10.36 mult=1 $X=59255 $Y=128755 $D=9
M353 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90007.3 a=1.26 p=14.36 mult=1 $X=59255 $Y=136860 $D=9
M354 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90007.3 a=1.26 p=14.36 mult=1 $X=59255 $Y=146860 $D=9
M355 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90007.3 a=1.26 p=14.36 mult=1 $X=59255 $Y=156860 $D=9
M356 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90007.3 a=1.26 p=14.36 mult=1 $X=59255 $Y=166860 $D=9
M357 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90006.6 a=1.26 p=14.36 mult=1 $X=59870 $Y=26860 $D=9
M358 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90006.6 a=1.26 p=14.36 mult=1 $X=59870 $Y=36860 $D=9
M359 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90006.6 a=1.26 p=14.36 mult=1 $X=59870 $Y=46860 $D=9
M360 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90006.6 a=1.26 p=14.36 mult=1 $X=59870 $Y=56860 $D=9
M361 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90006.6 a=0.9 p=10.36 mult=1 $X=59870 $Y=66860 $D=9
M362 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90006.6 a=1.26 p=14.36 mult=1 $X=59870 $Y=176860 $D=9
M363 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90006.6 a=1.26 p=14.36 mult=1 $X=59870 $Y=186860 $D=9
M364 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 r=27.7778 sa=90019.9 sb=90005.9 a=0.9 p=10.36 mult=1 $X=60605 $Y=128755 $D=9
M365 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90005.9 a=1.26 p=14.36 mult=1 $X=60605 $Y=136860 $D=9
M366 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90005.9 a=1.26 p=14.36 mult=1 $X=60605 $Y=146860 $D=9
M367 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90005.9 a=1.26 p=14.36 mult=1 $X=60605 $Y=156860 $D=9
M368 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90005.9 a=1.26 p=14.36 mult=1 $X=60605 $Y=166860 $D=9
M369 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90005.1 a=1.26 p=14.36 mult=1 $X=61450 $Y=26860 $D=9
M370 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90005.1 a=1.26 p=14.36 mult=1 $X=61450 $Y=36860 $D=9
M371 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90005.1 a=1.26 p=14.36 mult=1 $X=61450 $Y=46860 $D=9
M372 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90005.1 a=1.26 p=14.36 mult=1 $X=61450 $Y=56860 $D=9
M373 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90005.1 a=0.9 p=10.36 mult=1 $X=61450 $Y=66860 $D=9
M374 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90005.1 a=1.26 p=14.36 mult=1 $X=61450 $Y=176860 $D=9
M375 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90005.1 a=1.26 p=14.36 mult=1 $X=61450 $Y=186860 $D=9
M376 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90003.9 a=1.26 p=14.36 mult=1 $X=62640 $Y=26860 $D=9
M377 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90003.9 a=1.26 p=14.36 mult=1 $X=62640 $Y=36860 $D=9
M378 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90003.9 a=1.26 p=14.36 mult=1 $X=62640 $Y=46860 $D=9
M379 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90003.9 a=1.26 p=14.36 mult=1 $X=62640 $Y=56860 $D=9
M380 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90003.9 a=0.9 p=10.36 mult=1 $X=62640 $Y=66860 $D=9
M381 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90003.9 a=1.26 p=14.36 mult=1 $X=62640 $Y=176860 $D=9
M382 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90003.9 a=1.26 p=14.36 mult=1 $X=62640 $Y=186860 $D=9
M383 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 r=27.7778 sa=90019.9 sb=90003.1 a=0.9 p=10.36 mult=1 $X=63435 $Y=128755 $D=9
M384 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90003.1 a=1.26 p=14.36 mult=1 $X=63435 $Y=136860 $D=9
M385 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90003.1 a=1.26 p=14.36 mult=1 $X=63435 $Y=146860 $D=9
M386 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90003.1 a=1.26 p=14.36 mult=1 $X=63435 $Y=156860 $D=9
M387 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 r=38.8889 sa=90019.9 sb=90003.1 a=1.26 p=14.36 mult=1 $X=63435 $Y=166860 $D=9
M388 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90002.3 a=1.26 p=14.36 mult=1 $X=64220 $Y=26860 $D=9
M389 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90002.3 a=1.26 p=14.36 mult=1 $X=64220 $Y=36860 $D=9
M390 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90002.3 a=1.26 p=14.36 mult=1 $X=64220 $Y=46860 $D=9
M391 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90002.3 a=1.26 p=14.36 mult=1 $X=64220 $Y=56860 $D=9
M392 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 r=27.7778 sa=90019.9 sb=90002.3 a=0.9 p=10.36 mult=1 $X=64220 $Y=66860 $D=9
M393 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90002.3 a=1.26 p=14.36 mult=1 $X=64220 $Y=176860 $D=9
M394 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 r=38.8889 sa=90019.9 sb=90002.3 a=1.26 p=14.36 mult=1 $X=64220 $Y=186860 $D=9
M395 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 r=27.7778 sa=90019.9 sb=90001.7 a=0.9 p=10.36 mult=1 $X=64785 $Y=128755 $D=9
M396 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90001.7 a=1.26 p=14.36 mult=1 $X=64785 $Y=136860 $D=9
M397 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90001.7 a=1.26 p=14.36 mult=1 $X=64785 $Y=146860 $D=9
M398 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90001.7 a=1.26 p=14.36 mult=1 $X=64785 $Y=156860 $D=9
M399 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 r=38.8889 sa=90019.9 sb=90001.7 a=1.26 p=14.36 mult=1 $X=64785 $Y=166860 $D=9
M400 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90001.1 a=1.26 p=14.36 mult=1 $X=65410 $Y=26860 $D=9
M401 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90001.1 a=1.26 p=14.36 mult=1 $X=65410 $Y=36860 $D=9
M402 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90001.1 a=1.26 p=14.36 mult=1 $X=65410 $Y=46860 $D=9
M403 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90001.1 a=1.26 p=14.36 mult=1 $X=65410 $Y=56860 $D=9
M404 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 nshort L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 r=27.7778 sa=90019.9 sb=90001.1 a=0.9 p=10.36 mult=1 $X=65410 $Y=66860 $D=9
M405 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90001.1 a=1.26 p=14.36 mult=1 $X=65410 $Y=176860 $D=9
M406 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 nshort L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 r=38.8889 sa=90019.9 sb=90001.1 a=1.26 p=14.36 mult=1 $X=65410 $Y=186860 $D=9
M407 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 r=0.625 sa=4.00002e+06 sb=4e+06 a=40 p=26 mult=1 $X=58655 $Y=75805 $D=9
M408 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00002e+06 sb=4e+06 a=56 p=30 mult=1 $X=58655 $Y=82805 $D=9
M409 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 nshort L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00002e+06 sb=4e+06 a=56 p=30 mult=1 $X=58655 $Y=91300 $D=9
M410 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00002e+06 sb=4e+06 a=56 p=30 mult=1 $X=58655 $Y=101405 $D=9
M411 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00002e+06 sb=4e+06 a=56 p=30 mult=1 $X=58655 $Y=109900 $D=9
M412 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 nshort L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 r=0.875 sa=4.00002e+06 sb=4e+06 a=56 p=30 mult=1 $X=58655 $Y=118725 $D=9
X413 SRC_BDY_LVC1 VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=40185 $Y=114790 $D=150
X414 SRC_BDY_LVC2 VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=40605 $Y=34930 $D=150
X415 SRC_BDY_LVC1 VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=40640 $Y=196080 $D=150
X416 VSSD DRN_LVC1 Dpar a=108.41 p=46.58 m=1 $[nwdiode] $X=1015 $Y=685 $D=191
X417 VSSD DRN_LVC2 Dpar a=108.41 p=46.58 m=1 $[nwdiode] $X=67280 $Y=745 $D=191
X418 VSSD VDDIO Dpar a=10516.3 p=468.87 m=1 $[dnwdiode_psub] $X=9500 $Y=23605 $D=193
X419 SRC_BDY_LVC2 VDDIO Dpar a=4115.42 p=264.63 m=1 $[dnwdiode_pw] $X=10870 $Y=24975 $D=194
X420 SRC_BDY_LVC1 VDDIO Dpar a=5703.29 p=340.89 m=1 $[dnwdiode_pw] $X=10870 $Y=83485 $D=194
R421 DRN_LVC1 21 L=1950 W=0.33 m=1 mult=1 model="mrp1" $[mrp1] $X=240 $Y=19200 $D=257
R422 G_CORE G_PAD 0.01 m=1 $[short] $X=6670 $Y=103345 $D=286
X423 27 DRN_LVC2 sky130_fd_pr__res_bent_po__example_55959141808692 $T=70965 18130 0 90 $X=70615 $Y=17860
X424 DRN_LVC1 21 24 sky130_fd_pr__pfet_01v8__example_55959141808687 $T=2070 2020 0 0 $X=1610 $Y=1840
X425 DRN_LVC1 21 24 sky130_fd_pr__pfet_01v8__example_55959141808687 $T=2070 9670 0 0 $X=1610 $Y=9490
X426 DRN_LVC2 23 25 sky130_fd_pr__pfet_01v8__example_55959141808687 $T=68335 2080 0 0 $X=67875 $Y=1900
X427 DRN_LVC2 23 25 sky130_fd_pr__pfet_01v8__example_55959141808687 $T=68335 9730 0 0 $X=67875 $Y=9550
X616 23 26 sky130_fd_pr__res_bent_po__example_55959141808691 $T=66785 1745 1 90 $X=57045 $Y=1475
X622 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808704 $T=25815 136860 0 0 $X=23860 $Y=136700
X623 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808695 $T=25815 128755 0 0 $X=23860 $Y=128595
X630 VSSD BDY2_B2B SRC_BDY_LVC1 sky130_fd_io__gnd2gnd_120x2_lv_isosub $T=16525 18480 1 0 $X=16525 $Y=320
X631 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808701 $T=17130 176860 0 0 $X=15800 $Y=176700
X632 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808703 $T=17455 146860 0 0 $X=15500 $Y=146700
X633 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808703 $T=17455 156860 0 0 $X=15500 $Y=156700
X634 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808703 $T=17455 166860 0 0 $X=15500 $Y=166700
X635 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705 $T=14360 26860 0 0 $X=13030 $Y=26700
X636 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705 $T=14360 36860 0 0 $X=13030 $Y=36700
X637 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705 $T=14360 46860 0 0 $X=13030 $Y=46700
X638 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705 $T=14360 56860 0 0 $X=13030 $Y=56700
X639 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808705 $T=14360 186860 0 0 $X=13030 $Y=186700
X640 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808693 $T=14360 66860 0 0 $X=13030 $Y=66700
X642 22 26 sky130_fd_pr__res_bent_po__example_55959141808688 $T=11245 84330 0 90 $X=10895 $Y=84060
X643 27 22 sky130_fd_pr__res_bent_po__example_55959141808690 $T=69775 19510 0 180 $X=10025 $Y=19160
.ENDS
***************************************
.SUBCKT sky130_ef_io__vssd_lvc_clamped2_pad VSSD VSSA VSSIO VCCD VDDIO VSSD_PAD
** N=13 EP=6 IP=20 FDC=501
*.CALIBRE ISOLATED NETS: VCCHIB VDDA VSWITCH AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
X0 VSSD VSSD VSSIO VCCD VDDIO VCCD VSSA VSSD VSSD_PAD sky130_fd_io__top_ground_lvc_wpad $T=0 -35 0 0 $X=0 $Y=-35
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3 6 7 8 9 12 13 14 15 16
** N=17 EP=12 IP=52 FDC=1484
X0 1 9 6 8 15 sky130_ef_io__vdda_hvc_clamped_pad $T=197965 2415000 0 90 $X=0 $Y=2415000
X1 1 7 6 2 17 sky130_ef_io__vdda_hvc_clamped_pad $T=3390035 2594000 0 270 $X=3388000 $Y=2519000
X2 1 9 3 12 6 14 sky130_ef_io__vssd_lvc_clamped2_pad $T=197965 2204000 0 90 $X=0 $Y=2204000
X3 1 7 3 13 6 16 sky130_ef_io__vssd_lvc_clamped2_pad $T=3390035 2374000 0 270 $X=3379500 $Y=2287805
.ENDS
***************************************
.SUBCKT ICV_17 1 68 132 176 233 241
** N=329 EP=6 IP=25 FDC=482
X0 1 176 132 233 329 sky130_ef_io__vssa_hvc_clamped_pad $T=3390035 2153000 0 270 $X=3388000 $Y=2078000
X1 1 68 176 241 sky130_ef_io__vddio_hvc_clamped_pad $T=197965 551000 0 90 $X=0 $Y=551000
.ENDS
***************************************
.SUBCKT ICV_18 1 3 8 26 30 42 43
** N=88 EP=7 IP=38 FDC=723
X0 1 8 3 88 sky130_ef_io__vssio_hvc_clamped_pad $T=2920000 197965 0 180 $X=2845000 $Y=0
X1 1 8 26 30 42 sky130_ef_io__vssa_hvc_clamped_pad $T=469000 197965 0 180 $X=394000 $Y=0
X2 1 26 8 30 43 sky130_ef_io__vdda_hvc_clamped_pad $T=3189000 197965 0 180 $X=3114000 $Y=0
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em2o_cdns_55959141808653 2 3
** N=7 EP=2 IP=0 FDC=2
R0 2 6 0.01 m=1 $[short] $X=260 $Y=0 $D=283
R1 7 3 0.01 m=1 $[short] $X=1770 $Y=0 $D=283
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd2__example_55959141808202
** N=17 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808657
** N=5 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em2s_cdns_55959141808652 2 3
** N=6 EP=2 IP=0 FDC=2
R0 2 6 0.01 m=1 $[short] $X=260 $Y=0 $D=283
R1 6 3 0.01 m=1 $[short] $X=1770 $Y=0 $D=283
.ENDS
***************************************
.SUBCKT ICV_19
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_generic_po__example_5595914180838 2 3
** N=6 EP=2 IP=0 FDC=1
R0 2 3 L=10.2 W=0.5 m=1 mult=1 model="mrp1" $[mrp1] $X=0 $Y=0 $D=257
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_generic_po__example_5595914180864 2 3
** N=8 EP=2 IP=0 FDC=1
R0 2 3 L=1.5 W=0.8 m=1 mult=1 model="mrp1" $[mrp1] $X=0 $Y=0 $D=257
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em1s_cdns_5595914180859 2 3
** N=6 EP=2 IP=0 FDC=2
R0 2 6 0.01 m=1 $[short] $X=260 $Y=0 $D=282
R1 6 3 0.01 m=1 $[short] $X=1770 $Y=0 $D=282
.ENDS
***************************************
.SUBCKT sky130_fd_io__res250only_small PAD ROUT
** N=32 EP=2 IP=0 FDC=7
R0 PAD 6 L=0.17 W=2 m=1 mult=1 model="mrp1" $[mrp1] $X=300 $Y=10 $D=257
R1 6 7 L=10.07 W=2 m=1 mult=1 model="mrp1" $[mrp1] $X=640 $Y=10 $D=257
R2 7 ROUT L=0.17 W=2 m=1 mult=1 model="mrp1" $[mrp1] $X=10880 $Y=10 $D=257
R3 PAD 6 0.01 m=1 $[short] $X=380 $Y=0 $D=281
R4 7 ROUT 0.01 m=1 $[short] $X=10960 $Y=0 $D=281
R5 PAD 6 0.01 m=1 $[short] $X=380 $Y=5 $D=282
R6 7 ROUT 0.01 m=1 $[short] $X=10960 $Y=5 $D=282
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_5595914180862 2 3
** N=8 EP=2 IP=0 FDC=1
R0 2 3 L=6 W=0.8 m=1 mult=1 model="mrp1" $[mrp1] $X=0 $Y=0 $D=257
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_5595914180863 2 3
** N=8 EP=2 IP=0 FDC=1
R0 2 3 L=12 W=0.8 m=1 mult=1 model="mrp1" $[mrp1] $X=0 $Y=0 $D=257
.ENDS
***************************************
.SUBCKT sky130_fd_pr__model__pfet_highvoltage__example_55959141808616
** N=39 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_io__hvsbt_inv_x4
** N=74 EP=0 IP=44 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: IN OUT
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 2 3
** N=7 EP=2 IP=0 FDC=2
R0 2 6 0.01 m=1 $[short] $X=130 $Y=0 $D=282
R1 7 3 0.01 m=1 $[short] $X=280 $Y=0 $D=282
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_p_em1c_cdns_55959141808753 2
** N=6 EP=1 IP=0 FDC=2
R0 2 5 0.01 m=1 $[short] $X=160 $Y=0 $D=282
R1 2 6 0.01 m=1 $[short] $X=160 $Y=250 $D=282
.ENDS
***************************************
.SUBCKT ICV_20 2 3
** N=7 EP=2 IP=9 FDC=4
X0 2 3 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=0 0 0 0 $X=0 $Y=0
X1 2 sky130_fd_io__xres_p_em1c_cdns_55959141808753 $T=-10 -770 0 0 $X=-10 $Y=-770
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_generic_nd__example_55959141808754 2 3
** N=5 EP=2 IP=0 FDC=1
*.SEEDPROM
R0 2 3 L=14 W=0.5 m=1 $[mrdn] $X=0 $Y=0 $D=253
.ENDS
***************************************
.SUBCKT ICV_21 2 3 4 5
** N=9 EP=4 IP=10 FDC=2
*.SEEDPROM
X0 2 3 sky130_fd_pr__res_generic_nd__example_55959141808754 $T=14000 -770 1 180 $X=-340 $Y=-900
X1 4 5 sky130_fd_pr__res_generic_nd__example_55959141808754 $T=0 0 0 0 $X=-340 $Y=-130
.ENDS
***************************************
.SUBCKT ICV_22 2 3 4 5 6 7 8 9
** N=17 EP=8 IP=18 FDC=4
*.SEEDPROM
X0 4 2 3 5 ICV_21 $T=0 -1540 0 0 $X=-340 $Y=-2440
X1 8 6 7 9 ICV_21 $T=0 0 0 0 $X=-340 $Y=-900
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758 2 3
** N=7 EP=2 IP=0 FDC=2
R0 2 6 0.01 m=1 $[short] $X=130 $Y=0 $D=282
R1 7 3 0.01 m=1 $[short] $X=280 $Y=0 $D=282
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1c_cdns_55959141808760 2
** N=6 EP=1 IP=0 FDC=2
R0 2 5 0.01 m=1 $[short] $X=160 $Y=0 $D=282
R1 2 6 0.01 m=1 $[short] $X=160 $Y=640 $D=282
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1c_cdns_55959141808761 2
** N=6 EP=1 IP=0 FDC=2
R0 2 5 0.01 m=1 $[short] $X=160 $Y=0 $D=282
R1 2 6 0.01 m=1 $[short] $X=160 $Y=250 $D=282
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd__example_55959141808338
** N=22 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd2__example_55959141808337
** N=22 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__via_pol1__example_55959141808273
** N=13 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_23
** N=3 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_24
** N=5 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759 1
** N=5 EP=1 IP=0 FDC=2
R0 1 4 0.01 m=1 $[short] $X=160 $Y=0 $D=282
R1 1 5 0.01 m=1 $[short] $X=160 $Y=280 $D=282
.ENDS
***************************************
.SUBCKT ICV_25 2 3 4
** N=8 EP=3 IP=9 FDC=4
X0 2 3 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=0 0 0 0 $X=0 $Y=0
X1 4 sky130_fd_io__xres_p_em1c_cdns_55959141808753 $T=-10 770 0 0 $X=-10 $Y=770
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1o_cdns_55959141808756 1 2
** N=6 EP=2 IP=0 FDC=2
R0 2 5 0.01 m=1 $[short] $X=130 $Y=0 $D=282
R1 6 1 0.01 m=1 $[short] $X=280 $Y=0 $D=282
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_generic_nd__example_55959141808755 2 3
** N=5 EP=2 IP=0 FDC=1
*.SEEDPROM
R0 2 3 L=47 W=0.5 m=1 $[mrdn] $X=0 $Y=0 $D=253
.ENDS
***************************************
.SUBCKT ICV_26 2 3 4
** N=8 EP=3 IP=10 FDC=2
*.SEEDPROM
X0 2 3 sky130_fd_pr__res_generic_nd__example_55959141808754 $T=0 0 0 0 $X=-340 $Y=-130
X1 4 2 sky130_fd_pr__res_generic_nd__example_55959141808755 $T=-47510 0 0 0 $X=-47850 $Y=-130
.ENDS
***************************************
.SUBCKT ICV_27 2 3
** N=7 EP=2 IP=10 FDC=2
*.SEEDPROM
X0 2 2 sky130_fd_pr__res_generic_nd__example_55959141808754 $T=0 0 0 0 $X=-340 $Y=-130
X1 2 3 sky130_fd_pr__res_generic_nd__example_55959141808755 $T=14510 0 0 0 $X=14170 $Y=-130
.ENDS
***************************************
.SUBCKT ICV_28 2 3 4 5 6
** N=14 EP=5 IP=15 FDC=4
*.SEEDPROM
X0 3 4 2 ICV_26 $T=0 0 0 0 $X=-47850 $Y=-130
X1 5 6 ICV_27 $T=14000 770 1 180 $X=-47850 $Y=640
.ENDS
***************************************
.SUBCKT ICV_29 2 3 4 5 6 7 8 9 10 11
** N=27 EP=10 IP=28 FDC=8
*.SEEDPROM
X0 2 4 6 5 3 ICV_28 $T=0 0 0 0 $X=-47850 $Y=-130
X1 7 9 11 10 8 ICV_28 $T=0 1540 0 0 $X=-47850 $Y=1410
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres2v2_rcfilter_lpfv2 1 VCC_IO 3 4 5 6 7 8 9 10 11 12 13 IN
** N=5580 EP=14 IP=654 FDC=361
M0 1 3 1 1 nhv L=4 W=7 AD=0.98 AS=1.855 PD=7.28 PS=14.53 NRD=0 NRS=0 m=1 r=1.75 sa=2e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=2725 $Y=11605 $D=49
M1 1 4 1 1 nhv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=7005 $Y=11605 $D=49
M2 1 5 1 1 nhv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00001e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=11285 $Y=11605 $D=49
M3 1 6 1 1 nhv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00001e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=15565 $Y=11605 $D=49
M4 1 7 1 1 nhv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=19845 $Y=11605 $D=49
M5 1 8 1 1 nhv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=24125 $Y=11605 $D=49
M6 1 9 1 1 nhv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=28405 $Y=11605 $D=49
M7 1 10 1 1 nhv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=32685 $Y=11605 $D=49
M8 1 11 1 1 nhv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00001e+06 a=28 p=22 mult=1 $X=36965 $Y=11605 $D=49
M9 1 11 1 1 nhv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00001e+06 a=28 p=22 mult=1 $X=41245 $Y=11605 $D=49
M10 1 12 1 1 nhv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2e+06 a=28 p=22 mult=1 $X=45525 $Y=11605 $D=49
M11 1 13 1 1 nhv L=4 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2e+06 a=28 p=22 mult=1 $X=49805 $Y=11605 $D=49
M12 VCC_IO 3 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=1.855 PD=7.28 PS=14.53 NRD=0 NRS=0 m=1 r=1.75 sa=2e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=2625 $Y=21435 $D=109
M13 VCC_IO 4 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=6905 $Y=21435 $D=109
M14 VCC_IO 5 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00001e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=11185 $Y=21435 $D=109
M15 VCC_IO 6 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00001e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=15465 $Y=21435 $D=109
M16 VCC_IO 7 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=19745 $Y=21435 $D=109
M17 VCC_IO 8 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=24025 $Y=21435 $D=109
M18 VCC_IO 9 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=28305 $Y=21435 $D=109
M19 VCC_IO 10 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=32585 $Y=21435 $D=109
M20 VCC_IO 11 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00001e+06 a=28 p=22 mult=1 $X=36865 $Y=21435 $D=109
M21 VCC_IO 11 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00001e+06 a=28 p=22 mult=1 $X=41145 $Y=21435 $D=109
M22 VCC_IO 12 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2e+06 a=28 p=22 mult=1 $X=45425 $Y=21435 $D=109
M23 VCC_IO 13 VCC_IO VCC_IO phv L=4 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2e+06 a=28 p=22 mult=1 $X=49705 $Y=21435 $D=109
X24 1 8 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=815 $D=181
X25 1 7 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=2355 $D=181
X26 1 6 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=3895 $D=181
X27 1 5 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=5435 $D=181
X28 1 4 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=6975 $D=181
X29 1 3 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=8515 $D=181
X30 1 15 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=31330 $D=181
X31 1 16 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=32870 $D=181
X32 1 17 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=34410 $D=181
X33 1 18 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=35950 $D=181
X34 1 19 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=37490 $D=181
X35 1 20 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=39030 $D=181
X36 1 1 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=1585 $D=181
X37 1 1 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=3125 $D=181
X38 1 1 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=4665 $D=181
X39 1 1 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=6205 $D=181
X40 1 3 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=7745 $D=181
X41 1 9 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=9285 $D=181
X42 1 15 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=30560 $D=181
X43 1 16 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=32100 $D=181
X44 1 17 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=33640 $D=181
X45 1 18 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=35180 $D=181
X46 1 19 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=36720 $D=181
X47 1 20 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=38260 $D=181
X48 1 21 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=815 $D=181
X49 1 22 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=2355 $D=181
X50 1 23 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=3895 $D=181
X51 1 24 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=5435 $D=181
X52 1 25 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=6975 $D=181
X53 1 26 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=8515 $D=181
X54 1 27 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=31330 $D=181
X55 1 28 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=32870 $D=181
X56 1 29 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=34410 $D=181
X57 1 30 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=35950 $D=181
X58 1 31 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=37490 $D=181
X59 1 32 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=39030 $D=181
X60 1 1 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=1585 $D=181
X61 1 1 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=3125 $D=181
X62 1 1 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=4665 $D=181
X63 1 1 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=6205 $D=181
X64 1 3 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=7745 $D=181
X65 1 9 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=9285 $D=181
X66 1 15 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=30560 $D=181
X67 1 16 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=32100 $D=181
X68 1 17 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=33640 $D=181
X69 1 18 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=35180 $D=181
X70 1 19 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=36720 $D=181
X71 1 20 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=38260 $D=181
X72 1 38 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=815 $D=181
X73 1 39 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=1585 $D=181
X74 1 37 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=2355 $D=181
X75 1 40 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=3125 $D=181
X76 1 36 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=3895 $D=181
X77 1 41 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=4665 $D=181
X78 1 35 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=5435 $D=181
X79 1 42 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=6205 $D=181
X80 1 34 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=6975 $D=181
X81 1 43 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=7745 $D=181
X82 1 33 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=8515 $D=181
X83 1 44 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=9285 $D=181
X84 1 45 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=30560 $D=181
X85 1 10 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=31330 $D=181
X86 1 46 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=32100 $D=181
X87 1 11 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=32870 $D=181
X88 1 47 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=33640 $D=181
X89 1 11 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=34410 $D=181
X90 1 48 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=35180 $D=181
X91 1 12 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=35950 $D=181
X92 1 49 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=36720 $D=181
X93 1 13 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=37490 $D=181
X94 1 50 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=38260 $D=181
X95 1 IN Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=39030 $D=181
X96 1 33 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=10735 $D=181
X97 1 34 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=12275 $D=181
X98 1 35 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=13815 $D=181
X99 1 36 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=15355 $D=181
X100 1 37 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=16895 $D=181
X101 1 38 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=18435 $D=181
X102 1 13 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=21405 $D=181
X103 1 12 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=22945 $D=181
X104 1 11 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=24485 $D=181
X105 1 11 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=26025 $D=181
X106 1 10 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=27565 $D=181
X107 1 9 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=29105 $D=181
X108 1 33 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=11505 $D=181
X109 1 34 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=13045 $D=181
X110 1 35 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=14585 $D=181
X111 1 36 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=16125 $D=181
X112 1 37 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=17665 $D=181
X113 1 38 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=19205 $D=181
X114 1 IN Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=20635 $D=181
X115 1 13 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=22175 $D=181
X116 1 12 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=23715 $D=181
X117 1 11 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=25255 $D=181
X118 1 11 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=26795 $D=181
X119 1 10 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=28335 $D=181
X120 1 44 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=10735 $D=181
X121 1 33 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=11505 $D=181
X122 1 43 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=12275 $D=181
X123 1 34 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=13045 $D=181
X124 1 42 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=13815 $D=181
X125 1 35 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=14585 $D=181
X126 1 41 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=15355 $D=181
X127 1 36 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=16125 $D=181
X128 1 40 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=16895 $D=181
X129 1 37 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=17665 $D=181
X130 1 39 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=18435 $D=181
X131 1 38 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=19205 $D=181
X132 1 IN Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=20635 $D=181
X133 1 50 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=21405 $D=181
X134 1 13 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=22175 $D=181
X135 1 49 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=22945 $D=181
X136 1 12 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=23715 $D=181
X137 1 48 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=24485 $D=181
X138 1 11 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=25255 $D=181
X139 1 47 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=26025 $D=181
X140 1 11 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=26795 $D=181
X141 1 46 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=27565 $D=181
X142 1 10 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=28335 $D=181
X143 1 45 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=29105 $D=181
X144 1 VCC_IO Dpar a=501.44 p=125.96 m=1 $[nwdiode] $X=1350 $Y=20095 $D=191
X164 20 32 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=16535 39150 0 0 $X=16535 $Y=39150
X165 8 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=54510 935 0 0 $X=54510 $Y=935
X166 7 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=54510 2475 0 0 $X=54510 $Y=2475
X167 6 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=54510 4015 0 0 $X=54510 $Y=4015
X168 5 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=54510 5555 0 0 $X=54510 $Y=5555
X169 3 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=54510 8635 0 0 $X=54510 $Y=8635
X170 9 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=71780 29485 0 180 $X=71360 $Y=29225
X171 12 49 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=72265 23325 1 0 $X=72265 $Y=23065
X172 11 47 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=72265 26405 1 0 $X=72265 $Y=26145
X173 9 45 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=72265 29485 1 0 $X=72265 $Y=29225
X174 15 sky130_fd_io__xres_p_em1c_cdns_55959141808753 $T=16525 30680 0 0 $X=16525 $Y=30680
X175 IN sky130_fd_io__xres_p_em1c_cdns_55959141808753 $T=72255 21015 1 0 $X=72255 $Y=20755
X176 12 sky130_fd_io__xres_p_em1c_cdns_55959141808753 $T=72255 24095 1 0 $X=72255 $Y=23835
X177 11 sky130_fd_io__xres_p_em1c_cdns_55959141808753 $T=72255 27175 1 0 $X=72255 $Y=26915
X178 33 44 ICV_20 $T=72265 11115 1 0 $X=72255 $Y=10855
X179 34 43 ICV_20 $T=72265 12655 1 0 $X=72255 $Y=12395
X180 35 42 ICV_20 $T=72265 14195 1 0 $X=72255 $Y=13935
X181 36 41 ICV_20 $T=72265 15735 1 0 $X=72255 $Y=15475
X182 37 40 ICV_20 $T=72265 17275 1 0 $X=72255 $Y=17015
X183 38 39 ICV_20 $T=72265 18815 1 0 $X=72255 $Y=18555
X184 13 50 ICV_20 $T=72265 21785 1 0 $X=72255 $Y=21525
X185 11 48 ICV_20 $T=72265 24865 1 0 $X=72255 $Y=24605
X186 10 46 ICV_20 $T=72265 27945 1 0 $X=72255 $Y=27685
X187 34 43 34 34 33 44 33 33 ICV_22 $T=72640 11235 0 180 $X=58300 $Y=10605
X188 36 41 36 36 35 42 35 35 ICV_22 $T=72640 14315 0 180 $X=58300 $Y=13685
X189 38 39 38 38 37 40 37 37 ICV_22 $T=72640 17395 0 180 $X=58300 $Y=16765
X190 12 13 49 13 13 IN 50 IN ICV_22 $T=58640 21135 1 0 $X=58300 $Y=20505
X191 11 11 47 11 11 12 48 12 ICV_22 $T=58640 24215 1 0 $X=58300 $Y=23585
X192 9 10 45 10 10 11 46 11 ICV_22 $T=58640 27295 1 0 $X=58300 $Y=26665
X193 1 7 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758 $T=2980 2025 0 90 $X=2330 $Y=2025
X194 1 6 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758 $T=2980 3565 0 90 $X=2330 $Y=3565
X195 1 5 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758 $T=2980 5100 0 90 $X=2330 $Y=5100
X196 1 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758 $T=2980 6640 0 90 $X=2330 $Y=6640
X197 13 12 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758 $T=58060 22600 1 90 $X=58060 $Y=22600
X198 12 11 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758 $T=58060 24140 1 90 $X=58060 $Y=24140
X199 11 10 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758 $T=58060 27220 1 90 $X=58060 $Y=27220
X200 10 9 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758 $T=58060 28760 1 90 $X=58060 $Y=28760
X201 3 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808760 $T=2980 8155 0 90 $X=2330 $Y=8155
X202 11 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808760 $T=58060 25680 1 90 $X=58060 $Y=25680
X203 9 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808761 $T=29530 9405 0 0 $X=29530 $Y=9405
X204 4 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808761 $T=54470 7095 0 0 $X=54470 $Y=7095
X218 1 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759 $T=15570 6585 0 90 $X=15280 $Y=6585
X219 1 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759 $T=24130 5045 0 90 $X=23840 $Y=5045
X220 1 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759 $T=28410 3505 0 90 $X=28120 $Y=3505
X221 1 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759 $T=32690 1965 0 90 $X=32400 $Y=1965
X222 8 21 1 ICV_25 $T=16535 935 0 0 $X=16525 $Y=935
X223 7 22 1 ICV_25 $T=16535 2475 0 0 $X=16525 $Y=2475
X224 6 23 1 ICV_25 $T=16535 4015 0 0 $X=16525 $Y=4015
X225 5 24 1 ICV_25 $T=16535 5555 0 0 $X=16525 $Y=5555
X226 4 25 3 ICV_25 $T=16535 7095 0 0 $X=16525 $Y=7095
X227 3 26 9 ICV_25 $T=16535 8635 0 0 $X=16525 $Y=8635
X228 15 27 16 ICV_25 $T=16535 31450 0 0 $X=16525 $Y=31450
X229 16 28 17 ICV_25 $T=16535 32990 0 0 $X=16525 $Y=32990
X230 17 29 18 ICV_25 $T=16535 34530 0 0 $X=16525 $Y=34530
X231 18 30 19 ICV_25 $T=16535 36070 0 0 $X=16525 $Y=36070
X232 19 31 20 ICV_25 $T=16535 37610 0 0 $X=16525 $Y=37610
X233 1 9 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808756 $T=7010 9665 0 90 $X=6720 $Y=9665
X234 1 3 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808756 $T=11290 8125 0 90 $X=11000 $Y=8125
X235 32 20 IN ICV_26 $T=16910 39030 1 180 $X=2570 $Y=38900
X236 15 45 ICV_27 $T=2910 30560 0 0 $X=2570 $Y=30430
X237 13 31 19 20 50 ICV_28 $T=16910 37490 1 180 $X=2570 $Y=37360
X238 38 39 21 1 8 37 40 22 1 7 ICV_29 $T=16910 815 1 180 $X=2570 $Y=685
X239 36 41 23 1 6 35 42 24 1 5 ICV_29 $T=16910 3895 1 180 $X=2570 $Y=3765
X240 34 43 25 3 4 33 44 26 9 3 ICV_29 $T=16910 6975 1 180 $X=2570 $Y=6845
X241 10 46 27 16 15 11 47 28 17 16 ICV_29 $T=16910 31330 1 180 $X=2570 $Y=31200
X242 11 48 29 18 17 12 49 30 19 18 ICV_29 $T=16910 34410 1 180 $X=2570 $Y=34280
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_55959141808243
** N=5 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808723
** N=13 EP=0 IP=10 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd__example_5595914180848
** N=16 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_5595914180849
** N=17 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__model__pfet_highvoltage__example_55959141808371
** N=15 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_io__hvsbt_inv_x1
** N=31 EP=0 IP=24 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VGND VPWR OUT
.ENDS
***************************************
.SUBCKT sky130_fd_pr__model__pfet_highvoltage__example_55959141808421
** N=23 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_io__hvsbt_inv_x2
** N=44 EP=0 IP=28 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VGND VPWR IN OUT
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_55959141808719
** N=11 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808720
** N=24 EP=0 IP=22 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_5595914180829
** N=31 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808767 2 3 4 5
** N=26 EP=4 IP=22 FDC=1
*.SEEDPROM
M0 5 3 4 2 phv L=0.5 W=3 AD=0.84 AS=0.84 PD=6.56 PS=6.56 NRD=0 NRS=0 m=1 r=6 sa=250000 sb=250000 a=1.5 p=7 mult=1 $X=0 $Y=0 $D=109
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_tie_r_out_esd A B
** N=8 EP=2 IP=6 FDC=1
X0 A B sky130_fd_pr__res_generic_po__example_5595914180838 $T=1000 1095 0 0 $X=730 $Y=1095
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_55959141808765
** N=10 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808764 1 2 3 4
** N=9 EP=4 IP=4 FDC=1
M0 4 2 3 1 nhv L=0.5 W=3 AD=0.84 AS=0.84 PD=6.56 PS=6.56 NRD=0 NRS=0 m=1 r=6 sa=250000 sb=250000 a=1.5 p=7 mult=1 $X=0 $Y=0 $D=49
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808779 1 2 3 4
** N=15 EP=4 IP=10 FDC=1
M0 4 2 3 1 nhvnative L=0.9 W=1 AD=0.28 AS=0.28 PD=2.56 PS=2.56 NRD=0 NRS=0 m=1 r=1.11111 sa=450000 sb=450000 a=0.9 p=3.8 mult=1 $X=0 $Y=0 $D=59
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808777 1 2 3
** N=16 EP=3 IP=2 FDC=1
M0 3 2 1 1 nhv L=0.5 W=3 AD=0.84 AS=0.795 PD=6.56 PS=6.53 NRD=0 NRS=0 m=1 r=6 sa=250000 sb=250000 a=1.5 p=7 mult=1 $X=0 $Y=0 $D=49
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_5595914180827
** N=16 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd__example_55959141808233
** N=16 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808778
** N=53 EP=0 IP=48 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_55959141808449
** N=6 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808784 2 3 4
** N=9 EP=3 IP=6 FDC=1
*.SEEDPROM
M0 2 3 4 2 phv L=0.8 W=1 AD=0.28 AS=0.28 PD=2.56 PS=2.56 NRD=0 NRS=0 m=1 r=1.25 sa=400000 sb=400000 a=0.8 p=3.6 mult=1 $X=0 $Y=0 $D=109
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_559591418085
** N=16 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808783
** N=11 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd__example_55959141808782
** N=10 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808786
** N=35 EP=0 IP=33 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808787
** N=36 EP=0 IP=34 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__tpl1__example_55959141808151
** N=30 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__tpl1__example_55959141808148
** N=17 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__tpl1__example_55959141808150
** N=20 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__tpl1__example_55959141808149
** N=11 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1__example_55959141808158
** N=16 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_io__signal_5_sym_hv_local_5term NBODY NWELLRING GATE VGND IN 7
** N=101 EP=6 IP=102 FDC=3
*.SEEDPROM
M0 IN GATE VGND NBODY nhvesd L=0.6 W=5.4 AD=3.65486 AS=3.65486 PD=11.6192 PS=11.6192 NRD=8.436 NRS=9.2796 m=1 r=9 sa=300000 sb=300000 a=3.24 p=12 mult=1 $X=3675 $Y=3360 $D=129
R1 NWELLRING 7 0.01 m=1 $[short] $X=1015 $Y=330 $D=282
R2 NBODY 51 0.01 m=1 $[short] $X=2665 $Y=330 $D=282
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd__example_5595914180819
** N=10 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpio_buf_localesdv2 VGND VCC_IO VTRIP_SEL_H OUT_H 5
** N=179 EP=5 IP=209 FDC=25
*.SEEDPROM
M0 OUT_VT VTRIP_SEL_H OUT_H VGND nhv L=1 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 m=1 r=3 sa=500000 sb=500000 a=3 p=8 mult=1 $X=16175 $Y=17310 $D=49
X1 VGND VCC_IO Dpar a=8.5092 p=29.27 m=1 $[nwdiode] $X=1460 $Y=1770 $D=190
X2 VGND VCC_IO Dpar a=8.5092 p=29.27 m=1 $[nwdiode] $X=1460 $Y=12530 $D=190
X3 VGND VCC_IO Dpar a=8.5092 p=29.27 m=1 $[nwdiode] $X=8055 $Y=1770 $D=190
X4 VGND VCC_IO Dpar a=8.5092 p=29.27 m=1 $[nwdiode] $X=8055 $Y=12530 $D=190
X5 VGND VCC_IO Dpar a=5.1688 p=17.34 m=1 $[nwdiode] $X=14650 $Y=15810 $D=190
X6 5 OUT_H sky130_fd_io__res250only_small $T=17545 -185 0 90 $X=15525 $Y=-185
X7 VGND VCC_IO VGND VGND OUT_VT 8 sky130_fd_io__signal_5_sym_hv_local_5term $T=8335 690 1 180 $X=380 $Y=690
X8 VGND VCC_IO VGND VGND OUT_H 10 sky130_fd_io__signal_5_sym_hv_local_5term $T=8335 23570 0 180 $X=380 $Y=11450
X9 VGND VCC_IO VGND OUT_VT VCC_IO 7 sky130_fd_io__signal_5_sym_hv_local_5term $T=6975 690 0 0 $X=6975 $Y=690
X10 VGND VCC_IO VGND OUT_H VCC_IO 9 sky130_fd_io__signal_5_sym_hv_local_5term $T=6975 23570 1 0 $X=6975 $Y=11450
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpm1s2__example_55959141808659
** N=44 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808658
** N=36 EP=0 IP=26 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s__example_55959141808646
** N=31 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808647
** N=6 EP=0 IP=3 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpm1s2__example_55959141808649
** N=45 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_30
** N=4 EP=0 IP=8 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808650
** N=6 EP=0 IP=3 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2 1 2 VCC_IO 4 5 6 7 8 9 10 11 12 13 14
** N=3678 EP=14 IP=217 FDC=58
*.SEEDPROM
M0 14 4 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.425 PD=6.55 PS=11.37 NRD=10.374 NRS=8.7666 m=1 r=8.33333 sa=300002 sb=300020 a=3 p=11.2 mult=1 $X=4620 $Y=7285 $D=49
M1 14 4 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.425 PD=6.55 PS=11.37 NRD=10.374 NRS=8.7666 m=1 r=8.33333 sa=300002 sb=300020 a=3 p=11.2 mult=1 $X=4620 $Y=15290 $D=49
M2 2 4 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300004 sb=300020 a=3 p=11.2 mult=1 $X=6770 $Y=7285 $D=49
M3 2 4 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300004 sb=300020 a=3 p=11.2 mult=1 $X=6770 $Y=15290 $D=49
M4 14 4 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300007 sb=300020 a=3 p=11.2 mult=1 $X=9580 $Y=7285 $D=49
M5 14 4 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300007 sb=300020 a=3 p=11.2 mult=1 $X=9580 $Y=15290 $D=49
M6 2 4 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300009 sb=300020 a=3 p=11.2 mult=1 $X=11730 $Y=7285 $D=49
M7 2 4 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300009 sb=300020 a=3 p=11.2 mult=1 $X=11730 $Y=15290 $D=49
M8 14 5 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300011 sb=300020 a=3 p=11.2 mult=1 $X=14540 $Y=7285 $D=49
M9 14 5 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300011 sb=300020 a=3 p=11.2 mult=1 $X=14540 $Y=15290 $D=49
M10 2 5 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300014 sb=300020 a=3 p=11.2 mult=1 $X=16690 $Y=7285 $D=49
M11 2 5 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300014 sb=300020 a=3 p=11.2 mult=1 $X=16690 $Y=15290 $D=49
M12 14 5 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300016 sb=300020 a=3 p=11.2 mult=1 $X=19500 $Y=7285 $D=49
M13 14 5 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300016 sb=300020 a=3 p=11.2 mult=1 $X=19500 $Y=15290 $D=49
M14 2 6 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300019 sb=300020 a=3 p=11.2 mult=1 $X=21650 $Y=7285 $D=49
M15 2 6 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300019 sb=300020 a=3 p=11.2 mult=1 $X=21650 $Y=15290 $D=49
M16 14 6 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=24460 $Y=7285 $D=49
M17 14 6 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=24460 $Y=15290 $D=49
M18 2 6 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=26610 $Y=7285 $D=49
M19 2 6 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=26610 $Y=15290 $D=49
M20 14 7 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=29420 $Y=7285 $D=49
M21 14 7 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=29420 $Y=15290 $D=49
M22 2 7 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=31570 $Y=7285 $D=49
M23 2 7 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=31570 $Y=15290 $D=49
M24 14 7 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=34380 $Y=7285 $D=49
M25 14 7 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=34380 $Y=15290 $D=49
M26 2 8 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=36530 $Y=7285 $D=49
M27 2 8 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=36530 $Y=15290 $D=49
M28 14 9 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=39340 $Y=7285 $D=49
M29 14 9 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=39340 $Y=15290 $D=49
M30 2 9 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=41490 $Y=7285 $D=49
M31 2 9 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=41490 $Y=15290 $D=49
M32 14 9 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=44300 $Y=7285 $D=49
M33 14 9 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=44300 $Y=15290 $D=49
M34 2 10 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=46450 $Y=7285 $D=49
M35 2 10 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=46450 $Y=15290 $D=49
M36 14 10 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=49260 $Y=7285 $D=49
M37 14 10 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=49260 $Y=15290 $D=49
M38 2 10 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=51410 $Y=7285 $D=49
M39 2 10 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=51410 $Y=15290 $D=49
M40 14 10 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300018 a=3 p=11.2 mult=1 $X=54220 $Y=7285 $D=49
M41 14 10 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300018 a=3 p=11.2 mult=1 $X=54220 $Y=15290 $D=49
M42 2 10 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300016 a=3 p=11.2 mult=1 $X=56370 $Y=7285 $D=49
M43 2 10 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300016 a=3 p=11.2 mult=1 $X=56370 $Y=15290 $D=49
M44 14 10 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300013 a=3 p=11.2 mult=1 $X=59180 $Y=7285 $D=49
M45 14 10 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300013 a=3 p=11.2 mult=1 $X=59180 $Y=15290 $D=49
M46 2 11 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300011 a=3 p=11.2 mult=1 $X=61330 $Y=7285 $D=49
M47 2 11 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300011 a=3 p=11.2 mult=1 $X=61330 $Y=15290 $D=49
M48 14 12 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300008 a=3 p=11.2 mult=1 $X=64140 $Y=7285 $D=49
M49 14 12 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300008 a=3 p=11.2 mult=1 $X=64140 $Y=15290 $D=49
M50 2 13 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300006 a=3 p=11.2 mult=1 $X=66290 $Y=7285 $D=49
M51 2 13 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300006 a=3 p=11.2 mult=1 $X=66290 $Y=15290 $D=49
M52 14 13 2 2 nhv L=0.6 W=5 AD=2.975 AS=3.775 PD=6.19 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300003 a=3 p=11.2 mult=1 $X=69100 $Y=7285 $D=49
M53 14 13 2 2 nhv L=0.6 W=5 AD=2.975 AS=3.775 PD=6.19 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300003 a=3 p=11.2 mult=1 $X=69100 $Y=15290 $D=49
M54 2 13 14 2 nhv L=0.6 W=5 AD=3.425 AS=2.975 PD=11.37 PS=6.19 NRD=8.7666 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300002 a=3 p=11.2 mult=1 $X=70890 $Y=7285 $D=49
M55 2 13 14 2 nhv L=0.6 W=5 AD=3.425 AS=2.975 PD=11.37 PS=6.19 NRD=8.7666 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300002 a=3 p=11.2 mult=1 $X=70890 $Y=15290 $D=49
X56 1 VCC_IO Dpar a=1791.37 p=197.77 m=1 $[dnwdiode_psub] $X=440 $Y=2895 $D=193
X57 2 VCC_IO Dpar a=1558.74 p=186.49 m=1 $[dnwdiode_pw] $X=2345 $Y=3925 $D=194
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpio_pddrvr_strong_xres4v2 1 TIE_LO_ESD VGND_IO VCC_IO PD_H[2] PD_H[3] 7 8
** N=70 EP=8 IP=140 FDC=108
*.SEEDPROM
X0 VGND_IO VCC_IO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=6380 $Y=37555 $D=150
X1 PD_H[3] 7 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=3275 5230 1 90 $X=3275 $Y=5230
X2 PD_H[2] 7 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=4480 5230 1 90 $X=4480 $Y=5230
X3 PD_H[3] 15 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=8470 5230 0 90 $X=7820 $Y=5230
X4 TIE_LO_ESD 15 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=9885 5230 0 90 $X=9235 $Y=5230
X5 PD_H[3] 14 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=16120 5230 0 90 $X=15470 $Y=5230
X6 TIE_LO_ESD 14 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=17535 5230 0 90 $X=16885 $Y=5230
X7 PD_H[2] 13 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=34665 5230 0 90 $X=34015 $Y=5230
X8 TIE_LO_ESD 13 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=38965 5230 0 90 $X=38315 $Y=5230
X9 PD_H[2] 12 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=43175 5230 0 90 $X=42525 $Y=5230
X10 TIE_LO_ESD 12 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=47475 5230 0 90 $X=46825 $Y=5230
X11 PD_H[2] 11 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=50575 5230 0 90 $X=49925 $Y=5230
X12 TIE_LO_ESD 11 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=54875 5230 0 90 $X=54225 $Y=5230
X13 PD_H[2] 10 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=57290 5230 0 90 $X=56640 $Y=5230
X14 TIE_LO_ESD 10 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=61590 5230 0 90 $X=60940 $Y=5230
X15 PD_H[2] 9 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=64460 5230 0 90 $X=63810 $Y=5230
X16 PD_H[3] 9 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=66610 5230 0 90 $X=65960 $Y=5230
X17 TIE_LO_ESD 7 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=2065 5230 1 90 $X=2065 $Y=5230
X18 PD_H[2] 15 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=6950 5230 0 90 $X=6300 $Y=5230
X19 PD_H[2] 14 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=14600 5230 0 90 $X=13950 $Y=5230
X20 PD_H[3] 13 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=36815 5230 0 90 $X=36165 $Y=5230
X21 PD_H[3] 12 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=45325 5230 0 90 $X=44675 $Y=5230
X22 PD_H[3] 11 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=52725 5230 0 90 $X=52075 $Y=5230
X23 PD_H[3] 10 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=59440 5230 0 90 $X=58790 $Y=5230
X24 TIE_LO_ESD 9 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=68760 5230 0 90 $X=68110 $Y=5230
X25 TIE_LO_ESD VGND_IO sky130_fd_pr__res_generic_po__example_5595914180838 $T=2320 46835 0 0 $X=2050 $Y=46835
X26 1 VGND_IO VCC_IO 9 10 11 12 13 PD_H[2] PD_H[3] 14 15 7 8 sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2 $T=75440 42045 0 180 $X=-515 $Y=14600
.ENDS
***************************************
.SUBCKT ICV_1 VSSD VDDIO VCCHIB VDDIO_Q ENABLE_H EN_VDDIO_SIG_H INP_SEL_H ENABLE_VDDIO PAD PULLUP_H DISABLE_PULLUP_H PAD_A_ESD_H VSSIO FILT_IN_H XRES_H_N TIE_WEAK_HI_H
** N=38667 EP=16 IP=1572 FDC=776
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VCCD VDDA VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q
M0 VSSD ENABLE_VDDIO 36 VSSD nshort L=0.15 W=0.74 AD=0.2627 AS=0.2109 PD=2.19 PS=2.05 NRD=11.34 NRS=0 m=1 r=4.93333 sa=75000.2 sb=75000.3 a=0.111 p=1.78 mult=1 $X=16840 $Y=40175 $D=9
M1 61 34 VSSD VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=13.8396 NRS=0 m=1 r=1.16667 sa=300000 sb=300001 a=0.42 p=2.6 mult=1 $X=8460 $Y=7500 $D=49
M2 54 ENABLE_H 61 VSSD nhv L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=13.8396 m=1 r=1.16667 sa=300001 sb=300000 a=0.42 p=2.6 mult=1 $X=9340 $Y=7500 $D=49
M3 35 54 VSSD VSSD nhv L=0.6 W=0.7 AD=0.1855 AS=0.1855 PD=1.93 PS=1.93 NRD=0 NRS=0 m=1 r=1.16667 sa=300000 sb=300000 a=0.42 p=2.6 mult=1 $X=10845 $Y=7500 $D=49
M4 33 39 VSSD VSSD nhv L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 r=10 sa=250000 sb=250002 a=2.5 p=11 mult=1 $X=15285 $Y=20910 $D=49
M5 VSSD 39 33 VSSD nhv L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250001 sb=250002 a=2.5 p=11 mult=1 $X=15285 $Y=21690 $D=49
M6 32 37 VSSD VSSD nhv L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250002 sb=250001 a=2.5 p=11 mult=1 $X=15285 $Y=22470 $D=49
M7 VSSD 37 32 VSSD nhv L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250002 sb=250000 a=2.5 p=11 mult=1 $X=15285 $Y=23250 $D=49
M8 64 37 62 VSSD nhv L=0.8 W=5 AD=0.7 AS=1.4 PD=5.28 PS=10.56 NRD=0 NRS=0 m=1 r=6.25 sa=400000 sb=400007 a=4 p=11.6 mult=1 $X=15315 $Y=28245 $D=49
M9 62 37 64 VSSD nhv L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=6.25 sa=400001 sb=400006 a=4 p=11.6 mult=1 $X=15315 $Y=29325 $D=49
M10 64 37 62 VSSD nhv L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=6.25 sa=400002 sb=400005 a=4 p=11.6 mult=1 $X=15315 $Y=30405 $D=49
M11 62 37 64 VSSD nhv L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=6.25 sa=400003 sb=400004 a=4 p=11.6 mult=1 $X=15315 $Y=31485 $D=49
M12 VSSD 30 62 VSSD nhv L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=6.25 sa=400004 sb=400003 a=4 p=11.6 mult=1 $X=15315 $Y=32565 $D=49
M13 62 30 VSSD VSSD nhv L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=6.25 sa=400005 sb=400002 a=4 p=11.6 mult=1 $X=15315 $Y=33645 $D=49
M14 37 30 62 VSSD nhv L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=6.25 sa=400006 sb=400001 a=4 p=11.6 mult=1 $X=15315 $Y=34725 $D=49
M15 62 30 37 VSSD nhv L=0.8 W=5 AD=1.4 AS=0.7 PD=10.56 PS=5.28 NRD=0 NRS=0 m=1 r=6.25 sa=400007 sb=400000 a=4 p=11.6 mult=1 $X=15315 $Y=35805 $D=49
M16 62 37 57 VSSD nhv L=0.8 W=5 AD=1.4 AS=1.4 PD=10.56 PS=10.56 NRD=0 NRS=0 m=1 r=6.25 sa=400000 sb=400000 a=4 p=11.6 mult=1 $X=15315 $Y=37540 $D=49
M17 VSSD 31 52 VSSD nhv L=0.5 W=1 AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 m=1 r=2 sa=250000 sb=250002 a=0.5 p=3 mult=1 $X=21425 $Y=21690 $D=49
M18 52 31 VSSD VSSD nhv L=0.5 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=2 sa=250001 sb=250001 a=0.5 p=3 mult=1 $X=21425 $Y=22470 $D=49
M19 VSSD 31 52 VSSD nhv L=0.5 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 r=2 sa=250002 sb=250000 a=0.5 p=3 mult=1 $X=21425 $Y=23250 $D=49
M20 43 71 VSSD VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 r=1.16667 sa=300000 sb=300003 a=0.42 p=2.6 mult=1 $X=27755 $Y=29045 $D=49
M21 VSSD 71 43 VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300001 sb=300002 a=0.42 p=2.6 mult=1 $X=27755 $Y=29925 $D=49
M22 71 DISABLE_PULLUP_H VSSD VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300002 sb=300001 a=0.42 p=2.6 mult=1 $X=27755 $Y=30805 $D=49
M23 VSSD DISABLE_PULLUP_H 71 VSSD nhv L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300003 sb=300000 a=0.42 p=2.6 mult=1 $X=27755 $Y=31685 $D=49
M24 VSSD 41 63 VSSD nhv L=1 W=0.42 AD=0.1176 AS=0.1176 PD=1.4 PS=1.4 NRD=0 NRS=0 m=1 r=0.42 sa=500000 sb=500000 a=0.42 p=2.84 mult=1 $X=30440 $Y=14450 $D=49
M25 63 42 VSSD VSSD nhv L=1 W=1 AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 m=1 r=1 sa=500000 sb=500001 a=1 p=4 mult=1 $X=30720 $Y=9780 $D=49
M26 44 42 63 VSSD nhv L=1 W=1 AD=0.28 AS=0.14 PD=2.56 PS=1.28 NRD=0 NRS=0 m=1 r=1 sa=500001 sb=500000 a=1 p=4 mult=1 $X=30720 $Y=11060 $D=49
M27 41 44 VSSD VSSD nhv L=0.5 W=1 AD=0.28 AS=0.28 PD=2.56 PS=2.56 NRD=0 NRS=0 m=1 r=2 sa=250000 sb=250000 a=0.5 p=3 mult=1 $X=30720 $Y=12990 $D=49
M28 40 INP_SEL_H VSSD VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 r=1.16667 sa=300000 sb=300007 a=0.42 p=2.6 mult=1 $X=31240 $Y=17710 $D=49
M29 VSSD INP_SEL_H 40 VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300001 sb=300006 a=0.42 p=2.6 mult=1 $X=31240 $Y=18590 $D=49
M30 34 EN_VDDIO_SIG_H VSSD VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300002 sb=300005 a=0.42 p=2.6 mult=1 $X=31240 $Y=19470 $D=49
M31 VSSD EN_VDDIO_SIG_H 34 VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300003 sb=300004 a=0.42 p=2.6 mult=1 $X=31240 $Y=20350 $D=49
M32 XRES_H_N 72 VSSD VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300003 sb=300003 a=0.42 p=2.6 mult=1 $X=31240 $Y=21230 $D=49
M33 VSSD 72 XRES_H_N VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300004 sb=300003 a=0.42 p=2.6 mult=1 $X=31240 $Y=22110 $D=49
M34 XRES_H_N 72 VSSD VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300005 sb=300002 a=0.42 p=2.6 mult=1 $X=31240 $Y=22990 $D=49
M35 VSSD 72 XRES_H_N VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300006 sb=300001 a=0.42 p=2.6 mult=1 $X=31240 $Y=23870 $D=49
M36 72 41 VSSD VSSD nhv L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300007 sb=300000 a=0.42 p=2.6 mult=1 $X=31240 $Y=24750 $D=49
M37 XRES_H_N 72 VSSD VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 r=1.16667 sa=300000 sb=300003 a=0.42 p=2.6 mult=1 $X=35355 $Y=4770 $D=49
M38 VSSD 72 XRES_H_N VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300001 sb=300002 a=0.42 p=2.6 mult=1 $X=36235 $Y=4770 $D=49
M39 XRES_H_N 72 VSSD VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300002 sb=300001 a=0.42 p=2.6 mult=1 $X=37115 $Y=4770 $D=49
M40 VSSD 72 XRES_H_N VSSD nhv L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300003 sb=300000 a=0.42 p=2.6 mult=1 $X=37995 $Y=4770 $D=49
M41 24 35 60 VSSD nhvnative L=0.9 W=10 AD=2.8 AS=2.8 PD=20.56 PS=20.56 NRD=0 NRS=0 m=1 r=11.1111 sa=450000 sb=450000 a=9 p=21.8 mult=1 $X=21675 $Y=26745 $D=59
M42 VSSD VSSD VSSD VSSD nhvnative L=0.9 W=10 AD=2.8 AS=2.65 PD=20.56 PS=20.53 NRD=0 NRS=0 m=1 r=11.1111 sa=450000 sb=450000 a=9 p=21.8 mult=1 $X=23490 $Y=26745 $D=59
M43 VCCHIB ENABLE_VDDIO 36 VCCHIB phighvt L=0.15 W=1.12 AD=0.3864 AS=0.3304 PD=2.93 PS=2.83 NRD=10.5395 NRS=1.7533 m=1 r=7.46667 sa=75000.2 sb=75000.3 a=0.168 p=2.54 mult=1 $X=14990 $Y=40185 $D=89
M44 PAD 27 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=4.325 PD=6.55 PS=11.73 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300002 sb=300020 a=3 p=11.2 mult=1 $X=4065 $Y=107610 $D=109
M45 PAD 27 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=4.325 PD=6.55 PS=11.73 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300002 sb=300020 a=3 p=11.2 mult=1 $X=4065 $Y=115610 $D=109
M46 VDDIO 27 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300004 sb=300020 a=3 p=11.2 mult=1 $X=6215 $Y=107610 $D=109
M47 VDDIO 27 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300004 sb=300020 a=3 p=11.2 mult=1 $X=6215 $Y=115610 $D=109
M48 VDDIO_Q 32 33 VDDIO_Q phv L=0.5 W=0.42 AD=0.0588 AS=0.1176 PD=0.7 PS=1.4 NRD=0 NRS=0 m=1 r=0.84 sa=250000 sb=250001 a=0.21 p=1.84 mult=1 $X=7410 $Y=24400 $D=109
M49 32 33 VDDIO_Q VDDIO_Q phv L=0.5 W=0.42 AD=0.1176 AS=0.0588 PD=1.4 PS=0.7 NRD=0 NRS=0 m=1 r=0.84 sa=250001 sb=250000 a=0.21 p=1.84 mult=1 $X=7410 $Y=25180 $D=109
M50 54 34 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 r=1.66667 sa=300000 sb=300001 a=0.6 p=3.2 mult=1 $X=8460 $Y=4170 $D=109
M51 54 34 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 r=1.66667 sa=300000 sb=300001 a=0.6 p=3.2 mult=1 $X=8460 $Y=5510 $D=109
M52 PAD 27 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300007 sb=300020 a=3 p=11.2 mult=1 $X=9025 $Y=107610 $D=109
M53 PAD 27 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300007 sb=300020 a=3 p=11.2 mult=1 $X=9025 $Y=115610 $D=109
M54 VDDIO_Q ENABLE_H 54 VDDIO_Q phv L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300001 sb=300000 a=0.6 p=3.2 mult=1 $X=9340 $Y=4170 $D=109
M55 VDDIO_Q ENABLE_H 54 VDDIO_Q phv L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300001 sb=300000 a=0.6 p=3.2 mult=1 $X=9340 $Y=5510 $D=109
M56 VDDIO_Q 31 52 VDDIO_Q phv L=0.5 W=3 AD=0.42 AS=0.84 PD=3.28 PS=6.56 NRD=0 NRS=0 m=1 r=6 sa=250000 sb=250002 a=1.5 p=7 mult=1 $X=7095 $Y=19975 $D=109
M57 52 31 VDDIO_Q VDDIO_Q phv L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 r=6 sa=250001 sb=250001 a=1.5 p=7 mult=1 $X=7095 $Y=20755 $D=109
M58 VDDIO_Q 31 52 VDDIO_Q phv L=0.5 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 r=6 sa=250002 sb=250000 a=1.5 p=7 mult=1 $X=7095 $Y=21535 $D=109
M59 VDDIO_Q 32 31 VDDIO_Q phv L=0.5 W=3 AD=0.795 AS=0.84 PD=6.53 PS=6.56 NRD=0 NRS=0 m=1 r=6 sa=250000 sb=250000 a=1.5 p=7 mult=1 $X=7095 $Y=22950 $D=109
M60 35 54 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 r=1.66667 sa=300000 sb=300000 a=0.6 p=3.2 mult=1 $X=10845 $Y=4170 $D=109
M61 35 54 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 r=1.66667 sa=300000 sb=300000 a=0.6 p=3.2 mult=1 $X=10845 $Y=5510 $D=109
M62 VDDIO 27 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300009 sb=300020 a=3 p=11.2 mult=1 $X=11175 $Y=107610 $D=109
M63 VDDIO 27 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300009 sb=300020 a=3 p=11.2 mult=1 $X=11175 $Y=115610 $D=109
M64 VDDIO_Q ENABLE_H 55 VDDIO_Q phv L=0.5 W=5 AD=1.325 AS=1.4 PD=10.53 PS=10.56 NRD=0 NRS=0 m=1 r=10 sa=250000 sb=250000 a=2.5 p=11 mult=1 $X=6920 $Y=29660 $D=109
M65 51 30 37 VDDIO_Q phv L=0.5 W=5 AD=1.4 AS=1.4 PD=10.56 PS=10.56 NRD=0 NRS=0 m=1 r=10 sa=250000 sb=250000 a=2.5 p=11 mult=1 $X=6920 $Y=31460 $D=109
M66 56 35 VDDIO_Q VDDIO_Q phv L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 r=10 sa=250000 sb=250001 a=2.5 p=11 mult=1 $X=6920 $Y=32875 $D=109
M67 51 34 56 VDDIO_Q phv L=0.5 W=5 AD=1.4 AS=0.7 PD=10.56 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250001 sb=250000 a=2.5 p=11 mult=1 $X=6920 $Y=33655 $D=109
M68 VDDIO_Q 34 57 VDDIO_Q phv L=0.5 W=5 AD=0.7 AS=1.4 PD=5.28 PS=10.56 NRD=0 NRS=0 m=1 r=10 sa=250000 sb=250001 a=2.5 p=11 mult=1 $X=6920 $Y=35115 $D=109
M69 58 EN_VDDIO_SIG_H VDDIO_Q VDDIO_Q phv L=0.5 W=5 AD=1.4 AS=0.7 PD=10.56 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250001 sb=250000 a=2.5 p=11 mult=1 $X=6920 $Y=35895 $D=109
M70 VCCHIB 36 59 VCCHIB phv L=0.5 W=5 AD=0.7 AS=1.4 PD=5.28 PS=10.56 NRD=0 NRS=0 m=1 r=10 sa=250000 sb=250001 a=2.5 p=11 mult=1 $X=6920 $Y=39685 $D=109
M71 60 36 VCCHIB VCCHIB phv L=0.5 W=5 AD=1.4 AS=0.7 PD=10.56 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250001 sb=250000 a=2.5 p=11 mult=1 $X=6920 $Y=40465 $D=109
M72 25 37 39 25 phv L=0.5 W=5 AD=1.4 AS=1.4 PD=10.56 PS=10.56 NRD=0 NRS=0 m=1 r=10 sa=250000 sb=250000 a=2.5 p=11 mult=1 $X=7095 $Y=15515 $D=109
M73 45 37 39 VDDIO_Q phv L=0.5 W=5 AD=0.7 AS=1.4 PD=5.28 PS=10.56 NRD=0 NRS=0 m=1 r=10 sa=250000 sb=250002 a=2.5 p=11 mult=1 $X=7095 $Y=26635 $D=109
M74 26 34 45 VDDIO_Q phv L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250001 sb=250001 a=2.5 p=11 mult=1 $X=7095 $Y=27415 $D=109
M75 VDDIO_Q 35 26 VDDIO_Q phv L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250002 sb=250000 a=2.5 p=11 mult=1 $X=7095 $Y=28195 $D=109
M76 PAD 27 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300012 sb=300020 a=3 p=11.2 mult=1 $X=13985 $Y=107610 $D=109
M77 PAD 27 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300012 sb=300020 a=3 p=11.2 mult=1 $X=13985 $Y=115610 $D=109
M78 VDDIO 27 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300014 sb=300020 a=3 p=11.2 mult=1 $X=16135 $Y=107610 $D=109
M79 VDDIO 27 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300014 sb=300020 a=3 p=11.2 mult=1 $X=16135 $Y=115610 $D=109
M80 PAD 27 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300017 sb=300020 a=3 p=11.2 mult=1 $X=18945 $Y=107610 $D=109
M81 PAD 27 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300017 sb=300020 a=3 p=11.2 mult=1 $X=18945 $Y=115610 $D=109
M82 VDDIO 27 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300019 sb=300020 a=3 p=11.2 mult=1 $X=21095 $Y=107610 $D=109
M83 VDDIO 27 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300019 sb=300020 a=3 p=11.2 mult=1 $X=21095 $Y=115610 $D=109
M84 PAD 27 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=23905 $Y=107610 $D=109
M85 PAD 27 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=23905 $Y=115610 $D=109
M86 VDDIO 27 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=26055 $Y=107610 $D=109
M87 VDDIO 27 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=26055 $Y=115610 $D=109
M88 53 41 VDDIO_Q VDDIO_Q phv L=1 W=0.42 AD=0.1176 AS=0.1176 PD=1.4 PS=1.4 NRD=0 NRS=0 m=1 r=0.42 sa=500000 sb=500000 a=0.42 p=2.84 mult=1 $X=26705 $Y=14610 $D=109
M89 29 43 VDDIO VDDIO phv L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 r=10 sa=250000 sb=250002 a=2.5 p=11 mult=1 $X=27850 $Y=35625 $D=109
M90 40 INP_SEL_H VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 r=1.66667 sa=300000 sb=300007 a=0.6 p=3.2 mult=1 $X=27910 $Y=17710 $D=109
M91 VDDIO_Q INP_SEL_H 40 VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300001 sb=300006 a=0.6 p=3.2 mult=1 $X=27910 $Y=18590 $D=109
M92 34 EN_VDDIO_SIG_H VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300002 sb=300005 a=0.6 p=3.2 mult=1 $X=27910 $Y=19470 $D=109
M93 VDDIO_Q EN_VDDIO_SIG_H 34 VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300003 sb=300004 a=0.6 p=3.2 mult=1 $X=27910 $Y=20350 $D=109
M94 XRES_H_N 72 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300003 sb=300003 a=0.6 p=3.2 mult=1 $X=27910 $Y=21230 $D=109
M95 VDDIO_Q 72 XRES_H_N VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300004 sb=300003 a=0.6 p=3.2 mult=1 $X=27910 $Y=22110 $D=109
M96 XRES_H_N 72 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300005 sb=300002 a=0.6 p=3.2 mult=1 $X=27910 $Y=22990 $D=109
M97 VDDIO_Q 72 XRES_H_N VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300006 sb=300001 a=0.6 p=3.2 mult=1 $X=27910 $Y=23870 $D=109
M98 72 41 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300007 sb=300000 a=0.6 p=3.2 mult=1 $X=27910 $Y=24750 $D=109
M99 VDDIO 43 29 VDDIO phv L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250001 sb=250002 a=2.5 p=11 mult=1 $X=28630 $Y=35625 $D=109
M100 53 42 VDDIO_Q VDDIO_Q phv L=1 W=3 AD=0.42 AS=0.84 PD=3.28 PS=6.56 NRD=0 NRS=0 m=1 r=3 sa=500000 sb=500001 a=3 p=8 mult=1 $X=26420 $Y=9780 $D=109
M101 44 42 53 VDDIO_Q phv L=1 W=3 AD=0.84 AS=0.42 PD=6.56 PS=3.28 NRD=0 NRS=0 m=1 r=3 sa=500001 sb=500000 a=3 p=8 mult=1 $X=26420 $Y=11060 $D=109
M102 41 44 VDDIO_Q VDDIO_Q phv L=0.5 W=3 AD=0.84 AS=0.84 PD=6.56 PS=6.56 NRD=0 NRS=0 m=1 r=6 sa=250000 sb=250000 a=1.5 p=7 mult=1 $X=26420 $Y=12990 $D=109
M103 PAD 27 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=28865 $Y=107610 $D=109
M104 PAD 27 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=28865 $Y=115610 $D=109
M105 29 43 VDDIO VDDIO phv L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250002 sb=250001 a=2.5 p=11 mult=1 $X=29410 $Y=35625 $D=109
M106 40 INP_SEL_H VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 r=1.66667 sa=300000 sb=300007 a=0.6 p=3.2 mult=1 $X=29250 $Y=17710 $D=109
M107 VDDIO_Q INP_SEL_H 40 VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300001 sb=300006 a=0.6 p=3.2 mult=1 $X=29250 $Y=18590 $D=109
M108 34 EN_VDDIO_SIG_H VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300002 sb=300005 a=0.6 p=3.2 mult=1 $X=29250 $Y=19470 $D=109
M109 VDDIO_Q EN_VDDIO_SIG_H 34 VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300003 sb=300004 a=0.6 p=3.2 mult=1 $X=29250 $Y=20350 $D=109
M110 XRES_H_N 72 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300003 sb=300003 a=0.6 p=3.2 mult=1 $X=29250 $Y=21230 $D=109
M111 VDDIO_Q 72 XRES_H_N VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300004 sb=300003 a=0.6 p=3.2 mult=1 $X=29250 $Y=22110 $D=109
M112 XRES_H_N 72 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300005 sb=300002 a=0.6 p=3.2 mult=1 $X=29250 $Y=22990 $D=109
M113 VDDIO_Q 72 XRES_H_N VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300006 sb=300001 a=0.6 p=3.2 mult=1 $X=29250 $Y=23870 $D=109
M114 72 41 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300007 sb=300000 a=0.6 p=3.2 mult=1 $X=29250 $Y=24750 $D=109
M115 43 71 VDDIO VDDIO phv L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 r=1.66667 sa=300000 sb=300003 a=0.6 p=3.2 mult=1 $X=29445 $Y=29045 $D=109
M116 VDDIO 71 43 VDDIO phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300001 sb=300002 a=0.6 p=3.2 mult=1 $X=29445 $Y=29925 $D=109
M117 71 DISABLE_PULLUP_H VDDIO VDDIO phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300002 sb=300001 a=0.6 p=3.2 mult=1 $X=29445 $Y=30805 $D=109
M118 VDDIO DISABLE_PULLUP_H 71 VDDIO phv L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300003 sb=300000 a=0.6 p=3.2 mult=1 $X=29445 $Y=31685 $D=109
M119 VDDIO 43 29 VDDIO phv L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250002 sb=250000 a=2.5 p=11 mult=1 $X=30190 $Y=35625 $D=109
M120 VDDIO 27 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=31015 $Y=107610 $D=109
M121 VDDIO 27 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=31015 $Y=115610 $D=109
M122 43 71 VDDIO VDDIO phv L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 r=1.66667 sa=300000 sb=300003 a=0.6 p=3.2 mult=1 $X=30785 $Y=29045 $D=109
M123 VDDIO 71 43 VDDIO phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300001 sb=300002 a=0.6 p=3.2 mult=1 $X=30785 $Y=29925 $D=109
M124 71 DISABLE_PULLUP_H VDDIO VDDIO phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300002 sb=300001 a=0.6 p=3.2 mult=1 $X=30785 $Y=30805 $D=109
M125 VDDIO DISABLE_PULLUP_H 71 VDDIO phv L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300003 sb=300000 a=0.6 p=3.2 mult=1 $X=30785 $Y=31685 $D=109
M126 PAD 27 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=33825 $Y=107610 $D=109
M127 PAD 27 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=33825 $Y=115610 $D=109
M128 XRES_H_N 72 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 r=1.66667 sa=300000 sb=300003 a=0.6 p=3.2 mult=1 $X=35355 $Y=1440 $D=109
M129 XRES_H_N 72 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 r=1.66667 sa=300000 sb=300003 a=0.6 p=3.2 mult=1 $X=35355 $Y=2780 $D=109
M130 VDDIO 27 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=35975 $Y=107610 $D=109
M131 VDDIO 27 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=35975 $Y=115610 $D=109
M132 VDDIO_Q 72 XRES_H_N VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300001 sb=300002 a=0.6 p=3.2 mult=1 $X=36235 $Y=1440 $D=109
M133 VDDIO_Q 72 XRES_H_N VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300001 sb=300002 a=0.6 p=3.2 mult=1 $X=36235 $Y=2780 $D=109
M134 XRES_H_N 72 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300002 sb=300001 a=0.6 p=3.2 mult=1 $X=37115 $Y=1440 $D=109
M135 XRES_H_N 72 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300002 sb=300001 a=0.6 p=3.2 mult=1 $X=37115 $Y=2780 $D=109
M136 VDDIO_Q 72 XRES_H_N VDDIO_Q phv L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300003 sb=300000 a=0.6 p=3.2 mult=1 $X=37995 $Y=1440 $D=109
M137 VDDIO_Q 72 XRES_H_N VDDIO_Q phv L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300003 sb=300000 a=0.6 p=3.2 mult=1 $X=37995 $Y=2780 $D=109
M138 PAD 27 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=38785 $Y=107610 $D=109
M139 PAD 27 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=38785 $Y=115610 $D=109
M140 VDDIO 46 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=40935 $Y=107610 $D=109
M141 VDDIO 46 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=40935 $Y=115610 $D=109
M142 PAD 46 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=43745 $Y=107610 $D=109
M143 PAD 46 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=43745 $Y=115610 $D=109
M144 VDDIO 46 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=45895 $Y=107610 $D=109
M145 VDDIO 46 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=45895 $Y=115610 $D=109
M146 PAD 47 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=48705 $Y=107610 $D=109
M147 PAD 47 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=48705 $Y=115610 $D=109
M148 VDDIO 47 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=50855 $Y=107610 $D=109
M149 VDDIO 47 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=50855 $Y=115610 $D=109
M150 PAD 47 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300018 a=3 p=11.2 mult=1 $X=53665 $Y=107610 $D=109
M151 PAD 47 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300018 a=3 p=11.2 mult=1 $X=53665 $Y=115610 $D=109
M152 VDDIO 48 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300016 a=3 p=11.2 mult=1 $X=55815 $Y=107610 $D=109
M153 VDDIO 48 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300016 a=3 p=11.2 mult=1 $X=55815 $Y=115610 $D=109
M154 PAD 48 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300013 a=3 p=11.2 mult=1 $X=58625 $Y=107610 $D=109
M155 PAD 48 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300013 a=3 p=11.2 mult=1 $X=58625 $Y=115610 $D=109
M156 VDDIO 48 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300011 a=3 p=11.2 mult=1 $X=60775 $Y=107610 $D=109
M157 VDDIO 48 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300011 a=3 p=11.2 mult=1 $X=60775 $Y=115610 $D=109
M158 PAD 27 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300008 a=3 p=11.2 mult=1 $X=63585 $Y=107610 $D=109
M159 PAD 27 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300008 a=3 p=11.2 mult=1 $X=63585 $Y=115610 $D=109
M160 VDDIO 49 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300006 a=3 p=11.2 mult=1 $X=65735 $Y=107610 $D=109
M161 VDDIO 49 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300006 a=3 p=11.2 mult=1 $X=65735 $Y=115610 $D=109
M162 PAD 50 VDDIO VDDIO phv L=0.6 W=5 AD=2.975 AS=3.775 PD=6.19 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300003 a=3 p=11.2 mult=1 $X=68545 $Y=107610 $D=109
M163 PAD 50 VDDIO VDDIO phv L=0.6 W=5 AD=2.975 AS=3.775 PD=6.19 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300003 a=3 p=11.2 mult=1 $X=68545 $Y=115610 $D=109
M164 VDDIO 50 PAD VDDIO phv L=0.6 W=5 AD=4.3 AS=2.975 PD=11.72 PS=6.19 NRD=17.19 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300002 a=3 p=11.2 mult=1 $X=70335 $Y=107610 $D=109
M165 VDDIO 50 PAD VDDIO phv L=0.6 W=5 AD=4.3 AS=2.975 PD=11.72 PS=6.19 NRD=17.19 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300002 a=3 p=11.2 mult=1 $X=70335 $Y=115610 $D=109
X166 VSSD 56 Dpar a=156.97 p=1082.84 m=1 $[ndiode_h] $X=8720 $Y=183570 $D=182
X167 VSSD 51 Dpar a=156.981 p=1082.92 m=1 $[ndiode_h] $X=8720 $Y=189310 $D=182
X168 VSSD VDDIO_Q Dpar a=16.2631 p=16.27 m=1 $[nwdiode] $X=7655 $Y=3340 $D=191
X169 VSSD VCCHIB Dpar a=15.5 p=17.4 m=1 $[nwdiode] $X=6050 $Y=39075 $D=191
X170 VSSD VDDIO_Q Dpar a=96.7627 p=49.03 m=1 $[nwdiode] $X=6050 $Y=19410 $D=191
X171 VSSD 24 Dpar a=23.8226 p=21.54 m=1 $[nwdiode] $X=6220 $Y=9200 $D=191
X172 VSSD 25 Dpar a=21.9076 p=21.04 m=1 $[nwdiode] $X=6220 $Y=14310 $D=191
X173 VSSD VCCHIB Dpar a=4.2823 p=8.33 m=1 $[nwdiode] $X=14430 $Y=39555 $D=191
X174 VSSD VDDIO Dpar a=108.48 p=83.5 m=1 $[nwdiode] $X=5010 $Y=47395 $D=191
X175 VSSD VDDIO_Q Dpar a=40.2643 p=30.01 m=1 $[nwdiode] $X=20935 $Y=9430 $D=191
X176 VSSD VDDIO_Q Dpar a=32.0172 p=25.17 m=1 $[nwdiode] $X=27040 $Y=17115 $D=191
X177 VSSD VDDIO Dpar a=36.4812 p=24.46 m=1 $[nwdiode] $X=26670 $Y=34430 $D=191
X178 VSSD VDDIO Dpar a=15.7043 p=15.95 m=1 $[nwdiode] $X=29110 $Y=28450 $D=191
X179 VSSD VDDIO_Q Dpar a=16.8897 p=16.63 m=1 $[nwdiode] $X=34550 $Y=610 $D=191
X180 VSSD VDDIO Dpar a=1473.41 p=184.25 m=1 $[nwdiode] $X=1735 $Y=102850 $D=191
X181 VSSD VDDIO Dpar a=735.037 p=170.75 m=1 $[nwdiode] $X=-330 $Y=130665 $D=191
R182 56 51 L=1077.19 W=0.29 m=1 $[mrdn_hv] $X=8720 $Y=183570 $D=254
R183 28 29 L=50 W=0.8 m=1 mult=1 model="mrp1" $[mrp1] $X=5800 $Y=45140 $D=257
R184 VDDIO 38 L=50 W=0.8 m=1 mult=1 model="mrp1" $[mrp1] $X=13810 $Y=131810 $D=257
R185 45 26 L=713.695 W=0.4 m=1 mult=1 model="mrp1" $[mrp1] $X=3520 $Y=87005 $D=257
R186 65 91 0.01 m=1 $[short] $X=11385 $Y=43760 $D=282
R187 91 67 0.01 m=1 $[short] $X=11575 $Y=43760 $D=282
R188 67 93 0.01 m=1 $[short] $X=18125 $Y=43760 $D=282
R189 94 70 0.01 m=1 $[short] $X=18315 $Y=43760 $D=282
R190 73 97 0.01 m=1 $[short] $X=45905 $Y=129760 $D=282
R191 98 74 0.01 m=1 $[short] $X=47415 $Y=129760 $D=282
X192 27 46 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=44185 96810 1 90 $X=44185 $Y=96810
X193 27 46 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=45395 96810 1 90 $X=45395 $Y=96810
X194 27 47 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=52095 96810 1 90 $X=52095 $Y=96810
X195 27 47 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=54480 96810 1 90 $X=54480 $Y=96810
X196 27 48 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=59920 96455 1 90 $X=59920 $Y=96455
X197 27 48 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=61125 96455 1 90 $X=61125 $Y=96455
X198 27 49 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=65335 101140 1 90 $X=65335 $Y=101140
X199 27 49 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=67745 101140 1 90 $X=67745 $Y=101140
X200 27 50 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=70030 101140 1 90 $X=70030 $Y=101140
X201 27 50 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=71215 101140 1 90 $X=71215 $Y=101140
X210 27 46 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=46570 96810 1 90 $X=46570 $Y=96810
X211 27 47 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=53305 96810 1 90 $X=53305 $Y=96810
X212 27 48 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=58710 96455 1 90 $X=58710 $Y=96455
X213 27 49 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=66560 101140 1 90 $X=66560 $Y=101140
X214 27 50 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=68805 101140 1 90 $X=68805 $Y=101140
X241 27 VDDIO sky130_fd_pr__res_generic_po__example_5595914180838 $T=60050 98360 0 0 $X=59780 $Y=98360
X242 66 PULLUP_H sky130_fd_pr__res_generic_po__example_5595914180864 $T=8510 43145 0 180 $X=6740 $Y=42345
X243 68 66 sky130_fd_pr__res_generic_po__example_5595914180864 $T=11435 43145 0 180 $X=9665 $Y=42345
X244 69 68 sky130_fd_pr__res_generic_po__example_5595914180864 $T=14215 42335 1 180 $X=12445 $Y=42335
X245 65 69 sky130_fd_pr__res_generic_po__example_5595914180864 $T=17140 42335 1 180 $X=15370 $Y=42335
X246 78 75 sky130_fd_pr__res_generic_po__example_5595914180864 $T=57830 133080 1 180 $X=56060 $Y=133080
X247 76 77 sky130_fd_pr__res_generic_po__example_5595914180864 $T=56430 130495 1 0 $X=56160 $Y=129695
X248 79 78 sky130_fd_pr__res_generic_po__example_5595914180864 $T=60755 133080 1 180 $X=58985 $Y=133080
X249 77 79 sky130_fd_pr__res_generic_po__example_5595914180864 $T=59355 130495 1 0 $X=59085 $Y=129695
X250 66 PULLUP_H sky130_fd_io__tk_em1s_cdns_5595914180859 $T=8820 43070 0 180 $X=6780 $Y=42410
X251 68 66 sky130_fd_io__tk_em1s_cdns_5595914180859 $T=11620 43070 0 180 $X=9580 $Y=42410
X252 69 68 sky130_fd_io__tk_em1s_cdns_5595914180859 $T=14565 42410 1 180 $X=12525 $Y=42410
X253 65 69 sky130_fd_io__tk_em1s_cdns_5595914180859 $T=17470 42410 1 180 $X=15430 $Y=42410
X254 74 76 sky130_fd_io__tk_em1s_cdns_5595914180859 $T=52355 130420 1 0 $X=52355 $Y=129760
X255 78 75 sky130_fd_io__tk_em1s_cdns_5595914180859 $T=58180 133155 1 180 $X=56140 $Y=133155
X256 76 77 sky130_fd_io__tk_em1s_cdns_5595914180859 $T=56245 130420 1 0 $X=56245 $Y=129760
X257 77 79 sky130_fd_io__tk_em1s_cdns_5595914180859 $T=59045 130420 1 0 $X=59045 $Y=129760
X258 79 78 sky130_fd_io__tk_em1s_cdns_5595914180859 $T=61085 133155 1 180 $X=59045 $Y=133155
X259 PAD PAD_A_ESD_H sky130_fd_io__res250only_small $T=5710 1135 0 0 $X=5710 $Y=1135
X260 TIE_WEAK_HI_H 75 sky130_fd_io__res250only_small $T=66435 137450 0 180 $X=55085 $Y=135430
X261 67 65 sky130_fd_pr__res_bent_po__example_5595914180862 $T=11875 43685 1 180 $X=5605 $Y=43685
X262 70 67 sky130_fd_pr__res_bent_po__example_5595914180862 $T=18585 43685 1 180 $X=12315 $Y=43685
X263 74 73 sky130_fd_pr__res_bent_po__example_5595914180862 $T=49010 130505 0 180 $X=42740 $Y=129705
X264 76 74 sky130_fd_pr__res_bent_po__example_5595914180862 $T=55720 130505 0 180 $X=49450 $Y=129705
X265 70 28 sky130_fd_pr__res_bent_po__example_5595914180863 $T=19445 44485 1 0 $X=19175 $Y=43685
X266 73 38 sky130_fd_pr__res_bent_po__example_5595914180863 $T=52600 133880 0 180 $X=40330 $Y=133080
X269 VSSD VDDIO_Q 80 42 81 82 83 84 85 86 87 88 89 92 sky130_fd_io__xres2v2_rcfilter_lpfv2 $T=73595 4860 0 90 $X=33055 $Y=6020
X301 VDDIO_Q INP_SEL_H 52 92 sky130_fd_pr__pfet_01v8__example_55959141808767 $T=21265 10040 1 90 $X=20935 $Y=9430
X302 VDDIO_Q 40 92 FILT_IN_H sky130_fd_pr__pfet_01v8__example_55959141808767 $T=21265 11470 1 90 $X=20935 $Y=10860
X303 VSSIO TIE_LO_ESD sky130_fd_io__tk_tie_r_out_esd $T=17060 2635 0 0 $X=17450 $Y=3730
X304 VDDIO TIE_HI_ESD sky130_fd_io__tk_tie_r_out_esd $T=17060 3875 0 0 $X=17450 $Y=4970
X305 VSSD 40 52 92 sky130_fd_pr__nfet_01v8__example_55959141808764 $T=20005 10040 0 90 $X=16825 $Y=9580
X306 VSSD INP_SEL_H 92 FILT_IN_H sky130_fd_pr__nfet_01v8__example_55959141808764 $T=20005 11470 0 90 $X=16825 $Y=11010
X307 VSSD 30 64 58 sky130_fd_pr__nfet_01v8__example_55959141808779 $T=13635 35115 1 90 $X=13455 $Y=34655
X308 VSSD 35 59 25 sky130_fd_pr__nfet_01v8__example_55959141808779 $T=16525 17790 1 270 $X=15345 $Y=16430
X309 VSSD 32 31 sky130_fd_pr__nfet_01v8__example_55959141808777 $T=18315 20005 1 270 $X=15135 $Y=19045
X310 VSSD 37 39 sky130_fd_pr__nfet_01v8__example_55959141808777 $T=18390 25165 1 270 $X=15210 $Y=24205
X311 VSSD ENABLE_H 55 sky130_fd_pr__nfet_01v8__example_55959141808777 $T=18390 26580 1 270 $X=15210 $Y=25620
X327 24 24 24 sky130_fd_pr__pfet_01v8__example_55959141808784 $T=8380 11155 1 270 $X=7050 $Y=9745
X328 24 30 37 sky130_fd_pr__pfet_01v8__example_55959141808784 $T=10910 10355 0 90 $X=9580 $Y=9745
X348 VSSD VDDIO VSSD 30 PAD sky130_fd_io__gpio_buf_localesdv2 $T=4630 70965 1 0 $X=4923 $Y=47395
X351 VSSD 99 VSSIO VDDIO 99 99 90 PAD sky130_fd_io__gpio_pddrvr_strong_xres4v2 $T=0 184810 1 0 $X=-515 $Y=137270
.ENDS
***************************************
.SUBCKT ICV_2 VSSD VSSIO VCCD VDDIO VSSD_PAD
** N=13 EP=5 IP=20 FDC=501
*.CALIBRE ISOLATED NETS: VCCHIB VDDA VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
X0 VSSD VSSD VSSD VCCD VDDIO VCCD VSSIO VSSD VSSD_PAD sky130_fd_io__top_ground_lvc_wpad $T=0 -35 0 0 $X=0 $Y=-35
.ENDS
***************************************
.SUBCKT ICV_3 VSSD VSSIO VCCD VDDIO VCCD_PAD
** N=13 EP=5 IP=20 FDC=501
*.CALIBRE ISOLATED NETS: VCCHIB VDDA VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
X0 VSSD VSSD VSSD VCCD VDDIO VCCD VSSIO VCCD VCCD_PAD sky130_fd_io__top_power_lvc_wpad $T=0 -35 0 0 $X=0 $Y=-35
.ENDS
***************************************
.SUBCKT chip_io mprj_io_oeb[24] mprj_io_ib_mode_sel[24] mprj_io_vtrip_sel[24] mprj_io_out[24] mprj_io_holdover[24] mprj_io_dm[74] mprj_io_analog_sel[24] mprj_io_hldh_n[24] mprj_io_enh[24] mprj_io_inp_dis[24] mprj_io_analog_pol[24] mprj_io_dm[72] mprj_io_analog_en[24] mprj_io_dm[73] mprj_analog_io[17] mprj_io_slow_sel[24] mprj_io_in[24] porb_h mprj_io_oeb[23] mprj_io_ib_mode_sel[23]
+ mprj_io_vtrip_sel[23] mprj_io_out[23] mprj_io_holdover[23] mprj_io_dm[71] mprj_io_analog_sel[23] mprj_io_hldh_n[23] mprj_io_enh[23] mprj_io_inp_dis[23] mprj_io_analog_pol[23] mprj_io_dm[69] mprj_io_analog_en[23] mprj_io_dm[70] mprj_analog_io[16] mprj_io_slow_sel[23] mprj_io_in[23] mprj_io_oeb[22] mprj_io_ib_mode_sel[22] mprj_io_vtrip_sel[22] mprj_io_out[22] mprj_io_holdover[22]
+ mprj_io_dm[68] mprj_io_analog_sel[22] mprj_io_hldh_n[22] mprj_io_enh[22] mprj_io_inp_dis[22] mprj_io_analog_pol[22] mprj_io_dm[66] mprj_io_analog_en[22] mprj_io_dm[67] mprj_analog_io[15] mprj_io_slow_sel[22] mprj_io_in[22] mprj_io_oeb[21] mprj_io_ib_mode_sel[21] mprj_io_vtrip_sel[21] mprj_io_out[21] mprj_io_holdover[21] mprj_io_dm[65] mprj_io_analog_sel[21] mprj_io_hldh_n[21]
+ mprj_io_enh[21] mprj_io_inp_dis[21] mprj_io_analog_pol[21] mprj_io_dm[63] mprj_io_analog_en[21] mprj_io_dm[64] mprj_analog_io[14] mprj_io_slow_sel[21] mprj_io_in[21] mprj_io_oeb[20] mprj_io_ib_mode_sel[20] mprj_io_vtrip_sel[20] mprj_io_out[20] mprj_io_holdover[20] mprj_io_dm[62] mprj_io_analog_sel[20] mprj_io_hldh_n[20] mprj_io_enh[20] mprj_io_inp_dis[20] mprj_io_analog_pol[20]
+ mprj_io_dm[60] mprj_io_analog_en[20] mprj_io_dm[61] mprj_analog_io[13] mprj_io_slow_sel[20] mprj_io_in[20] mprj_io_oeb[19] mprj_io_ib_mode_sel[19] mprj_io_vtrip_sel[19] mprj_io_out[19] mprj_io_holdover[19] mprj_io_dm[59] mprj_io_analog_sel[19] mprj_io_hldh_n[19] mprj_io_enh[19] mprj_io_inp_dis[19] mprj_io_analog_pol[19] mprj_io_dm[57] mprj_io_analog_en[19] mprj_io_dm[58]
+ mprj_analog_io[12] mprj_io_slow_sel[19] mprj_io_in[19] mprj_io_oeb[18] mprj_io_ib_mode_sel[18] mprj_io_vtrip_sel[18] mprj_io_out[18] mprj_io_holdover[18] mprj_io_dm[56] mprj_io_analog_sel[18] mprj_io_hldh_n[18] mprj_io_enh[18] mprj_io_inp_dis[18] mprj_io_analog_pol[18] mprj_io_dm[54] mprj_io_analog_en[18] mprj_io_dm[55] mprj_analog_io[11] mprj_io_slow_sel[18] mprj_io_in[18]
+ mprj_io_oeb[17] mprj_io_ib_mode_sel[17] mprj_io_vtrip_sel[17] mprj_io_out[17] mprj_io_holdover[17] mprj_io_dm[53] mprj_io_analog_sel[17] mprj_io_hldh_n[17] mprj_io_enh[17] mprj_io_inp_dis[17] mprj_io_analog_pol[17] mprj_io_dm[51] mprj_io_analog_en[17] mprj_io_dm[52] mprj_analog_io[10] mprj_io_slow_sel[17] mprj_io_in[17] mprj_io_oeb[16] mprj_io_ib_mode_sel[16] mprj_io_vtrip_sel[16]
+ mprj_io_out[16] mprj_io_holdover[16] mprj_io_dm[50] mprj_io_analog_sel[16] mprj_io_hldh_n[16] mprj_io_enh[16] mprj_io_inp_dis[16] mprj_io_analog_pol[16] mprj_io_dm[48] mprj_io_analog_en[16] mprj_io_dm[49] mprj_analog_io[9] mprj_io_slow_sel[16] mprj_io_in[16] mprj_io_oeb[15] mprj_io_ib_mode_sel[15] mprj_io_vtrip_sel[15] mprj_io_out[15] mprj_io_holdover[15] mprj_io_dm[47]
+ mprj_io_analog_sel[15] mprj_io_hldh_n[15] mprj_io_enh[15] mprj_io_inp_dis[15] mprj_io_analog_pol[15] mprj_io_dm[45] mprj_io_analog_en[15] mprj_io_dm[46] mprj_analog_io[8] mprj_io_slow_sel[15] mprj_io_in[15] mprj_io_in[14] mprj_io_slow_sel[14] mprj_analog_io[7] mprj_io_dm[43] mprj_io_analog_en[14] mprj_io_dm[42] mprj_io_analog_pol[14] mprj_io_inp_dis[14] mprj_io_enh[14]
+ mprj_io_hldh_n[14] mprj_io_analog_sel[14] mprj_io_dm[44] mprj_io_holdover[14] mprj_io_out[14] mprj_io_vtrip_sel[14] mprj_io_ib_mode_sel[14] mprj_io_oeb[14] mprj_io_in[13] mprj_io_slow_sel[13] mprj_analog_io[6] mprj_io_dm[40] mprj_io_analog_en[13] mprj_io_dm[39] mprj_io_analog_pol[13] mprj_io_inp_dis[13] mprj_io_enh[13] mprj_io_hldh_n[13] mprj_io_analog_sel[13] mprj_io_dm[41]
+ mprj_io_holdover[13] mprj_io_out[13] mprj_io_vtrip_sel[13] mprj_io_ib_mode_sel[13] mprj_io_oeb[13] mprj_io_oeb[31] mprj_io_ib_mode_sel[31] mprj_io_vtrip_sel[31] mprj_io_out[31] mprj_io_holdover[31] mprj_io_dm[95] mprj_io_analog_sel[31] mprj_io_hldh_n[31] mprj_io_enh[31] mprj_io_inp_dis[31] mprj_io_analog_pol[31] mprj_io_dm[93] mprj_io_analog_en[31] mprj_io_dm[94] mprj_analog_io[24]
+ mprj_io_slow_sel[31] mprj_io_in[31] mprj_io_oeb[30] mprj_io_ib_mode_sel[30] mprj_io_vtrip_sel[30] mprj_io_out[30] mprj_io_holdover[30] mprj_io_dm[92] mprj_io_analog_sel[30] mprj_io_hldh_n[30] mprj_io_enh[30] mprj_io_inp_dis[30] mprj_io_analog_pol[30] mprj_io_dm[90] mprj_io_analog_en[30] mprj_io_dm[91] mprj_analog_io[23] mprj_io_slow_sel[30] mprj_io_in[30] mprj_io_oeb[29]
+ mprj_io_ib_mode_sel[29] mprj_io_vtrip_sel[29] mprj_io_out[29] mprj_io_holdover[29] mprj_io_dm[89] mprj_io_analog_sel[29] mprj_io_hldh_n[29] mprj_io_enh[29] mprj_io_inp_dis[29] mprj_io_analog_pol[29] mprj_io_dm[87] mprj_io_analog_en[29] mprj_io_dm[88] mprj_analog_io[22] mprj_io_slow_sel[29] mprj_io_in[29] mprj_io_oeb[28] mprj_io_ib_mode_sel[28] mprj_io_vtrip_sel[28] mprj_io_out[28]
+ mprj_io_holdover[28] mprj_io_dm[86] mprj_io_analog_sel[28] mprj_io_hldh_n[28] mprj_io_enh[28] mprj_io_inp_dis[28] mprj_io_analog_pol[28] mprj_io_dm[84] mprj_io_analog_en[28] mprj_io_dm[85] mprj_analog_io[21] mprj_io_slow_sel[28] mprj_io_in[28] mprj_io_oeb[27] mprj_io_ib_mode_sel[27] mprj_io_vtrip_sel[27] mprj_io_out[27] mprj_io_holdover[27] mprj_io_dm[83] mprj_io_analog_sel[27]
+ mprj_io_hldh_n[27] mprj_io_enh[27] mprj_io_inp_dis[27] mprj_io_analog_pol[27] mprj_io_dm[81] mprj_io_analog_en[27] mprj_io_dm[82] mprj_analog_io[20] mprj_io_slow_sel[27] mprj_io_in[27] mprj_io_oeb[26] mprj_io_ib_mode_sel[26] mprj_io_vtrip_sel[26] mprj_io_out[26] mprj_io_holdover[26] mprj_io_dm[80] mprj_io_analog_sel[26] mprj_io_hldh_n[26] mprj_io_enh[26] mprj_io_inp_dis[26]
+ mprj_io_analog_pol[26] mprj_io_dm[78] mprj_io_analog_en[26] mprj_io_dm[79] mprj_analog_io[19] mprj_io_slow_sel[26] mprj_io_in[26] mprj_io_oeb[25] mprj_io_ib_mode_sel[25] mprj_io_vtrip_sel[25] mprj_io_out[25] mprj_io_holdover[25] mprj_io_dm[77] mprj_io_analog_sel[25] mprj_io_hldh_n[25] mprj_io_enh[25] mprj_io_inp_dis[25] mprj_io_analog_pol[25] mprj_io_dm[75] mprj_io_analog_en[25]
+ mprj_io_dm[76] mprj_analog_io[18] mprj_io_slow_sel[25] mprj_io_in[25] mprj_io_in[7] mprj_io_slow_sel[7] mprj_analog_io[0] mprj_io_dm[22] mprj_io_analog_en[7] mprj_io_dm[21] mprj_io_analog_pol[7] mprj_io_inp_dis[7] mprj_io_enh[7] mprj_io_hldh_n[7] mprj_io_analog_sel[7] mprj_io_dm[23] mprj_io_holdover[7] mprj_io_out[7] mprj_io_vtrip_sel[7] mprj_io_ib_mode_sel[7]
+ mprj_io_oeb[7] mprj_io_in[8] mprj_io_slow_sel[8] mprj_analog_io[1] mprj_io_dm[25] mprj_io_analog_en[8] mprj_io_dm[24] mprj_io_analog_pol[8] mprj_io_inp_dis[8] mprj_io_enh[8] mprj_io_hldh_n[8] mprj_io_analog_sel[8] mprj_io_dm[26] mprj_io_holdover[8] mprj_io_out[8] mprj_io_vtrip_sel[8] mprj_io_ib_mode_sel[8] mprj_io_oeb[8] mprj_io_in[9] mprj_io_slow_sel[9]
+ mprj_analog_io[2] mprj_io_dm[28] mprj_io_analog_en[9] mprj_io_dm[27] mprj_io_analog_pol[9] mprj_io_inp_dis[9] mprj_io_enh[9] mprj_io_hldh_n[9] mprj_io_analog_sel[9] mprj_io_dm[29] mprj_io_holdover[9] mprj_io_out[9] mprj_io_vtrip_sel[9] mprj_io_ib_mode_sel[9] mprj_io_oeb[9] mprj_io_in[10] mprj_io_slow_sel[10] mprj_analog_io[3] mprj_io_dm[31] mprj_io_analog_en[10]
+ mprj_io_dm[30] mprj_io_analog_pol[10] mprj_io_inp_dis[10] mprj_io_enh[10] mprj_io_hldh_n[10] mprj_io_analog_sel[10] mprj_io_dm[32] mprj_io_holdover[10] mprj_io_out[10] mprj_io_vtrip_sel[10] mprj_io_ib_mode_sel[10] mprj_io_oeb[10] mprj_io_in[11] mprj_io_slow_sel[11] mprj_analog_io[4] mprj_io_dm[34] mprj_io_analog_en[11] mprj_io_dm[33] mprj_io_analog_pol[11] mprj_io_inp_dis[11]
+ mprj_io_enh[11] mprj_io_hldh_n[11] mprj_io_analog_sel[11] mprj_io_dm[35] mprj_io_holdover[11] mprj_io_out[11] mprj_io_vtrip_sel[11] mprj_io_ib_mode_sel[11] mprj_io_oeb[11] mprj_io_in[12] mprj_io_slow_sel[12] mprj_analog_io[5] mprj_io_dm[37] mprj_io_analog_en[12] mprj_io_dm[36] mprj_io_analog_pol[12] mprj_io_inp_dis[12] mprj_io_enh[12] mprj_io_hldh_n[12] mprj_io_analog_sel[12]
+ mprj_io_dm[38] mprj_io_holdover[12] mprj_io_out[12] mprj_io_vtrip_sel[12] mprj_io_ib_mode_sel[12] mprj_io_oeb[12] mprj_io_oeb[37] mprj_io_ib_mode_sel[37] mprj_io_vtrip_sel[37] mprj_io_out[37] mprj_io_holdover[37] mprj_io_dm[113] mprj_io_analog_sel[37] mprj_io_hldh_n[37] mprj_io_enh[37] mprj_io_inp_dis[37] mprj_io_analog_pol[37] mprj_io_dm[111] mprj_io_analog_en[37] mprj_io_dm[112]
+ mprj_io_slow_sel[37] mprj_io_in[37] mprj_io_oeb[36] mprj_io_ib_mode_sel[36] mprj_io_vtrip_sel[36] mprj_io_out[36] mprj_io_holdover[36] mprj_io_dm[110] mprj_io_analog_sel[36] mprj_io_hldh_n[36] mprj_io_enh[36] mprj_io_inp_dis[36] mprj_io_analog_pol[36] mprj_io_dm[108] mprj_io_analog_en[36] mprj_io_dm[109] mprj_io_slow_sel[36] mprj_io_in[36] mprj_io_oeb[35] mprj_io_ib_mode_sel[35]
+ mprj_io_vtrip_sel[35] mprj_io_out[35] mprj_io_holdover[35] mprj_io_dm[107] mprj_io_analog_sel[35] mprj_io_hldh_n[35] mprj_io_enh[35] mprj_io_inp_dis[35] mprj_io_analog_pol[35] mprj_io_dm[105] mprj_io_analog_en[35] mprj_io_dm[106] mprj_analog_io[28] mprj_io_slow_sel[35] mprj_io_in[35] mprj_io_oeb[34] mprj_io_ib_mode_sel[34] mprj_io_vtrip_sel[34] mprj_io_out[34] mprj_io_holdover[34]
+ mprj_io_dm[104] mprj_io_analog_sel[34] mprj_io_hldh_n[34] mprj_io_enh[34] mprj_io_inp_dis[34] mprj_io_analog_pol[34] mprj_io_dm[102] mprj_io_analog_en[34] mprj_io_dm[103] mprj_analog_io[27] mprj_io_slow_sel[34] mprj_io_in[34] mprj_io_oeb[33] mprj_io_ib_mode_sel[33] mprj_io_vtrip_sel[33] mprj_io_out[33] mprj_io_holdover[33] mprj_io_dm[101] mprj_io_analog_sel[33] mprj_io_hldh_n[33]
+ mprj_io_enh[33] mprj_io_inp_dis[33] mprj_io_analog_pol[33] mprj_io_dm[99] mprj_io_analog_en[33] mprj_io_dm[100] mprj_analog_io[26] mprj_io_slow_sel[33] mprj_io_in[33] mprj_io_oeb[32] mprj_io_ib_mode_sel[32] mprj_io_vtrip_sel[32] mprj_io_out[32] mprj_io_holdover[32] mprj_io_dm[98] mprj_io_analog_sel[32] mprj_io_hldh_n[32] mprj_io_enh[32] mprj_io_inp_dis[32] mprj_io_analog_pol[32]
+ mprj_io_dm[96] mprj_io_analog_en[32] mprj_io_dm[97] mprj_analog_io[25] mprj_io_slow_sel[32] mprj_io_in[32] mprj_io_in[0] mprj_io_slow_sel[0] mprj_io_dm[1] mprj_io_analog_en[0] mprj_io_dm[0] mprj_io_analog_pol[0] mprj_io_inp_dis[0] mprj_io_enh[0] mprj_io_hldh_n[0] mprj_io_analog_sel[0] mprj_io_dm[2] mprj_io_holdover[0] mprj_io_out[0] mprj_io_vtrip_sel[0]
+ mprj_io_ib_mode_sel[0] mprj_io_oeb[0] mprj_io_in[1] mprj_io_slow_sel[1] mprj_io_dm[4] mprj_io_analog_en[1] mprj_io_dm[3] mprj_io_analog_pol[1] mprj_io_inp_dis[1] mprj_io_enh[1] mprj_io_hldh_n[1] mprj_io_analog_sel[1] mprj_io_dm[5] mprj_io_holdover[1] mprj_io_out[1] mprj_io_vtrip_sel[1] mprj_io_ib_mode_sel[1] mprj_io_oeb[1] mprj_io_in[2] mprj_io_slow_sel[2]
+ mprj_io_dm[7] mprj_io_analog_en[2] mprj_io_dm[6] mprj_io_analog_pol[2] mprj_io_inp_dis[2] mprj_io_enh[2] mprj_io_hldh_n[2] mprj_io_analog_sel[2] mprj_io_dm[8] mprj_io_holdover[2] mprj_io_out[2] mprj_io_vtrip_sel[2] mprj_io_ib_mode_sel[2] mprj_io_oeb[2] mprj_io_in[3] mprj_io_slow_sel[3] mprj_io_dm[10] mprj_io_analog_en[3] mprj_io_dm[9] mprj_io_analog_pol[3]
+ mprj_io_inp_dis[3] mprj_io_enh[3] mprj_io_hldh_n[3] mprj_io_analog_sel[3] mprj_io_dm[11] mprj_io_holdover[3] mprj_io_out[3] mprj_io_vtrip_sel[3] mprj_io_ib_mode_sel[3] mprj_io_oeb[3] mprj_io_in[4] mprj_io_slow_sel[4] mprj_io_dm[13] mprj_io_analog_en[4] mprj_io_dm[12] mprj_io_analog_pol[4] mprj_io_inp_dis[4] mprj_io_enh[4] mprj_io_hldh_n[4] mprj_io_analog_sel[4]
+ mprj_io_dm[14] mprj_io_holdover[4] mprj_io_out[4] mprj_io_vtrip_sel[4] mprj_io_ib_mode_sel[4] mprj_io_oeb[4] mprj_io_in[5] mprj_io_slow_sel[5] mprj_io_dm[16] mprj_io_analog_en[5] mprj_io_dm[15] mprj_io_analog_pol[5] mprj_io_inp_dis[5] mprj_io_enh[5] mprj_io_hldh_n[5] mprj_io_analog_sel[5] mprj_io_dm[17] mprj_io_holdover[5] mprj_io_out[5] mprj_io_vtrip_sel[5]
+ mprj_io_ib_mode_sel[5] mprj_io_oeb[5] mprj_io_in[6] mprj_io_slow_sel[6] mprj_io_dm[19] mprj_io_analog_en[6] mprj_io_dm[18] mprj_io_analog_pol[6] mprj_io_inp_dis[6] mprj_io_enh[6] mprj_io_hldh_n[6] mprj_io_analog_sel[6] mprj_io_dm[20] mprj_io_holdover[6] mprj_io_out[6] mprj_io_vtrip_sel[6] mprj_io_ib_mode_sel[6] mprj_io_oeb[6] clock_core por
+ flash_csb_ieb_core flash_csb_core flash_csb_oeb_core flash_clk_ieb_core flash_clk_core flash_clk_oeb_core flash_io0_di_core flash_io0_ieb_core flash_io0_do_core flash_io0_oeb_core flash_io1_di_core flash_io1_ieb_core flash_io1_do_core flash_io1_oeb_core gpio_in_core gpio_mode0_core gpio_inenb_core gpio_mode1_core gpio_out_core gpio_outenb_core
+ resetb_core_h mprj_io[24] vccd2_pad mprj_io[23] mprj_io[22] mprj_io[21] mprj_io[20] mprj_io[19] vssio_pad mprj_io[18] mprj_io[17] mprj_io[16] vssa1_pad mprj_io[15] vccd1_pad mprj_io[14] mprj_io[13] mprj_io[31] mprj_io[30] mprj_io[29]
+ mprj_io[28] mprj_io[27] mprj_io[26] mprj_io[25] vssa2_pad vdda1_pad mprj_io[7] mprj_io[8] mprj_io[9] mprj_io[10] mprj_io[11] mprj_io[12] vssd2_pad vdda2_pad vssd1_pad mprj_io[37] mprj_io[36] mprj_io[35] mprj_io[34] mprj_io[33]
+ mprj_io[32] vddio_pad mprj_io[0] mprj_io[1] mprj_io[2] mprj_io[3] mprj_io[4] mprj_io[5] mprj_io[6] vssa_pad clock flash_csb flash_clk flash_io0 flash_io1 gpio vdda_pad resetb vssd_pad vccd_pad
** N=735 EP=720 IP=844 FDC=6675
X0 1 193 Dpar a=57.3765 p=0 m=1 $[nwdiode] $X=662380 $Y=29790 $D=189
X1 1 2 175 669 193 673 330 674 vccd2_pad vssio_pad vssa1_pad vccd1_pad ICV_13 $T=0 0 0 0 $X=0 $Y=4526800
X2 1 2 193 ICV_14 $T=0 0 0 0 $X=0 $Y=4213000
X3 1 330 193 175 669 672 vssa2_pad vdda1_pad ICV_15 $T=0 0 0 0 $X=0 $Y=2594000
X4 1 330 2 193 175 672 669 673 674 vssd2_pad vdda2_pad vssd1_pad ICV_16 $T=0 0 0 0 $X=0 $Y=2204000
X5 1 2 175 193 330 vddio_pad ICV_17 $T=0 0 0 0 $X=0 $Y=426200
X6 1 2 193 675 676 vssa_pad vdda_pad ICV_18 $T=0 0 0 0 $X=0 $Y=0
X7 1 193 174 193 porb_h 2 2 174 resetb 2 2 645 2 2 resetb_core_h 645 ICV_1 $T=738000 200000 0 180 $X=662380 $Y=0
X8 1 2 174 193 vssd_pad ICV_2 $T=1281000 197965 0 180 $X=1194860 $Y=0
X9 1 2 174 193 vccd_pad ICV_3 $T=197965 340000 0 90 $X=0 $Y=329025
.ENDS
***************************************
