VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_protect
  CLASS BLOCK ;
  FOREIGN mgmt_protect ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 90.000 ;
  PIN caravel_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 15.000 0.300 15.600 ;
    END
  END caravel_clk
  PIN caravel_clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 44.920 0.300 45.520 ;
    END
  END caravel_clk2
  PIN caravel_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 74.840 0.300 75.440 ;
    END
  END caravel_rstn
  PIN la_data_in_core[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 89.700 9.570 92.000 ;
    END
  END la_data_in_core[0]
  PIN la_data_in_core[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 89.700 227.610 92.000 ;
    END
  END la_data_in_core[100]
  PIN la_data_in_core[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 89.700 229.910 92.000 ;
    END
  END la_data_in_core[101]
  PIN la_data_in_core[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 89.700 232.210 92.000 ;
    END
  END la_data_in_core[102]
  PIN la_data_in_core[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 89.700 234.050 92.000 ;
    END
  END la_data_in_core[103]
  PIN la_data_in_core[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 89.700 236.350 92.000 ;
    END
  END la_data_in_core[104]
  PIN la_data_in_core[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 89.700 238.650 92.000 ;
    END
  END la_data_in_core[105]
  PIN la_data_in_core[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 89.700 240.950 92.000 ;
    END
  END la_data_in_core[106]
  PIN la_data_in_core[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 89.700 242.790 92.000 ;
    END
  END la_data_in_core[107]
  PIN la_data_in_core[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 89.700 245.090 92.000 ;
    END
  END la_data_in_core[108]
  PIN la_data_in_core[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 89.700 247.390 92.000 ;
    END
  END la_data_in_core[109]
  PIN la_data_in_core[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 89.700 31.650 92.000 ;
    END
  END la_data_in_core[10]
  PIN la_data_in_core[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 89.700 249.230 92.000 ;
    END
  END la_data_in_core[110]
  PIN la_data_in_core[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 89.700 251.530 92.000 ;
    END
  END la_data_in_core[111]
  PIN la_data_in_core[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 89.700 253.830 92.000 ;
    END
  END la_data_in_core[112]
  PIN la_data_in_core[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 89.700 256.130 92.000 ;
    END
  END la_data_in_core[113]
  PIN la_data_in_core[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 89.700 257.970 92.000 ;
    END
  END la_data_in_core[114]
  PIN la_data_in_core[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 89.700 260.270 92.000 ;
    END
  END la_data_in_core[115]
  PIN la_data_in_core[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 89.700 262.570 92.000 ;
    END
  END la_data_in_core[116]
  PIN la_data_in_core[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 89.700 264.870 92.000 ;
    END
  END la_data_in_core[117]
  PIN la_data_in_core[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 89.700 266.710 92.000 ;
    END
  END la_data_in_core[118]
  PIN la_data_in_core[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 89.700 269.010 92.000 ;
    END
  END la_data_in_core[119]
  PIN la_data_in_core[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 89.700 33.950 92.000 ;
    END
  END la_data_in_core[11]
  PIN la_data_in_core[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 89.700 271.310 92.000 ;
    END
  END la_data_in_core[120]
  PIN la_data_in_core[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 89.700 273.610 92.000 ;
    END
  END la_data_in_core[121]
  PIN la_data_in_core[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 89.700 275.450 92.000 ;
    END
  END la_data_in_core[122]
  PIN la_data_in_core[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 89.700 277.750 92.000 ;
    END
  END la_data_in_core[123]
  PIN la_data_in_core[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 89.700 280.050 92.000 ;
    END
  END la_data_in_core[124]
  PIN la_data_in_core[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 89.700 281.890 92.000 ;
    END
  END la_data_in_core[125]
  PIN la_data_in_core[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 89.700 284.190 92.000 ;
    END
  END la_data_in_core[126]
  PIN la_data_in_core[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 89.700 286.490 92.000 ;
    END
  END la_data_in_core[127]
  PIN la_data_in_core[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 89.700 35.790 92.000 ;
    END
  END la_data_in_core[12]
  PIN la_data_in_core[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 89.700 38.090 92.000 ;
    END
  END la_data_in_core[13]
  PIN la_data_in_core[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 89.700 40.390 92.000 ;
    END
  END la_data_in_core[14]
  PIN la_data_in_core[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 89.700 42.230 92.000 ;
    END
  END la_data_in_core[15]
  PIN la_data_in_core[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 89.700 44.530 92.000 ;
    END
  END la_data_in_core[16]
  PIN la_data_in_core[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 89.700 46.830 92.000 ;
    END
  END la_data_in_core[17]
  PIN la_data_in_core[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 89.700 49.130 92.000 ;
    END
  END la_data_in_core[18]
  PIN la_data_in_core[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 89.700 50.970 92.000 ;
    END
  END la_data_in_core[19]
  PIN la_data_in_core[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 89.700 11.870 92.000 ;
    END
  END la_data_in_core[1]
  PIN la_data_in_core[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 89.700 53.270 92.000 ;
    END
  END la_data_in_core[20]
  PIN la_data_in_core[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 89.700 55.570 92.000 ;
    END
  END la_data_in_core[21]
  PIN la_data_in_core[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 89.700 57.870 92.000 ;
    END
  END la_data_in_core[22]
  PIN la_data_in_core[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 89.700 59.710 92.000 ;
    END
  END la_data_in_core[23]
  PIN la_data_in_core[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 89.700 62.010 92.000 ;
    END
  END la_data_in_core[24]
  PIN la_data_in_core[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 89.700 64.310 92.000 ;
    END
  END la_data_in_core[25]
  PIN la_data_in_core[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 89.700 66.610 92.000 ;
    END
  END la_data_in_core[26]
  PIN la_data_in_core[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 89.700 68.450 92.000 ;
    END
  END la_data_in_core[27]
  PIN la_data_in_core[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 89.700 70.750 92.000 ;
    END
  END la_data_in_core[28]
  PIN la_data_in_core[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 89.700 73.050 92.000 ;
    END
  END la_data_in_core[29]
  PIN la_data_in_core[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 89.700 14.170 92.000 ;
    END
  END la_data_in_core[2]
  PIN la_data_in_core[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 89.700 75.350 92.000 ;
    END
  END la_data_in_core[30]
  PIN la_data_in_core[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 89.700 77.190 92.000 ;
    END
  END la_data_in_core[31]
  PIN la_data_in_core[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 89.700 79.490 92.000 ;
    END
  END la_data_in_core[32]
  PIN la_data_in_core[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 89.700 81.790 92.000 ;
    END
  END la_data_in_core[33]
  PIN la_data_in_core[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 89.700 83.630 92.000 ;
    END
  END la_data_in_core[34]
  PIN la_data_in_core[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 89.700 85.930 92.000 ;
    END
  END la_data_in_core[35]
  PIN la_data_in_core[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 89.700 88.230 92.000 ;
    END
  END la_data_in_core[36]
  PIN la_data_in_core[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 89.700 90.530 92.000 ;
    END
  END la_data_in_core[37]
  PIN la_data_in_core[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 89.700 92.370 92.000 ;
    END
  END la_data_in_core[38]
  PIN la_data_in_core[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 89.700 94.670 92.000 ;
    END
  END la_data_in_core[39]
  PIN la_data_in_core[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 89.700 16.470 92.000 ;
    END
  END la_data_in_core[3]
  PIN la_data_in_core[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 89.700 96.970 92.000 ;
    END
  END la_data_in_core[40]
  PIN la_data_in_core[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 89.700 99.270 92.000 ;
    END
  END la_data_in_core[41]
  PIN la_data_in_core[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 89.700 101.110 92.000 ;
    END
  END la_data_in_core[42]
  PIN la_data_in_core[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 89.700 103.410 92.000 ;
    END
  END la_data_in_core[43]
  PIN la_data_in_core[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 89.700 105.710 92.000 ;
    END
  END la_data_in_core[44]
  PIN la_data_in_core[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 89.700 108.010 92.000 ;
    END
  END la_data_in_core[45]
  PIN la_data_in_core[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 89.700 109.850 92.000 ;
    END
  END la_data_in_core[46]
  PIN la_data_in_core[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 89.700 112.150 92.000 ;
    END
  END la_data_in_core[47]
  PIN la_data_in_core[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 89.700 114.450 92.000 ;
    END
  END la_data_in_core[48]
  PIN la_data_in_core[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 89.700 116.750 92.000 ;
    END
  END la_data_in_core[49]
  PIN la_data_in_core[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 89.700 18.310 92.000 ;
    END
  END la_data_in_core[4]
  PIN la_data_in_core[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 89.700 118.590 92.000 ;
    END
  END la_data_in_core[50]
  PIN la_data_in_core[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 89.700 120.890 92.000 ;
    END
  END la_data_in_core[51]
  PIN la_data_in_core[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 89.700 123.190 92.000 ;
    END
  END la_data_in_core[52]
  PIN la_data_in_core[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 89.700 125.030 92.000 ;
    END
  END la_data_in_core[53]
  PIN la_data_in_core[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 89.700 127.330 92.000 ;
    END
  END la_data_in_core[54]
  PIN la_data_in_core[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 89.700 129.630 92.000 ;
    END
  END la_data_in_core[55]
  PIN la_data_in_core[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 89.700 131.930 92.000 ;
    END
  END la_data_in_core[56]
  PIN la_data_in_core[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 89.700 133.770 92.000 ;
    END
  END la_data_in_core[57]
  PIN la_data_in_core[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 89.700 136.070 92.000 ;
    END
  END la_data_in_core[58]
  PIN la_data_in_core[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 89.700 138.370 92.000 ;
    END
  END la_data_in_core[59]
  PIN la_data_in_core[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 89.700 20.610 92.000 ;
    END
  END la_data_in_core[5]
  PIN la_data_in_core[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 89.700 140.670 92.000 ;
    END
  END la_data_in_core[60]
  PIN la_data_in_core[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 89.700 142.510 92.000 ;
    END
  END la_data_in_core[61]
  PIN la_data_in_core[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 89.700 144.810 92.000 ;
    END
  END la_data_in_core[62]
  PIN la_data_in_core[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 89.700 147.110 92.000 ;
    END
  END la_data_in_core[63]
  PIN la_data_in_core[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 89.700 149.410 92.000 ;
    END
  END la_data_in_core[64]
  PIN la_data_in_core[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 89.700 151.250 92.000 ;
    END
  END la_data_in_core[65]
  PIN la_data_in_core[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 89.700 153.550 92.000 ;
    END
  END la_data_in_core[66]
  PIN la_data_in_core[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 89.700 155.850 92.000 ;
    END
  END la_data_in_core[67]
  PIN la_data_in_core[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 89.700 158.150 92.000 ;
    END
  END la_data_in_core[68]
  PIN la_data_in_core[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 89.700 159.990 92.000 ;
    END
  END la_data_in_core[69]
  PIN la_data_in_core[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 89.700 22.910 92.000 ;
    END
  END la_data_in_core[6]
  PIN la_data_in_core[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 89.700 162.290 92.000 ;
    END
  END la_data_in_core[70]
  PIN la_data_in_core[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 89.700 164.590 92.000 ;
    END
  END la_data_in_core[71]
  PIN la_data_in_core[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 89.700 166.430 92.000 ;
    END
  END la_data_in_core[72]
  PIN la_data_in_core[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 89.700 168.730 92.000 ;
    END
  END la_data_in_core[73]
  PIN la_data_in_core[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 89.700 171.030 92.000 ;
    END
  END la_data_in_core[74]
  PIN la_data_in_core[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 89.700 173.330 92.000 ;
    END
  END la_data_in_core[75]
  PIN la_data_in_core[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 89.700 175.170 92.000 ;
    END
  END la_data_in_core[76]
  PIN la_data_in_core[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 89.700 177.470 92.000 ;
    END
  END la_data_in_core[77]
  PIN la_data_in_core[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 89.700 179.770 92.000 ;
    END
  END la_data_in_core[78]
  PIN la_data_in_core[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 89.700 182.070 92.000 ;
    END
  END la_data_in_core[79]
  PIN la_data_in_core[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 89.700 25.210 92.000 ;
    END
  END la_data_in_core[7]
  PIN la_data_in_core[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 89.700 183.910 92.000 ;
    END
  END la_data_in_core[80]
  PIN la_data_in_core[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 89.700 186.210 92.000 ;
    END
  END la_data_in_core[81]
  PIN la_data_in_core[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 89.700 188.510 92.000 ;
    END
  END la_data_in_core[82]
  PIN la_data_in_core[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 89.700 190.810 92.000 ;
    END
  END la_data_in_core[83]
  PIN la_data_in_core[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 89.700 192.650 92.000 ;
    END
  END la_data_in_core[84]
  PIN la_data_in_core[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 89.700 194.950 92.000 ;
    END
  END la_data_in_core[85]
  PIN la_data_in_core[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 89.700 197.250 92.000 ;
    END
  END la_data_in_core[86]
  PIN la_data_in_core[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 89.700 199.550 92.000 ;
    END
  END la_data_in_core[87]
  PIN la_data_in_core[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 89.700 201.390 92.000 ;
    END
  END la_data_in_core[88]
  PIN la_data_in_core[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 89.700 203.690 92.000 ;
    END
  END la_data_in_core[89]
  PIN la_data_in_core[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 89.700 27.050 92.000 ;
    END
  END la_data_in_core[8]
  PIN la_data_in_core[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 89.700 205.990 92.000 ;
    END
  END la_data_in_core[90]
  PIN la_data_in_core[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 89.700 207.830 92.000 ;
    END
  END la_data_in_core[91]
  PIN la_data_in_core[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 89.700 210.130 92.000 ;
    END
  END la_data_in_core[92]
  PIN la_data_in_core[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 89.700 212.430 92.000 ;
    END
  END la_data_in_core[93]
  PIN la_data_in_core[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 89.700 214.730 92.000 ;
    END
  END la_data_in_core[94]
  PIN la_data_in_core[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 89.700 216.570 92.000 ;
    END
  END la_data_in_core[95]
  PIN la_data_in_core[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 89.700 218.870 92.000 ;
    END
  END la_data_in_core[96]
  PIN la_data_in_core[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 89.700 221.170 92.000 ;
    END
  END la_data_in_core[97]
  PIN la_data_in_core[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 89.700 223.470 92.000 ;
    END
  END la_data_in_core[98]
  PIN la_data_in_core[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 89.700 225.310 92.000 ;
    END
  END la_data_in_core[99]
  PIN la_data_in_core[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 89.700 29.350 92.000 ;
    END
  END la_data_in_core[9]
  PIN la_data_in_mprj[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 -2.000 280.050 0.300 ;
    END
  END la_data_in_mprj[0]
  PIN la_data_in_mprj[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 -2.000 497.630 0.300 ;
    END
  END la_data_in_mprj[100]
  PIN la_data_in_mprj[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 -2.000 499.930 0.300 ;
    END
  END la_data_in_mprj[101]
  PIN la_data_in_mprj[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 -2.000 502.230 0.300 ;
    END
  END la_data_in_mprj[102]
  PIN la_data_in_mprj[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 -2.000 504.530 0.300 ;
    END
  END la_data_in_mprj[103]
  PIN la_data_in_mprj[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 -2.000 506.370 0.300 ;
    END
  END la_data_in_mprj[104]
  PIN la_data_in_mprj[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 -2.000 508.670 0.300 ;
    END
  END la_data_in_mprj[105]
  PIN la_data_in_mprj[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 -2.000 510.970 0.300 ;
    END
  END la_data_in_mprj[106]
  PIN la_data_in_mprj[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 -2.000 513.270 0.300 ;
    END
  END la_data_in_mprj[107]
  PIN la_data_in_mprj[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 -2.000 515.110 0.300 ;
    END
  END la_data_in_mprj[108]
  PIN la_data_in_mprj[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 -2.000 517.410 0.300 ;
    END
  END la_data_in_mprj[109]
  PIN la_data_in_mprj[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 -2.000 301.670 0.300 ;
    END
  END la_data_in_mprj[10]
  PIN la_data_in_mprj[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 -2.000 519.710 0.300 ;
    END
  END la_data_in_mprj[110]
  PIN la_data_in_mprj[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 -2.000 521.550 0.300 ;
    END
  END la_data_in_mprj[111]
  PIN la_data_in_mprj[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.570 -2.000 523.850 0.300 ;
    END
  END la_data_in_mprj[112]
  PIN la_data_in_mprj[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.870 -2.000 526.150 0.300 ;
    END
  END la_data_in_mprj[113]
  PIN la_data_in_mprj[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 -2.000 528.450 0.300 ;
    END
  END la_data_in_mprj[114]
  PIN la_data_in_mprj[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 -2.000 530.290 0.300 ;
    END
  END la_data_in_mprj[115]
  PIN la_data_in_mprj[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 -2.000 532.590 0.300 ;
    END
  END la_data_in_mprj[116]
  PIN la_data_in_mprj[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 -2.000 534.890 0.300 ;
    END
  END la_data_in_mprj[117]
  PIN la_data_in_mprj[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 -2.000 537.190 0.300 ;
    END
  END la_data_in_mprj[118]
  PIN la_data_in_mprj[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 -2.000 539.030 0.300 ;
    END
  END la_data_in_mprj[119]
  PIN la_data_in_mprj[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 -2.000 303.970 0.300 ;
    END
  END la_data_in_mprj[11]
  PIN la_data_in_mprj[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 -2.000 541.330 0.300 ;
    END
  END la_data_in_mprj[120]
  PIN la_data_in_mprj[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 -2.000 543.630 0.300 ;
    END
  END la_data_in_mprj[121]
  PIN la_data_in_mprj[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 -2.000 545.930 0.300 ;
    END
  END la_data_in_mprj[122]
  PIN la_data_in_mprj[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 -2.000 547.770 0.300 ;
    END
  END la_data_in_mprj[123]
  PIN la_data_in_mprj[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 -2.000 550.070 0.300 ;
    END
  END la_data_in_mprj[124]
  PIN la_data_in_mprj[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 -2.000 552.370 0.300 ;
    END
  END la_data_in_mprj[125]
  PIN la_data_in_mprj[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 -2.000 554.670 0.300 ;
    END
  END la_data_in_mprj[126]
  PIN la_data_in_mprj[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 -2.000 556.510 0.300 ;
    END
  END la_data_in_mprj[127]
  PIN la_data_in_mprj[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 -2.000 306.270 0.300 ;
    END
  END la_data_in_mprj[12]
  PIN la_data_in_mprj[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 -2.000 308.110 0.300 ;
    END
  END la_data_in_mprj[13]
  PIN la_data_in_mprj[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 -2.000 310.410 0.300 ;
    END
  END la_data_in_mprj[14]
  PIN la_data_in_mprj[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 -2.000 312.710 0.300 ;
    END
  END la_data_in_mprj[15]
  PIN la_data_in_mprj[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 -2.000 315.010 0.300 ;
    END
  END la_data_in_mprj[16]
  PIN la_data_in_mprj[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 -2.000 316.850 0.300 ;
    END
  END la_data_in_mprj[17]
  PIN la_data_in_mprj[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 -2.000 319.150 0.300 ;
    END
  END la_data_in_mprj[18]
  PIN la_data_in_mprj[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 -2.000 321.450 0.300 ;
    END
  END la_data_in_mprj[19]
  PIN la_data_in_mprj[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 -2.000 281.890 0.300 ;
    END
  END la_data_in_mprj[1]
  PIN la_data_in_mprj[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 -2.000 323.290 0.300 ;
    END
  END la_data_in_mprj[20]
  PIN la_data_in_mprj[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 -2.000 325.590 0.300 ;
    END
  END la_data_in_mprj[21]
  PIN la_data_in_mprj[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 -2.000 327.890 0.300 ;
    END
  END la_data_in_mprj[22]
  PIN la_data_in_mprj[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 -2.000 330.190 0.300 ;
    END
  END la_data_in_mprj[23]
  PIN la_data_in_mprj[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 -2.000 332.030 0.300 ;
    END
  END la_data_in_mprj[24]
  PIN la_data_in_mprj[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 -2.000 334.330 0.300 ;
    END
  END la_data_in_mprj[25]
  PIN la_data_in_mprj[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 -2.000 336.630 0.300 ;
    END
  END la_data_in_mprj[26]
  PIN la_data_in_mprj[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 -2.000 338.930 0.300 ;
    END
  END la_data_in_mprj[27]
  PIN la_data_in_mprj[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 -2.000 340.770 0.300 ;
    END
  END la_data_in_mprj[28]
  PIN la_data_in_mprj[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 -2.000 343.070 0.300 ;
    END
  END la_data_in_mprj[29]
  PIN la_data_in_mprj[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 -2.000 284.190 0.300 ;
    END
  END la_data_in_mprj[2]
  PIN la_data_in_mprj[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 -2.000 345.370 0.300 ;
    END
  END la_data_in_mprj[30]
  PIN la_data_in_mprj[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 -2.000 347.670 0.300 ;
    END
  END la_data_in_mprj[31]
  PIN la_data_in_mprj[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 -2.000 349.510 0.300 ;
    END
  END la_data_in_mprj[32]
  PIN la_data_in_mprj[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 -2.000 351.810 0.300 ;
    END
  END la_data_in_mprj[33]
  PIN la_data_in_mprj[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 -2.000 354.110 0.300 ;
    END
  END la_data_in_mprj[34]
  PIN la_data_in_mprj[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 -2.000 356.410 0.300 ;
    END
  END la_data_in_mprj[35]
  PIN la_data_in_mprj[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 -2.000 358.250 0.300 ;
    END
  END la_data_in_mprj[36]
  PIN la_data_in_mprj[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 -2.000 360.550 0.300 ;
    END
  END la_data_in_mprj[37]
  PIN la_data_in_mprj[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 -2.000 362.850 0.300 ;
    END
  END la_data_in_mprj[38]
  PIN la_data_in_mprj[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 -2.000 364.690 0.300 ;
    END
  END la_data_in_mprj[39]
  PIN la_data_in_mprj[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 -2.000 286.490 0.300 ;
    END
  END la_data_in_mprj[3]
  PIN la_data_in_mprj[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 -2.000 366.990 0.300 ;
    END
  END la_data_in_mprj[40]
  PIN la_data_in_mprj[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 -2.000 369.290 0.300 ;
    END
  END la_data_in_mprj[41]
  PIN la_data_in_mprj[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 -2.000 371.590 0.300 ;
    END
  END la_data_in_mprj[42]
  PIN la_data_in_mprj[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 -2.000 373.430 0.300 ;
    END
  END la_data_in_mprj[43]
  PIN la_data_in_mprj[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 -2.000 375.730 0.300 ;
    END
  END la_data_in_mprj[44]
  PIN la_data_in_mprj[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 -2.000 378.030 0.300 ;
    END
  END la_data_in_mprj[45]
  PIN la_data_in_mprj[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 -2.000 380.330 0.300 ;
    END
  END la_data_in_mprj[46]
  PIN la_data_in_mprj[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 -2.000 382.170 0.300 ;
    END
  END la_data_in_mprj[47]
  PIN la_data_in_mprj[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 -2.000 384.470 0.300 ;
    END
  END la_data_in_mprj[48]
  PIN la_data_in_mprj[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 -2.000 386.770 0.300 ;
    END
  END la_data_in_mprj[49]
  PIN la_data_in_mprj[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 -2.000 288.790 0.300 ;
    END
  END la_data_in_mprj[4]
  PIN la_data_in_mprj[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 -2.000 389.070 0.300 ;
    END
  END la_data_in_mprj[50]
  PIN la_data_in_mprj[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 -2.000 390.910 0.300 ;
    END
  END la_data_in_mprj[51]
  PIN la_data_in_mprj[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 -2.000 393.210 0.300 ;
    END
  END la_data_in_mprj[52]
  PIN la_data_in_mprj[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 -2.000 395.510 0.300 ;
    END
  END la_data_in_mprj[53]
  PIN la_data_in_mprj[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 -2.000 397.810 0.300 ;
    END
  END la_data_in_mprj[54]
  PIN la_data_in_mprj[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 -2.000 399.650 0.300 ;
    END
  END la_data_in_mprj[55]
  PIN la_data_in_mprj[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 -2.000 401.950 0.300 ;
    END
  END la_data_in_mprj[56]
  PIN la_data_in_mprj[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 -2.000 404.250 0.300 ;
    END
  END la_data_in_mprj[57]
  PIN la_data_in_mprj[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 -2.000 406.090 0.300 ;
    END
  END la_data_in_mprj[58]
  PIN la_data_in_mprj[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 -2.000 408.390 0.300 ;
    END
  END la_data_in_mprj[59]
  PIN la_data_in_mprj[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 -2.000 290.630 0.300 ;
    END
  END la_data_in_mprj[5]
  PIN la_data_in_mprj[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 -2.000 410.690 0.300 ;
    END
  END la_data_in_mprj[60]
  PIN la_data_in_mprj[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 -2.000 412.990 0.300 ;
    END
  END la_data_in_mprj[61]
  PIN la_data_in_mprj[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 -2.000 414.830 0.300 ;
    END
  END la_data_in_mprj[62]
  PIN la_data_in_mprj[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 -2.000 417.130 0.300 ;
    END
  END la_data_in_mprj[63]
  PIN la_data_in_mprj[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 -2.000 419.430 0.300 ;
    END
  END la_data_in_mprj[64]
  PIN la_data_in_mprj[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 -2.000 421.730 0.300 ;
    END
  END la_data_in_mprj[65]
  PIN la_data_in_mprj[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 -2.000 423.570 0.300 ;
    END
  END la_data_in_mprj[66]
  PIN la_data_in_mprj[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 -2.000 425.870 0.300 ;
    END
  END la_data_in_mprj[67]
  PIN la_data_in_mprj[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 -2.000 428.170 0.300 ;
    END
  END la_data_in_mprj[68]
  PIN la_data_in_mprj[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 -2.000 430.470 0.300 ;
    END
  END la_data_in_mprj[69]
  PIN la_data_in_mprj[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 -2.000 292.930 0.300 ;
    END
  END la_data_in_mprj[6]
  PIN la_data_in_mprj[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 -2.000 432.310 0.300 ;
    END
  END la_data_in_mprj[70]
  PIN la_data_in_mprj[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 -2.000 434.610 0.300 ;
    END
  END la_data_in_mprj[71]
  PIN la_data_in_mprj[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 -2.000 436.910 0.300 ;
    END
  END la_data_in_mprj[72]
  PIN la_data_in_mprj[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 -2.000 439.210 0.300 ;
    END
  END la_data_in_mprj[73]
  PIN la_data_in_mprj[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 -2.000 441.050 0.300 ;
    END
  END la_data_in_mprj[74]
  PIN la_data_in_mprj[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 -2.000 443.350 0.300 ;
    END
  END la_data_in_mprj[75]
  PIN la_data_in_mprj[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 -2.000 445.650 0.300 ;
    END
  END la_data_in_mprj[76]
  PIN la_data_in_mprj[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 -2.000 447.490 0.300 ;
    END
  END la_data_in_mprj[77]
  PIN la_data_in_mprj[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 -2.000 449.790 0.300 ;
    END
  END la_data_in_mprj[78]
  PIN la_data_in_mprj[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 -2.000 452.090 0.300 ;
    END
  END la_data_in_mprj[79]
  PIN la_data_in_mprj[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 -2.000 295.230 0.300 ;
    END
  END la_data_in_mprj[7]
  PIN la_data_in_mprj[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 -2.000 454.390 0.300 ;
    END
  END la_data_in_mprj[80]
  PIN la_data_in_mprj[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 -2.000 456.230 0.300 ;
    END
  END la_data_in_mprj[81]
  PIN la_data_in_mprj[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 -2.000 458.530 0.300 ;
    END
  END la_data_in_mprj[82]
  PIN la_data_in_mprj[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 -2.000 460.830 0.300 ;
    END
  END la_data_in_mprj[83]
  PIN la_data_in_mprj[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 -2.000 463.130 0.300 ;
    END
  END la_data_in_mprj[84]
  PIN la_data_in_mprj[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 -2.000 464.970 0.300 ;
    END
  END la_data_in_mprj[85]
  PIN la_data_in_mprj[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 -2.000 467.270 0.300 ;
    END
  END la_data_in_mprj[86]
  PIN la_data_in_mprj[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 -2.000 469.570 0.300 ;
    END
  END la_data_in_mprj[87]
  PIN la_data_in_mprj[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 -2.000 471.870 0.300 ;
    END
  END la_data_in_mprj[88]
  PIN la_data_in_mprj[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 -2.000 473.710 0.300 ;
    END
  END la_data_in_mprj[89]
  PIN la_data_in_mprj[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 -2.000 297.530 0.300 ;
    END
  END la_data_in_mprj[8]
  PIN la_data_in_mprj[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 -2.000 476.010 0.300 ;
    END
  END la_data_in_mprj[90]
  PIN la_data_in_mprj[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 -2.000 478.310 0.300 ;
    END
  END la_data_in_mprj[91]
  PIN la_data_in_mprj[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 -2.000 480.610 0.300 ;
    END
  END la_data_in_mprj[92]
  PIN la_data_in_mprj[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 -2.000 482.450 0.300 ;
    END
  END la_data_in_mprj[93]
  PIN la_data_in_mprj[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 -2.000 484.750 0.300 ;
    END
  END la_data_in_mprj[94]
  PIN la_data_in_mprj[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 -2.000 487.050 0.300 ;
    END
  END la_data_in_mprj[95]
  PIN la_data_in_mprj[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 -2.000 488.890 0.300 ;
    END
  END la_data_in_mprj[96]
  PIN la_data_in_mprj[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 -2.000 491.190 0.300 ;
    END
  END la_data_in_mprj[97]
  PIN la_data_in_mprj[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 -2.000 493.490 0.300 ;
    END
  END la_data_in_mprj[98]
  PIN la_data_in_mprj[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 -2.000 495.790 0.300 ;
    END
  END la_data_in_mprj[99]
  PIN la_data_in_mprj[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 -2.000 299.370 0.300 ;
    END
  END la_data_in_mprj[9]
  PIN la_data_out_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 89.700 288.790 92.000 ;
    END
  END la_data_out_core[0]
  PIN la_data_out_core[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 89.700 506.370 92.000 ;
    END
  END la_data_out_core[100]
  PIN la_data_out_core[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 89.700 508.670 92.000 ;
    END
  END la_data_out_core[101]
  PIN la_data_out_core[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 89.700 510.970 92.000 ;
    END
  END la_data_out_core[102]
  PIN la_data_out_core[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 89.700 513.270 92.000 ;
    END
  END la_data_out_core[103]
  PIN la_data_out_core[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 89.700 515.110 92.000 ;
    END
  END la_data_out_core[104]
  PIN la_data_out_core[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 89.700 517.410 92.000 ;
    END
  END la_data_out_core[105]
  PIN la_data_out_core[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 89.700 519.710 92.000 ;
    END
  END la_data_out_core[106]
  PIN la_data_out_core[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 89.700 521.550 92.000 ;
    END
  END la_data_out_core[107]
  PIN la_data_out_core[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.570 89.700 523.850 92.000 ;
    END
  END la_data_out_core[108]
  PIN la_data_out_core[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.870 89.700 526.150 92.000 ;
    END
  END la_data_out_core[109]
  PIN la_data_out_core[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 89.700 310.410 92.000 ;
    END
  END la_data_out_core[10]
  PIN la_data_out_core[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 89.700 528.450 92.000 ;
    END
  END la_data_out_core[110]
  PIN la_data_out_core[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 89.700 530.290 92.000 ;
    END
  END la_data_out_core[111]
  PIN la_data_out_core[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 89.700 532.590 92.000 ;
    END
  END la_data_out_core[112]
  PIN la_data_out_core[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 89.700 534.890 92.000 ;
    END
  END la_data_out_core[113]
  PIN la_data_out_core[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 89.700 537.190 92.000 ;
    END
  END la_data_out_core[114]
  PIN la_data_out_core[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 89.700 539.030 92.000 ;
    END
  END la_data_out_core[115]
  PIN la_data_out_core[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 89.700 541.330 92.000 ;
    END
  END la_data_out_core[116]
  PIN la_data_out_core[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 89.700 543.630 92.000 ;
    END
  END la_data_out_core[117]
  PIN la_data_out_core[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 89.700 545.930 92.000 ;
    END
  END la_data_out_core[118]
  PIN la_data_out_core[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 89.700 547.770 92.000 ;
    END
  END la_data_out_core[119]
  PIN la_data_out_core[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 89.700 312.710 92.000 ;
    END
  END la_data_out_core[11]
  PIN la_data_out_core[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 89.700 550.070 92.000 ;
    END
  END la_data_out_core[120]
  PIN la_data_out_core[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 89.700 552.370 92.000 ;
    END
  END la_data_out_core[121]
  PIN la_data_out_core[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 89.700 554.670 92.000 ;
    END
  END la_data_out_core[122]
  PIN la_data_out_core[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 89.700 556.510 92.000 ;
    END
  END la_data_out_core[123]
  PIN la_data_out_core[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 89.700 558.810 92.000 ;
    END
  END la_data_out_core[124]
  PIN la_data_out_core[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 89.700 561.110 92.000 ;
    END
  END la_data_out_core[125]
  PIN la_data_out_core[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 89.700 562.950 92.000 ;
    END
  END la_data_out_core[126]
  PIN la_data_out_core[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 89.700 565.250 92.000 ;
    END
  END la_data_out_core[127]
  PIN la_data_out_core[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 89.700 315.010 92.000 ;
    END
  END la_data_out_core[12]
  PIN la_data_out_core[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 89.700 316.850 92.000 ;
    END
  END la_data_out_core[13]
  PIN la_data_out_core[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 89.700 319.150 92.000 ;
    END
  END la_data_out_core[14]
  PIN la_data_out_core[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 89.700 321.450 92.000 ;
    END
  END la_data_out_core[15]
  PIN la_data_out_core[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 89.700 323.290 92.000 ;
    END
  END la_data_out_core[16]
  PIN la_data_out_core[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 89.700 325.590 92.000 ;
    END
  END la_data_out_core[17]
  PIN la_data_out_core[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 89.700 327.890 92.000 ;
    END
  END la_data_out_core[18]
  PIN la_data_out_core[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 89.700 330.190 92.000 ;
    END
  END la_data_out_core[19]
  PIN la_data_out_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 89.700 290.630 92.000 ;
    END
  END la_data_out_core[1]
  PIN la_data_out_core[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 89.700 332.030 92.000 ;
    END
  END la_data_out_core[20]
  PIN la_data_out_core[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 89.700 334.330 92.000 ;
    END
  END la_data_out_core[21]
  PIN la_data_out_core[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 89.700 336.630 92.000 ;
    END
  END la_data_out_core[22]
  PIN la_data_out_core[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 89.700 338.930 92.000 ;
    END
  END la_data_out_core[23]
  PIN la_data_out_core[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 89.700 340.770 92.000 ;
    END
  END la_data_out_core[24]
  PIN la_data_out_core[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 89.700 343.070 92.000 ;
    END
  END la_data_out_core[25]
  PIN la_data_out_core[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 89.700 345.370 92.000 ;
    END
  END la_data_out_core[26]
  PIN la_data_out_core[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 89.700 347.670 92.000 ;
    END
  END la_data_out_core[27]
  PIN la_data_out_core[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 89.700 349.510 92.000 ;
    END
  END la_data_out_core[28]
  PIN la_data_out_core[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 89.700 351.810 92.000 ;
    END
  END la_data_out_core[29]
  PIN la_data_out_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 89.700 292.930 92.000 ;
    END
  END la_data_out_core[2]
  PIN la_data_out_core[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 89.700 354.110 92.000 ;
    END
  END la_data_out_core[30]
  PIN la_data_out_core[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 89.700 356.410 92.000 ;
    END
  END la_data_out_core[31]
  PIN la_data_out_core[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 89.700 358.250 92.000 ;
    END
  END la_data_out_core[32]
  PIN la_data_out_core[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 89.700 360.550 92.000 ;
    END
  END la_data_out_core[33]
  PIN la_data_out_core[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 89.700 362.850 92.000 ;
    END
  END la_data_out_core[34]
  PIN la_data_out_core[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 89.700 364.690 92.000 ;
    END
  END la_data_out_core[35]
  PIN la_data_out_core[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 89.700 366.990 92.000 ;
    END
  END la_data_out_core[36]
  PIN la_data_out_core[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 89.700 369.290 92.000 ;
    END
  END la_data_out_core[37]
  PIN la_data_out_core[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 89.700 371.590 92.000 ;
    END
  END la_data_out_core[38]
  PIN la_data_out_core[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 89.700 373.430 92.000 ;
    END
  END la_data_out_core[39]
  PIN la_data_out_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 89.700 295.230 92.000 ;
    END
  END la_data_out_core[3]
  PIN la_data_out_core[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 89.700 375.730 92.000 ;
    END
  END la_data_out_core[40]
  PIN la_data_out_core[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 89.700 378.030 92.000 ;
    END
  END la_data_out_core[41]
  PIN la_data_out_core[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 89.700 380.330 92.000 ;
    END
  END la_data_out_core[42]
  PIN la_data_out_core[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 89.700 382.170 92.000 ;
    END
  END la_data_out_core[43]
  PIN la_data_out_core[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 89.700 384.470 92.000 ;
    END
  END la_data_out_core[44]
  PIN la_data_out_core[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 89.700 386.770 92.000 ;
    END
  END la_data_out_core[45]
  PIN la_data_out_core[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 89.700 389.070 92.000 ;
    END
  END la_data_out_core[46]
  PIN la_data_out_core[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 89.700 390.910 92.000 ;
    END
  END la_data_out_core[47]
  PIN la_data_out_core[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 89.700 393.210 92.000 ;
    END
  END la_data_out_core[48]
  PIN la_data_out_core[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 89.700 395.510 92.000 ;
    END
  END la_data_out_core[49]
  PIN la_data_out_core[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 89.700 297.530 92.000 ;
    END
  END la_data_out_core[4]
  PIN la_data_out_core[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 89.700 397.810 92.000 ;
    END
  END la_data_out_core[50]
  PIN la_data_out_core[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 89.700 399.650 92.000 ;
    END
  END la_data_out_core[51]
  PIN la_data_out_core[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 89.700 401.950 92.000 ;
    END
  END la_data_out_core[52]
  PIN la_data_out_core[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 89.700 404.250 92.000 ;
    END
  END la_data_out_core[53]
  PIN la_data_out_core[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 89.700 406.090 92.000 ;
    END
  END la_data_out_core[54]
  PIN la_data_out_core[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 89.700 408.390 92.000 ;
    END
  END la_data_out_core[55]
  PIN la_data_out_core[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 89.700 410.690 92.000 ;
    END
  END la_data_out_core[56]
  PIN la_data_out_core[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 89.700 412.990 92.000 ;
    END
  END la_data_out_core[57]
  PIN la_data_out_core[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 89.700 414.830 92.000 ;
    END
  END la_data_out_core[58]
  PIN la_data_out_core[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 89.700 417.130 92.000 ;
    END
  END la_data_out_core[59]
  PIN la_data_out_core[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 89.700 299.370 92.000 ;
    END
  END la_data_out_core[5]
  PIN la_data_out_core[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 89.700 419.430 92.000 ;
    END
  END la_data_out_core[60]
  PIN la_data_out_core[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 89.700 421.730 92.000 ;
    END
  END la_data_out_core[61]
  PIN la_data_out_core[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 89.700 423.570 92.000 ;
    END
  END la_data_out_core[62]
  PIN la_data_out_core[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 89.700 425.870 92.000 ;
    END
  END la_data_out_core[63]
  PIN la_data_out_core[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 89.700 428.170 92.000 ;
    END
  END la_data_out_core[64]
  PIN la_data_out_core[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 89.700 430.470 92.000 ;
    END
  END la_data_out_core[65]
  PIN la_data_out_core[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 89.700 432.310 92.000 ;
    END
  END la_data_out_core[66]
  PIN la_data_out_core[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 89.700 434.610 92.000 ;
    END
  END la_data_out_core[67]
  PIN la_data_out_core[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 89.700 436.910 92.000 ;
    END
  END la_data_out_core[68]
  PIN la_data_out_core[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 89.700 439.210 92.000 ;
    END
  END la_data_out_core[69]
  PIN la_data_out_core[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 89.700 301.670 92.000 ;
    END
  END la_data_out_core[6]
  PIN la_data_out_core[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 89.700 441.050 92.000 ;
    END
  END la_data_out_core[70]
  PIN la_data_out_core[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 89.700 443.350 92.000 ;
    END
  END la_data_out_core[71]
  PIN la_data_out_core[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 89.700 445.650 92.000 ;
    END
  END la_data_out_core[72]
  PIN la_data_out_core[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 89.700 447.490 92.000 ;
    END
  END la_data_out_core[73]
  PIN la_data_out_core[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 89.700 449.790 92.000 ;
    END
  END la_data_out_core[74]
  PIN la_data_out_core[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 89.700 452.090 92.000 ;
    END
  END la_data_out_core[75]
  PIN la_data_out_core[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 89.700 454.390 92.000 ;
    END
  END la_data_out_core[76]
  PIN la_data_out_core[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 89.700 456.230 92.000 ;
    END
  END la_data_out_core[77]
  PIN la_data_out_core[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 89.700 458.530 92.000 ;
    END
  END la_data_out_core[78]
  PIN la_data_out_core[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 89.700 460.830 92.000 ;
    END
  END la_data_out_core[79]
  PIN la_data_out_core[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 89.700 303.970 92.000 ;
    END
  END la_data_out_core[7]
  PIN la_data_out_core[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 89.700 463.130 92.000 ;
    END
  END la_data_out_core[80]
  PIN la_data_out_core[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 89.700 464.970 92.000 ;
    END
  END la_data_out_core[81]
  PIN la_data_out_core[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 89.700 467.270 92.000 ;
    END
  END la_data_out_core[82]
  PIN la_data_out_core[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 89.700 469.570 92.000 ;
    END
  END la_data_out_core[83]
  PIN la_data_out_core[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 89.700 471.870 92.000 ;
    END
  END la_data_out_core[84]
  PIN la_data_out_core[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 89.700 473.710 92.000 ;
    END
  END la_data_out_core[85]
  PIN la_data_out_core[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 89.700 476.010 92.000 ;
    END
  END la_data_out_core[86]
  PIN la_data_out_core[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 89.700 478.310 92.000 ;
    END
  END la_data_out_core[87]
  PIN la_data_out_core[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 89.700 480.610 92.000 ;
    END
  END la_data_out_core[88]
  PIN la_data_out_core[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 89.700 482.450 92.000 ;
    END
  END la_data_out_core[89]
  PIN la_data_out_core[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 89.700 306.270 92.000 ;
    END
  END la_data_out_core[8]
  PIN la_data_out_core[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 89.700 484.750 92.000 ;
    END
  END la_data_out_core[90]
  PIN la_data_out_core[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 89.700 487.050 92.000 ;
    END
  END la_data_out_core[91]
  PIN la_data_out_core[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 89.700 488.890 92.000 ;
    END
  END la_data_out_core[92]
  PIN la_data_out_core[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 89.700 491.190 92.000 ;
    END
  END la_data_out_core[93]
  PIN la_data_out_core[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 89.700 493.490 92.000 ;
    END
  END la_data_out_core[94]
  PIN la_data_out_core[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 89.700 495.790 92.000 ;
    END
  END la_data_out_core[95]
  PIN la_data_out_core[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 89.700 497.630 92.000 ;
    END
  END la_data_out_core[96]
  PIN la_data_out_core[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 89.700 499.930 92.000 ;
    END
  END la_data_out_core[97]
  PIN la_data_out_core[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 89.700 502.230 92.000 ;
    END
  END la_data_out_core[98]
  PIN la_data_out_core[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 89.700 504.530 92.000 ;
    END
  END la_data_out_core[99]
  PIN la_data_out_core[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 89.700 308.110 92.000 ;
    END
  END la_data_out_core[9]
  PIN la_data_out_mprj[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 -2.000 1.290 0.300 ;
    END
  END la_data_out_mprj[0]
  PIN la_data_out_mprj[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 -2.000 218.870 0.300 ;
    END
  END la_data_out_mprj[100]
  PIN la_data_out_mprj[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 -2.000 221.170 0.300 ;
    END
  END la_data_out_mprj[101]
  PIN la_data_out_mprj[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 -2.000 223.470 0.300 ;
    END
  END la_data_out_mprj[102]
  PIN la_data_out_mprj[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 -2.000 225.310 0.300 ;
    END
  END la_data_out_mprj[103]
  PIN la_data_out_mprj[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 -2.000 227.610 0.300 ;
    END
  END la_data_out_mprj[104]
  PIN la_data_out_mprj[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 -2.000 229.910 0.300 ;
    END
  END la_data_out_mprj[105]
  PIN la_data_out_mprj[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 -2.000 232.210 0.300 ;
    END
  END la_data_out_mprj[106]
  PIN la_data_out_mprj[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 -2.000 234.050 0.300 ;
    END
  END la_data_out_mprj[107]
  PIN la_data_out_mprj[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 -2.000 236.350 0.300 ;
    END
  END la_data_out_mprj[108]
  PIN la_data_out_mprj[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 -2.000 238.650 0.300 ;
    END
  END la_data_out_mprj[109]
  PIN la_data_out_mprj[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 -2.000 22.910 0.300 ;
    END
  END la_data_out_mprj[10]
  PIN la_data_out_mprj[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 -2.000 240.950 0.300 ;
    END
  END la_data_out_mprj[110]
  PIN la_data_out_mprj[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 -2.000 242.790 0.300 ;
    END
  END la_data_out_mprj[111]
  PIN la_data_out_mprj[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 -2.000 245.090 0.300 ;
    END
  END la_data_out_mprj[112]
  PIN la_data_out_mprj[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 -2.000 247.390 0.300 ;
    END
  END la_data_out_mprj[113]
  PIN la_data_out_mprj[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 -2.000 249.230 0.300 ;
    END
  END la_data_out_mprj[114]
  PIN la_data_out_mprj[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 -2.000 251.530 0.300 ;
    END
  END la_data_out_mprj[115]
  PIN la_data_out_mprj[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 -2.000 253.830 0.300 ;
    END
  END la_data_out_mprj[116]
  PIN la_data_out_mprj[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 -2.000 256.130 0.300 ;
    END
  END la_data_out_mprj[117]
  PIN la_data_out_mprj[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 -2.000 257.970 0.300 ;
    END
  END la_data_out_mprj[118]
  PIN la_data_out_mprj[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 -2.000 260.270 0.300 ;
    END
  END la_data_out_mprj[119]
  PIN la_data_out_mprj[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 -2.000 25.210 0.300 ;
    END
  END la_data_out_mprj[11]
  PIN la_data_out_mprj[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 -2.000 262.570 0.300 ;
    END
  END la_data_out_mprj[120]
  PIN la_data_out_mprj[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 -2.000 264.870 0.300 ;
    END
  END la_data_out_mprj[121]
  PIN la_data_out_mprj[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 -2.000 266.710 0.300 ;
    END
  END la_data_out_mprj[122]
  PIN la_data_out_mprj[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 -2.000 269.010 0.300 ;
    END
  END la_data_out_mprj[123]
  PIN la_data_out_mprj[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 -2.000 271.310 0.300 ;
    END
  END la_data_out_mprj[124]
  PIN la_data_out_mprj[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 -2.000 273.610 0.300 ;
    END
  END la_data_out_mprj[125]
  PIN la_data_out_mprj[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 -2.000 275.450 0.300 ;
    END
  END la_data_out_mprj[126]
  PIN la_data_out_mprj[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 -2.000 277.750 0.300 ;
    END
  END la_data_out_mprj[127]
  PIN la_data_out_mprj[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 -2.000 27.050 0.300 ;
    END
  END la_data_out_mprj[12]
  PIN la_data_out_mprj[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 -2.000 29.350 0.300 ;
    END
  END la_data_out_mprj[13]
  PIN la_data_out_mprj[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 -2.000 31.650 0.300 ;
    END
  END la_data_out_mprj[14]
  PIN la_data_out_mprj[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 -2.000 33.950 0.300 ;
    END
  END la_data_out_mprj[15]
  PIN la_data_out_mprj[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 -2.000 35.790 0.300 ;
    END
  END la_data_out_mprj[16]
  PIN la_data_out_mprj[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 -2.000 38.090 0.300 ;
    END
  END la_data_out_mprj[17]
  PIN la_data_out_mprj[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 -2.000 40.390 0.300 ;
    END
  END la_data_out_mprj[18]
  PIN la_data_out_mprj[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 -2.000 42.230 0.300 ;
    END
  END la_data_out_mprj[19]
  PIN la_data_out_mprj[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 -2.000 3.130 0.300 ;
    END
  END la_data_out_mprj[1]
  PIN la_data_out_mprj[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 -2.000 44.530 0.300 ;
    END
  END la_data_out_mprj[20]
  PIN la_data_out_mprj[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 -2.000 46.830 0.300 ;
    END
  END la_data_out_mprj[21]
  PIN la_data_out_mprj[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 -2.000 49.130 0.300 ;
    END
  END la_data_out_mprj[22]
  PIN la_data_out_mprj[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 -2.000 50.970 0.300 ;
    END
  END la_data_out_mprj[23]
  PIN la_data_out_mprj[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 -2.000 53.270 0.300 ;
    END
  END la_data_out_mprj[24]
  PIN la_data_out_mprj[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 -2.000 55.570 0.300 ;
    END
  END la_data_out_mprj[25]
  PIN la_data_out_mprj[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 -2.000 57.870 0.300 ;
    END
  END la_data_out_mprj[26]
  PIN la_data_out_mprj[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 -2.000 59.710 0.300 ;
    END
  END la_data_out_mprj[27]
  PIN la_data_out_mprj[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 -2.000 62.010 0.300 ;
    END
  END la_data_out_mprj[28]
  PIN la_data_out_mprj[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 -2.000 64.310 0.300 ;
    END
  END la_data_out_mprj[29]
  PIN la_data_out_mprj[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 -2.000 5.430 0.300 ;
    END
  END la_data_out_mprj[2]
  PIN la_data_out_mprj[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 -2.000 66.610 0.300 ;
    END
  END la_data_out_mprj[30]
  PIN la_data_out_mprj[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 -2.000 68.450 0.300 ;
    END
  END la_data_out_mprj[31]
  PIN la_data_out_mprj[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 -2.000 70.750 0.300 ;
    END
  END la_data_out_mprj[32]
  PIN la_data_out_mprj[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 -2.000 73.050 0.300 ;
    END
  END la_data_out_mprj[33]
  PIN la_data_out_mprj[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 -2.000 75.350 0.300 ;
    END
  END la_data_out_mprj[34]
  PIN la_data_out_mprj[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 -2.000 77.190 0.300 ;
    END
  END la_data_out_mprj[35]
  PIN la_data_out_mprj[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 -2.000 79.490 0.300 ;
    END
  END la_data_out_mprj[36]
  PIN la_data_out_mprj[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 -2.000 81.790 0.300 ;
    END
  END la_data_out_mprj[37]
  PIN la_data_out_mprj[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 -2.000 83.630 0.300 ;
    END
  END la_data_out_mprj[38]
  PIN la_data_out_mprj[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 -2.000 85.930 0.300 ;
    END
  END la_data_out_mprj[39]
  PIN la_data_out_mprj[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 -2.000 7.730 0.300 ;
    END
  END la_data_out_mprj[3]
  PIN la_data_out_mprj[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 -2.000 88.230 0.300 ;
    END
  END la_data_out_mprj[40]
  PIN la_data_out_mprj[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 -2.000 90.530 0.300 ;
    END
  END la_data_out_mprj[41]
  PIN la_data_out_mprj[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 -2.000 92.370 0.300 ;
    END
  END la_data_out_mprj[42]
  PIN la_data_out_mprj[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 -2.000 94.670 0.300 ;
    END
  END la_data_out_mprj[43]
  PIN la_data_out_mprj[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 -2.000 96.970 0.300 ;
    END
  END la_data_out_mprj[44]
  PIN la_data_out_mprj[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 -2.000 99.270 0.300 ;
    END
  END la_data_out_mprj[45]
  PIN la_data_out_mprj[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 -2.000 101.110 0.300 ;
    END
  END la_data_out_mprj[46]
  PIN la_data_out_mprj[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 -2.000 103.410 0.300 ;
    END
  END la_data_out_mprj[47]
  PIN la_data_out_mprj[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 -2.000 105.710 0.300 ;
    END
  END la_data_out_mprj[48]
  PIN la_data_out_mprj[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 -2.000 108.010 0.300 ;
    END
  END la_data_out_mprj[49]
  PIN la_data_out_mprj[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 -2.000 9.570 0.300 ;
    END
  END la_data_out_mprj[4]
  PIN la_data_out_mprj[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 -2.000 109.850 0.300 ;
    END
  END la_data_out_mprj[50]
  PIN la_data_out_mprj[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 -2.000 112.150 0.300 ;
    END
  END la_data_out_mprj[51]
  PIN la_data_out_mprj[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 -2.000 114.450 0.300 ;
    END
  END la_data_out_mprj[52]
  PIN la_data_out_mprj[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 -2.000 116.750 0.300 ;
    END
  END la_data_out_mprj[53]
  PIN la_data_out_mprj[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 -2.000 118.590 0.300 ;
    END
  END la_data_out_mprj[54]
  PIN la_data_out_mprj[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 -2.000 120.890 0.300 ;
    END
  END la_data_out_mprj[55]
  PIN la_data_out_mprj[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 -2.000 123.190 0.300 ;
    END
  END la_data_out_mprj[56]
  PIN la_data_out_mprj[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 -2.000 125.030 0.300 ;
    END
  END la_data_out_mprj[57]
  PIN la_data_out_mprj[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 -2.000 127.330 0.300 ;
    END
  END la_data_out_mprj[58]
  PIN la_data_out_mprj[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 -2.000 129.630 0.300 ;
    END
  END la_data_out_mprj[59]
  PIN la_data_out_mprj[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 -2.000 11.870 0.300 ;
    END
  END la_data_out_mprj[5]
  PIN la_data_out_mprj[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 -2.000 131.930 0.300 ;
    END
  END la_data_out_mprj[60]
  PIN la_data_out_mprj[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 -2.000 133.770 0.300 ;
    END
  END la_data_out_mprj[61]
  PIN la_data_out_mprj[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 -2.000 136.070 0.300 ;
    END
  END la_data_out_mprj[62]
  PIN la_data_out_mprj[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 -2.000 138.370 0.300 ;
    END
  END la_data_out_mprj[63]
  PIN la_data_out_mprj[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 -2.000 140.670 0.300 ;
    END
  END la_data_out_mprj[64]
  PIN la_data_out_mprj[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 -2.000 142.510 0.300 ;
    END
  END la_data_out_mprj[65]
  PIN la_data_out_mprj[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 -2.000 144.810 0.300 ;
    END
  END la_data_out_mprj[66]
  PIN la_data_out_mprj[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 -2.000 147.110 0.300 ;
    END
  END la_data_out_mprj[67]
  PIN la_data_out_mprj[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 -2.000 149.410 0.300 ;
    END
  END la_data_out_mprj[68]
  PIN la_data_out_mprj[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 -2.000 151.250 0.300 ;
    END
  END la_data_out_mprj[69]
  PIN la_data_out_mprj[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 -2.000 14.170 0.300 ;
    END
  END la_data_out_mprj[6]
  PIN la_data_out_mprj[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 -2.000 153.550 0.300 ;
    END
  END la_data_out_mprj[70]
  PIN la_data_out_mprj[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 -2.000 155.850 0.300 ;
    END
  END la_data_out_mprj[71]
  PIN la_data_out_mprj[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 -2.000 158.150 0.300 ;
    END
  END la_data_out_mprj[72]
  PIN la_data_out_mprj[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 -2.000 159.990 0.300 ;
    END
  END la_data_out_mprj[73]
  PIN la_data_out_mprj[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 -2.000 162.290 0.300 ;
    END
  END la_data_out_mprj[74]
  PIN la_data_out_mprj[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 -2.000 164.590 0.300 ;
    END
  END la_data_out_mprj[75]
  PIN la_data_out_mprj[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 -2.000 166.430 0.300 ;
    END
  END la_data_out_mprj[76]
  PIN la_data_out_mprj[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 -2.000 168.730 0.300 ;
    END
  END la_data_out_mprj[77]
  PIN la_data_out_mprj[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 -2.000 171.030 0.300 ;
    END
  END la_data_out_mprj[78]
  PIN la_data_out_mprj[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 -2.000 173.330 0.300 ;
    END
  END la_data_out_mprj[79]
  PIN la_data_out_mprj[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 -2.000 16.470 0.300 ;
    END
  END la_data_out_mprj[7]
  PIN la_data_out_mprj[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 -2.000 175.170 0.300 ;
    END
  END la_data_out_mprj[80]
  PIN la_data_out_mprj[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 -2.000 177.470 0.300 ;
    END
  END la_data_out_mprj[81]
  PIN la_data_out_mprj[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 -2.000 179.770 0.300 ;
    END
  END la_data_out_mprj[82]
  PIN la_data_out_mprj[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 -2.000 182.070 0.300 ;
    END
  END la_data_out_mprj[83]
  PIN la_data_out_mprj[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 -2.000 183.910 0.300 ;
    END
  END la_data_out_mprj[84]
  PIN la_data_out_mprj[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 -2.000 186.210 0.300 ;
    END
  END la_data_out_mprj[85]
  PIN la_data_out_mprj[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 -2.000 188.510 0.300 ;
    END
  END la_data_out_mprj[86]
  PIN la_data_out_mprj[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 -2.000 190.810 0.300 ;
    END
  END la_data_out_mprj[87]
  PIN la_data_out_mprj[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 -2.000 192.650 0.300 ;
    END
  END la_data_out_mprj[88]
  PIN la_data_out_mprj[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 -2.000 194.950 0.300 ;
    END
  END la_data_out_mprj[89]
  PIN la_data_out_mprj[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 -2.000 18.310 0.300 ;
    END
  END la_data_out_mprj[8]
  PIN la_data_out_mprj[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 -2.000 197.250 0.300 ;
    END
  END la_data_out_mprj[90]
  PIN la_data_out_mprj[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 -2.000 199.550 0.300 ;
    END
  END la_data_out_mprj[91]
  PIN la_data_out_mprj[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 -2.000 201.390 0.300 ;
    END
  END la_data_out_mprj[92]
  PIN la_data_out_mprj[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 -2.000 203.690 0.300 ;
    END
  END la_data_out_mprj[93]
  PIN la_data_out_mprj[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 -2.000 205.990 0.300 ;
    END
  END la_data_out_mprj[94]
  PIN la_data_out_mprj[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 -2.000 207.830 0.300 ;
    END
  END la_data_out_mprj[95]
  PIN la_data_out_mprj[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 -2.000 210.130 0.300 ;
    END
  END la_data_out_mprj[96]
  PIN la_data_out_mprj[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 -2.000 212.430 0.300 ;
    END
  END la_data_out_mprj[97]
  PIN la_data_out_mprj[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 -2.000 214.730 0.300 ;
    END
  END la_data_out_mprj[98]
  PIN la_data_out_mprj[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 -2.000 216.570 0.300 ;
    END
  END la_data_out_mprj[99]
  PIN la_data_out_mprj[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 -2.000 20.610 0.300 ;
    END
  END la_data_out_mprj[9]
  PIN la_oen_core[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 89.700 567.550 92.000 ;
    END
  END la_oen_core[0]
  PIN la_oen_core[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 89.700 785.590 92.000 ;
    END
  END la_oen_core[100]
  PIN la_oen_core[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 89.700 787.430 92.000 ;
    END
  END la_oen_core[101]
  PIN la_oen_core[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 89.700 789.730 92.000 ;
    END
  END la_oen_core[102]
  PIN la_oen_core[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.750 89.700 792.030 92.000 ;
    END
  END la_oen_core[103]
  PIN la_oen_core[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 89.700 794.330 92.000 ;
    END
  END la_oen_core[104]
  PIN la_oen_core[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 89.700 796.170 92.000 ;
    END
  END la_oen_core[105]
  PIN la_oen_core[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 89.700 798.470 92.000 ;
    END
  END la_oen_core[106]
  PIN la_oen_core[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.490 89.700 800.770 92.000 ;
    END
  END la_oen_core[107]
  PIN la_oen_core[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.330 89.700 802.610 92.000 ;
    END
  END la_oen_core[108]
  PIN la_oen_core[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.630 89.700 804.910 92.000 ;
    END
  END la_oen_core[109]
  PIN la_oen_core[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 89.700 589.170 92.000 ;
    END
  END la_oen_core[10]
  PIN la_oen_core[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.930 89.700 807.210 92.000 ;
    END
  END la_oen_core[110]
  PIN la_oen_core[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.230 89.700 809.510 92.000 ;
    END
  END la_oen_core[111]
  PIN la_oen_core[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.070 89.700 811.350 92.000 ;
    END
  END la_oen_core[112]
  PIN la_oen_core[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.370 89.700 813.650 92.000 ;
    END
  END la_oen_core[113]
  PIN la_oen_core[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.670 89.700 815.950 92.000 ;
    END
  END la_oen_core[114]
  PIN la_oen_core[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 89.700 818.250 92.000 ;
    END
  END la_oen_core[115]
  PIN la_oen_core[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 89.700 820.090 92.000 ;
    END
  END la_oen_core[116]
  PIN la_oen_core[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.110 89.700 822.390 92.000 ;
    END
  END la_oen_core[117]
  PIN la_oen_core[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 89.700 824.690 92.000 ;
    END
  END la_oen_core[118]
  PIN la_oen_core[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.710 89.700 826.990 92.000 ;
    END
  END la_oen_core[119]
  PIN la_oen_core[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 89.700 591.470 92.000 ;
    END
  END la_oen_core[11]
  PIN la_oen_core[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.550 89.700 828.830 92.000 ;
    END
  END la_oen_core[120]
  PIN la_oen_core[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 89.700 831.130 92.000 ;
    END
  END la_oen_core[121]
  PIN la_oen_core[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 89.700 833.430 92.000 ;
    END
  END la_oen_core[122]
  PIN la_oen_core[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.450 89.700 835.730 92.000 ;
    END
  END la_oen_core[123]
  PIN la_oen_core[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 89.700 837.570 92.000 ;
    END
  END la_oen_core[124]
  PIN la_oen_core[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.590 89.700 839.870 92.000 ;
    END
  END la_oen_core[125]
  PIN la_oen_core[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.890 89.700 842.170 92.000 ;
    END
  END la_oen_core[126]
  PIN la_oen_core[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 89.700 844.010 92.000 ;
    END
  END la_oen_core[127]
  PIN la_oen_core[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 89.700 593.770 92.000 ;
    END
  END la_oen_core[12]
  PIN la_oen_core[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 89.700 596.070 92.000 ;
    END
  END la_oen_core[13]
  PIN la_oen_core[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 89.700 597.910 92.000 ;
    END
  END la_oen_core[14]
  PIN la_oen_core[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 89.700 600.210 92.000 ;
    END
  END la_oen_core[15]
  PIN la_oen_core[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 89.700 602.510 92.000 ;
    END
  END la_oen_core[16]
  PIN la_oen_core[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 89.700 604.350 92.000 ;
    END
  END la_oen_core[17]
  PIN la_oen_core[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 89.700 606.650 92.000 ;
    END
  END la_oen_core[18]
  PIN la_oen_core[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 89.700 608.950 92.000 ;
    END
  END la_oen_core[19]
  PIN la_oen_core[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 89.700 569.850 92.000 ;
    END
  END la_oen_core[1]
  PIN la_oen_core[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 89.700 611.250 92.000 ;
    END
  END la_oen_core[20]
  PIN la_oen_core[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 89.700 613.090 92.000 ;
    END
  END la_oen_core[21]
  PIN la_oen_core[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 89.700 615.390 92.000 ;
    END
  END la_oen_core[22]
  PIN la_oen_core[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 89.700 617.690 92.000 ;
    END
  END la_oen_core[23]
  PIN la_oen_core[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 89.700 619.990 92.000 ;
    END
  END la_oen_core[24]
  PIN la_oen_core[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 89.700 621.830 92.000 ;
    END
  END la_oen_core[25]
  PIN la_oen_core[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 89.700 624.130 92.000 ;
    END
  END la_oen_core[26]
  PIN la_oen_core[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.150 89.700 626.430 92.000 ;
    END
  END la_oen_core[27]
  PIN la_oen_core[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 89.700 628.730 92.000 ;
    END
  END la_oen_core[28]
  PIN la_oen_core[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 89.700 630.570 92.000 ;
    END
  END la_oen_core[29]
  PIN la_oen_core[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 89.700 571.690 92.000 ;
    END
  END la_oen_core[2]
  PIN la_oen_core[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.590 89.700 632.870 92.000 ;
    END
  END la_oen_core[30]
  PIN la_oen_core[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 89.700 635.170 92.000 ;
    END
  END la_oen_core[31]
  PIN la_oen_core[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 89.700 637.470 92.000 ;
    END
  END la_oen_core[32]
  PIN la_oen_core[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 89.700 639.310 92.000 ;
    END
  END la_oen_core[33]
  PIN la_oen_core[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 89.700 641.610 92.000 ;
    END
  END la_oen_core[34]
  PIN la_oen_core[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.630 89.700 643.910 92.000 ;
    END
  END la_oen_core[35]
  PIN la_oen_core[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.470 89.700 645.750 92.000 ;
    END
  END la_oen_core[36]
  PIN la_oen_core[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.770 89.700 648.050 92.000 ;
    END
  END la_oen_core[37]
  PIN la_oen_core[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 89.700 650.350 92.000 ;
    END
  END la_oen_core[38]
  PIN la_oen_core[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 89.700 652.650 92.000 ;
    END
  END la_oen_core[39]
  PIN la_oen_core[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.710 89.700 573.990 92.000 ;
    END
  END la_oen_core[3]
  PIN la_oen_core[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 89.700 654.490 92.000 ;
    END
  END la_oen_core[40]
  PIN la_oen_core[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 89.700 656.790 92.000 ;
    END
  END la_oen_core[41]
  PIN la_oen_core[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.810 89.700 659.090 92.000 ;
    END
  END la_oen_core[42]
  PIN la_oen_core[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 89.700 661.390 92.000 ;
    END
  END la_oen_core[43]
  PIN la_oen_core[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.950 89.700 663.230 92.000 ;
    END
  END la_oen_core[44]
  PIN la_oen_core[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.250 89.700 665.530 92.000 ;
    END
  END la_oen_core[45]
  PIN la_oen_core[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 89.700 667.830 92.000 ;
    END
  END la_oen_core[46]
  PIN la_oen_core[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 89.700 670.130 92.000 ;
    END
  END la_oen_core[47]
  PIN la_oen_core[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.690 89.700 671.970 92.000 ;
    END
  END la_oen_core[48]
  PIN la_oen_core[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 89.700 674.270 92.000 ;
    END
  END la_oen_core[49]
  PIN la_oen_core[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 89.700 576.290 92.000 ;
    END
  END la_oen_core[4]
  PIN la_oen_core[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 89.700 676.570 92.000 ;
    END
  END la_oen_core[50]
  PIN la_oen_core[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.590 89.700 678.870 92.000 ;
    END
  END la_oen_core[51]
  PIN la_oen_core[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 89.700 680.710 92.000 ;
    END
  END la_oen_core[52]
  PIN la_oen_core[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 89.700 683.010 92.000 ;
    END
  END la_oen_core[53]
  PIN la_oen_core[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 89.700 685.310 92.000 ;
    END
  END la_oen_core[54]
  PIN la_oen_core[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.870 89.700 687.150 92.000 ;
    END
  END la_oen_core[55]
  PIN la_oen_core[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 89.700 689.450 92.000 ;
    END
  END la_oen_core[56]
  PIN la_oen_core[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.470 89.700 691.750 92.000 ;
    END
  END la_oen_core[57]
  PIN la_oen_core[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 89.700 694.050 92.000 ;
    END
  END la_oen_core[58]
  PIN la_oen_core[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 89.700 695.890 92.000 ;
    END
  END la_oen_core[59]
  PIN la_oen_core[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 89.700 578.590 92.000 ;
    END
  END la_oen_core[5]
  PIN la_oen_core[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.910 89.700 698.190 92.000 ;
    END
  END la_oen_core[60]
  PIN la_oen_core[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 89.700 700.490 92.000 ;
    END
  END la_oen_core[61]
  PIN la_oen_core[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 89.700 702.790 92.000 ;
    END
  END la_oen_core[62]
  PIN la_oen_core[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.350 89.700 704.630 92.000 ;
    END
  END la_oen_core[63]
  PIN la_oen_core[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.650 89.700 706.930 92.000 ;
    END
  END la_oen_core[64]
  PIN la_oen_core[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.950 89.700 709.230 92.000 ;
    END
  END la_oen_core[65]
  PIN la_oen_core[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 89.700 711.530 92.000 ;
    END
  END la_oen_core[66]
  PIN la_oen_core[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 89.700 713.370 92.000 ;
    END
  END la_oen_core[67]
  PIN la_oen_core[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 89.700 715.670 92.000 ;
    END
  END la_oen_core[68]
  PIN la_oen_core[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 89.700 717.970 92.000 ;
    END
  END la_oen_core[69]
  PIN la_oen_core[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 89.700 580.430 92.000 ;
    END
  END la_oen_core[6]
  PIN la_oen_core[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.990 89.700 720.270 92.000 ;
    END
  END la_oen_core[70]
  PIN la_oen_core[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.830 89.700 722.110 92.000 ;
    END
  END la_oen_core[71]
  PIN la_oen_core[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 89.700 724.410 92.000 ;
    END
  END la_oen_core[72]
  PIN la_oen_core[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.430 89.700 726.710 92.000 ;
    END
  END la_oen_core[73]
  PIN la_oen_core[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.270 89.700 728.550 92.000 ;
    END
  END la_oen_core[74]
  PIN la_oen_core[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.570 89.700 730.850 92.000 ;
    END
  END la_oen_core[75]
  PIN la_oen_core[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 89.700 733.150 92.000 ;
    END
  END la_oen_core[76]
  PIN la_oen_core[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 89.700 735.450 92.000 ;
    END
  END la_oen_core[77]
  PIN la_oen_core[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 89.700 737.290 92.000 ;
    END
  END la_oen_core[78]
  PIN la_oen_core[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.310 89.700 739.590 92.000 ;
    END
  END la_oen_core[79]
  PIN la_oen_core[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 89.700 582.730 92.000 ;
    END
  END la_oen_core[7]
  PIN la_oen_core[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 89.700 741.890 92.000 ;
    END
  END la_oen_core[80]
  PIN la_oen_core[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 89.700 744.190 92.000 ;
    END
  END la_oen_core[81]
  PIN la_oen_core[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.750 89.700 746.030 92.000 ;
    END
  END la_oen_core[82]
  PIN la_oen_core[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 89.700 748.330 92.000 ;
    END
  END la_oen_core[83]
  PIN la_oen_core[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 89.700 750.630 92.000 ;
    END
  END la_oen_core[84]
  PIN la_oen_core[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 89.700 752.930 92.000 ;
    END
  END la_oen_core[85]
  PIN la_oen_core[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 89.700 754.770 92.000 ;
    END
  END la_oen_core[86]
  PIN la_oen_core[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 89.700 757.070 92.000 ;
    END
  END la_oen_core[87]
  PIN la_oen_core[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 89.700 759.370 92.000 ;
    END
  END la_oen_core[88]
  PIN la_oen_core[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.930 89.700 761.210 92.000 ;
    END
  END la_oen_core[89]
  PIN la_oen_core[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.750 89.700 585.030 92.000 ;
    END
  END la_oen_core[8]
  PIN la_oen_core[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 89.700 763.510 92.000 ;
    END
  END la_oen_core[90]
  PIN la_oen_core[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.530 89.700 765.810 92.000 ;
    END
  END la_oen_core[91]
  PIN la_oen_core[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 89.700 768.110 92.000 ;
    END
  END la_oen_core[92]
  PIN la_oen_core[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 89.700 769.950 92.000 ;
    END
  END la_oen_core[93]
  PIN la_oen_core[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 89.700 772.250 92.000 ;
    END
  END la_oen_core[94]
  PIN la_oen_core[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.270 89.700 774.550 92.000 ;
    END
  END la_oen_core[95]
  PIN la_oen_core[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 89.700 776.850 92.000 ;
    END
  END la_oen_core[96]
  PIN la_oen_core[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.410 89.700 778.690 92.000 ;
    END
  END la_oen_core[97]
  PIN la_oen_core[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.710 89.700 780.990 92.000 ;
    END
  END la_oen_core[98]
  PIN la_oen_core[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 89.700 783.290 92.000 ;
    END
  END la_oen_core[99]
  PIN la_oen_core[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 89.700 587.330 92.000 ;
    END
  END la_oen_core[9]
  PIN la_oen_mprj[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 -2.000 558.810 0.300 ;
    END
  END la_oen_mprj[0]
  PIN la_oen_mprj[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 -2.000 776.850 0.300 ;
    END
  END la_oen_mprj[100]
  PIN la_oen_mprj[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.410 -2.000 778.690 0.300 ;
    END
  END la_oen_mprj[101]
  PIN la_oen_mprj[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.710 -2.000 780.990 0.300 ;
    END
  END la_oen_mprj[102]
  PIN la_oen_mprj[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 -2.000 783.290 0.300 ;
    END
  END la_oen_mprj[103]
  PIN la_oen_mprj[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 -2.000 785.590 0.300 ;
    END
  END la_oen_mprj[104]
  PIN la_oen_mprj[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 -2.000 787.430 0.300 ;
    END
  END la_oen_mprj[105]
  PIN la_oen_mprj[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 -2.000 789.730 0.300 ;
    END
  END la_oen_mprj[106]
  PIN la_oen_mprj[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.750 -2.000 792.030 0.300 ;
    END
  END la_oen_mprj[107]
  PIN la_oen_mprj[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 -2.000 794.330 0.300 ;
    END
  END la_oen_mprj[108]
  PIN la_oen_mprj[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 -2.000 796.170 0.300 ;
    END
  END la_oen_mprj[109]
  PIN la_oen_mprj[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 -2.000 580.430 0.300 ;
    END
  END la_oen_mprj[10]
  PIN la_oen_mprj[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 -2.000 798.470 0.300 ;
    END
  END la_oen_mprj[110]
  PIN la_oen_mprj[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.490 -2.000 800.770 0.300 ;
    END
  END la_oen_mprj[111]
  PIN la_oen_mprj[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.330 -2.000 802.610 0.300 ;
    END
  END la_oen_mprj[112]
  PIN la_oen_mprj[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.630 -2.000 804.910 0.300 ;
    END
  END la_oen_mprj[113]
  PIN la_oen_mprj[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.930 -2.000 807.210 0.300 ;
    END
  END la_oen_mprj[114]
  PIN la_oen_mprj[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.230 -2.000 809.510 0.300 ;
    END
  END la_oen_mprj[115]
  PIN la_oen_mprj[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.070 -2.000 811.350 0.300 ;
    END
  END la_oen_mprj[116]
  PIN la_oen_mprj[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.370 -2.000 813.650 0.300 ;
    END
  END la_oen_mprj[117]
  PIN la_oen_mprj[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.670 -2.000 815.950 0.300 ;
    END
  END la_oen_mprj[118]
  PIN la_oen_mprj[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 -2.000 818.250 0.300 ;
    END
  END la_oen_mprj[119]
  PIN la_oen_mprj[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 -2.000 582.730 0.300 ;
    END
  END la_oen_mprj[11]
  PIN la_oen_mprj[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 -2.000 820.090 0.300 ;
    END
  END la_oen_mprj[120]
  PIN la_oen_mprj[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.110 -2.000 822.390 0.300 ;
    END
  END la_oen_mprj[121]
  PIN la_oen_mprj[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 -2.000 824.690 0.300 ;
    END
  END la_oen_mprj[122]
  PIN la_oen_mprj[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.710 -2.000 826.990 0.300 ;
    END
  END la_oen_mprj[123]
  PIN la_oen_mprj[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.550 -2.000 828.830 0.300 ;
    END
  END la_oen_mprj[124]
  PIN la_oen_mprj[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 -2.000 831.130 0.300 ;
    END
  END la_oen_mprj[125]
  PIN la_oen_mprj[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 -2.000 833.430 0.300 ;
    END
  END la_oen_mprj[126]
  PIN la_oen_mprj[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.450 -2.000 835.730 0.300 ;
    END
  END la_oen_mprj[127]
  PIN la_oen_mprj[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.750 -2.000 585.030 0.300 ;
    END
  END la_oen_mprj[12]
  PIN la_oen_mprj[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 -2.000 587.330 0.300 ;
    END
  END la_oen_mprj[13]
  PIN la_oen_mprj[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 -2.000 589.170 0.300 ;
    END
  END la_oen_mprj[14]
  PIN la_oen_mprj[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 -2.000 591.470 0.300 ;
    END
  END la_oen_mprj[15]
  PIN la_oen_mprj[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 -2.000 593.770 0.300 ;
    END
  END la_oen_mprj[16]
  PIN la_oen_mprj[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 -2.000 596.070 0.300 ;
    END
  END la_oen_mprj[17]
  PIN la_oen_mprj[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 -2.000 597.910 0.300 ;
    END
  END la_oen_mprj[18]
  PIN la_oen_mprj[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 -2.000 600.210 0.300 ;
    END
  END la_oen_mprj[19]
  PIN la_oen_mprj[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 -2.000 561.110 0.300 ;
    END
  END la_oen_mprj[1]
  PIN la_oen_mprj[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 -2.000 602.510 0.300 ;
    END
  END la_oen_mprj[20]
  PIN la_oen_mprj[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 -2.000 604.350 0.300 ;
    END
  END la_oen_mprj[21]
  PIN la_oen_mprj[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 -2.000 606.650 0.300 ;
    END
  END la_oen_mprj[22]
  PIN la_oen_mprj[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 -2.000 608.950 0.300 ;
    END
  END la_oen_mprj[23]
  PIN la_oen_mprj[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 -2.000 611.250 0.300 ;
    END
  END la_oen_mprj[24]
  PIN la_oen_mprj[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 -2.000 613.090 0.300 ;
    END
  END la_oen_mprj[25]
  PIN la_oen_mprj[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 -2.000 615.390 0.300 ;
    END
  END la_oen_mprj[26]
  PIN la_oen_mprj[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 -2.000 617.690 0.300 ;
    END
  END la_oen_mprj[27]
  PIN la_oen_mprj[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 -2.000 619.990 0.300 ;
    END
  END la_oen_mprj[28]
  PIN la_oen_mprj[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 -2.000 621.830 0.300 ;
    END
  END la_oen_mprj[29]
  PIN la_oen_mprj[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 -2.000 562.950 0.300 ;
    END
  END la_oen_mprj[2]
  PIN la_oen_mprj[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 -2.000 624.130 0.300 ;
    END
  END la_oen_mprj[30]
  PIN la_oen_mprj[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.150 -2.000 626.430 0.300 ;
    END
  END la_oen_mprj[31]
  PIN la_oen_mprj[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 -2.000 628.730 0.300 ;
    END
  END la_oen_mprj[32]
  PIN la_oen_mprj[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 -2.000 630.570 0.300 ;
    END
  END la_oen_mprj[33]
  PIN la_oen_mprj[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.590 -2.000 632.870 0.300 ;
    END
  END la_oen_mprj[34]
  PIN la_oen_mprj[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 -2.000 635.170 0.300 ;
    END
  END la_oen_mprj[35]
  PIN la_oen_mprj[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 -2.000 637.470 0.300 ;
    END
  END la_oen_mprj[36]
  PIN la_oen_mprj[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 -2.000 639.310 0.300 ;
    END
  END la_oen_mprj[37]
  PIN la_oen_mprj[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 -2.000 641.610 0.300 ;
    END
  END la_oen_mprj[38]
  PIN la_oen_mprj[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.630 -2.000 643.910 0.300 ;
    END
  END la_oen_mprj[39]
  PIN la_oen_mprj[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 -2.000 565.250 0.300 ;
    END
  END la_oen_mprj[3]
  PIN la_oen_mprj[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.470 -2.000 645.750 0.300 ;
    END
  END la_oen_mprj[40]
  PIN la_oen_mprj[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.770 -2.000 648.050 0.300 ;
    END
  END la_oen_mprj[41]
  PIN la_oen_mprj[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 -2.000 650.350 0.300 ;
    END
  END la_oen_mprj[42]
  PIN la_oen_mprj[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 -2.000 652.650 0.300 ;
    END
  END la_oen_mprj[43]
  PIN la_oen_mprj[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 -2.000 654.490 0.300 ;
    END
  END la_oen_mprj[44]
  PIN la_oen_mprj[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 -2.000 656.790 0.300 ;
    END
  END la_oen_mprj[45]
  PIN la_oen_mprj[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.810 -2.000 659.090 0.300 ;
    END
  END la_oen_mprj[46]
  PIN la_oen_mprj[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 -2.000 661.390 0.300 ;
    END
  END la_oen_mprj[47]
  PIN la_oen_mprj[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.950 -2.000 663.230 0.300 ;
    END
  END la_oen_mprj[48]
  PIN la_oen_mprj[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.250 -2.000 665.530 0.300 ;
    END
  END la_oen_mprj[49]
  PIN la_oen_mprj[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 -2.000 567.550 0.300 ;
    END
  END la_oen_mprj[4]
  PIN la_oen_mprj[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 -2.000 667.830 0.300 ;
    END
  END la_oen_mprj[50]
  PIN la_oen_mprj[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 -2.000 670.130 0.300 ;
    END
  END la_oen_mprj[51]
  PIN la_oen_mprj[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.690 -2.000 671.970 0.300 ;
    END
  END la_oen_mprj[52]
  PIN la_oen_mprj[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 -2.000 674.270 0.300 ;
    END
  END la_oen_mprj[53]
  PIN la_oen_mprj[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 -2.000 676.570 0.300 ;
    END
  END la_oen_mprj[54]
  PIN la_oen_mprj[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.590 -2.000 678.870 0.300 ;
    END
  END la_oen_mprj[55]
  PIN la_oen_mprj[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 -2.000 680.710 0.300 ;
    END
  END la_oen_mprj[56]
  PIN la_oen_mprj[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 -2.000 683.010 0.300 ;
    END
  END la_oen_mprj[57]
  PIN la_oen_mprj[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 -2.000 685.310 0.300 ;
    END
  END la_oen_mprj[58]
  PIN la_oen_mprj[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.870 -2.000 687.150 0.300 ;
    END
  END la_oen_mprj[59]
  PIN la_oen_mprj[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 -2.000 569.850 0.300 ;
    END
  END la_oen_mprj[5]
  PIN la_oen_mprj[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 -2.000 689.450 0.300 ;
    END
  END la_oen_mprj[60]
  PIN la_oen_mprj[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.470 -2.000 691.750 0.300 ;
    END
  END la_oen_mprj[61]
  PIN la_oen_mprj[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 -2.000 694.050 0.300 ;
    END
  END la_oen_mprj[62]
  PIN la_oen_mprj[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 -2.000 695.890 0.300 ;
    END
  END la_oen_mprj[63]
  PIN la_oen_mprj[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.910 -2.000 698.190 0.300 ;
    END
  END la_oen_mprj[64]
  PIN la_oen_mprj[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 -2.000 700.490 0.300 ;
    END
  END la_oen_mprj[65]
  PIN la_oen_mprj[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 -2.000 702.790 0.300 ;
    END
  END la_oen_mprj[66]
  PIN la_oen_mprj[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.350 -2.000 704.630 0.300 ;
    END
  END la_oen_mprj[67]
  PIN la_oen_mprj[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.650 -2.000 706.930 0.300 ;
    END
  END la_oen_mprj[68]
  PIN la_oen_mprj[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.950 -2.000 709.230 0.300 ;
    END
  END la_oen_mprj[69]
  PIN la_oen_mprj[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 -2.000 571.690 0.300 ;
    END
  END la_oen_mprj[6]
  PIN la_oen_mprj[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 -2.000 711.530 0.300 ;
    END
  END la_oen_mprj[70]
  PIN la_oen_mprj[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 -2.000 713.370 0.300 ;
    END
  END la_oen_mprj[71]
  PIN la_oen_mprj[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 -2.000 715.670 0.300 ;
    END
  END la_oen_mprj[72]
  PIN la_oen_mprj[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 -2.000 717.970 0.300 ;
    END
  END la_oen_mprj[73]
  PIN la_oen_mprj[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.990 -2.000 720.270 0.300 ;
    END
  END la_oen_mprj[74]
  PIN la_oen_mprj[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.830 -2.000 722.110 0.300 ;
    END
  END la_oen_mprj[75]
  PIN la_oen_mprj[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 -2.000 724.410 0.300 ;
    END
  END la_oen_mprj[76]
  PIN la_oen_mprj[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.430 -2.000 726.710 0.300 ;
    END
  END la_oen_mprj[77]
  PIN la_oen_mprj[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.270 -2.000 728.550 0.300 ;
    END
  END la_oen_mprj[78]
  PIN la_oen_mprj[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.570 -2.000 730.850 0.300 ;
    END
  END la_oen_mprj[79]
  PIN la_oen_mprj[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.710 -2.000 573.990 0.300 ;
    END
  END la_oen_mprj[7]
  PIN la_oen_mprj[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 -2.000 733.150 0.300 ;
    END
  END la_oen_mprj[80]
  PIN la_oen_mprj[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 -2.000 735.450 0.300 ;
    END
  END la_oen_mprj[81]
  PIN la_oen_mprj[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 -2.000 737.290 0.300 ;
    END
  END la_oen_mprj[82]
  PIN la_oen_mprj[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.310 -2.000 739.590 0.300 ;
    END
  END la_oen_mprj[83]
  PIN la_oen_mprj[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 -2.000 741.890 0.300 ;
    END
  END la_oen_mprj[84]
  PIN la_oen_mprj[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 -2.000 744.190 0.300 ;
    END
  END la_oen_mprj[85]
  PIN la_oen_mprj[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.750 -2.000 746.030 0.300 ;
    END
  END la_oen_mprj[86]
  PIN la_oen_mprj[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 -2.000 748.330 0.300 ;
    END
  END la_oen_mprj[87]
  PIN la_oen_mprj[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 -2.000 750.630 0.300 ;
    END
  END la_oen_mprj[88]
  PIN la_oen_mprj[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 -2.000 752.930 0.300 ;
    END
  END la_oen_mprj[89]
  PIN la_oen_mprj[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 -2.000 576.290 0.300 ;
    END
  END la_oen_mprj[8]
  PIN la_oen_mprj[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 -2.000 754.770 0.300 ;
    END
  END la_oen_mprj[90]
  PIN la_oen_mprj[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 -2.000 757.070 0.300 ;
    END
  END la_oen_mprj[91]
  PIN la_oen_mprj[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 -2.000 759.370 0.300 ;
    END
  END la_oen_mprj[92]
  PIN la_oen_mprj[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.930 -2.000 761.210 0.300 ;
    END
  END la_oen_mprj[93]
  PIN la_oen_mprj[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 -2.000 763.510 0.300 ;
    END
  END la_oen_mprj[94]
  PIN la_oen_mprj[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.530 -2.000 765.810 0.300 ;
    END
  END la_oen_mprj[95]
  PIN la_oen_mprj[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 -2.000 768.110 0.300 ;
    END
  END la_oen_mprj[96]
  PIN la_oen_mprj[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 -2.000 769.950 0.300 ;
    END
  END la_oen_mprj[97]
  PIN la_oen_mprj[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 -2.000 772.250 0.300 ;
    END
  END la_oen_mprj[98]
  PIN la_oen_mprj[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.270 -2.000 774.550 0.300 ;
    END
  END la_oen_mprj[99]
  PIN la_oen_mprj[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 -2.000 578.590 0.300 ;
    END
  END la_oen_mprj[9]
  PIN mprj_adr_o_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 -2.000 844.010 0.300 ;
    END
  END mprj_adr_o_core[0]
  PIN mprj_adr_o_core[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.170 -2.000 896.450 0.300 ;
    END
  END mprj_adr_o_core[10]
  PIN mprj_adr_o_core[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.770 -2.000 901.050 0.300 ;
    END
  END mprj_adr_o_core[11]
  PIN mprj_adr_o_core[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 -2.000 905.190 0.300 ;
    END
  END mprj_adr_o_core[12]
  PIN mprj_adr_o_core[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 -2.000 909.790 0.300 ;
    END
  END mprj_adr_o_core[13]
  PIN mprj_adr_o_core[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.650 -2.000 913.930 0.300 ;
    END
  END mprj_adr_o_core[14]
  PIN mprj_adr_o_core[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.250 -2.000 918.530 0.300 ;
    END
  END mprj_adr_o_core[15]
  PIN mprj_adr_o_core[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.390 -2.000 922.670 0.300 ;
    END
  END mprj_adr_o_core[16]
  PIN mprj_adr_o_core[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.530 -2.000 926.810 0.300 ;
    END
  END mprj_adr_o_core[17]
  PIN mprj_adr_o_core[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.130 -2.000 931.410 0.300 ;
    END
  END mprj_adr_o_core[18]
  PIN mprj_adr_o_core[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.270 -2.000 935.550 0.300 ;
    END
  END mprj_adr_o_core[19]
  PIN mprj_adr_o_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.630 -2.000 850.910 0.300 ;
    END
  END mprj_adr_o_core[1]
  PIN mprj_adr_o_core[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.870 -2.000 940.150 0.300 ;
    END
  END mprj_adr_o_core[20]
  PIN mprj_adr_o_core[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.010 -2.000 944.290 0.300 ;
    END
  END mprj_adr_o_core[21]
  PIN mprj_adr_o_core[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.610 -2.000 948.890 0.300 ;
    END
  END mprj_adr_o_core[22]
  PIN mprj_adr_o_core[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.750 -2.000 953.030 0.300 ;
    END
  END mprj_adr_o_core[23]
  PIN mprj_adr_o_core[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.350 -2.000 957.630 0.300 ;
    END
  END mprj_adr_o_core[24]
  PIN mprj_adr_o_core[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.490 -2.000 961.770 0.300 ;
    END
  END mprj_adr_o_core[25]
  PIN mprj_adr_o_core[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 -2.000 966.370 0.300 ;
    END
  END mprj_adr_o_core[26]
  PIN mprj_adr_o_core[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.230 -2.000 970.510 0.300 ;
    END
  END mprj_adr_o_core[27]
  PIN mprj_adr_o_core[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.830 -2.000 975.110 0.300 ;
    END
  END mprj_adr_o_core[28]
  PIN mprj_adr_o_core[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 -2.000 979.250 0.300 ;
    END
  END mprj_adr_o_core[29]
  PIN mprj_adr_o_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.070 -2.000 857.350 0.300 ;
    END
  END mprj_adr_o_core[2]
  PIN mprj_adr_o_core[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.570 -2.000 983.850 0.300 ;
    END
  END mprj_adr_o_core[30]
  PIN mprj_adr_o_core[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.710 -2.000 987.990 0.300 ;
    END
  END mprj_adr_o_core[31]
  PIN mprj_adr_o_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.510 -2.000 863.790 0.300 ;
    END
  END mprj_adr_o_core[3]
  PIN mprj_adr_o_core[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.950 -2.000 870.230 0.300 ;
    END
  END mprj_adr_o_core[4]
  PIN mprj_adr_o_core[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.550 -2.000 874.830 0.300 ;
    END
  END mprj_adr_o_core[5]
  PIN mprj_adr_o_core[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.690 -2.000 878.970 0.300 ;
    END
  END mprj_adr_o_core[6]
  PIN mprj_adr_o_core[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.290 -2.000 883.570 0.300 ;
    END
  END mprj_adr_o_core[7]
  PIN mprj_adr_o_core[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.430 -2.000 887.710 0.300 ;
    END
  END mprj_adr_o_core[8]
  PIN mprj_adr_o_core[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 -2.000 892.310 0.300 ;
    END
  END mprj_adr_o_core[9]
  PIN mprj_adr_o_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.470 89.700 852.750 92.000 ;
    END
  END mprj_adr_o_user[0]
  PIN mprj_adr_o_user[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 89.700 905.190 92.000 ;
    END
  END mprj_adr_o_user[10]
  PIN mprj_adr_o_user[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 89.700 909.790 92.000 ;
    END
  END mprj_adr_o_user[11]
  PIN mprj_adr_o_user[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.650 89.700 913.930 92.000 ;
    END
  END mprj_adr_o_user[12]
  PIN mprj_adr_o_user[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.250 89.700 918.530 92.000 ;
    END
  END mprj_adr_o_user[13]
  PIN mprj_adr_o_user[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.390 89.700 922.670 92.000 ;
    END
  END mprj_adr_o_user[14]
  PIN mprj_adr_o_user[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.530 89.700 926.810 92.000 ;
    END
  END mprj_adr_o_user[15]
  PIN mprj_adr_o_user[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.130 89.700 931.410 92.000 ;
    END
  END mprj_adr_o_user[16]
  PIN mprj_adr_o_user[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.270 89.700 935.550 92.000 ;
    END
  END mprj_adr_o_user[17]
  PIN mprj_adr_o_user[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.870 89.700 940.150 92.000 ;
    END
  END mprj_adr_o_user[18]
  PIN mprj_adr_o_user[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.010 89.700 944.290 92.000 ;
    END
  END mprj_adr_o_user[19]
  PIN mprj_adr_o_user[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.370 89.700 859.650 92.000 ;
    END
  END mprj_adr_o_user[1]
  PIN mprj_adr_o_user[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.610 89.700 948.890 92.000 ;
    END
  END mprj_adr_o_user[20]
  PIN mprj_adr_o_user[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.750 89.700 953.030 92.000 ;
    END
  END mprj_adr_o_user[21]
  PIN mprj_adr_o_user[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.350 89.700 957.630 92.000 ;
    END
  END mprj_adr_o_user[22]
  PIN mprj_adr_o_user[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.490 89.700 961.770 92.000 ;
    END
  END mprj_adr_o_user[23]
  PIN mprj_adr_o_user[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 89.700 966.370 92.000 ;
    END
  END mprj_adr_o_user[24]
  PIN mprj_adr_o_user[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.230 89.700 970.510 92.000 ;
    END
  END mprj_adr_o_user[25]
  PIN mprj_adr_o_user[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.830 89.700 975.110 92.000 ;
    END
  END mprj_adr_o_user[26]
  PIN mprj_adr_o_user[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 89.700 979.250 92.000 ;
    END
  END mprj_adr_o_user[27]
  PIN mprj_adr_o_user[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.570 89.700 983.850 92.000 ;
    END
  END mprj_adr_o_user[28]
  PIN mprj_adr_o_user[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.710 89.700 987.990 92.000 ;
    END
  END mprj_adr_o_user[29]
  PIN mprj_adr_o_user[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.810 89.700 866.090 92.000 ;
    END
  END mprj_adr_o_user[2]
  PIN mprj_adr_o_user[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.310 89.700 992.590 92.000 ;
    END
  END mprj_adr_o_user[30]
  PIN mprj_adr_o_user[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.450 89.700 996.730 92.000 ;
    END
  END mprj_adr_o_user[31]
  PIN mprj_adr_o_user[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 89.700 872.530 92.000 ;
    END
  END mprj_adr_o_user[3]
  PIN mprj_adr_o_user[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.690 89.700 878.970 92.000 ;
    END
  END mprj_adr_o_user[4]
  PIN mprj_adr_o_user[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.290 89.700 883.570 92.000 ;
    END
  END mprj_adr_o_user[5]
  PIN mprj_adr_o_user[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.430 89.700 887.710 92.000 ;
    END
  END mprj_adr_o_user[6]
  PIN mprj_adr_o_user[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 89.700 892.310 92.000 ;
    END
  END mprj_adr_o_user[7]
  PIN mprj_adr_o_user[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.170 89.700 896.450 92.000 ;
    END
  END mprj_adr_o_user[8]
  PIN mprj_adr_o_user[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.770 89.700 901.050 92.000 ;
    END
  END mprj_adr_o_user[9]
  PIN mprj_cyc_o_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 -2.000 837.570 0.300 ;
    END
  END mprj_cyc_o_core
  PIN mprj_cyc_o_user
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.030 89.700 846.310 92.000 ;
    END
  END mprj_cyc_o_user
  PIN mprj_dat_o_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.030 -2.000 846.310 0.300 ;
    END
  END mprj_dat_o_core[0]
  PIN mprj_dat_o_core[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 -2.000 898.750 0.300 ;
    END
  END mprj_dat_o_core[10]
  PIN mprj_dat_o_core[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.610 -2.000 902.890 0.300 ;
    END
  END mprj_dat_o_core[11]
  PIN mprj_dat_o_core[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.210 -2.000 907.490 0.300 ;
    END
  END mprj_dat_o_core[12]
  PIN mprj_dat_o_core[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 -2.000 911.630 0.300 ;
    END
  END mprj_dat_o_core[13]
  PIN mprj_dat_o_core[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.950 -2.000 916.230 0.300 ;
    END
  END mprj_dat_o_core[14]
  PIN mprj_dat_o_core[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.090 -2.000 920.370 0.300 ;
    END
  END mprj_dat_o_core[15]
  PIN mprj_dat_o_core[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.690 -2.000 924.970 0.300 ;
    END
  END mprj_dat_o_core[16]
  PIN mprj_dat_o_core[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.830 -2.000 929.110 0.300 ;
    END
  END mprj_dat_o_core[17]
  PIN mprj_dat_o_core[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.430 -2.000 933.710 0.300 ;
    END
  END mprj_dat_o_core[18]
  PIN mprj_dat_o_core[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.570 -2.000 937.850 0.300 ;
    END
  END mprj_dat_o_core[19]
  PIN mprj_dat_o_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.470 -2.000 852.750 0.300 ;
    END
  END mprj_dat_o_core[1]
  PIN mprj_dat_o_core[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.170 -2.000 942.450 0.300 ;
    END
  END mprj_dat_o_core[20]
  PIN mprj_dat_o_core[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.310 -2.000 946.590 0.300 ;
    END
  END mprj_dat_o_core[21]
  PIN mprj_dat_o_core[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.910 -2.000 951.190 0.300 ;
    END
  END mprj_dat_o_core[22]
  PIN mprj_dat_o_core[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 -2.000 955.330 0.300 ;
    END
  END mprj_dat_o_core[23]
  PIN mprj_dat_o_core[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 -2.000 959.930 0.300 ;
    END
  END mprj_dat_o_core[24]
  PIN mprj_dat_o_core[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.790 -2.000 964.070 0.300 ;
    END
  END mprj_dat_o_core[25]
  PIN mprj_dat_o_core[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.930 -2.000 968.210 0.300 ;
    END
  END mprj_dat_o_core[26]
  PIN mprj_dat_o_core[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 -2.000 972.810 0.300 ;
    END
  END mprj_dat_o_core[27]
  PIN mprj_dat_o_core[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.670 -2.000 976.950 0.300 ;
    END
  END mprj_dat_o_core[28]
  PIN mprj_dat_o_core[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.270 -2.000 981.550 0.300 ;
    END
  END mprj_dat_o_core[29]
  PIN mprj_dat_o_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.370 -2.000 859.650 0.300 ;
    END
  END mprj_dat_o_core[2]
  PIN mprj_dat_o_core[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 -2.000 985.690 0.300 ;
    END
  END mprj_dat_o_core[30]
  PIN mprj_dat_o_core[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.010 -2.000 990.290 0.300 ;
    END
  END mprj_dat_o_core[31]
  PIN mprj_dat_o_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.810 -2.000 866.090 0.300 ;
    END
  END mprj_dat_o_core[3]
  PIN mprj_dat_o_core[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 -2.000 872.530 0.300 ;
    END
  END mprj_dat_o_core[4]
  PIN mprj_dat_o_core[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.850 -2.000 877.130 0.300 ;
    END
  END mprj_dat_o_core[5]
  PIN mprj_dat_o_core[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.990 -2.000 881.270 0.300 ;
    END
  END mprj_dat_o_core[6]
  PIN mprj_dat_o_core[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.130 -2.000 885.410 0.300 ;
    END
  END mprj_dat_o_core[7]
  PIN mprj_dat_o_core[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.730 -2.000 890.010 0.300 ;
    END
  END mprj_dat_o_core[8]
  PIN mprj_dat_o_core[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.870 -2.000 894.150 0.300 ;
    END
  END mprj_dat_o_core[9]
  PIN mprj_dat_o_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.770 89.700 855.050 92.000 ;
    END
  END mprj_dat_o_user[0]
  PIN mprj_dat_o_user[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.210 89.700 907.490 92.000 ;
    END
  END mprj_dat_o_user[10]
  PIN mprj_dat_o_user[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 89.700 911.630 92.000 ;
    END
  END mprj_dat_o_user[11]
  PIN mprj_dat_o_user[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.950 89.700 916.230 92.000 ;
    END
  END mprj_dat_o_user[12]
  PIN mprj_dat_o_user[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.090 89.700 920.370 92.000 ;
    END
  END mprj_dat_o_user[13]
  PIN mprj_dat_o_user[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.690 89.700 924.970 92.000 ;
    END
  END mprj_dat_o_user[14]
  PIN mprj_dat_o_user[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.830 89.700 929.110 92.000 ;
    END
  END mprj_dat_o_user[15]
  PIN mprj_dat_o_user[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.430 89.700 933.710 92.000 ;
    END
  END mprj_dat_o_user[16]
  PIN mprj_dat_o_user[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.570 89.700 937.850 92.000 ;
    END
  END mprj_dat_o_user[17]
  PIN mprj_dat_o_user[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.170 89.700 942.450 92.000 ;
    END
  END mprj_dat_o_user[18]
  PIN mprj_dat_o_user[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.310 89.700 946.590 92.000 ;
    END
  END mprj_dat_o_user[19]
  PIN mprj_dat_o_user[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.210 89.700 861.490 92.000 ;
    END
  END mprj_dat_o_user[1]
  PIN mprj_dat_o_user[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.910 89.700 951.190 92.000 ;
    END
  END mprj_dat_o_user[20]
  PIN mprj_dat_o_user[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 89.700 955.330 92.000 ;
    END
  END mprj_dat_o_user[21]
  PIN mprj_dat_o_user[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 89.700 959.930 92.000 ;
    END
  END mprj_dat_o_user[22]
  PIN mprj_dat_o_user[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.790 89.700 964.070 92.000 ;
    END
  END mprj_dat_o_user[23]
  PIN mprj_dat_o_user[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.930 89.700 968.210 92.000 ;
    END
  END mprj_dat_o_user[24]
  PIN mprj_dat_o_user[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 89.700 972.810 92.000 ;
    END
  END mprj_dat_o_user[25]
  PIN mprj_dat_o_user[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.670 89.700 976.950 92.000 ;
    END
  END mprj_dat_o_user[26]
  PIN mprj_dat_o_user[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.270 89.700 981.550 92.000 ;
    END
  END mprj_dat_o_user[27]
  PIN mprj_dat_o_user[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 89.700 985.690 92.000 ;
    END
  END mprj_dat_o_user[28]
  PIN mprj_dat_o_user[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.010 89.700 990.290 92.000 ;
    END
  END mprj_dat_o_user[29]
  PIN mprj_dat_o_user[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.110 89.700 868.390 92.000 ;
    END
  END mprj_dat_o_user[2]
  PIN mprj_dat_o_user[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.150 89.700 994.430 92.000 ;
    END
  END mprj_dat_o_user[30]
  PIN mprj_dat_o_user[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 89.700 999.030 92.000 ;
    END
  END mprj_dat_o_user[31]
  PIN mprj_dat_o_user[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.550 89.700 874.830 92.000 ;
    END
  END mprj_dat_o_user[3]
  PIN mprj_dat_o_user[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.990 89.700 881.270 92.000 ;
    END
  END mprj_dat_o_user[4]
  PIN mprj_dat_o_user[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.130 89.700 885.410 92.000 ;
    END
  END mprj_dat_o_user[5]
  PIN mprj_dat_o_user[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.730 89.700 890.010 92.000 ;
    END
  END mprj_dat_o_user[6]
  PIN mprj_dat_o_user[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.870 89.700 894.150 92.000 ;
    END
  END mprj_dat_o_user[7]
  PIN mprj_dat_o_user[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 89.700 898.750 92.000 ;
    END
  END mprj_dat_o_user[8]
  PIN mprj_dat_o_user[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.610 89.700 902.890 92.000 ;
    END
  END mprj_dat_o_user[9]
  PIN mprj_sel_o_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.330 -2.000 848.610 0.300 ;
    END
  END mprj_sel_o_core[0]
  PIN mprj_sel_o_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.770 -2.000 855.050 0.300 ;
    END
  END mprj_sel_o_core[1]
  PIN mprj_sel_o_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.210 -2.000 861.490 0.300 ;
    END
  END mprj_sel_o_core[2]
  PIN mprj_sel_o_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.110 -2.000 868.390 0.300 ;
    END
  END mprj_sel_o_core[3]
  PIN mprj_sel_o_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.070 89.700 857.350 92.000 ;
    END
  END mprj_sel_o_user[0]
  PIN mprj_sel_o_user[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.510 89.700 863.790 92.000 ;
    END
  END mprj_sel_o_user[1]
  PIN mprj_sel_o_user[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.950 89.700 870.230 92.000 ;
    END
  END mprj_sel_o_user[2]
  PIN mprj_sel_o_user[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.850 89.700 877.130 92.000 ;
    END
  END mprj_sel_o_user[3]
  PIN mprj_stb_o_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.590 -2.000 839.870 0.300 ;
    END
  END mprj_stb_o_core
  PIN mprj_stb_o_user
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.330 89.700 848.610 92.000 ;
    END
  END mprj_stb_o_user
  PIN mprj_we_o_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.890 -2.000 842.170 0.300 ;
    END
  END mprj_we_o_core
  PIN mprj_we_o_user
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.630 89.700 850.910 92.000 ;
    END
  END mprj_we_o_user
  PIN user1_vcc_powergood
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.310 -2.000 992.590 0.300 ;
    END
  END user1_vcc_powergood
  PIN user1_vdd_powergood
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.150 -2.000 994.430 0.300 ;
    END
  END user1_vdd_powergood
  PIN user2_vcc_powergood
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.450 -2.000 996.730 0.300 ;
    END
  END user2_vcc_powergood
  PIN user2_vdd_powergood
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 -2.000 999.030 0.300 ;
    END
  END user2_vdd_powergood
  PIN user_clock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 89.700 1.290 92.000 ;
    END
  END user_clock
  PIN user_clock2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 89.700 3.130 92.000 ;
    END
  END user_clock2
  PIN user_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 89.700 5.430 92.000 ;
    END
  END user_reset
  PIN user_resetn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 89.700 7.730 92.000 ;
    END
  END user_resetn
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 19.920 91.470 21.120 91.480 ;
        RECT 169.920 91.470 171.120 91.480 ;
        RECT 319.920 91.470 321.120 91.480 ;
        RECT 469.920 91.470 471.120 91.480 ;
        RECT 619.920 91.470 621.120 91.480 ;
        RECT 769.920 91.470 771.120 91.480 ;
        RECT 919.920 91.470 921.120 91.480 ;
        RECT -1.630 91.170 1001.210 91.470 ;
        RECT 19.920 91.160 21.120 91.170 ;
        RECT 169.920 91.160 171.120 91.170 ;
        RECT 319.920 91.160 321.120 91.170 ;
        RECT 469.920 91.160 471.120 91.170 ;
        RECT 619.920 91.160 621.120 91.170 ;
        RECT 769.920 91.160 771.120 91.170 ;
        RECT 919.920 91.160 921.120 91.170 ;
        RECT 19.920 -1.410 21.120 -1.400 ;
        RECT 169.920 -1.410 171.120 -1.400 ;
        RECT 319.920 -1.410 321.120 -1.400 ;
        RECT 469.920 -1.410 471.120 -1.400 ;
        RECT 619.920 -1.410 621.120 -1.400 ;
        RECT 769.920 -1.410 771.120 -1.400 ;
        RECT 919.920 -1.410 921.120 -1.400 ;
        RECT -1.630 -1.710 1001.210 -1.410 ;
        RECT 19.920 -1.720 21.120 -1.710 ;
        RECT 169.920 -1.720 171.120 -1.710 ;
        RECT 319.920 -1.720 321.120 -1.710 ;
        RECT 469.920 -1.720 471.120 -1.710 ;
        RECT 619.920 -1.720 621.120 -1.710 ;
        RECT 769.920 -1.720 771.120 -1.710 ;
        RECT 919.920 -1.720 921.120 -1.710 ;
      LAYER via3 ;
        RECT 19.960 91.160 20.280 91.480 ;
        RECT 20.360 91.160 20.680 91.480 ;
        RECT 20.760 91.160 21.080 91.480 ;
        RECT 169.960 91.160 170.280 91.480 ;
        RECT 170.360 91.160 170.680 91.480 ;
        RECT 170.760 91.160 171.080 91.480 ;
        RECT 319.960 91.160 320.280 91.480 ;
        RECT 320.360 91.160 320.680 91.480 ;
        RECT 320.760 91.160 321.080 91.480 ;
        RECT 469.960 91.160 470.280 91.480 ;
        RECT 470.360 91.160 470.680 91.480 ;
        RECT 470.760 91.160 471.080 91.480 ;
        RECT 619.960 91.160 620.280 91.480 ;
        RECT 620.360 91.160 620.680 91.480 ;
        RECT 620.760 91.160 621.080 91.480 ;
        RECT 769.960 91.160 770.280 91.480 ;
        RECT 770.360 91.160 770.680 91.480 ;
        RECT 770.760 91.160 771.080 91.480 ;
        RECT 919.960 91.160 920.280 91.480 ;
        RECT 920.360 91.160 920.680 91.480 ;
        RECT 920.760 91.160 921.080 91.480 ;
        RECT 19.960 -1.720 20.280 -1.400 ;
        RECT 20.360 -1.720 20.680 -1.400 ;
        RECT 20.760 -1.720 21.080 -1.400 ;
        RECT 169.960 -1.720 170.280 -1.400 ;
        RECT 170.360 -1.720 170.680 -1.400 ;
        RECT 170.760 -1.720 171.080 -1.400 ;
        RECT 319.960 -1.720 320.280 -1.400 ;
        RECT 320.360 -1.720 320.680 -1.400 ;
        RECT 320.760 -1.720 321.080 -1.400 ;
        RECT 469.960 -1.720 470.280 -1.400 ;
        RECT 470.360 -1.720 470.680 -1.400 ;
        RECT 470.760 -1.720 471.080 -1.400 ;
        RECT 619.960 -1.720 620.280 -1.400 ;
        RECT 620.360 -1.720 620.680 -1.400 ;
        RECT 620.760 -1.720 621.080 -1.400 ;
        RECT 769.960 -1.720 770.280 -1.400 ;
        RECT 770.360 -1.720 770.680 -1.400 ;
        RECT 770.760 -1.720 771.080 -1.400 ;
        RECT 919.960 -1.720 920.280 -1.400 ;
        RECT 920.360 -1.720 920.680 -1.400 ;
        RECT 920.760 -1.720 921.080 -1.400 ;
      LAYER met4 ;
        RECT 19.920 89.700 21.120 92.170 ;
        RECT 169.920 89.700 171.120 92.170 ;
        RECT 319.920 89.700 321.120 92.170 ;
        RECT 469.920 89.700 471.120 92.170 ;
        RECT 619.920 89.700 621.120 92.170 ;
        RECT 769.920 89.700 771.120 92.170 ;
        RECT 919.920 89.700 921.120 92.170 ;
        RECT 19.920 -2.410 21.120 0.300 ;
        RECT 169.920 -2.410 171.120 0.300 ;
        RECT 319.920 -2.410 321.120 0.300 ;
        RECT 469.920 -2.410 471.120 0.300 ;
        RECT 619.920 -2.410 621.120 0.300 ;
        RECT 769.920 -2.410 771.120 0.300 ;
        RECT 919.920 -2.410 921.120 0.300 ;
    END
  END vccd
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1000.910 -1.710 1001.210 91.470 ;
    END
  END vccd
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -1.630 -1.710 -1.330 91.470 ;
    END
  END vccd
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 94.920 92.170 96.120 92.180 ;
        RECT 244.920 92.170 246.120 92.180 ;
        RECT 394.920 92.170 396.120 92.180 ;
        RECT 544.920 92.170 546.120 92.180 ;
        RECT 694.920 92.170 696.120 92.180 ;
        RECT 844.920 92.170 846.120 92.180 ;
        RECT -2.330 91.870 1001.910 92.170 ;
        RECT 94.920 91.860 96.120 91.870 ;
        RECT 244.920 91.860 246.120 91.870 ;
        RECT 394.920 91.860 396.120 91.870 ;
        RECT 544.920 91.860 546.120 91.870 ;
        RECT 694.920 91.860 696.120 91.870 ;
        RECT 844.920 91.860 846.120 91.870 ;
        RECT 94.920 -2.110 96.120 -2.100 ;
        RECT 244.920 -2.110 246.120 -2.100 ;
        RECT 394.920 -2.110 396.120 -2.100 ;
        RECT 544.920 -2.110 546.120 -2.100 ;
        RECT 694.920 -2.110 696.120 -2.100 ;
        RECT 844.920 -2.110 846.120 -2.100 ;
        RECT -2.330 -2.410 1001.910 -2.110 ;
        RECT 94.920 -2.420 96.120 -2.410 ;
        RECT 244.920 -2.420 246.120 -2.410 ;
        RECT 394.920 -2.420 396.120 -2.410 ;
        RECT 544.920 -2.420 546.120 -2.410 ;
        RECT 694.920 -2.420 696.120 -2.410 ;
        RECT 844.920 -2.420 846.120 -2.410 ;
      LAYER via3 ;
        RECT 94.960 91.860 95.280 92.180 ;
        RECT 95.360 91.860 95.680 92.180 ;
        RECT 95.760 91.860 96.080 92.180 ;
        RECT 244.960 91.860 245.280 92.180 ;
        RECT 245.360 91.860 245.680 92.180 ;
        RECT 245.760 91.860 246.080 92.180 ;
        RECT 394.960 91.860 395.280 92.180 ;
        RECT 395.360 91.860 395.680 92.180 ;
        RECT 395.760 91.860 396.080 92.180 ;
        RECT 544.960 91.860 545.280 92.180 ;
        RECT 545.360 91.860 545.680 92.180 ;
        RECT 545.760 91.860 546.080 92.180 ;
        RECT 694.960 91.860 695.280 92.180 ;
        RECT 695.360 91.860 695.680 92.180 ;
        RECT 695.760 91.860 696.080 92.180 ;
        RECT 844.960 91.860 845.280 92.180 ;
        RECT 845.360 91.860 845.680 92.180 ;
        RECT 845.760 91.860 846.080 92.180 ;
        RECT 94.960 -2.420 95.280 -2.100 ;
        RECT 95.360 -2.420 95.680 -2.100 ;
        RECT 95.760 -2.420 96.080 -2.100 ;
        RECT 244.960 -2.420 245.280 -2.100 ;
        RECT 245.360 -2.420 245.680 -2.100 ;
        RECT 245.760 -2.420 246.080 -2.100 ;
        RECT 394.960 -2.420 395.280 -2.100 ;
        RECT 395.360 -2.420 395.680 -2.100 ;
        RECT 395.760 -2.420 396.080 -2.100 ;
        RECT 544.960 -2.420 545.280 -2.100 ;
        RECT 545.360 -2.420 545.680 -2.100 ;
        RECT 545.760 -2.420 546.080 -2.100 ;
        RECT 694.960 -2.420 695.280 -2.100 ;
        RECT 695.360 -2.420 695.680 -2.100 ;
        RECT 695.760 -2.420 696.080 -2.100 ;
        RECT 844.960 -2.420 845.280 -2.100 ;
        RECT 845.360 -2.420 845.680 -2.100 ;
        RECT 845.760 -2.420 846.080 -2.100 ;
      LAYER met4 ;
        RECT 94.920 89.700 96.120 92.185 ;
        RECT 244.920 89.700 246.120 92.185 ;
        RECT 394.920 89.700 396.120 92.185 ;
        RECT 544.920 89.700 546.120 92.185 ;
        RECT 694.920 89.700 696.120 92.185 ;
        RECT 844.920 89.700 846.120 92.185 ;
        RECT 94.920 -2.425 96.120 0.300 ;
        RECT 244.920 -2.425 246.120 0.300 ;
        RECT 394.920 -2.425 396.120 0.300 ;
        RECT 544.920 -2.425 546.120 0.300 ;
        RECT 694.920 -2.425 696.120 0.300 ;
        RECT 844.920 -2.425 846.120 0.300 ;
    END
  END vssd
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1001.610 -2.410 1001.910 92.170 ;
    END
  END vssd
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -2.330 -2.410 -2.030 92.170 ;
    END
  END vssd
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 24.320 92.870 25.520 92.880 ;
        RECT 174.320 92.870 175.520 92.880 ;
        RECT 324.320 92.870 325.520 92.880 ;
        RECT 474.320 92.870 475.520 92.880 ;
        RECT 624.320 92.870 625.520 92.880 ;
        RECT 774.320 92.870 775.520 92.880 ;
        RECT 924.320 92.870 925.520 92.880 ;
        RECT -3.030 92.570 1002.610 92.870 ;
        RECT 24.320 92.560 25.520 92.570 ;
        RECT 174.320 92.560 175.520 92.570 ;
        RECT 324.320 92.560 325.520 92.570 ;
        RECT 474.320 92.560 475.520 92.570 ;
        RECT 624.320 92.560 625.520 92.570 ;
        RECT 774.320 92.560 775.520 92.570 ;
        RECT 924.320 92.560 925.520 92.570 ;
        RECT 24.320 -2.810 25.520 -2.800 ;
        RECT 174.320 -2.810 175.520 -2.800 ;
        RECT 324.320 -2.810 325.520 -2.800 ;
        RECT 474.320 -2.810 475.520 -2.800 ;
        RECT 624.320 -2.810 625.520 -2.800 ;
        RECT 774.320 -2.810 775.520 -2.800 ;
        RECT 924.320 -2.810 925.520 -2.800 ;
        RECT -3.030 -3.110 1002.610 -2.810 ;
        RECT 24.320 -3.120 25.520 -3.110 ;
        RECT 174.320 -3.120 175.520 -3.110 ;
        RECT 324.320 -3.120 325.520 -3.110 ;
        RECT 474.320 -3.120 475.520 -3.110 ;
        RECT 624.320 -3.120 625.520 -3.110 ;
        RECT 774.320 -3.120 775.520 -3.110 ;
        RECT 924.320 -3.120 925.520 -3.110 ;
      LAYER via3 ;
        RECT 24.360 92.560 24.680 92.880 ;
        RECT 24.760 92.560 25.080 92.880 ;
        RECT 25.160 92.560 25.480 92.880 ;
        RECT 174.360 92.560 174.680 92.880 ;
        RECT 174.760 92.560 175.080 92.880 ;
        RECT 175.160 92.560 175.480 92.880 ;
        RECT 324.360 92.560 324.680 92.880 ;
        RECT 324.760 92.560 325.080 92.880 ;
        RECT 325.160 92.560 325.480 92.880 ;
        RECT 474.360 92.560 474.680 92.880 ;
        RECT 474.760 92.560 475.080 92.880 ;
        RECT 475.160 92.560 475.480 92.880 ;
        RECT 624.360 92.560 624.680 92.880 ;
        RECT 624.760 92.560 625.080 92.880 ;
        RECT 625.160 92.560 625.480 92.880 ;
        RECT 774.360 92.560 774.680 92.880 ;
        RECT 774.760 92.560 775.080 92.880 ;
        RECT 775.160 92.560 775.480 92.880 ;
        RECT 924.360 92.560 924.680 92.880 ;
        RECT 924.760 92.560 925.080 92.880 ;
        RECT 925.160 92.560 925.480 92.880 ;
        RECT 24.360 -3.120 24.680 -2.800 ;
        RECT 24.760 -3.120 25.080 -2.800 ;
        RECT 25.160 -3.120 25.480 -2.800 ;
        RECT 174.360 -3.120 174.680 -2.800 ;
        RECT 174.760 -3.120 175.080 -2.800 ;
        RECT 175.160 -3.120 175.480 -2.800 ;
        RECT 324.360 -3.120 324.680 -2.800 ;
        RECT 324.760 -3.120 325.080 -2.800 ;
        RECT 325.160 -3.120 325.480 -2.800 ;
        RECT 474.360 -3.120 474.680 -2.800 ;
        RECT 474.760 -3.120 475.080 -2.800 ;
        RECT 475.160 -3.120 475.480 -2.800 ;
        RECT 624.360 -3.120 624.680 -2.800 ;
        RECT 624.760 -3.120 625.080 -2.800 ;
        RECT 625.160 -3.120 625.480 -2.800 ;
        RECT 774.360 -3.120 774.680 -2.800 ;
        RECT 774.760 -3.120 775.080 -2.800 ;
        RECT 775.160 -3.120 775.480 -2.800 ;
        RECT 924.360 -3.120 924.680 -2.800 ;
        RECT 924.760 -3.120 925.080 -2.800 ;
        RECT 925.160 -3.120 925.480 -2.800 ;
      LAYER met4 ;
        RECT 24.320 89.700 25.520 93.570 ;
        RECT 174.320 89.700 175.520 93.570 ;
        RECT 324.320 89.700 325.520 93.570 ;
        RECT 474.320 89.700 475.520 93.570 ;
        RECT 624.320 89.700 625.520 93.570 ;
        RECT 774.320 89.700 775.520 93.570 ;
        RECT 924.320 89.700 925.520 93.570 ;
        RECT 24.320 -3.810 25.520 0.300 ;
        RECT 174.320 -3.810 175.520 0.300 ;
        RECT 324.320 -3.810 325.520 0.300 ;
        RECT 474.320 -3.810 475.520 0.300 ;
        RECT 624.320 -3.810 625.520 0.300 ;
        RECT 774.320 -3.810 775.520 0.300 ;
        RECT 924.320 -3.810 925.520 0.300 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1002.310 -3.110 1002.610 92.870 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -3.030 -3.110 -2.730 92.870 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 99.320 93.570 100.520 93.580 ;
        RECT 249.320 93.570 250.520 93.580 ;
        RECT 399.320 93.570 400.520 93.580 ;
        RECT 549.320 93.570 550.520 93.580 ;
        RECT 699.320 93.570 700.520 93.580 ;
        RECT 849.320 93.570 850.520 93.580 ;
        RECT -3.730 93.270 1003.310 93.570 ;
        RECT 99.320 93.260 100.520 93.270 ;
        RECT 249.320 93.260 250.520 93.270 ;
        RECT 399.320 93.260 400.520 93.270 ;
        RECT 549.320 93.260 550.520 93.270 ;
        RECT 699.320 93.260 700.520 93.270 ;
        RECT 849.320 93.260 850.520 93.270 ;
        RECT 99.320 -3.510 100.520 -3.500 ;
        RECT 249.320 -3.510 250.520 -3.500 ;
        RECT 399.320 -3.510 400.520 -3.500 ;
        RECT 549.320 -3.510 550.520 -3.500 ;
        RECT 699.320 -3.510 700.520 -3.500 ;
        RECT 849.320 -3.510 850.520 -3.500 ;
        RECT -3.730 -3.810 1003.310 -3.510 ;
        RECT 99.320 -3.820 100.520 -3.810 ;
        RECT 249.320 -3.820 250.520 -3.810 ;
        RECT 399.320 -3.820 400.520 -3.810 ;
        RECT 549.320 -3.820 550.520 -3.810 ;
        RECT 699.320 -3.820 700.520 -3.810 ;
        RECT 849.320 -3.820 850.520 -3.810 ;
      LAYER via3 ;
        RECT 99.360 93.260 99.680 93.580 ;
        RECT 99.760 93.260 100.080 93.580 ;
        RECT 100.160 93.260 100.480 93.580 ;
        RECT 249.360 93.260 249.680 93.580 ;
        RECT 249.760 93.260 250.080 93.580 ;
        RECT 250.160 93.260 250.480 93.580 ;
        RECT 399.360 93.260 399.680 93.580 ;
        RECT 399.760 93.260 400.080 93.580 ;
        RECT 400.160 93.260 400.480 93.580 ;
        RECT 549.360 93.260 549.680 93.580 ;
        RECT 549.760 93.260 550.080 93.580 ;
        RECT 550.160 93.260 550.480 93.580 ;
        RECT 699.360 93.260 699.680 93.580 ;
        RECT 699.760 93.260 700.080 93.580 ;
        RECT 700.160 93.260 700.480 93.580 ;
        RECT 849.360 93.260 849.680 93.580 ;
        RECT 849.760 93.260 850.080 93.580 ;
        RECT 850.160 93.260 850.480 93.580 ;
        RECT 99.360 -3.820 99.680 -3.500 ;
        RECT 99.760 -3.820 100.080 -3.500 ;
        RECT 100.160 -3.820 100.480 -3.500 ;
        RECT 249.360 -3.820 249.680 -3.500 ;
        RECT 249.760 -3.820 250.080 -3.500 ;
        RECT 250.160 -3.820 250.480 -3.500 ;
        RECT 399.360 -3.820 399.680 -3.500 ;
        RECT 399.760 -3.820 400.080 -3.500 ;
        RECT 400.160 -3.820 400.480 -3.500 ;
        RECT 549.360 -3.820 549.680 -3.500 ;
        RECT 549.760 -3.820 550.080 -3.500 ;
        RECT 550.160 -3.820 550.480 -3.500 ;
        RECT 699.360 -3.820 699.680 -3.500 ;
        RECT 699.760 -3.820 700.080 -3.500 ;
        RECT 700.160 -3.820 700.480 -3.500 ;
        RECT 849.360 -3.820 849.680 -3.500 ;
        RECT 849.760 -3.820 850.080 -3.500 ;
        RECT 850.160 -3.820 850.480 -3.500 ;
      LAYER met4 ;
        RECT 99.320 89.700 100.520 93.585 ;
        RECT 249.320 89.700 250.520 93.585 ;
        RECT 399.320 89.700 400.520 93.585 ;
        RECT 549.320 89.700 550.520 93.585 ;
        RECT 699.320 89.700 700.520 93.585 ;
        RECT 849.320 89.700 850.520 93.585 ;
        RECT 99.320 -3.825 100.520 0.300 ;
        RECT 249.320 -3.825 250.520 0.300 ;
        RECT 399.320 -3.825 400.520 0.300 ;
        RECT 549.320 -3.825 550.520 0.300 ;
        RECT 699.320 -3.825 700.520 0.300 ;
        RECT 849.320 -3.825 850.520 0.300 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1003.010 -3.810 1003.310 93.570 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -3.730 -3.810 -3.430 93.570 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 28.720 94.270 29.920 94.280 ;
        RECT 178.720 94.270 179.920 94.280 ;
        RECT 328.720 94.270 329.920 94.280 ;
        RECT 478.720 94.270 479.920 94.280 ;
        RECT 628.720 94.270 629.920 94.280 ;
        RECT 778.720 94.270 779.920 94.280 ;
        RECT 928.720 94.270 929.920 94.280 ;
        RECT -4.430 93.970 1004.010 94.270 ;
        RECT 28.720 93.960 29.920 93.970 ;
        RECT 178.720 93.960 179.920 93.970 ;
        RECT 328.720 93.960 329.920 93.970 ;
        RECT 478.720 93.960 479.920 93.970 ;
        RECT 628.720 93.960 629.920 93.970 ;
        RECT 778.720 93.960 779.920 93.970 ;
        RECT 928.720 93.960 929.920 93.970 ;
        RECT 28.720 -4.210 29.920 -4.200 ;
        RECT 178.720 -4.210 179.920 -4.200 ;
        RECT 328.720 -4.210 329.920 -4.200 ;
        RECT 478.720 -4.210 479.920 -4.200 ;
        RECT 628.720 -4.210 629.920 -4.200 ;
        RECT 778.720 -4.210 779.920 -4.200 ;
        RECT 928.720 -4.210 929.920 -4.200 ;
        RECT -4.430 -4.510 1004.010 -4.210 ;
        RECT 28.720 -4.520 29.920 -4.510 ;
        RECT 178.720 -4.520 179.920 -4.510 ;
        RECT 328.720 -4.520 329.920 -4.510 ;
        RECT 478.720 -4.520 479.920 -4.510 ;
        RECT 628.720 -4.520 629.920 -4.510 ;
        RECT 778.720 -4.520 779.920 -4.510 ;
        RECT 928.720 -4.520 929.920 -4.510 ;
      LAYER via3 ;
        RECT 28.760 93.960 29.080 94.280 ;
        RECT 29.160 93.960 29.480 94.280 ;
        RECT 29.560 93.960 29.880 94.280 ;
        RECT 178.760 93.960 179.080 94.280 ;
        RECT 179.160 93.960 179.480 94.280 ;
        RECT 179.560 93.960 179.880 94.280 ;
        RECT 328.760 93.960 329.080 94.280 ;
        RECT 329.160 93.960 329.480 94.280 ;
        RECT 329.560 93.960 329.880 94.280 ;
        RECT 478.760 93.960 479.080 94.280 ;
        RECT 479.160 93.960 479.480 94.280 ;
        RECT 479.560 93.960 479.880 94.280 ;
        RECT 628.760 93.960 629.080 94.280 ;
        RECT 629.160 93.960 629.480 94.280 ;
        RECT 629.560 93.960 629.880 94.280 ;
        RECT 778.760 93.960 779.080 94.280 ;
        RECT 779.160 93.960 779.480 94.280 ;
        RECT 779.560 93.960 779.880 94.280 ;
        RECT 928.760 93.960 929.080 94.280 ;
        RECT 929.160 93.960 929.480 94.280 ;
        RECT 929.560 93.960 929.880 94.280 ;
        RECT 28.760 -4.520 29.080 -4.200 ;
        RECT 29.160 -4.520 29.480 -4.200 ;
        RECT 29.560 -4.520 29.880 -4.200 ;
        RECT 178.760 -4.520 179.080 -4.200 ;
        RECT 179.160 -4.520 179.480 -4.200 ;
        RECT 179.560 -4.520 179.880 -4.200 ;
        RECT 328.760 -4.520 329.080 -4.200 ;
        RECT 329.160 -4.520 329.480 -4.200 ;
        RECT 329.560 -4.520 329.880 -4.200 ;
        RECT 478.760 -4.520 479.080 -4.200 ;
        RECT 479.160 -4.520 479.480 -4.200 ;
        RECT 479.560 -4.520 479.880 -4.200 ;
        RECT 628.760 -4.520 629.080 -4.200 ;
        RECT 629.160 -4.520 629.480 -4.200 ;
        RECT 629.560 -4.520 629.880 -4.200 ;
        RECT 778.760 -4.520 779.080 -4.200 ;
        RECT 779.160 -4.520 779.480 -4.200 ;
        RECT 779.560 -4.520 779.880 -4.200 ;
        RECT 928.760 -4.520 929.080 -4.200 ;
        RECT 929.160 -4.520 929.480 -4.200 ;
        RECT 929.560 -4.520 929.880 -4.200 ;
      LAYER met4 ;
        RECT 28.720 89.700 29.920 94.970 ;
        RECT 178.720 89.700 179.920 94.970 ;
        RECT 328.720 89.700 329.920 94.970 ;
        RECT 478.720 89.700 479.920 94.970 ;
        RECT 628.720 89.700 629.920 94.970 ;
        RECT 778.720 89.700 779.920 94.970 ;
        RECT 928.720 89.700 929.920 94.970 ;
        RECT 28.720 -5.210 29.920 0.300 ;
        RECT 178.720 -5.210 179.920 0.300 ;
        RECT 328.720 -5.210 329.920 0.300 ;
        RECT 478.720 -5.210 479.920 0.300 ;
        RECT 628.720 -5.210 629.920 0.300 ;
        RECT 778.720 -5.210 779.920 0.300 ;
        RECT 928.720 -5.210 929.920 0.300 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1003.710 -4.510 1004.010 94.270 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -4.430 -4.510 -4.130 94.270 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 103.720 94.970 104.920 94.980 ;
        RECT 253.720 94.970 254.920 94.980 ;
        RECT 403.720 94.970 404.920 94.980 ;
        RECT 553.720 94.970 554.920 94.980 ;
        RECT 703.720 94.970 704.920 94.980 ;
        RECT 853.720 94.970 854.920 94.980 ;
        RECT -5.130 94.670 1004.710 94.970 ;
        RECT 103.720 94.660 104.920 94.670 ;
        RECT 253.720 94.660 254.920 94.670 ;
        RECT 403.720 94.660 404.920 94.670 ;
        RECT 553.720 94.660 554.920 94.670 ;
        RECT 703.720 94.660 704.920 94.670 ;
        RECT 853.720 94.660 854.920 94.670 ;
        RECT 103.720 -4.910 104.920 -4.900 ;
        RECT 253.720 -4.910 254.920 -4.900 ;
        RECT 403.720 -4.910 404.920 -4.900 ;
        RECT 553.720 -4.910 554.920 -4.900 ;
        RECT 703.720 -4.910 704.920 -4.900 ;
        RECT 853.720 -4.910 854.920 -4.900 ;
        RECT -5.130 -5.210 1004.710 -4.910 ;
        RECT 103.720 -5.220 104.920 -5.210 ;
        RECT 253.720 -5.220 254.920 -5.210 ;
        RECT 403.720 -5.220 404.920 -5.210 ;
        RECT 553.720 -5.220 554.920 -5.210 ;
        RECT 703.720 -5.220 704.920 -5.210 ;
        RECT 853.720 -5.220 854.920 -5.210 ;
      LAYER via3 ;
        RECT 103.760 94.660 104.080 94.980 ;
        RECT 104.160 94.660 104.480 94.980 ;
        RECT 104.560 94.660 104.880 94.980 ;
        RECT 253.760 94.660 254.080 94.980 ;
        RECT 254.160 94.660 254.480 94.980 ;
        RECT 254.560 94.660 254.880 94.980 ;
        RECT 403.760 94.660 404.080 94.980 ;
        RECT 404.160 94.660 404.480 94.980 ;
        RECT 404.560 94.660 404.880 94.980 ;
        RECT 553.760 94.660 554.080 94.980 ;
        RECT 554.160 94.660 554.480 94.980 ;
        RECT 554.560 94.660 554.880 94.980 ;
        RECT 703.760 94.660 704.080 94.980 ;
        RECT 704.160 94.660 704.480 94.980 ;
        RECT 704.560 94.660 704.880 94.980 ;
        RECT 853.760 94.660 854.080 94.980 ;
        RECT 854.160 94.660 854.480 94.980 ;
        RECT 854.560 94.660 854.880 94.980 ;
        RECT 103.760 -5.220 104.080 -4.900 ;
        RECT 104.160 -5.220 104.480 -4.900 ;
        RECT 104.560 -5.220 104.880 -4.900 ;
        RECT 253.760 -5.220 254.080 -4.900 ;
        RECT 254.160 -5.220 254.480 -4.900 ;
        RECT 254.560 -5.220 254.880 -4.900 ;
        RECT 403.760 -5.220 404.080 -4.900 ;
        RECT 404.160 -5.220 404.480 -4.900 ;
        RECT 404.560 -5.220 404.880 -4.900 ;
        RECT 553.760 -5.220 554.080 -4.900 ;
        RECT 554.160 -5.220 554.480 -4.900 ;
        RECT 554.560 -5.220 554.880 -4.900 ;
        RECT 703.760 -5.220 704.080 -4.900 ;
        RECT 704.160 -5.220 704.480 -4.900 ;
        RECT 704.560 -5.220 704.880 -4.900 ;
        RECT 853.760 -5.220 854.080 -4.900 ;
        RECT 854.160 -5.220 854.480 -4.900 ;
        RECT 854.560 -5.220 854.880 -4.900 ;
      LAYER met4 ;
        RECT 103.720 89.700 104.920 94.985 ;
        RECT 253.720 89.700 254.920 94.985 ;
        RECT 403.720 89.700 404.920 94.985 ;
        RECT 553.720 89.700 554.920 94.985 ;
        RECT 703.720 89.700 704.920 94.985 ;
        RECT 853.720 89.700 854.920 94.985 ;
        RECT 103.720 -5.225 104.920 0.300 ;
        RECT 253.720 -5.225 254.920 0.300 ;
        RECT 403.720 -5.225 404.920 0.300 ;
        RECT 553.720 -5.225 554.920 0.300 ;
        RECT 703.720 -5.225 704.920 0.300 ;
        RECT 853.720 -5.225 854.920 0.300 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1004.410 -5.210 1004.710 94.970 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -5.130 -5.210 -4.830 94.970 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 33.120 95.670 34.320 95.680 ;
        RECT 183.120 95.670 184.320 95.680 ;
        RECT 333.120 95.670 334.320 95.680 ;
        RECT 483.120 95.670 484.320 95.680 ;
        RECT 633.120 95.670 634.320 95.680 ;
        RECT 783.120 95.670 784.320 95.680 ;
        RECT 933.120 95.670 934.320 95.680 ;
        RECT -5.830 95.370 1005.410 95.670 ;
        RECT 33.120 95.360 34.320 95.370 ;
        RECT 183.120 95.360 184.320 95.370 ;
        RECT 333.120 95.360 334.320 95.370 ;
        RECT 483.120 95.360 484.320 95.370 ;
        RECT 633.120 95.360 634.320 95.370 ;
        RECT 783.120 95.360 784.320 95.370 ;
        RECT 933.120 95.360 934.320 95.370 ;
        RECT 33.120 -5.610 34.320 -5.600 ;
        RECT 183.120 -5.610 184.320 -5.600 ;
        RECT 333.120 -5.610 334.320 -5.600 ;
        RECT 483.120 -5.610 484.320 -5.600 ;
        RECT 633.120 -5.610 634.320 -5.600 ;
        RECT 783.120 -5.610 784.320 -5.600 ;
        RECT 933.120 -5.610 934.320 -5.600 ;
        RECT -5.830 -5.910 1005.410 -5.610 ;
        RECT 33.120 -5.920 34.320 -5.910 ;
        RECT 183.120 -5.920 184.320 -5.910 ;
        RECT 333.120 -5.920 334.320 -5.910 ;
        RECT 483.120 -5.920 484.320 -5.910 ;
        RECT 633.120 -5.920 634.320 -5.910 ;
        RECT 783.120 -5.920 784.320 -5.910 ;
        RECT 933.120 -5.920 934.320 -5.910 ;
      LAYER via3 ;
        RECT 33.160 95.360 33.480 95.680 ;
        RECT 33.560 95.360 33.880 95.680 ;
        RECT 33.960 95.360 34.280 95.680 ;
        RECT 183.160 95.360 183.480 95.680 ;
        RECT 183.560 95.360 183.880 95.680 ;
        RECT 183.960 95.360 184.280 95.680 ;
        RECT 333.160 95.360 333.480 95.680 ;
        RECT 333.560 95.360 333.880 95.680 ;
        RECT 333.960 95.360 334.280 95.680 ;
        RECT 483.160 95.360 483.480 95.680 ;
        RECT 483.560 95.360 483.880 95.680 ;
        RECT 483.960 95.360 484.280 95.680 ;
        RECT 633.160 95.360 633.480 95.680 ;
        RECT 633.560 95.360 633.880 95.680 ;
        RECT 633.960 95.360 634.280 95.680 ;
        RECT 783.160 95.360 783.480 95.680 ;
        RECT 783.560 95.360 783.880 95.680 ;
        RECT 783.960 95.360 784.280 95.680 ;
        RECT 933.160 95.360 933.480 95.680 ;
        RECT 933.560 95.360 933.880 95.680 ;
        RECT 933.960 95.360 934.280 95.680 ;
        RECT 33.160 -5.920 33.480 -5.600 ;
        RECT 33.560 -5.920 33.880 -5.600 ;
        RECT 33.960 -5.920 34.280 -5.600 ;
        RECT 183.160 -5.920 183.480 -5.600 ;
        RECT 183.560 -5.920 183.880 -5.600 ;
        RECT 183.960 -5.920 184.280 -5.600 ;
        RECT 333.160 -5.920 333.480 -5.600 ;
        RECT 333.560 -5.920 333.880 -5.600 ;
        RECT 333.960 -5.920 334.280 -5.600 ;
        RECT 483.160 -5.920 483.480 -5.600 ;
        RECT 483.560 -5.920 483.880 -5.600 ;
        RECT 483.960 -5.920 484.280 -5.600 ;
        RECT 633.160 -5.920 633.480 -5.600 ;
        RECT 633.560 -5.920 633.880 -5.600 ;
        RECT 633.960 -5.920 634.280 -5.600 ;
        RECT 783.160 -5.920 783.480 -5.600 ;
        RECT 783.560 -5.920 783.880 -5.600 ;
        RECT 783.960 -5.920 784.280 -5.600 ;
        RECT 933.160 -5.920 933.480 -5.600 ;
        RECT 933.560 -5.920 933.880 -5.600 ;
        RECT 933.960 -5.920 934.280 -5.600 ;
      LAYER met4 ;
        RECT 33.120 89.700 34.320 96.370 ;
        RECT 183.120 89.700 184.320 96.370 ;
        RECT 333.120 89.700 334.320 96.370 ;
        RECT 483.120 89.700 484.320 96.370 ;
        RECT 633.120 89.700 634.320 96.370 ;
        RECT 783.120 89.700 784.320 96.370 ;
        RECT 933.120 89.700 934.320 96.370 ;
        RECT 33.120 -6.610 34.320 0.300 ;
        RECT 183.120 -6.610 184.320 0.300 ;
        RECT 333.120 -6.610 334.320 0.300 ;
        RECT 483.120 -6.610 484.320 0.300 ;
        RECT 633.120 -6.610 634.320 0.300 ;
        RECT 783.120 -6.610 784.320 0.300 ;
        RECT 933.120 -6.610 934.320 0.300 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1005.110 -5.910 1005.410 95.670 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -5.830 -5.910 -5.530 95.670 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 108.120 96.370 109.320 96.380 ;
        RECT 258.120 96.370 259.320 96.380 ;
        RECT 408.120 96.370 409.320 96.380 ;
        RECT 558.120 96.370 559.320 96.380 ;
        RECT 708.120 96.370 709.320 96.380 ;
        RECT 858.120 96.370 859.320 96.380 ;
        RECT -6.530 96.070 1006.110 96.370 ;
        RECT 108.120 96.060 109.320 96.070 ;
        RECT 258.120 96.060 259.320 96.070 ;
        RECT 408.120 96.060 409.320 96.070 ;
        RECT 558.120 96.060 559.320 96.070 ;
        RECT 708.120 96.060 709.320 96.070 ;
        RECT 858.120 96.060 859.320 96.070 ;
        RECT 108.120 -6.310 109.320 -6.300 ;
        RECT 258.120 -6.310 259.320 -6.300 ;
        RECT 408.120 -6.310 409.320 -6.300 ;
        RECT 558.120 -6.310 559.320 -6.300 ;
        RECT 708.120 -6.310 709.320 -6.300 ;
        RECT 858.120 -6.310 859.320 -6.300 ;
        RECT -6.530 -6.610 1006.110 -6.310 ;
        RECT 108.120 -6.620 109.320 -6.610 ;
        RECT 258.120 -6.620 259.320 -6.610 ;
        RECT 408.120 -6.620 409.320 -6.610 ;
        RECT 558.120 -6.620 559.320 -6.610 ;
        RECT 708.120 -6.620 709.320 -6.610 ;
        RECT 858.120 -6.620 859.320 -6.610 ;
      LAYER via3 ;
        RECT 108.160 96.060 108.480 96.380 ;
        RECT 108.560 96.060 108.880 96.380 ;
        RECT 108.960 96.060 109.280 96.380 ;
        RECT 258.160 96.060 258.480 96.380 ;
        RECT 258.560 96.060 258.880 96.380 ;
        RECT 258.960 96.060 259.280 96.380 ;
        RECT 408.160 96.060 408.480 96.380 ;
        RECT 408.560 96.060 408.880 96.380 ;
        RECT 408.960 96.060 409.280 96.380 ;
        RECT 558.160 96.060 558.480 96.380 ;
        RECT 558.560 96.060 558.880 96.380 ;
        RECT 558.960 96.060 559.280 96.380 ;
        RECT 708.160 96.060 708.480 96.380 ;
        RECT 708.560 96.060 708.880 96.380 ;
        RECT 708.960 96.060 709.280 96.380 ;
        RECT 858.160 96.060 858.480 96.380 ;
        RECT 858.560 96.060 858.880 96.380 ;
        RECT 858.960 96.060 859.280 96.380 ;
        RECT 108.160 -6.620 108.480 -6.300 ;
        RECT 108.560 -6.620 108.880 -6.300 ;
        RECT 108.960 -6.620 109.280 -6.300 ;
        RECT 258.160 -6.620 258.480 -6.300 ;
        RECT 258.560 -6.620 258.880 -6.300 ;
        RECT 258.960 -6.620 259.280 -6.300 ;
        RECT 408.160 -6.620 408.480 -6.300 ;
        RECT 408.560 -6.620 408.880 -6.300 ;
        RECT 408.960 -6.620 409.280 -6.300 ;
        RECT 558.160 -6.620 558.480 -6.300 ;
        RECT 558.560 -6.620 558.880 -6.300 ;
        RECT 558.960 -6.620 559.280 -6.300 ;
        RECT 708.160 -6.620 708.480 -6.300 ;
        RECT 708.560 -6.620 708.880 -6.300 ;
        RECT 708.960 -6.620 709.280 -6.300 ;
        RECT 858.160 -6.620 858.480 -6.300 ;
        RECT 858.560 -6.620 858.880 -6.300 ;
        RECT 858.960 -6.620 859.280 -6.300 ;
      LAYER met4 ;
        RECT 108.120 89.700 109.320 96.385 ;
        RECT 258.120 89.700 259.320 96.385 ;
        RECT 408.120 89.700 409.320 96.385 ;
        RECT 558.120 89.700 559.320 96.385 ;
        RECT 708.120 89.700 709.320 96.385 ;
        RECT 858.120 89.700 859.320 96.385 ;
        RECT 108.120 -6.625 109.320 0.300 ;
        RECT 258.120 -6.625 259.320 0.300 ;
        RECT 408.120 -6.625 409.320 0.300 ;
        RECT 558.120 -6.625 559.320 0.300 ;
        RECT 708.120 -6.625 709.320 0.300 ;
        RECT 858.120 -6.625 859.320 0.300 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1005.810 -6.610 1006.110 96.370 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -6.530 -6.610 -6.230 96.370 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 37.520 97.070 38.720 97.080 ;
        RECT 187.520 97.070 188.720 97.080 ;
        RECT 337.520 97.070 338.720 97.080 ;
        RECT 487.520 97.070 488.720 97.080 ;
        RECT 637.520 97.070 638.720 97.080 ;
        RECT 787.520 97.070 788.720 97.080 ;
        RECT 937.520 97.070 938.720 97.080 ;
        RECT -7.230 96.770 1006.810 97.070 ;
        RECT 37.520 96.760 38.720 96.770 ;
        RECT 187.520 96.760 188.720 96.770 ;
        RECT 337.520 96.760 338.720 96.770 ;
        RECT 487.520 96.760 488.720 96.770 ;
        RECT 637.520 96.760 638.720 96.770 ;
        RECT 787.520 96.760 788.720 96.770 ;
        RECT 937.520 96.760 938.720 96.770 ;
        RECT 37.520 -7.010 38.720 -7.000 ;
        RECT 187.520 -7.010 188.720 -7.000 ;
        RECT 337.520 -7.010 338.720 -7.000 ;
        RECT 487.520 -7.010 488.720 -7.000 ;
        RECT 637.520 -7.010 638.720 -7.000 ;
        RECT 787.520 -7.010 788.720 -7.000 ;
        RECT 937.520 -7.010 938.720 -7.000 ;
        RECT -7.230 -7.310 1006.810 -7.010 ;
        RECT 37.520 -7.320 38.720 -7.310 ;
        RECT 187.520 -7.320 188.720 -7.310 ;
        RECT 337.520 -7.320 338.720 -7.310 ;
        RECT 487.520 -7.320 488.720 -7.310 ;
        RECT 637.520 -7.320 638.720 -7.310 ;
        RECT 787.520 -7.320 788.720 -7.310 ;
        RECT 937.520 -7.320 938.720 -7.310 ;
      LAYER via3 ;
        RECT 37.560 96.760 37.880 97.080 ;
        RECT 37.960 96.760 38.280 97.080 ;
        RECT 38.360 96.760 38.680 97.080 ;
        RECT 187.560 96.760 187.880 97.080 ;
        RECT 187.960 96.760 188.280 97.080 ;
        RECT 188.360 96.760 188.680 97.080 ;
        RECT 337.560 96.760 337.880 97.080 ;
        RECT 337.960 96.760 338.280 97.080 ;
        RECT 338.360 96.760 338.680 97.080 ;
        RECT 487.560 96.760 487.880 97.080 ;
        RECT 487.960 96.760 488.280 97.080 ;
        RECT 488.360 96.760 488.680 97.080 ;
        RECT 637.560 96.760 637.880 97.080 ;
        RECT 637.960 96.760 638.280 97.080 ;
        RECT 638.360 96.760 638.680 97.080 ;
        RECT 787.560 96.760 787.880 97.080 ;
        RECT 787.960 96.760 788.280 97.080 ;
        RECT 788.360 96.760 788.680 97.080 ;
        RECT 937.560 96.760 937.880 97.080 ;
        RECT 937.960 96.760 938.280 97.080 ;
        RECT 938.360 96.760 938.680 97.080 ;
        RECT 37.560 -7.320 37.880 -7.000 ;
        RECT 37.960 -7.320 38.280 -7.000 ;
        RECT 38.360 -7.320 38.680 -7.000 ;
        RECT 187.560 -7.320 187.880 -7.000 ;
        RECT 187.960 -7.320 188.280 -7.000 ;
        RECT 188.360 -7.320 188.680 -7.000 ;
        RECT 337.560 -7.320 337.880 -7.000 ;
        RECT 337.960 -7.320 338.280 -7.000 ;
        RECT 338.360 -7.320 338.680 -7.000 ;
        RECT 487.560 -7.320 487.880 -7.000 ;
        RECT 487.960 -7.320 488.280 -7.000 ;
        RECT 488.360 -7.320 488.680 -7.000 ;
        RECT 637.560 -7.320 637.880 -7.000 ;
        RECT 637.960 -7.320 638.280 -7.000 ;
        RECT 638.360 -7.320 638.680 -7.000 ;
        RECT 787.560 -7.320 787.880 -7.000 ;
        RECT 787.960 -7.320 788.280 -7.000 ;
        RECT 788.360 -7.320 788.680 -7.000 ;
        RECT 937.560 -7.320 937.880 -7.000 ;
        RECT 937.960 -7.320 938.280 -7.000 ;
        RECT 938.360 -7.320 938.680 -7.000 ;
      LAYER met4 ;
        RECT 37.520 89.700 38.720 97.770 ;
        RECT 187.520 89.700 188.720 97.770 ;
        RECT 337.520 89.700 338.720 97.770 ;
        RECT 487.520 89.700 488.720 97.770 ;
        RECT 637.520 89.700 638.720 97.770 ;
        RECT 787.520 89.700 788.720 97.770 ;
        RECT 937.520 89.700 938.720 97.770 ;
        RECT 37.520 -8.010 38.720 0.300 ;
        RECT 187.520 -8.010 188.720 0.300 ;
        RECT 337.520 -8.010 338.720 0.300 ;
        RECT 487.520 -8.010 488.720 0.300 ;
        RECT 637.520 -8.010 638.720 0.300 ;
        RECT 787.520 -8.010 788.720 0.300 ;
        RECT 937.520 -8.010 938.720 0.300 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1006.510 -7.310 1006.810 97.070 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -7.230 -7.310 -6.930 97.070 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 112.520 97.770 113.720 97.780 ;
        RECT 262.520 97.770 263.720 97.780 ;
        RECT 412.520 97.770 413.720 97.780 ;
        RECT 562.520 97.770 563.720 97.780 ;
        RECT 712.520 97.770 713.720 97.780 ;
        RECT 862.520 97.770 863.720 97.780 ;
        RECT -7.930 97.470 1007.510 97.770 ;
        RECT 112.520 97.460 113.720 97.470 ;
        RECT 262.520 97.460 263.720 97.470 ;
        RECT 412.520 97.460 413.720 97.470 ;
        RECT 562.520 97.460 563.720 97.470 ;
        RECT 712.520 97.460 713.720 97.470 ;
        RECT 862.520 97.460 863.720 97.470 ;
        RECT 112.520 -7.710 113.720 -7.700 ;
        RECT 262.520 -7.710 263.720 -7.700 ;
        RECT 412.520 -7.710 413.720 -7.700 ;
        RECT 562.520 -7.710 563.720 -7.700 ;
        RECT 712.520 -7.710 713.720 -7.700 ;
        RECT 862.520 -7.710 863.720 -7.700 ;
        RECT -7.930 -8.010 1007.510 -7.710 ;
        RECT 112.520 -8.020 113.720 -8.010 ;
        RECT 262.520 -8.020 263.720 -8.010 ;
        RECT 412.520 -8.020 413.720 -8.010 ;
        RECT 562.520 -8.020 563.720 -8.010 ;
        RECT 712.520 -8.020 713.720 -8.010 ;
        RECT 862.520 -8.020 863.720 -8.010 ;
      LAYER via3 ;
        RECT 112.560 97.460 112.880 97.780 ;
        RECT 112.960 97.460 113.280 97.780 ;
        RECT 113.360 97.460 113.680 97.780 ;
        RECT 262.560 97.460 262.880 97.780 ;
        RECT 262.960 97.460 263.280 97.780 ;
        RECT 263.360 97.460 263.680 97.780 ;
        RECT 412.560 97.460 412.880 97.780 ;
        RECT 412.960 97.460 413.280 97.780 ;
        RECT 413.360 97.460 413.680 97.780 ;
        RECT 562.560 97.460 562.880 97.780 ;
        RECT 562.960 97.460 563.280 97.780 ;
        RECT 563.360 97.460 563.680 97.780 ;
        RECT 712.560 97.460 712.880 97.780 ;
        RECT 712.960 97.460 713.280 97.780 ;
        RECT 713.360 97.460 713.680 97.780 ;
        RECT 862.560 97.460 862.880 97.780 ;
        RECT 862.960 97.460 863.280 97.780 ;
        RECT 863.360 97.460 863.680 97.780 ;
        RECT 112.560 -8.020 112.880 -7.700 ;
        RECT 112.960 -8.020 113.280 -7.700 ;
        RECT 113.360 -8.020 113.680 -7.700 ;
        RECT 262.560 -8.020 262.880 -7.700 ;
        RECT 262.960 -8.020 263.280 -7.700 ;
        RECT 263.360 -8.020 263.680 -7.700 ;
        RECT 412.560 -8.020 412.880 -7.700 ;
        RECT 412.960 -8.020 413.280 -7.700 ;
        RECT 413.360 -8.020 413.680 -7.700 ;
        RECT 562.560 -8.020 562.880 -7.700 ;
        RECT 562.960 -8.020 563.280 -7.700 ;
        RECT 563.360 -8.020 563.680 -7.700 ;
        RECT 712.560 -8.020 712.880 -7.700 ;
        RECT 712.960 -8.020 713.280 -7.700 ;
        RECT 713.360 -8.020 713.680 -7.700 ;
        RECT 862.560 -8.020 862.880 -7.700 ;
        RECT 862.960 -8.020 863.280 -7.700 ;
        RECT 863.360 -8.020 863.680 -7.700 ;
      LAYER met4 ;
        RECT 112.520 89.700 113.720 97.785 ;
        RECT 262.520 89.700 263.720 97.785 ;
        RECT 412.520 89.700 413.720 97.785 ;
        RECT 562.520 89.700 563.720 97.785 ;
        RECT 712.520 89.700 713.720 97.785 ;
        RECT 862.520 89.700 863.720 97.785 ;
        RECT 112.520 -8.025 113.720 0.300 ;
        RECT 262.520 -8.025 263.720 0.300 ;
        RECT 412.520 -8.025 413.720 0.300 ;
        RECT 562.520 -8.025 563.720 0.300 ;
        RECT 712.520 -8.025 713.720 0.300 ;
        RECT 862.520 -8.025 863.720 0.300 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1007.210 -8.010 1007.510 97.770 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -7.930 -8.010 -7.630 97.770 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 326.285 89.845 328.295 90.015 ;
        RECT 328.125 89.700 328.295 89.845 ;
        RECT 453.245 89.845 473.195 90.015 ;
        RECT 453.245 89.700 453.415 89.845 ;
        RECT 473.025 89.700 473.195 89.845 ;
        RECT 5.520 5.355 994.060 89.700 ;
      LAYER met1 ;
        RECT 296.310 90.000 296.630 90.060 ;
        RECT 326.225 90.000 326.515 90.045 ;
        RECT 296.310 89.860 326.515 90.000 ;
        RECT 296.310 89.800 296.630 89.860 ;
        RECT 326.225 89.815 326.515 89.860 ;
        RECT 326.670 90.000 326.990 90.060 ;
        RECT 600.830 90.000 601.150 90.060 ;
        RECT 326.670 89.860 601.150 90.000 ;
        RECT 326.670 89.800 326.990 89.860 ;
        RECT 600.830 89.800 601.150 89.860 ;
        RECT 132.550 89.700 132.870 89.720 ;
        RECT 472.505 89.700 472.795 89.705 ;
        RECT 472.965 89.700 473.255 89.705 ;
        RECT 475.725 89.700 476.015 89.705 ;
        RECT 476.170 89.700 476.490 89.720 ;
        RECT 754.010 89.700 754.330 89.720 ;
        RECT 0.990 3.100 999.050 89.700 ;
      LAYER via ;
        RECT 296.340 89.800 296.600 90.060 ;
        RECT 326.700 89.800 326.960 90.060 ;
        RECT 600.860 89.800 601.120 90.060 ;
        RECT 132.580 89.460 132.840 89.720 ;
        RECT 476.200 89.460 476.460 89.720 ;
        RECT 754.040 89.460 754.300 89.720 ;
      LAYER met2 ;
        RECT 296.340 89.770 296.600 90.090 ;
        RECT 326.700 89.770 326.960 90.090 ;
        RECT 600.860 89.770 601.120 90.090 ;
        RECT 132.580 89.700 132.840 89.750 ;
        RECT 296.400 89.700 296.540 89.770 ;
        RECT 326.760 89.700 326.900 89.770 ;
        RECT 476.200 89.700 476.460 89.750 ;
        RECT 600.920 89.700 601.060 89.770 ;
        RECT 754.040 89.700 754.300 89.750 ;
        RECT 1.010 0.300 999.030 89.700 ;
      LAYER met3 ;
        RECT 0.300 4.255 973.295 89.585 ;
      LAYER met4 ;
        RECT 19.920 0.300 938.720 89.700 ;
  END
END mgmt_protect
END LIBRARY

