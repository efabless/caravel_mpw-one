* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param
+ sky130_fd_pr__pfet_01v8_mvt__noia_mult = 100.0
.param sky130_fd_pr__pfet_01v8_mvt__toxe_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_mvt__vth0_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_mvt__voff_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_mvt__nfactor_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__pfet_01v8_mvt__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_mvt__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_mvt__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_mvt__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__pfet_01v8_mvt d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1 
msky130_fd_pr__pfet_01v8_mvt d g s b sky130_fd_pr__pfet_01v8_mvt__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} 
.model sky130_fd_pr__pfet_01v8_mvt__model.0 pmos
* Model Flag Parameters
+ lmin = 1.45e-007 lmax = 1.55e-007 wmin = 1.675e-006 wmax = 1.685e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_mvt__toxe_mult}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1*sky130_fd_pr__pfet_01v8_mvt__rshp_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {7.304e-009+sky130_fd_pr__pfet_01v8_mvt__wint_diff}
+ lint = {-1.399e-008+sky130_fd_pr__pfet_01v8_mvt__lint_diff}
+ vth0 = {-0.7375+sky130_fd_pr__pfet_01v8_mvt__vth0_diff_0}
+ k1 = 0.2078
+ k2 = {0.09904+sky130_fd_pr__pfet_01v8_mvt__k2_diff_0}
+ k3 = -15.85
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.496
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.977
+ dvt1w = 1147000.0
+ dvt2w = -0.00896
+ dsub = 0.26
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.02472
+ cdscb = 0.003175
+ cdscd = 0.0
+ cit = 0.0001462
+ voff = {-0.4483+sky130_fd_pr__pfet_01v8_mvt__voff_diff_0}
+ nfactor = {4.228+sky130_fd_pr__pfet_01v8_mvt__nfactor_diff_0}
+ eta0 = {0.5735+sky130_fd_pr__pfet_01v8_mvt__eta0_diff_0}
+ etab = -0.03063
+ u0 = {0.002233+sky130_fd_pr__pfet_01v8_mvt__u0_diff_0}
+ ua = {-2.832e-009+sky130_fd_pr__pfet_01v8_mvt__ua_diff_0}
+ ub = {2.789e-018+sky130_fd_pr__pfet_01v8_mvt__ub_diff_0}
+ uc = -1.076e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {47470+sky130_fd_pr__pfet_01v8_mvt__vsat_diff_0}
+ a0 = {1.047+sky130_fd_pr__pfet_01v8_mvt__a0_diff_0}
+ ags = {0.5789+sky130_fd_pr__pfet_01v8_mvt__ags_diff_0}
+ a1 = 0.0
+ a2 = 0.9995
+ b0 = {0+sky130_fd_pr__pfet_01v8_mvt__b0_diff_0}
+ b1 = {0+sky130_fd_pr__pfet_01v8_mvt__b1_diff_0}
+ keta = {0.09663+sky130_fd_pr__pfet_01v8_mvt__keta_diff_0}
+ dwg = -5.722e-9
+ dwb = -1.786e-8
+ pclm = {0.2853+sky130_fd_pr__pfet_01v8_mvt__pclm_diff_0}
+ pdiblc1 = 0.0195
+ pdiblc2 = 0.00043
+ pdiblcb = -2.441e-5
+ drout = 1.0
+ pscbe1 = 7.69e+8
+ pscbe2 = 8.801e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_mvt__pdits_diff_0}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_mvt__pditsd_diff_0}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {547.9+sky130_fd_pr__pfet_01v8_mvt__rdsw_diff_0}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.3235
+ prwg = 0.1376
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.261
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {2.214e-010+sky130_fd_pr__pfet_01v8_mvt__agidl_diff_0}
+ bgidl = {1e+009+sky130_fd_pr__pfet_01v8_mvt__bgidl_diff_0}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_mvt__cgidl_diff_0}
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {1.536e-008+sky130_fd_pr__pfet_01v8_mvt__dlc_diff}
+ dwc = {0+sky130_fd_pr__pfet_01v8_mvt__dwc_diff}
+ xpart = 0.0
+ cgso = {7.17e-011*sky130_fd_pr__pfet_01v8_mvt__overlap_mult}
+ cgdo = {8.17e-011*sky130_fd_pr__pfet_01v8_mvt__overlap_mult}
+ cgbo = 0.0
+ cgdl = {5.5e-013*sky130_fd_pr__pfet_01v8_mvt__overlap_mult}
+ cgsl = {5.5e-013*sky130_fd_pr__pfet_01v8_mvt__overlap_mult}
+ clc = 0.0
+ cle = 1.0
+ cf = 6.0e-12
+ ckappas = 0.6
+ vfbcv = -0.1447
+ acde = 0.3136
+ moin = 25.0
+ noff = 3.9
+ voffcv = 0.1462
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 1.0
+ noia = {2.7e+042*sky130_fd_pr__pfet_01v8_mvt__noia_mult}
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ ntnoi = 1.0
+ lintnoi = -2.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 2.5e+7
+ tnoib = 0.0
+ rnoia = 0.69
+ rnoib = 0.34
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.148e-5
+ jsws = 8.04e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.69
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = {0.000738*sky130_fd_pr__pfet_01v8_mvt__ajunction_mult}
+ mjs = 0.3463
+ pbsws = 0.7418
+ cjsws = {9.889e-011*sky130_fd_pr__pfet_01v8_mvt__pjunction_mult}
+ mjsws = 0.2978
+ pbswgs = 1.434
+ cjswgs = {2.232e-010*sky130_fd_pr__pfet_01v8_mvt__pjunction_mult}
+ mjswgs = 0.9274
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.5434+sky130_fd_pr__pfet_01v8_mvt__kt1_diff_0}
+ kt2 = -0.1167
+ at = 21110.0
+ ute = -0.2531
+ ua1 = -8.749e-10
+ ub1 = 2.358e-18
+ uc1 = 7.088e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_mvt__tvoff_diff_0}
+ njs = 1.363
+ tpb = 0.002039
+ tcj = 0.001241
+ tpbsw = 0.001246
+ tcjsw = 0.0003736
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 5.2
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 3.29e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.5
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_mvt__model.1 pmos
* Model Flag Parameters
+ lmin = 1.45e-007 lmax = 1.55e-007 wmin = 8.35e-007 wmax = 8.45e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_mvt__toxe_mult}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1*sky130_fd_pr__pfet_01v8_mvt__rshp_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {7.304e-009+sky130_fd_pr__pfet_01v8_mvt__wint_diff}
+ lint = {-1.399e-008+sky130_fd_pr__pfet_01v8_mvt__lint_diff}
+ vth0 = {-0.7375+sky130_fd_pr__pfet_01v8_mvt__vth0_diff_1}
+ k1 = 0.2078
+ k2 = {0.107+sky130_fd_pr__pfet_01v8_mvt__k2_diff_1}
+ k3 = -15.85
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.496
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.977
+ dvt1w = 1147000.0
+ dvt2w = -0.00896
+ dsub = 0.26
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.02522
+ cdscb = 0.004958
+ cdscd = 0.0
+ cit = 0.0001462
+ voff = {-0.4483+sky130_fd_pr__pfet_01v8_mvt__voff_diff_1}
+ nfactor = {4.228+sky130_fd_pr__pfet_01v8_mvt__nfactor_diff_1}
+ eta0 = {0.6128+sky130_fd_pr__pfet_01v8_mvt__eta0_diff_1}
+ etab = -0.04874
+ u0 = {0.002175+sky130_fd_pr__pfet_01v8_mvt__u0_diff_1}
+ ua = {-2.801e-009+sky130_fd_pr__pfet_01v8_mvt__ua_diff_1}
+ ub = {2.717e-018+sky130_fd_pr__pfet_01v8_mvt__ub_diff_1}
+ uc = -2.128e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {45410+sky130_fd_pr__pfet_01v8_mvt__vsat_diff_1}
+ a0 = {1.047+sky130_fd_pr__pfet_01v8_mvt__a0_diff_1}
+ ags = {0.5789+sky130_fd_pr__pfet_01v8_mvt__ags_diff_1}
+ a1 = 0.0
+ a2 = 0.9995
+ b0 = {0+sky130_fd_pr__pfet_01v8_mvt__b0_diff_1}
+ b1 = {0+sky130_fd_pr__pfet_01v8_mvt__b1_diff_1}
+ keta = {0.09663+sky130_fd_pr__pfet_01v8_mvt__keta_diff_1}
+ dwg = -5.722e-9
+ dwb = -1.786e-8
+ pclm = {0.2853+sky130_fd_pr__pfet_01v8_mvt__pclm_diff_1}
+ pdiblc1 = 0.0195
+ pdiblc2 = 0.00043
+ pdiblcb = -2.441e-5
+ drout = 1.0
+ pscbe1 = 7.69e+8
+ pscbe2 = 8.801e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_mvt__pdits_diff_1}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_mvt__pditsd_diff_1}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {547.9+sky130_fd_pr__pfet_01v8_mvt__rdsw_diff_1}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.3235
+ prwg = 0.1376
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.261
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {2.214e-010+sky130_fd_pr__pfet_01v8_mvt__agidl_diff_1}
+ bgidl = {1e+009+sky130_fd_pr__pfet_01v8_mvt__bgidl_diff_1}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_mvt__cgidl_diff_1}
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {3.536e-008+sky130_fd_pr__pfet_01v8_mvt__dlc_diff}
+ dwc = {0+sky130_fd_pr__pfet_01v8_mvt__dwc_diff}
+ xpart = 0.0
+ cgso = {1e-013*sky130_fd_pr__pfet_01v8_mvt__overlap_mult}
+ cgdo = {1.857e-010*sky130_fd_pr__pfet_01v8_mvt__overlap_mult}
+ cgbo = 0.0
+ cgdl = {9.55e-012*sky130_fd_pr__pfet_01v8_mvt__overlap_mult}
+ cgsl = {9.55e-012*sky130_fd_pr__pfet_01v8_mvt__overlap_mult}
+ clc = 0.0
+ cle = 1.0
+ cf = 1.2e-13
+ ckappas = 0.6
+ vfbcv = -0.1447
+ acde = 0.3136
+ moin = 25.0
+ noff = 3.9
+ voffcv = 0.1462
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 1.0
+ noia = {2.7e+042*sky130_fd_pr__pfet_01v8_mvt__noia_mult}
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ ntnoi = 1.0
+ lintnoi = -2.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 2.5e+7
+ tnoib = 0.0
+ rnoia = 0.69
+ rnoib = 0.34
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.148e-5
+ jsws = 8.04e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.69
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = {0.000738*sky130_fd_pr__pfet_01v8_mvt__ajunction_mult}
+ mjs = 0.3463
+ pbsws = 0.7418
+ cjsws = {9.889e-011*sky130_fd_pr__pfet_01v8_mvt__pjunction_mult}
+ mjsws = 0.2978
+ pbswgs = 1.434
+ cjswgs = {2.232e-010*sky130_fd_pr__pfet_01v8_mvt__pjunction_mult}
+ mjswgs = 0.9274
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.7955+sky130_fd_pr__pfet_01v8_mvt__kt1_diff_1}
+ kt2 = -0.1319
+ at = 21110.0
+ ute = -0.1462
+ ua1 = -1.988e-10
+ ub1 = 1.323e-18
+ uc1 = 5.411e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_mvt__tvoff_diff_1}
+ njs = 1.363
+ tpb = 0.002039
+ tcj = 0.001241
+ tpbsw = 0.001246
+ tcjsw = 0.0003736
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 5.2
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 3.29e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.5
+ steta0 = 0.0
.ends sky130_fd_pr__pfet_01v8_mvt
* Well Proximity Effect Parameters
