* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__special_pfet_pass__tox_slope_spectre = 0.0
.param sky130_fd_pr__special_pfet_pass__vth0_slope_spectre = 0.0
.param sky130_fd_pr__special_pfet_pass__voff_slope_spectre = 0.0
.param sky130_fd_pr__special_pfet_pass__nfactor_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__special_pfet_pass__tox_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__special_pfet_pass__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__special_pfet_pass__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__special_pfet_pass__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__special_pfet_pass d g s b
+
.param  l = 1 w = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 mult = 1 sa = 0 sb = 0 sd = 0.0
msky130_fd_pr__special_pfet_pass d g s b sky130_fd_pr__special_pfet_pass__model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs}
.model sky130_fd_pr__special_pfet_pass__model.0 pmos
+ lmin = 1.495e-007 lmax = 1.505e-007 wmin = 1.395e-007 wmax = 1.405e-7
+ level = 49.0
+
+ tnom = 30.0
+ version = 3.2
+ tox = {4.214e-009*sky130_fd_pr__special_pfet_pass__tox_mult}
+ toxm = 4.214e-9
+ xj = 1.15e-7
+ nch = 7.919257e+17
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {0+sky130_fd_pr__special_pfet_pass__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {0+sky130_fd_pr__special_pfet_pass__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ mobmod = 1.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* Diode Parameters
+
*+ ldif = 0.0
*+ hdif = 0.0
*+ rd = 0.0
*+ rs = 0.0
*+ rsc = 0.0
*+ rdc = 0.0
+
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.8866+sky130_fd_pr__special_pfet_pass__vth0_diff_0}
+ k1 = 0.48313
+ k2 = {-0.086211+sky130_fd_pr__special_pfet_pass__k2_diff_0}
+ k3 = {0+sky130_fd_pr__special_pfet_pass__k3_diff}
+ dvt0 = {0+sky130_fd_pr__special_pfet_pass__dvt0_diff}
+ dvt1 = 1.0e-10
+ dvt2 = 0.0
+ dvt0w = 0.0
+ dvt1w = 10001.0
+ dvt2w = 0.0
+ nlx = 0.0
+ w0 = 1.0e-10
+ k3b = 0.0
+ ngate = 1.0e+23
+ vfb = -0.3872688
* Mobility Parameters
+ vsat = {100410+sky130_fd_pr__special_pfet_pass__vsat_diff_0}
+ ua = -1.5724e-9
+ ub = 1.0206e-18
+ uc = -2.1234e-11
+ rdsw = {659.8838+sky130_fd_pr__special_pfet_pass__rdsw_diff_0}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.0038566+sky130_fd_pr__special_pfet_pass__u0_diff_0}
+ a0 = 1.6572
+ keta = 0.032965
+ a1 = 0.0
+ a2 = 0.4
+ ags = 0.01944
+ b0 = 0.0
+ b1 = 0.0
* Subthreshold Current Parameters
+ voff = {-0.17082+sky130_fd_pr__special_pfet_pass__voff_diff_0}
+ nfactor = {2+sky130_fd_pr__special_pfet_pass__nfactor_diff_0}
+ cit = {-0.002+sky130_fd_pr__special_pfet_pass__cit_diff}
+ cdsc = {0+sky130_fd_pr__special_pfet_pass__cdsc_diff}
+ cdscb = {0.0005+sky130_fd_pr__special_pfet_pass__cdscb_diff}
+ cdscd = {0+sky130_fd_pr__special_pfet_pass__cdscd_diff}
+ eta0 = 0.001
+ etab = 0.0
+ dsub = 1.0e-10
* Rout Parameters
+ pclm = 2.4129
+ pdiblc1 = 0.0
+ pdiblc2 = 0.023805348
+ pdiblcb = -0.5
+ drout = 1.0e-10
+ pscbe1 = 7.0054e+8
+ pscbe2 = 1.0e-20
+ pvag = 0.0
+ delta = 0.071729
+ alpha0 = 1.3735e-6
+ alpha1 = 0.0
+ beta0 = 23.765
* Temperature Effects Parameters
+ kt1 = {-0.50219+sky130_fd_pr__special_pfet_pass__kt1_diff_0}
+ kt2 = {-0.048934+sky130_fd_pr__special_pfet_pass__kt2_diff}
+ at = 3000.3
+ ute = -0.8
+ ua1 = -4.1272e-11
+ ub1 = 4.0968e-19
+ uc1 = 1.2689e-11
+ kt1l = {0+sky130_fd_pr__special_pfet_pass__kt1l_diff}
+ prt = 0.49191
* Capacitance Parameters
+ cj = {0.00074079*sky130_fd_pr__special_pfet_pass__ajunction_mult}
+ mj = 0.34629
+ pb = 0.6587
+ cjsw = {9.88e-011*sky130_fd_pr__special_pfet_pass__pjunction_mult}
+ mjsw = 0.29781
+ pbsw = 0.7418
+ cjswg = 2.3894e-10
+ mjswg = 0.9274
+ pbswg = 1.4338
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ js = 2.1483e-5
+ jsw = 8.040000000000001e-10
+ nj = 1.3632
+ xti = 5.2
+ cgdo = {1.4045e-010*sky130_fd_pr__special_pfet_pass__overlap_mult}
+ cgso = {1.4045e-010*sky130_fd_pr__special_pfet_pass__overlap_mult}
+ cgbo = 0.0
+ capmod = 3.0
*+ nqsmod = 0.0
+ elm = 0.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__special_pfet_pass__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__special_pfet_pass__overlap_mult}
+ ckappa = 0.6
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {5.67e-009+sky130_fd_pr__special_pfet_pass__dlc_diff+sky130_fd_pr__special_pfet_pass__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__special_pfet_pass__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.401
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
.model sky130_fd_pr__special_pfet_pass__model.1 pmos
+ lmin = 0.25e-007 lmax = 0.5e-007 wmin = 1.395e-007 wmax = 1.405e-7
+ level = 49.0
+
+ tnom = 30.0
+ version = 3.2
+ tox = {4.214e-009*sky130_fd_pr__special_pfet_pass__tox_mult}
+ toxm = 4.214e-9
+ xj = 1.15e-7
+ nch = 7.919257e+17
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-2.4825e-8+sky130_fd_pr__special_pfet_pass__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {-5.522e-8+sky130_fd_pr__special_pfet_pass__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ mobmod = 1.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* Diode Parameters
+
+ ldif = 0.0
+ hdif = 0.0
+ rd = 0.0
+ rs = 0.0
+ rsc = 0.0
+ rdc = 0.0
+
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.8866+sky130_fd_pr__special_pfet_pass__vth0_diff_0}
+ k1 = 0.48313
+ k2 = {-0.086211+sky130_fd_pr__special_pfet_pass__k2_diff_0}
+ k3 = {0+sky130_fd_pr__special_pfet_pass__k3_diff}
+ dvt0 = {0+sky130_fd_pr__special_pfet_pass__dvt0_diff}
+ dvt1 = 1.0e-10
+ dvt2 = 0.0
+ dvt0w = 0.0
+ dvt1w = 10001.0
+ dvt2w = 0.0
+ nlx = 0.0
+ w0 = 1.0e-10
+ k3b = 0.0
+ ngate = 1.0e+23
+ vfb = -0.3872688
* Mobility Parameters
+ vsat = {100410+sky130_fd_pr__special_pfet_pass__vsat_diff_0}
+ ua = -1.5724e-9
+ ub = 1.0206e-18
+ uc = -2.1234e-11
+ rdsw = {659.8838+sky130_fd_pr__special_pfet_pass__rdsw_diff_0}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.0038566+sky130_fd_pr__special_pfet_pass__u0_diff_0}
+ a0 = 1.6572
+ keta = 0.032965
+ a1 = 0.0
+ a2 = 0.4
+ ags = 0.01944
+ b0 = 0.0
+ b1 = 0.0
* Subthreshold Current Parameters
+ voff = {-0.17082+sky130_fd_pr__special_pfet_pass__voff_diff_0}
+ nfactor = {2+sky130_fd_pr__special_pfet_pass__nfactor_diff_0}
+ cit = {-0.002+sky130_fd_pr__special_pfet_pass__cit_diff}
+ cdsc = {0+sky130_fd_pr__special_pfet_pass__cdsc_diff}
+ cdscb = {0.0005+sky130_fd_pr__special_pfet_pass__cdscb_diff}
+ cdscd = {0+sky130_fd_pr__special_pfet_pass__cdscd_diff}
+ eta0 = 0.001
+ etab = 0.0
+ dsub = 1.0e-10
* Rout Parameters
+ pclm = 2.4129
+ pdiblc1 = 0.0
+ pdiblc2 = 0.023805348
+ pdiblcb = -0.5
+ drout = 1.0e-10
+ pscbe1 = 7.0054e+8
+ pscbe2 = 1.0e-20
+ pvag = 0.0
+ delta = 0.071729
+ alpha0 = 1.3735e-6
+ alpha1 = 0.0
+ beta0 = 23.765
* Temperature Effects Parameters
+ kt1 = {-0.50219+sky130_fd_pr__special_pfet_pass__kt1_diff_0}
+ kt2 = {-0.048934+sky130_fd_pr__special_pfet_pass__kt2_diff}
+ at = 3000.3
+ ute = -0.8
+ ua1 = -4.1272e-11
+ ub1 = 4.0968e-19
+ uc1 = 1.2689e-11
+ kt1l = {0+sky130_fd_pr__special_pfet_pass__kt1l_diff}
+ prt = 0.49191
* Capacitance Parameters
+ cj = {0.00074079*sky130_fd_pr__special_pfet_pass__ajunction_mult}
+ mj = 0.34629
+ pb = 0.6587
+ cjsw = {9.88e-011*sky130_fd_pr__special_pfet_pass__pjunction_mult}
+ mjsw = 0.29781
+ pbsw = 0.7418
+ cjswg = 2.3894e-10
+ mjswg = 0.9274
+ pbswg = 1.4338
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ js = 2.1483e-5
+ jsw = 8.040000000000001e-10
+ nj = 1.3632
+ xti = 5.2
+ cgdo = {1.4045e-010*sky130_fd_pr__special_pfet_pass__overlap_mult}
+ cgso = {1.4045e-010*sky130_fd_pr__special_pfet_pass__overlap_mult}
+ cgbo = 0.0
+ capmod = 3.0
+ nqsmod = 0.0
+ elm = 0.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__special_pfet_pass__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__special_pfet_pass__overlap_mult}
+ ckappa = 0.6
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.4825e-8+sky130_fd_pr__special_pfet_pass__dlc_diff+sky130_fd_pr__special_pfet_pass__dlc_rotweak}
+ dwc = {3.622e-8+sky130_fd_pr__special_pfet_pass__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.401
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
+ noimod = 2.0
+ noia = {5.3000000E+40*1.6e-21}
+ noib = {5.6400000E+22*1.6e-21}
+ noic = {6.0700000E+07*1.6e-21}
+ em = 4.1000000e+7
+ ef = 0.88
.ends sky130_fd_pr__special_pfet_pass
