// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

/* Generated by Yosys 0.9+3621 (git sha1 84e9fa7, gcc 8.3.1 -fPIC -Os) */

module mgmt_protect_hv(mprj2_vdd_logic1, mprj_vdd_logic1, vccd, vssd, vdda1, vssa1, vdda2, vssa2);
  output mprj2_vdd_logic1;
  wire mprj2_vdd_logic1_h;
  output mprj_vdd_logic1;
  wire mprj_vdd_logic1_h;
  input vccd;
  input vdda1;
  input vdda2;
  input vssa1;
  input vssa2;
  input vssd;
  sky130_fd_sc_hvl__decap_8 FILLER_0_0 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_104 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_112 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_120 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_128 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_136 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_144 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_152 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_16 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_160 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_168 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_176 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_184 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_192 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_200 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_208 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_216 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_224 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_232 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_24 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_240 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_248 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_256 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_264 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_272 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_280 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_288 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_296 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_304 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_312 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_32 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_320 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_328 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_336 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_344 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_352 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_360 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_368 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_376 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_384 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_392 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_40 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_4 FILLER_0_400 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__fill_2 FILLER_0_404 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_48 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_56 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_64 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_72 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_8 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_80 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_88 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_0_96 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_0 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_114 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_122 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_130 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_138 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_146 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_154 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_16 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_162 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_170 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_178 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_186 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_194 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_202 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_210 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_218 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_226 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_234 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_24 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_242 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_250 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_258 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_266 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_274 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_282 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_290 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_298 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_306 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_314 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_32 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_322 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_330 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_338 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_346 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_354 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_362 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__fill_2 FILLER_1_370 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_389 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_397 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_40 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__fill_1 FILLER_1_405 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_48 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_56 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_64 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_72 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_8 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_80 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_1_88 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__fill_1 FILLER_1_96 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_0 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_114 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_122 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_130 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_138 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_146 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_154 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_16 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_162 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_170 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_178 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_186 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_194 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_202 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_210 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_218 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_226 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_234 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_24 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_242 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_250 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_258 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_266 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_274 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_282 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_290 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_298 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_306 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_314 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_32 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_322 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_330 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_338 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_346 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_354 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_362 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__fill_2 FILLER_2_370 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_389 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_397 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_40 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__fill_1 FILLER_2_405 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_48 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_56 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_64 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_72 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_8 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_80 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_2_88 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__fill_1 FILLER_2_96 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_0 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_104 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_112 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_120 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__fill_1 FILLER_3_128 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_134 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__fill_1 FILLER_3_142 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_148 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_156 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_16 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_164 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_172 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_180 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_188 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_196 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_204 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_212 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_220 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_228 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_236 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_24 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_244 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_252 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_260 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_268 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_276 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_284 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_292 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_300 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_308 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_316 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_32 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_324 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_332 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_340 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_348 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_356 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_364 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_372 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_380 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_388 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_396 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_40 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__fill_2 FILLER_3_404 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_48 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_56 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_64 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_72 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_8 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_80 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_88 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_3_96 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_0 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_104 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_112 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_120 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_128 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_136 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_144 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_152 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_16 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_160 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_168 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_176 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_184 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_192 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_200 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_208 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_216 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_224 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_232 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_24 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_240 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_248 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_256 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_264 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_272 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_280 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_288 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_296 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_304 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_312 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_32 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_320 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_328 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_336 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_344 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_352 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_360 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_368 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_376 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_384 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_392 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_40 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_4 FILLER_4_400 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__fill_2 FILLER_4_404 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_48 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_56 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_64 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_72 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_8 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_80 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_88 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__decap_8 FILLER_4_96 (
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__conb_1 mprj2_logic_high_hvl (
    .HI(mprj2_vdd_logic1_h),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__lsbufhv2lv_1 mprj2_logic_high_lv (
    .A(mprj2_vdd_logic1_h),
    .LVPWR(vdda2),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .X(mprj2_vdd_logic1)
  );
  sky130_fd_sc_hvl__conb_1 mprj_logic_high_hvl (
    .HI(mprj_vdd_logic1_h),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2)
  );
  sky130_fd_sc_hvl__lsbufhv2lv_1 mprj_logic_high_lv (
    .A(mprj_vdd_logic1_h),
    .LVPWR(vdda2),
    .VGND(vssa2),
    .VNB(vssa2),
    .VPB(vdda2),
    .VPWR(vdda2),
    .X(mprj_vdd_logic1)
  );
endmodule
