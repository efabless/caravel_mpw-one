VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_core
  CLASS BLOCK ;
  FOREIGN mgmt_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 2150.000 BY 860.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END clock
  PIN core_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 856.000 1.750 860.000 ;
    END
  END core_clk
  PIN core_rstn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 856.000 4.970 860.000 ;
    END
  END core_rstn
  PIN flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.870 0.000 1124.150 4.000 ;
    END
  END flash_clk
  PIN flash_clk_ieb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.390 0.000 1221.670 4.000 ;
    END
  END flash_clk_ieb
  PIN flash_clk_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1318.910 0.000 1319.190 4.000 ;
    END
  END flash_clk_oeb
  PIN flash_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.390 0.000 830.670 4.000 ;
    END
  END flash_csb
  PIN flash_csb_ieb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.370 0.000 928.650 4.000 ;
    END
  END flash_csb_ieb
  PIN flash_csb_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.890 0.000 1026.170 4.000 ;
    END
  END flash_csb_oeb
  PIN flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.890 0.000 1417.170 4.000 ;
    END
  END flash_io0_di
  PIN flash_io0_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1514.410 0.000 1514.690 4.000 ;
    END
  END flash_io0_do
  PIN flash_io0_ieb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1612.390 0.000 1612.670 4.000 ;
    END
  END flash_io0_ieb
  PIN flash_io0_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.910 0.000 1710.190 4.000 ;
    END
  END flash_io0_oeb
  PIN flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1807.890 0.000 1808.170 4.000 ;
    END
  END flash_io1_di
  PIN flash_io1_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.410 0.000 1905.690 4.000 ;
    END
  END flash_io1_do
  PIN flash_io1_ieb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2003.390 0.000 2003.670 4.000 ;
    END
  END flash_io1_ieb
  PIN flash_io1_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.910 0.000 2101.190 4.000 ;
    END
  END flash_io1_oeb
  PIN flash_io2_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 845.960 4.000 846.560 ;
    END
  END flash_io2_do
  PIN flash_io2_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 845.280 2150.000 845.880 ;
    END
  END flash_io2_oeb
  PIN flash_io3_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 854.800 2150.000 855.400 ;
    END
  END flash_io3_do
  PIN flash_io3_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 851.400 4.000 852.000 ;
    END
  END flash_io3_oeb
  PIN gpio_in_pad
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END gpio_in_pad
  PIN gpio_inenb_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 4.000 ;
    END
  END gpio_inenb_pad
  PIN gpio_mode0_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 0.000 439.670 4.000 ;
    END
  END gpio_mode0_pad
  PIN gpio_mode1_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 0.000 537.650 4.000 ;
    END
  END gpio_mode1_pad
  PIN gpio_out_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 0.000 635.170 4.000 ;
    END
  END gpio_out_pad
  PIN gpio_outenb_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 0.000 733.150 4.000 ;
    END
  END gpio_outenb_pad
  PIN jtag_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 323.720 2150.000 324.320 ;
    END
  END jtag_out
  PIN jtag_outenb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 333.240 2150.000 333.840 ;
    END
  END jtag_outenb
  PIN la_iena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 856.000 440.130 860.000 ;
    END
  END la_iena[0]
  PIN la_iena[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.610 856.000 764.890 860.000 ;
    END
  END la_iena[100]
  PIN la_iena[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 856.000 768.110 860.000 ;
    END
  END la_iena[101]
  PIN la_iena[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.050 856.000 771.330 860.000 ;
    END
  END la_iena[102]
  PIN la_iena[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.270 856.000 774.550 860.000 ;
    END
  END la_iena[103]
  PIN la_iena[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.490 856.000 777.770 860.000 ;
    END
  END la_iena[104]
  PIN la_iena[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.710 856.000 780.990 860.000 ;
    END
  END la_iena[105]
  PIN la_iena[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.930 856.000 784.210 860.000 ;
    END
  END la_iena[106]
  PIN la_iena[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 856.000 787.430 860.000 ;
    END
  END la_iena[107]
  PIN la_iena[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.370 856.000 790.650 860.000 ;
    END
  END la_iena[108]
  PIN la_iena[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 856.000 793.870 860.000 ;
    END
  END la_iena[109]
  PIN la_iena[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 856.000 472.330 860.000 ;
    END
  END la_iena[10]
  PIN la_iena[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.810 856.000 797.090 860.000 ;
    END
  END la_iena[110]
  PIN la_iena[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.030 856.000 800.310 860.000 ;
    END
  END la_iena[111]
  PIN la_iena[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.250 856.000 803.530 860.000 ;
    END
  END la_iena[112]
  PIN la_iena[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.470 856.000 806.750 860.000 ;
    END
  END la_iena[113]
  PIN la_iena[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.150 856.000 810.430 860.000 ;
    END
  END la_iena[114]
  PIN la_iena[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.370 856.000 813.650 860.000 ;
    END
  END la_iena[115]
  PIN la_iena[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.590 856.000 816.870 860.000 ;
    END
  END la_iena[116]
  PIN la_iena[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 856.000 820.090 860.000 ;
    END
  END la_iena[117]
  PIN la_iena[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.030 856.000 823.310 860.000 ;
    END
  END la_iena[118]
  PIN la_iena[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.250 856.000 826.530 860.000 ;
    END
  END la_iena[119]
  PIN la_iena[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 856.000 475.550 860.000 ;
    END
  END la_iena[11]
  PIN la_iena[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.470 856.000 829.750 860.000 ;
    END
  END la_iena[120]
  PIN la_iena[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.690 856.000 832.970 860.000 ;
    END
  END la_iena[121]
  PIN la_iena[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.910 856.000 836.190 860.000 ;
    END
  END la_iena[122]
  PIN la_iena[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.130 856.000 839.410 860.000 ;
    END
  END la_iena[123]
  PIN la_iena[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.350 856.000 842.630 860.000 ;
    END
  END la_iena[124]
  PIN la_iena[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.570 856.000 845.850 860.000 ;
    END
  END la_iena[125]
  PIN la_iena[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 856.000 849.070 860.000 ;
    END
  END la_iena[126]
  PIN la_iena[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.010 856.000 852.290 860.000 ;
    END
  END la_iena[127]
  PIN la_iena[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 856.000 478.770 860.000 ;
    END
  END la_iena[12]
  PIN la_iena[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 856.000 481.990 860.000 ;
    END
  END la_iena[13]
  PIN la_iena[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 856.000 485.670 860.000 ;
    END
  END la_iena[14]
  PIN la_iena[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 856.000 488.890 860.000 ;
    END
  END la_iena[15]
  PIN la_iena[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 856.000 492.110 860.000 ;
    END
  END la_iena[16]
  PIN la_iena[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 856.000 495.330 860.000 ;
    END
  END la_iena[17]
  PIN la_iena[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.270 856.000 498.550 860.000 ;
    END
  END la_iena[18]
  PIN la_iena[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.490 856.000 501.770 860.000 ;
    END
  END la_iena[19]
  PIN la_iena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 856.000 443.350 860.000 ;
    END
  END la_iena[1]
  PIN la_iena[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 856.000 504.990 860.000 ;
    END
  END la_iena[20]
  PIN la_iena[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 856.000 508.210 860.000 ;
    END
  END la_iena[21]
  PIN la_iena[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.150 856.000 511.430 860.000 ;
    END
  END la_iena[22]
  PIN la_iena[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.370 856.000 514.650 860.000 ;
    END
  END la_iena[23]
  PIN la_iena[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 856.000 517.870 860.000 ;
    END
  END la_iena[24]
  PIN la_iena[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 856.000 521.090 860.000 ;
    END
  END la_iena[25]
  PIN la_iena[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 856.000 524.310 860.000 ;
    END
  END la_iena[26]
  PIN la_iena[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.250 856.000 527.530 860.000 ;
    END
  END la_iena[27]
  PIN la_iena[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 856.000 530.750 860.000 ;
    END
  END la_iena[28]
  PIN la_iena[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 856.000 533.970 860.000 ;
    END
  END la_iena[29]
  PIN la_iena[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 856.000 446.570 860.000 ;
    END
  END la_iena[2]
  PIN la_iena[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 856.000 537.190 860.000 ;
    END
  END la_iena[30]
  PIN la_iena[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 856.000 540.870 860.000 ;
    END
  END la_iena[31]
  PIN la_iena[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 856.000 544.090 860.000 ;
    END
  END la_iena[32]
  PIN la_iena[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 856.000 547.310 860.000 ;
    END
  END la_iena[33]
  PIN la_iena[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 856.000 550.530 860.000 ;
    END
  END la_iena[34]
  PIN la_iena[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 856.000 553.750 860.000 ;
    END
  END la_iena[35]
  PIN la_iena[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 856.000 556.970 860.000 ;
    END
  END la_iena[36]
  PIN la_iena[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 856.000 560.190 860.000 ;
    END
  END la_iena[37]
  PIN la_iena[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.130 856.000 563.410 860.000 ;
    END
  END la_iena[38]
  PIN la_iena[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 856.000 566.630 860.000 ;
    END
  END la_iena[39]
  PIN la_iena[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 856.000 449.790 860.000 ;
    END
  END la_iena[3]
  PIN la_iena[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 856.000 569.850 860.000 ;
    END
  END la_iena[40]
  PIN la_iena[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 856.000 573.070 860.000 ;
    END
  END la_iena[41]
  PIN la_iena[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 856.000 576.290 860.000 ;
    END
  END la_iena[42]
  PIN la_iena[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 856.000 579.510 860.000 ;
    END
  END la_iena[43]
  PIN la_iena[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 856.000 582.730 860.000 ;
    END
  END la_iena[44]
  PIN la_iena[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 856.000 585.950 860.000 ;
    END
  END la_iena[45]
  PIN la_iena[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 856.000 589.170 860.000 ;
    END
  END la_iena[46]
  PIN la_iena[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 856.000 592.390 860.000 ;
    END
  END la_iena[47]
  PIN la_iena[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 856.000 596.070 860.000 ;
    END
  END la_iena[48]
  PIN la_iena[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 856.000 599.290 860.000 ;
    END
  END la_iena[49]
  PIN la_iena[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 856.000 453.010 860.000 ;
    END
  END la_iena[4]
  PIN la_iena[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 856.000 602.510 860.000 ;
    END
  END la_iena[50]
  PIN la_iena[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 856.000 605.730 860.000 ;
    END
  END la_iena[51]
  PIN la_iena[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 856.000 608.950 860.000 ;
    END
  END la_iena[52]
  PIN la_iena[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 856.000 612.170 860.000 ;
    END
  END la_iena[53]
  PIN la_iena[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 856.000 615.390 860.000 ;
    END
  END la_iena[54]
  PIN la_iena[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 856.000 618.610 860.000 ;
    END
  END la_iena[55]
  PIN la_iena[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 856.000 621.830 860.000 ;
    END
  END la_iena[56]
  PIN la_iena[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 856.000 625.050 860.000 ;
    END
  END la_iena[57]
  PIN la_iena[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 856.000 628.270 860.000 ;
    END
  END la_iena[58]
  PIN la_iena[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 856.000 631.490 860.000 ;
    END
  END la_iena[59]
  PIN la_iena[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 856.000 456.230 860.000 ;
    END
  END la_iena[5]
  PIN la_iena[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 856.000 634.710 860.000 ;
    END
  END la_iena[60]
  PIN la_iena[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 856.000 637.930 860.000 ;
    END
  END la_iena[61]
  PIN la_iena[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 856.000 641.150 860.000 ;
    END
  END la_iena[62]
  PIN la_iena[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 856.000 644.370 860.000 ;
    END
  END la_iena[63]
  PIN la_iena[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.770 856.000 648.050 860.000 ;
    END
  END la_iena[64]
  PIN la_iena[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.990 856.000 651.270 860.000 ;
    END
  END la_iena[65]
  PIN la_iena[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 856.000 654.490 860.000 ;
    END
  END la_iena[66]
  PIN la_iena[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 856.000 657.710 860.000 ;
    END
  END la_iena[67]
  PIN la_iena[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 856.000 660.930 860.000 ;
    END
  END la_iena[68]
  PIN la_iena[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 856.000 664.150 860.000 ;
    END
  END la_iena[69]
  PIN la_iena[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 856.000 459.450 860.000 ;
    END
  END la_iena[6]
  PIN la_iena[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 856.000 667.370 860.000 ;
    END
  END la_iena[70]
  PIN la_iena[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 856.000 670.590 860.000 ;
    END
  END la_iena[71]
  PIN la_iena[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 856.000 673.810 860.000 ;
    END
  END la_iena[72]
  PIN la_iena[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 856.000 677.030 860.000 ;
    END
  END la_iena[73]
  PIN la_iena[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 856.000 680.250 860.000 ;
    END
  END la_iena[74]
  PIN la_iena[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 856.000 683.470 860.000 ;
    END
  END la_iena[75]
  PIN la_iena[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 856.000 686.690 860.000 ;
    END
  END la_iena[76]
  PIN la_iena[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.630 856.000 689.910 860.000 ;
    END
  END la_iena[77]
  PIN la_iena[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.850 856.000 693.130 860.000 ;
    END
  END la_iena[78]
  PIN la_iena[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 856.000 696.350 860.000 ;
    END
  END la_iena[79]
  PIN la_iena[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 856.000 462.670 860.000 ;
    END
  END la_iena[7]
  PIN la_iena[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 856.000 699.570 860.000 ;
    END
  END la_iena[80]
  PIN la_iena[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.970 856.000 703.250 860.000 ;
    END
  END la_iena[81]
  PIN la_iena[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.190 856.000 706.470 860.000 ;
    END
  END la_iena[82]
  PIN la_iena[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 856.000 709.690 860.000 ;
    END
  END la_iena[83]
  PIN la_iena[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 856.000 712.910 860.000 ;
    END
  END la_iena[84]
  PIN la_iena[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 856.000 716.130 860.000 ;
    END
  END la_iena[85]
  PIN la_iena[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.070 856.000 719.350 860.000 ;
    END
  END la_iena[86]
  PIN la_iena[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.290 856.000 722.570 860.000 ;
    END
  END la_iena[87]
  PIN la_iena[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.510 856.000 725.790 860.000 ;
    END
  END la_iena[88]
  PIN la_iena[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.730 856.000 729.010 860.000 ;
    END
  END la_iena[89]
  PIN la_iena[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 856.000 465.890 860.000 ;
    END
  END la_iena[8]
  PIN la_iena[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.950 856.000 732.230 860.000 ;
    END
  END la_iena[90]
  PIN la_iena[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 856.000 735.450 860.000 ;
    END
  END la_iena[91]
  PIN la_iena[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.390 856.000 738.670 860.000 ;
    END
  END la_iena[92]
  PIN la_iena[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 856.000 741.890 860.000 ;
    END
  END la_iena[93]
  PIN la_iena[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.830 856.000 745.110 860.000 ;
    END
  END la_iena[94]
  PIN la_iena[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 856.000 748.330 860.000 ;
    END
  END la_iena[95]
  PIN la_iena[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.270 856.000 751.550 860.000 ;
    END
  END la_iena[96]
  PIN la_iena[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.950 856.000 755.230 860.000 ;
    END
  END la_iena[97]
  PIN la_iena[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 856.000 758.450 860.000 ;
    END
  END la_iena[98]
  PIN la_iena[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.390 856.000 761.670 860.000 ;
    END
  END la_iena[99]
  PIN la_iena[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.830 856.000 469.110 860.000 ;
    END
  END la_iena[9]
  PIN la_input[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.230 856.000 855.510 860.000 ;
    END
  END la_input[0]
  PIN la_input[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.990 856.000 1180.270 860.000 ;
    END
  END la_input[100]
  PIN la_input[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.210 856.000 1183.490 860.000 ;
    END
  END la_input[101]
  PIN la_input[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1186.890 856.000 1187.170 860.000 ;
    END
  END la_input[102]
  PIN la_input[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.110 856.000 1190.390 860.000 ;
    END
  END la_input[103]
  PIN la_input[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1193.330 856.000 1193.610 860.000 ;
    END
  END la_input[104]
  PIN la_input[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.550 856.000 1196.830 860.000 ;
    END
  END la_input[105]
  PIN la_input[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1199.770 856.000 1200.050 860.000 ;
    END
  END la_input[106]
  PIN la_input[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.990 856.000 1203.270 860.000 ;
    END
  END la_input[107]
  PIN la_input[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1206.210 856.000 1206.490 860.000 ;
    END
  END la_input[108]
  PIN la_input[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1209.430 856.000 1209.710 860.000 ;
    END
  END la_input[109]
  PIN la_input[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.890 856.000 888.170 860.000 ;
    END
  END la_input[10]
  PIN la_input[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1212.650 856.000 1212.930 860.000 ;
    END
  END la_input[110]
  PIN la_input[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.870 856.000 1216.150 860.000 ;
    END
  END la_input[111]
  PIN la_input[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1219.090 856.000 1219.370 860.000 ;
    END
  END la_input[112]
  PIN la_input[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1222.310 856.000 1222.590 860.000 ;
    END
  END la_input[113]
  PIN la_input[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.530 856.000 1225.810 860.000 ;
    END
  END la_input[114]
  PIN la_input[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1228.750 856.000 1229.030 860.000 ;
    END
  END la_input[115]
  PIN la_input[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.970 856.000 1232.250 860.000 ;
    END
  END la_input[116]
  PIN la_input[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1235.190 856.000 1235.470 860.000 ;
    END
  END la_input[117]
  PIN la_input[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.870 856.000 1239.150 860.000 ;
    END
  END la_input[118]
  PIN la_input[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.090 856.000 1242.370 860.000 ;
    END
  END la_input[119]
  PIN la_input[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.110 856.000 891.390 860.000 ;
    END
  END la_input[11]
  PIN la_input[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1245.310 856.000 1245.590 860.000 ;
    END
  END la_input[120]
  PIN la_input[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1248.530 856.000 1248.810 860.000 ;
    END
  END la_input[121]
  PIN la_input[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1251.750 856.000 1252.030 860.000 ;
    END
  END la_input[122]
  PIN la_input[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1254.970 856.000 1255.250 860.000 ;
    END
  END la_input[123]
  PIN la_input[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.190 856.000 1258.470 860.000 ;
    END
  END la_input[124]
  PIN la_input[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.410 856.000 1261.690 860.000 ;
    END
  END la_input[125]
  PIN la_input[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.630 856.000 1264.910 860.000 ;
    END
  END la_input[126]
  PIN la_input[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.850 856.000 1268.130 860.000 ;
    END
  END la_input[127]
  PIN la_input[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.330 856.000 894.610 860.000 ;
    END
  END la_input[12]
  PIN la_input[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.550 856.000 897.830 860.000 ;
    END
  END la_input[13]
  PIN la_input[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.770 856.000 901.050 860.000 ;
    END
  END la_input[14]
  PIN la_input[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.990 856.000 904.270 860.000 ;
    END
  END la_input[15]
  PIN la_input[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.210 856.000 907.490 860.000 ;
    END
  END la_input[16]
  PIN la_input[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.430 856.000 910.710 860.000 ;
    END
  END la_input[17]
  PIN la_input[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.650 856.000 913.930 860.000 ;
    END
  END la_input[18]
  PIN la_input[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.330 856.000 917.610 860.000 ;
    END
  END la_input[19]
  PIN la_input[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.450 856.000 858.730 860.000 ;
    END
  END la_input[1]
  PIN la_input[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.550 856.000 920.830 860.000 ;
    END
  END la_input[20]
  PIN la_input[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.770 856.000 924.050 860.000 ;
    END
  END la_input[21]
  PIN la_input[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.990 856.000 927.270 860.000 ;
    END
  END la_input[22]
  PIN la_input[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.210 856.000 930.490 860.000 ;
    END
  END la_input[23]
  PIN la_input[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.430 856.000 933.710 860.000 ;
    END
  END la_input[24]
  PIN la_input[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.650 856.000 936.930 860.000 ;
    END
  END la_input[25]
  PIN la_input[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.870 856.000 940.150 860.000 ;
    END
  END la_input[26]
  PIN la_input[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.090 856.000 943.370 860.000 ;
    END
  END la_input[27]
  PIN la_input[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.310 856.000 946.590 860.000 ;
    END
  END la_input[28]
  PIN la_input[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.530 856.000 949.810 860.000 ;
    END
  END la_input[29]
  PIN la_input[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.130 856.000 862.410 860.000 ;
    END
  END la_input[2]
  PIN la_input[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.750 856.000 953.030 860.000 ;
    END
  END la_input[30]
  PIN la_input[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.970 856.000 956.250 860.000 ;
    END
  END la_input[31]
  PIN la_input[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.190 856.000 959.470 860.000 ;
    END
  END la_input[32]
  PIN la_input[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.410 856.000 962.690 860.000 ;
    END
  END la_input[33]
  PIN la_input[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.630 856.000 965.910 860.000 ;
    END
  END la_input[34]
  PIN la_input[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 856.000 969.590 860.000 ;
    END
  END la_input[35]
  PIN la_input[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 856.000 972.810 860.000 ;
    END
  END la_input[36]
  PIN la_input[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 856.000 976.030 860.000 ;
    END
  END la_input[37]
  PIN la_input[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 856.000 979.250 860.000 ;
    END
  END la_input[38]
  PIN la_input[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.190 856.000 982.470 860.000 ;
    END
  END la_input[39]
  PIN la_input[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.350 856.000 865.630 860.000 ;
    END
  END la_input[3]
  PIN la_input[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 856.000 985.690 860.000 ;
    END
  END la_input[40]
  PIN la_input[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.630 856.000 988.910 860.000 ;
    END
  END la_input[41]
  PIN la_input[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 856.000 992.130 860.000 ;
    END
  END la_input[42]
  PIN la_input[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.070 856.000 995.350 860.000 ;
    END
  END la_input[43]
  PIN la_input[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 856.000 998.570 860.000 ;
    END
  END la_input[44]
  PIN la_input[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 856.000 1001.790 860.000 ;
    END
  END la_input[45]
  PIN la_input[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.730 856.000 1005.010 860.000 ;
    END
  END la_input[46]
  PIN la_input[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 856.000 1008.230 860.000 ;
    END
  END la_input[47]
  PIN la_input[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.170 856.000 1011.450 860.000 ;
    END
  END la_input[48]
  PIN la_input[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 856.000 1014.670 860.000 ;
    END
  END la_input[49]
  PIN la_input[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.570 856.000 868.850 860.000 ;
    END
  END la_input[4]
  PIN la_input[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.610 856.000 1017.890 860.000 ;
    END
  END la_input[50]
  PIN la_input[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 856.000 1021.110 860.000 ;
    END
  END la_input[51]
  PIN la_input[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.510 856.000 1024.790 860.000 ;
    END
  END la_input[52]
  PIN la_input[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.730 856.000 1028.010 860.000 ;
    END
  END la_input[53]
  PIN la_input[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.950 856.000 1031.230 860.000 ;
    END
  END la_input[54]
  PIN la_input[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.170 856.000 1034.450 860.000 ;
    END
  END la_input[55]
  PIN la_input[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.390 856.000 1037.670 860.000 ;
    END
  END la_input[56]
  PIN la_input[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.610 856.000 1040.890 860.000 ;
    END
  END la_input[57]
  PIN la_input[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.830 856.000 1044.110 860.000 ;
    END
  END la_input[58]
  PIN la_input[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.050 856.000 1047.330 860.000 ;
    END
  END la_input[59]
  PIN la_input[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.790 856.000 872.070 860.000 ;
    END
  END la_input[5]
  PIN la_input[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.270 856.000 1050.550 860.000 ;
    END
  END la_input[60]
  PIN la_input[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.490 856.000 1053.770 860.000 ;
    END
  END la_input[61]
  PIN la_input[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.710 856.000 1056.990 860.000 ;
    END
  END la_input[62]
  PIN la_input[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.930 856.000 1060.210 860.000 ;
    END
  END la_input[63]
  PIN la_input[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.150 856.000 1063.430 860.000 ;
    END
  END la_input[64]
  PIN la_input[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.370 856.000 1066.650 860.000 ;
    END
  END la_input[65]
  PIN la_input[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.590 856.000 1069.870 860.000 ;
    END
  END la_input[66]
  PIN la_input[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.810 856.000 1073.090 860.000 ;
    END
  END la_input[67]
  PIN la_input[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.490 856.000 1076.770 860.000 ;
    END
  END la_input[68]
  PIN la_input[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.710 856.000 1079.990 860.000 ;
    END
  END la_input[69]
  PIN la_input[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.010 856.000 875.290 860.000 ;
    END
  END la_input[6]
  PIN la_input[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.930 856.000 1083.210 860.000 ;
    END
  END la_input[70]
  PIN la_input[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.150 856.000 1086.430 860.000 ;
    END
  END la_input[71]
  PIN la_input[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1089.370 856.000 1089.650 860.000 ;
    END
  END la_input[72]
  PIN la_input[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.590 856.000 1092.870 860.000 ;
    END
  END la_input[73]
  PIN la_input[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.810 856.000 1096.090 860.000 ;
    END
  END la_input[74]
  PIN la_input[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.030 856.000 1099.310 860.000 ;
    END
  END la_input[75]
  PIN la_input[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.250 856.000 1102.530 860.000 ;
    END
  END la_input[76]
  PIN la_input[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.470 856.000 1105.750 860.000 ;
    END
  END la_input[77]
  PIN la_input[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.690 856.000 1108.970 860.000 ;
    END
  END la_input[78]
  PIN la_input[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.910 856.000 1112.190 860.000 ;
    END
  END la_input[79]
  PIN la_input[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.230 856.000 878.510 860.000 ;
    END
  END la_input[7]
  PIN la_input[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1115.130 856.000 1115.410 860.000 ;
    END
  END la_input[80]
  PIN la_input[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1118.350 856.000 1118.630 860.000 ;
    END
  END la_input[81]
  PIN la_input[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.570 856.000 1121.850 860.000 ;
    END
  END la_input[82]
  PIN la_input[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.790 856.000 1125.070 860.000 ;
    END
  END la_input[83]
  PIN la_input[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.010 856.000 1128.290 860.000 ;
    END
  END la_input[84]
  PIN la_input[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.690 856.000 1131.970 860.000 ;
    END
  END la_input[85]
  PIN la_input[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.910 856.000 1135.190 860.000 ;
    END
  END la_input[86]
  PIN la_input[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.130 856.000 1138.410 860.000 ;
    END
  END la_input[87]
  PIN la_input[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.350 856.000 1141.630 860.000 ;
    END
  END la_input[88]
  PIN la_input[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1144.570 856.000 1144.850 860.000 ;
    END
  END la_input[89]
  PIN la_input[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.450 856.000 881.730 860.000 ;
    END
  END la_input[8]
  PIN la_input[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.790 856.000 1148.070 860.000 ;
    END
  END la_input[90]
  PIN la_input[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.010 856.000 1151.290 860.000 ;
    END
  END la_input[91]
  PIN la_input[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.230 856.000 1154.510 860.000 ;
    END
  END la_input[92]
  PIN la_input[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.450 856.000 1157.730 860.000 ;
    END
  END la_input[93]
  PIN la_input[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.670 856.000 1160.950 860.000 ;
    END
  END la_input[94]
  PIN la_input[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1163.890 856.000 1164.170 860.000 ;
    END
  END la_input[95]
  PIN la_input[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1167.110 856.000 1167.390 860.000 ;
    END
  END la_input[96]
  PIN la_input[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1170.330 856.000 1170.610 860.000 ;
    END
  END la_input[97]
  PIN la_input[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.550 856.000 1173.830 860.000 ;
    END
  END la_input[98]
  PIN la_input[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.770 856.000 1177.050 860.000 ;
    END
  END la_input[99]
  PIN la_input[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.670 856.000 884.950 860.000 ;
    END
  END la_input[9]
  PIN la_oenb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.070 856.000 1271.350 860.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1595.830 856.000 1596.110 860.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1599.050 856.000 1599.330 860.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1602.270 856.000 1602.550 860.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1605.490 856.000 1605.770 860.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1608.710 856.000 1608.990 860.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.930 856.000 1612.210 860.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1615.610 856.000 1615.890 860.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1618.830 856.000 1619.110 860.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.050 856.000 1622.330 860.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1625.270 856.000 1625.550 860.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.730 856.000 1304.010 860.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1628.490 856.000 1628.770 860.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1631.710 856.000 1631.990 860.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.930 856.000 1635.210 860.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1638.150 856.000 1638.430 860.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1641.370 856.000 1641.650 860.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1644.590 856.000 1644.870 860.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1647.810 856.000 1648.090 860.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.030 856.000 1651.310 860.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1654.250 856.000 1654.530 860.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.470 856.000 1657.750 860.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1306.950 856.000 1307.230 860.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1660.690 856.000 1660.970 860.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.910 856.000 1664.190 860.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.130 856.000 1667.410 860.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1670.810 856.000 1671.090 860.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.030 856.000 1674.310 860.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1677.250 856.000 1677.530 860.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.470 856.000 1680.750 860.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1683.690 856.000 1683.970 860.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.170 856.000 1310.450 860.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.390 856.000 1313.670 860.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.610 856.000 1316.890 860.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1319.830 856.000 1320.110 860.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.050 856.000 1323.330 860.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.270 856.000 1326.550 860.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.490 856.000 1329.770 860.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.710 856.000 1332.990 860.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.290 856.000 1274.570 860.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.930 856.000 1336.210 860.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1339.150 856.000 1339.430 860.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.370 856.000 1342.650 860.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.050 856.000 1346.330 860.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.270 856.000 1349.550 860.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.490 856.000 1352.770 860.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.710 856.000 1355.990 860.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.930 856.000 1359.210 860.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.150 856.000 1362.430 860.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1365.370 856.000 1365.650 860.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.510 856.000 1277.790 860.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.590 856.000 1368.870 860.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.810 856.000 1372.090 860.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.030 856.000 1375.310 860.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.250 856.000 1378.530 860.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.470 856.000 1381.750 860.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1384.690 856.000 1384.970 860.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.910 856.000 1388.190 860.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.130 856.000 1391.410 860.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.350 856.000 1394.630 860.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.570 856.000 1397.850 860.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.730 856.000 1281.010 860.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1401.250 856.000 1401.530 860.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.470 856.000 1404.750 860.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.690 856.000 1407.970 860.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.910 856.000 1411.190 860.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1414.130 856.000 1414.410 860.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.350 856.000 1417.630 860.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.570 856.000 1420.850 860.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.790 856.000 1424.070 860.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.010 856.000 1427.290 860.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1430.230 856.000 1430.510 860.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.950 856.000 1284.230 860.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1433.450 856.000 1433.730 860.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.670 856.000 1436.950 860.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.890 856.000 1440.170 860.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1443.110 856.000 1443.390 860.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1446.330 856.000 1446.610 860.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.550 856.000 1449.830 860.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.230 856.000 1453.510 860.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.450 856.000 1456.730 860.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.670 856.000 1459.950 860.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.890 856.000 1463.170 860.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.170 856.000 1287.450 860.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1466.110 856.000 1466.390 860.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1469.330 856.000 1469.610 860.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.550 856.000 1472.830 860.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.770 856.000 1476.050 860.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.990 856.000 1479.270 860.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1482.210 856.000 1482.490 860.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1485.430 856.000 1485.710 860.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1488.650 856.000 1488.930 860.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1491.870 856.000 1492.150 860.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1495.090 856.000 1495.370 860.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1290.390 856.000 1290.670 860.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.310 856.000 1498.590 860.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1501.530 856.000 1501.810 860.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1504.750 856.000 1505.030 860.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1508.430 856.000 1508.710 860.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1511.650 856.000 1511.930 860.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1514.870 856.000 1515.150 860.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.090 856.000 1518.370 860.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.310 856.000 1521.590 860.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1524.530 856.000 1524.810 860.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.750 856.000 1528.030 860.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.070 856.000 1294.350 860.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.970 856.000 1531.250 860.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.190 856.000 1534.470 860.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1537.410 856.000 1537.690 860.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1540.630 856.000 1540.910 860.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1543.850 856.000 1544.130 860.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1547.070 856.000 1547.350 860.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1550.290 856.000 1550.570 860.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1553.510 856.000 1553.790 860.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1556.730 856.000 1557.010 860.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1560.410 856.000 1560.690 860.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.290 856.000 1297.570 860.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.630 856.000 1563.910 860.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1566.850 856.000 1567.130 860.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1570.070 856.000 1570.350 860.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1573.290 856.000 1573.570 860.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.510 856.000 1576.790 860.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1579.730 856.000 1580.010 860.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1582.950 856.000 1583.230 860.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.170 856.000 1586.450 860.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.390 856.000 1589.670 860.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.610 856.000 1592.890 860.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1300.510 856.000 1300.790 860.000 ;
    END
  END la_oenb[9]
  PIN la_output[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1686.910 856.000 1687.190 860.000 ;
    END
  END la_output[0]
  PIN la_output[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2011.670 856.000 2011.950 860.000 ;
    END
  END la_output[100]
  PIN la_output[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2014.890 856.000 2015.170 860.000 ;
    END
  END la_output[101]
  PIN la_output[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2018.110 856.000 2018.390 860.000 ;
    END
  END la_output[102]
  PIN la_output[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2021.330 856.000 2021.610 860.000 ;
    END
  END la_output[103]
  PIN la_output[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2024.550 856.000 2024.830 860.000 ;
    END
  END la_output[104]
  PIN la_output[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2027.770 856.000 2028.050 860.000 ;
    END
  END la_output[105]
  PIN la_output[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.990 856.000 2031.270 860.000 ;
    END
  END la_output[106]
  PIN la_output[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2034.210 856.000 2034.490 860.000 ;
    END
  END la_output[107]
  PIN la_output[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2037.430 856.000 2037.710 860.000 ;
    END
  END la_output[108]
  PIN la_output[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2040.650 856.000 2040.930 860.000 ;
    END
  END la_output[109]
  PIN la_output[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1719.110 856.000 1719.390 860.000 ;
    END
  END la_output[10]
  PIN la_output[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2044.330 856.000 2044.610 860.000 ;
    END
  END la_output[110]
  PIN la_output[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.550 856.000 2047.830 860.000 ;
    END
  END la_output[111]
  PIN la_output[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2050.770 856.000 2051.050 860.000 ;
    END
  END la_output[112]
  PIN la_output[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.990 856.000 2054.270 860.000 ;
    END
  END la_output[113]
  PIN la_output[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2057.210 856.000 2057.490 860.000 ;
    END
  END la_output[114]
  PIN la_output[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2060.430 856.000 2060.710 860.000 ;
    END
  END la_output[115]
  PIN la_output[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2063.650 856.000 2063.930 860.000 ;
    END
  END la_output[116]
  PIN la_output[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2066.870 856.000 2067.150 860.000 ;
    END
  END la_output[117]
  PIN la_output[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2070.090 856.000 2070.370 860.000 ;
    END
  END la_output[118]
  PIN la_output[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2073.310 856.000 2073.590 860.000 ;
    END
  END la_output[119]
  PIN la_output[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.790 856.000 1723.070 860.000 ;
    END
  END la_output[11]
  PIN la_output[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2076.530 856.000 2076.810 860.000 ;
    END
  END la_output[120]
  PIN la_output[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2079.750 856.000 2080.030 860.000 ;
    END
  END la_output[121]
  PIN la_output[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2082.970 856.000 2083.250 860.000 ;
    END
  END la_output[122]
  PIN la_output[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2086.190 856.000 2086.470 860.000 ;
    END
  END la_output[123]
  PIN la_output[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.410 856.000 2089.690 860.000 ;
    END
  END la_output[124]
  PIN la_output[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2092.630 856.000 2092.910 860.000 ;
    END
  END la_output[125]
  PIN la_output[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2095.850 856.000 2096.130 860.000 ;
    END
  END la_output[126]
  PIN la_output[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2099.530 856.000 2099.810 860.000 ;
    END
  END la_output[127]
  PIN la_output[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.010 856.000 1726.290 860.000 ;
    END
  END la_output[12]
  PIN la_output[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.230 856.000 1729.510 860.000 ;
    END
  END la_output[13]
  PIN la_output[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.450 856.000 1732.730 860.000 ;
    END
  END la_output[14]
  PIN la_output[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1735.670 856.000 1735.950 860.000 ;
    END
  END la_output[15]
  PIN la_output[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.890 856.000 1739.170 860.000 ;
    END
  END la_output[16]
  PIN la_output[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.110 856.000 1742.390 860.000 ;
    END
  END la_output[17]
  PIN la_output[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.330 856.000 1745.610 860.000 ;
    END
  END la_output[18]
  PIN la_output[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1748.550 856.000 1748.830 860.000 ;
    END
  END la_output[19]
  PIN la_output[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1690.130 856.000 1690.410 860.000 ;
    END
  END la_output[1]
  PIN la_output[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.770 856.000 1752.050 860.000 ;
    END
  END la_output[20]
  PIN la_output[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.990 856.000 1755.270 860.000 ;
    END
  END la_output[21]
  PIN la_output[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.210 856.000 1758.490 860.000 ;
    END
  END la_output[22]
  PIN la_output[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.430 856.000 1761.710 860.000 ;
    END
  END la_output[23]
  PIN la_output[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.650 856.000 1764.930 860.000 ;
    END
  END la_output[24]
  PIN la_output[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1767.870 856.000 1768.150 860.000 ;
    END
  END la_output[25]
  PIN la_output[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1771.090 856.000 1771.370 860.000 ;
    END
  END la_output[26]
  PIN la_output[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.310 856.000 1774.590 860.000 ;
    END
  END la_output[27]
  PIN la_output[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.990 856.000 1778.270 860.000 ;
    END
  END la_output[28]
  PIN la_output[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.210 856.000 1781.490 860.000 ;
    END
  END la_output[29]
  PIN la_output[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.350 856.000 1693.630 860.000 ;
    END
  END la_output[2]
  PIN la_output[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1784.430 856.000 1784.710 860.000 ;
    END
  END la_output[30]
  PIN la_output[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.650 856.000 1787.930 860.000 ;
    END
  END la_output[31]
  PIN la_output[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1790.870 856.000 1791.150 860.000 ;
    END
  END la_output[32]
  PIN la_output[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1794.090 856.000 1794.370 860.000 ;
    END
  END la_output[33]
  PIN la_output[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1797.310 856.000 1797.590 860.000 ;
    END
  END la_output[34]
  PIN la_output[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1800.530 856.000 1800.810 860.000 ;
    END
  END la_output[35]
  PIN la_output[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1803.750 856.000 1804.030 860.000 ;
    END
  END la_output[36]
  PIN la_output[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1806.970 856.000 1807.250 860.000 ;
    END
  END la_output[37]
  PIN la_output[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.190 856.000 1810.470 860.000 ;
    END
  END la_output[38]
  PIN la_output[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1813.410 856.000 1813.690 860.000 ;
    END
  END la_output[39]
  PIN la_output[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1696.570 856.000 1696.850 860.000 ;
    END
  END la_output[3]
  PIN la_output[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.630 856.000 1816.910 860.000 ;
    END
  END la_output[40]
  PIN la_output[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1819.850 856.000 1820.130 860.000 ;
    END
  END la_output[41]
  PIN la_output[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1823.070 856.000 1823.350 860.000 ;
    END
  END la_output[42]
  PIN la_output[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1826.290 856.000 1826.570 860.000 ;
    END
  END la_output[43]
  PIN la_output[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1829.970 856.000 1830.250 860.000 ;
    END
  END la_output[44]
  PIN la_output[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1833.190 856.000 1833.470 860.000 ;
    END
  END la_output[45]
  PIN la_output[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1836.410 856.000 1836.690 860.000 ;
    END
  END la_output[46]
  PIN la_output[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1839.630 856.000 1839.910 860.000 ;
    END
  END la_output[47]
  PIN la_output[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1842.850 856.000 1843.130 860.000 ;
    END
  END la_output[48]
  PIN la_output[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.070 856.000 1846.350 860.000 ;
    END
  END la_output[49]
  PIN la_output[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.790 856.000 1700.070 860.000 ;
    END
  END la_output[4]
  PIN la_output[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1849.290 856.000 1849.570 860.000 ;
    END
  END la_output[50]
  PIN la_output[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.510 856.000 1852.790 860.000 ;
    END
  END la_output[51]
  PIN la_output[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1855.730 856.000 1856.010 860.000 ;
    END
  END la_output[52]
  PIN la_output[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.950 856.000 1859.230 860.000 ;
    END
  END la_output[53]
  PIN la_output[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1862.170 856.000 1862.450 860.000 ;
    END
  END la_output[54]
  PIN la_output[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1865.390 856.000 1865.670 860.000 ;
    END
  END la_output[55]
  PIN la_output[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1868.610 856.000 1868.890 860.000 ;
    END
  END la_output[56]
  PIN la_output[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1871.830 856.000 1872.110 860.000 ;
    END
  END la_output[57]
  PIN la_output[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1875.050 856.000 1875.330 860.000 ;
    END
  END la_output[58]
  PIN la_output[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1878.270 856.000 1878.550 860.000 ;
    END
  END la_output[59]
  PIN la_output[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.010 856.000 1703.290 860.000 ;
    END
  END la_output[5]
  PIN la_output[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.490 856.000 1881.770 860.000 ;
    END
  END la_output[60]
  PIN la_output[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1885.170 856.000 1885.450 860.000 ;
    END
  END la_output[61]
  PIN la_output[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.390 856.000 1888.670 860.000 ;
    END
  END la_output[62]
  PIN la_output[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1891.610 856.000 1891.890 860.000 ;
    END
  END la_output[63]
  PIN la_output[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1894.830 856.000 1895.110 860.000 ;
    END
  END la_output[64]
  PIN la_output[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1898.050 856.000 1898.330 860.000 ;
    END
  END la_output[65]
  PIN la_output[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1901.270 856.000 1901.550 860.000 ;
    END
  END la_output[66]
  PIN la_output[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.490 856.000 1904.770 860.000 ;
    END
  END la_output[67]
  PIN la_output[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1907.710 856.000 1907.990 860.000 ;
    END
  END la_output[68]
  PIN la_output[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1910.930 856.000 1911.210 860.000 ;
    END
  END la_output[69]
  PIN la_output[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.230 856.000 1706.510 860.000 ;
    END
  END la_output[6]
  PIN la_output[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1914.150 856.000 1914.430 860.000 ;
    END
  END la_output[70]
  PIN la_output[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.370 856.000 1917.650 860.000 ;
    END
  END la_output[71]
  PIN la_output[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1920.590 856.000 1920.870 860.000 ;
    END
  END la_output[72]
  PIN la_output[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.810 856.000 1924.090 860.000 ;
    END
  END la_output[73]
  PIN la_output[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1927.030 856.000 1927.310 860.000 ;
    END
  END la_output[74]
  PIN la_output[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1930.250 856.000 1930.530 860.000 ;
    END
  END la_output[75]
  PIN la_output[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1933.470 856.000 1933.750 860.000 ;
    END
  END la_output[76]
  PIN la_output[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1937.150 856.000 1937.430 860.000 ;
    END
  END la_output[77]
  PIN la_output[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1940.370 856.000 1940.650 860.000 ;
    END
  END la_output[78]
  PIN la_output[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1943.590 856.000 1943.870 860.000 ;
    END
  END la_output[79]
  PIN la_output[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.450 856.000 1709.730 860.000 ;
    END
  END la_output[7]
  PIN la_output[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1946.810 856.000 1947.090 860.000 ;
    END
  END la_output[80]
  PIN la_output[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1950.030 856.000 1950.310 860.000 ;
    END
  END la_output[81]
  PIN la_output[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.250 856.000 1953.530 860.000 ;
    END
  END la_output[82]
  PIN la_output[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1956.470 856.000 1956.750 860.000 ;
    END
  END la_output[83]
  PIN la_output[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.690 856.000 1959.970 860.000 ;
    END
  END la_output[84]
  PIN la_output[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1962.910 856.000 1963.190 860.000 ;
    END
  END la_output[85]
  PIN la_output[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1966.130 856.000 1966.410 860.000 ;
    END
  END la_output[86]
  PIN la_output[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1969.350 856.000 1969.630 860.000 ;
    END
  END la_output[87]
  PIN la_output[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1972.570 856.000 1972.850 860.000 ;
    END
  END la_output[88]
  PIN la_output[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1975.790 856.000 1976.070 860.000 ;
    END
  END la_output[89]
  PIN la_output[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1712.670 856.000 1712.950 860.000 ;
    END
  END la_output[8]
  PIN la_output[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1979.010 856.000 1979.290 860.000 ;
    END
  END la_output[90]
  PIN la_output[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1982.230 856.000 1982.510 860.000 ;
    END
  END la_output[91]
  PIN la_output[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1985.450 856.000 1985.730 860.000 ;
    END
  END la_output[92]
  PIN la_output[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.670 856.000 1988.950 860.000 ;
    END
  END la_output[93]
  PIN la_output[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1992.350 856.000 1992.630 860.000 ;
    END
  END la_output[94]
  PIN la_output[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1995.570 856.000 1995.850 860.000 ;
    END
  END la_output[95]
  PIN la_output[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1998.790 856.000 1999.070 860.000 ;
    END
  END la_output[96]
  PIN la_output[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2002.010 856.000 2002.290 860.000 ;
    END
  END la_output[97]
  PIN la_output[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2005.230 856.000 2005.510 860.000 ;
    END
  END la_output[98]
  PIN la_output[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2008.450 856.000 2008.730 860.000 ;
    END
  END la_output[99]
  PIN la_output[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.890 856.000 1716.170 860.000 ;
    END
  END la_output[9]
  PIN mask_rev[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 4.800 2150.000 5.400 ;
    END
  END mask_rev[0]
  PIN mask_rev[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 101.360 2150.000 101.960 ;
    END
  END mask_rev[10]
  PIN mask_rev[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 110.880 2150.000 111.480 ;
    END
  END mask_rev[11]
  PIN mask_rev[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 120.400 2150.000 121.000 ;
    END
  END mask_rev[12]
  PIN mask_rev[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 129.920 2150.000 130.520 ;
    END
  END mask_rev[13]
  PIN mask_rev[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 139.440 2150.000 140.040 ;
    END
  END mask_rev[14]
  PIN mask_rev[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 149.640 2150.000 150.240 ;
    END
  END mask_rev[15]
  PIN mask_rev[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 159.160 2150.000 159.760 ;
    END
  END mask_rev[16]
  PIN mask_rev[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 168.680 2150.000 169.280 ;
    END
  END mask_rev[17]
  PIN mask_rev[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 178.200 2150.000 178.800 ;
    END
  END mask_rev[18]
  PIN mask_rev[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 188.400 2150.000 189.000 ;
    END
  END mask_rev[19]
  PIN mask_rev[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 14.320 2150.000 14.920 ;
    END
  END mask_rev[1]
  PIN mask_rev[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 197.920 2150.000 198.520 ;
    END
  END mask_rev[20]
  PIN mask_rev[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 207.440 2150.000 208.040 ;
    END
  END mask_rev[21]
  PIN mask_rev[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 216.960 2150.000 217.560 ;
    END
  END mask_rev[22]
  PIN mask_rev[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 226.480 2150.000 227.080 ;
    END
  END mask_rev[23]
  PIN mask_rev[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 236.680 2150.000 237.280 ;
    END
  END mask_rev[24]
  PIN mask_rev[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 246.200 2150.000 246.800 ;
    END
  END mask_rev[25]
  PIN mask_rev[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 255.720 2150.000 256.320 ;
    END
  END mask_rev[26]
  PIN mask_rev[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 265.240 2150.000 265.840 ;
    END
  END mask_rev[27]
  PIN mask_rev[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 274.760 2150.000 275.360 ;
    END
  END mask_rev[28]
  PIN mask_rev[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 284.960 2150.000 285.560 ;
    END
  END mask_rev[29]
  PIN mask_rev[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 23.840 2150.000 24.440 ;
    END
  END mask_rev[2]
  PIN mask_rev[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 294.480 2150.000 295.080 ;
    END
  END mask_rev[30]
  PIN mask_rev[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 304.000 2150.000 304.600 ;
    END
  END mask_rev[31]
  PIN mask_rev[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 33.360 2150.000 33.960 ;
    END
  END mask_rev[3]
  PIN mask_rev[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 42.880 2150.000 43.480 ;
    END
  END mask_rev[4]
  PIN mask_rev[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 53.080 2150.000 53.680 ;
    END
  END mask_rev[5]
  PIN mask_rev[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 62.600 2150.000 63.200 ;
    END
  END mask_rev[6]
  PIN mask_rev[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 72.120 2150.000 72.720 ;
    END
  END mask_rev[7]
  PIN mask_rev[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 81.640 2150.000 82.240 ;
    END
  END mask_rev[8]
  PIN mask_rev[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 91.160 2150.000 91.760 ;
    END
  END mask_rev[9]
  PIN mgmt_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END mgmt_addr[0]
  PIN mgmt_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END mgmt_addr[1]
  PIN mgmt_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END mgmt_addr[2]
  PIN mgmt_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END mgmt_addr[3]
  PIN mgmt_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END mgmt_addr[4]
  PIN mgmt_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END mgmt_addr[5]
  PIN mgmt_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END mgmt_addr[6]
  PIN mgmt_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END mgmt_addr[7]
  PIN mgmt_addr_ro[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END mgmt_addr_ro[0]
  PIN mgmt_addr_ro[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END mgmt_addr_ro[1]
  PIN mgmt_addr_ro[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END mgmt_addr_ro[2]
  PIN mgmt_addr_ro[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END mgmt_addr_ro[3]
  PIN mgmt_addr_ro[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END mgmt_addr_ro[4]
  PIN mgmt_addr_ro[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END mgmt_addr_ro[5]
  PIN mgmt_addr_ro[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END mgmt_addr_ro[6]
  PIN mgmt_addr_ro[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END mgmt_addr_ro[7]
  PIN mgmt_ena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END mgmt_ena[0]
  PIN mgmt_ena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END mgmt_ena[1]
  PIN mgmt_ena_ro
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END mgmt_ena_ro
  PIN mgmt_in_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 381.520 2150.000 382.120 ;
    END
  END mgmt_in_data[0]
  PIN mgmt_in_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 574.640 2150.000 575.240 ;
    END
  END mgmt_in_data[10]
  PIN mgmt_in_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 594.360 2150.000 594.960 ;
    END
  END mgmt_in_data[11]
  PIN mgmt_in_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 613.400 2150.000 614.000 ;
    END
  END mgmt_in_data[12]
  PIN mgmt_in_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 632.440 2150.000 633.040 ;
    END
  END mgmt_in_data[13]
  PIN mgmt_in_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 652.160 2150.000 652.760 ;
    END
  END mgmt_in_data[14]
  PIN mgmt_in_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 671.200 2150.000 671.800 ;
    END
  END mgmt_in_data[15]
  PIN mgmt_in_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 690.920 2150.000 691.520 ;
    END
  END mgmt_in_data[16]
  PIN mgmt_in_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 709.960 2150.000 710.560 ;
    END
  END mgmt_in_data[17]
  PIN mgmt_in_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 729.680 2150.000 730.280 ;
    END
  END mgmt_in_data[18]
  PIN mgmt_in_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 748.720 2150.000 749.320 ;
    END
  END mgmt_in_data[19]
  PIN mgmt_in_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 400.560 2150.000 401.160 ;
    END
  END mgmt_in_data[1]
  PIN mgmt_in_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 767.760 2150.000 768.360 ;
    END
  END mgmt_in_data[20]
  PIN mgmt_in_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 787.480 2150.000 788.080 ;
    END
  END mgmt_in_data[21]
  PIN mgmt_in_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 806.520 2150.000 807.120 ;
    END
  END mgmt_in_data[22]
  PIN mgmt_in_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 826.240 2150.000 826.840 ;
    END
  END mgmt_in_data[23]
  PIN mgmt_in_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 856.000 95.590 860.000 ;
    END
  END mgmt_in_data[24]
  PIN mgmt_in_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 856.000 89.150 860.000 ;
    END
  END mgmt_in_data[25]
  PIN mgmt_in_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 856.000 82.710 860.000 ;
    END
  END mgmt_in_data[26]
  PIN mgmt_in_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 856.000 76.270 860.000 ;
    END
  END mgmt_in_data[27]
  PIN mgmt_in_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 856.000 69.830 860.000 ;
    END
  END mgmt_in_data[28]
  PIN mgmt_in_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 856.000 63.390 860.000 ;
    END
  END mgmt_in_data[29]
  PIN mgmt_in_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 420.280 2150.000 420.880 ;
    END
  END mgmt_in_data[2]
  PIN mgmt_in_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 856.000 56.950 860.000 ;
    END
  END mgmt_in_data[30]
  PIN mgmt_in_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 856.000 50.050 860.000 ;
    END
  END mgmt_in_data[31]
  PIN mgmt_in_data[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 856.000 43.610 860.000 ;
    END
  END mgmt_in_data[32]
  PIN mgmt_in_data[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 856.000 37.170 860.000 ;
    END
  END mgmt_in_data[33]
  PIN mgmt_in_data[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 856.000 30.730 860.000 ;
    END
  END mgmt_in_data[34]
  PIN mgmt_in_data[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 856.000 24.290 860.000 ;
    END
  END mgmt_in_data[35]
  PIN mgmt_in_data[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 856.000 17.850 860.000 ;
    END
  END mgmt_in_data[36]
  PIN mgmt_in_data[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 856.000 11.410 860.000 ;
    END
  END mgmt_in_data[37]
  PIN mgmt_in_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 439.320 2150.000 439.920 ;
    END
  END mgmt_in_data[3]
  PIN mgmt_in_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 459.040 2150.000 459.640 ;
    END
  END mgmt_in_data[4]
  PIN mgmt_in_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 478.080 2150.000 478.680 ;
    END
  END mgmt_in_data[5]
  PIN mgmt_in_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 497.120 2150.000 497.720 ;
    END
  END mgmt_in_data[6]
  PIN mgmt_in_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 516.840 2150.000 517.440 ;
    END
  END mgmt_in_data[7]
  PIN mgmt_in_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 535.880 2150.000 536.480 ;
    END
  END mgmt_in_data[8]
  PIN mgmt_in_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 555.600 2150.000 556.200 ;
    END
  END mgmt_in_data[9]
  PIN mgmt_out_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 391.040 2150.000 391.640 ;
    END
  END mgmt_out_data[0]
  PIN mgmt_out_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 584.160 2150.000 584.760 ;
    END
  END mgmt_out_data[10]
  PIN mgmt_out_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 603.880 2150.000 604.480 ;
    END
  END mgmt_out_data[11]
  PIN mgmt_out_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 622.920 2150.000 623.520 ;
    END
  END mgmt_out_data[12]
  PIN mgmt_out_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 642.640 2150.000 643.240 ;
    END
  END mgmt_out_data[13]
  PIN mgmt_out_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 661.680 2150.000 662.280 ;
    END
  END mgmt_out_data[14]
  PIN mgmt_out_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 680.720 2150.000 681.320 ;
    END
  END mgmt_out_data[15]
  PIN mgmt_out_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 700.440 2150.000 701.040 ;
    END
  END mgmt_out_data[16]
  PIN mgmt_out_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 719.480 2150.000 720.080 ;
    END
  END mgmt_out_data[17]
  PIN mgmt_out_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 739.200 2150.000 739.800 ;
    END
  END mgmt_out_data[18]
  PIN mgmt_out_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 758.240 2150.000 758.840 ;
    END
  END mgmt_out_data[19]
  PIN mgmt_out_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 410.080 2150.000 410.680 ;
    END
  END mgmt_out_data[1]
  PIN mgmt_out_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 777.960 2150.000 778.560 ;
    END
  END mgmt_out_data[20]
  PIN mgmt_out_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 797.000 2150.000 797.600 ;
    END
  END mgmt_out_data[21]
  PIN mgmt_out_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 816.040 2150.000 816.640 ;
    END
  END mgmt_out_data[22]
  PIN mgmt_out_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 835.760 2150.000 836.360 ;
    END
  END mgmt_out_data[23]
  PIN mgmt_out_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 856.000 98.810 860.000 ;
    END
  END mgmt_out_data[24]
  PIN mgmt_out_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 856.000 92.370 860.000 ;
    END
  END mgmt_out_data[25]
  PIN mgmt_out_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 856.000 85.930 860.000 ;
    END
  END mgmt_out_data[26]
  PIN mgmt_out_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 856.000 79.490 860.000 ;
    END
  END mgmt_out_data[27]
  PIN mgmt_out_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 856.000 73.050 860.000 ;
    END
  END mgmt_out_data[28]
  PIN mgmt_out_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 856.000 66.610 860.000 ;
    END
  END mgmt_out_data[29]
  PIN mgmt_out_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 429.800 2150.000 430.400 ;
    END
  END mgmt_out_data[2]
  PIN mgmt_out_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 856.000 60.170 860.000 ;
    END
  END mgmt_out_data[30]
  PIN mgmt_out_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 856.000 53.270 860.000 ;
    END
  END mgmt_out_data[31]
  PIN mgmt_out_data[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 856.000 46.830 860.000 ;
    END
  END mgmt_out_data[32]
  PIN mgmt_out_data[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 856.000 40.390 860.000 ;
    END
  END mgmt_out_data[33]
  PIN mgmt_out_data[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 856.000 33.950 860.000 ;
    END
  END mgmt_out_data[34]
  PIN mgmt_out_data[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 856.000 27.510 860.000 ;
    END
  END mgmt_out_data[35]
  PIN mgmt_out_data[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 856.000 21.070 860.000 ;
    END
  END mgmt_out_data[36]
  PIN mgmt_out_data[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 856.000 14.630 860.000 ;
    END
  END mgmt_out_data[37]
  PIN mgmt_out_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 448.840 2150.000 449.440 ;
    END
  END mgmt_out_data[3]
  PIN mgmt_out_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 468.560 2150.000 469.160 ;
    END
  END mgmt_out_data[4]
  PIN mgmt_out_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 487.600 2150.000 488.200 ;
    END
  END mgmt_out_data[5]
  PIN mgmt_out_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 507.320 2150.000 507.920 ;
    END
  END mgmt_out_data[6]
  PIN mgmt_out_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 526.360 2150.000 526.960 ;
    END
  END mgmt_out_data[7]
  PIN mgmt_out_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 545.400 2150.000 546.000 ;
    END
  END mgmt_out_data[8]
  PIN mgmt_out_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 565.120 2150.000 565.720 ;
    END
  END mgmt_out_data[9]
  PIN mgmt_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 4.000 104.680 ;
    END
  END mgmt_rdata[0]
  PIN mgmt_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END mgmt_rdata[10]
  PIN mgmt_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END mgmt_rdata[11]
  PIN mgmt_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END mgmt_rdata[12]
  PIN mgmt_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END mgmt_rdata[13]
  PIN mgmt_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END mgmt_rdata[14]
  PIN mgmt_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END mgmt_rdata[15]
  PIN mgmt_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.760 4.000 190.360 ;
    END
  END mgmt_rdata[16]
  PIN mgmt_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.200 4.000 195.800 ;
    END
  END mgmt_rdata[17]
  PIN mgmt_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END mgmt_rdata[18]
  PIN mgmt_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END mgmt_rdata[19]
  PIN mgmt_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END mgmt_rdata[1]
  PIN mgmt_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.520 4.000 212.120 ;
    END
  END mgmt_rdata[20]
  PIN mgmt_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END mgmt_rdata[21]
  PIN mgmt_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.400 4.000 223.000 ;
    END
  END mgmt_rdata[22]
  PIN mgmt_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END mgmt_rdata[23]
  PIN mgmt_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END mgmt_rdata[24]
  PIN mgmt_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END mgmt_rdata[25]
  PIN mgmt_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END mgmt_rdata[26]
  PIN mgmt_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END mgmt_rdata[27]
  PIN mgmt_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END mgmt_rdata[28]
  PIN mgmt_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END mgmt_rdata[29]
  PIN mgmt_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END mgmt_rdata[2]
  PIN mgmt_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END mgmt_rdata[30]
  PIN mgmt_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END mgmt_rdata[31]
  PIN mgmt_rdata[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END mgmt_rdata[32]
  PIN mgmt_rdata[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END mgmt_rdata[33]
  PIN mgmt_rdata[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END mgmt_rdata[34]
  PIN mgmt_rdata[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.760 4.000 292.360 ;
    END
  END mgmt_rdata[35]
  PIN mgmt_rdata[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.200 4.000 297.800 ;
    END
  END mgmt_rdata[36]
  PIN mgmt_rdata[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END mgmt_rdata[37]
  PIN mgmt_rdata[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.080 4.000 308.680 ;
    END
  END mgmt_rdata[38]
  PIN mgmt_rdata[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 313.520 4.000 314.120 ;
    END
  END mgmt_rdata[39]
  PIN mgmt_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END mgmt_rdata[3]
  PIN mgmt_rdata[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.960 4.000 319.560 ;
    END
  END mgmt_rdata[40]
  PIN mgmt_rdata[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 324.400 4.000 325.000 ;
    END
  END mgmt_rdata[41]
  PIN mgmt_rdata[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END mgmt_rdata[42]
  PIN mgmt_rdata[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.280 4.000 335.880 ;
    END
  END mgmt_rdata[43]
  PIN mgmt_rdata[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END mgmt_rdata[44]
  PIN mgmt_rdata[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 4.000 346.760 ;
    END
  END mgmt_rdata[45]
  PIN mgmt_rdata[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END mgmt_rdata[46]
  PIN mgmt_rdata[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END mgmt_rdata[47]
  PIN mgmt_rdata[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END mgmt_rdata[48]
  PIN mgmt_rdata[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END mgmt_rdata[49]
  PIN mgmt_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END mgmt_rdata[4]
  PIN mgmt_rdata[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END mgmt_rdata[50]
  PIN mgmt_rdata[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END mgmt_rdata[51]
  PIN mgmt_rdata[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END mgmt_rdata[52]
  PIN mgmt_rdata[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END mgmt_rdata[53]
  PIN mgmt_rdata[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END mgmt_rdata[54]
  PIN mgmt_rdata[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 4.000 400.480 ;
    END
  END mgmt_rdata[55]
  PIN mgmt_rdata[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END mgmt_rdata[56]
  PIN mgmt_rdata[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.080 4.000 410.680 ;
    END
  END mgmt_rdata[57]
  PIN mgmt_rdata[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 415.520 4.000 416.120 ;
    END
  END mgmt_rdata[58]
  PIN mgmt_rdata[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.960 4.000 421.560 ;
    END
  END mgmt_rdata[59]
  PIN mgmt_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END mgmt_rdata[5]
  PIN mgmt_rdata[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 426.400 4.000 427.000 ;
    END
  END mgmt_rdata[60]
  PIN mgmt_rdata[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END mgmt_rdata[61]
  PIN mgmt_rdata[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.280 4.000 437.880 ;
    END
  END mgmt_rdata[62]
  PIN mgmt_rdata[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.720 4.000 443.320 ;
    END
  END mgmt_rdata[63]
  PIN mgmt_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END mgmt_rdata[6]
  PIN mgmt_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END mgmt_rdata[7]
  PIN mgmt_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END mgmt_rdata[8]
  PIN mgmt_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END mgmt_rdata[9]
  PIN mgmt_rdata_ro[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.160 4.000 448.760 ;
    END
  END mgmt_rdata_ro[0]
  PIN mgmt_rdata_ro[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END mgmt_rdata_ro[10]
  PIN mgmt_rdata_ro[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END mgmt_rdata_ro[11]
  PIN mgmt_rdata_ro[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END mgmt_rdata_ro[12]
  PIN mgmt_rdata_ro[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END mgmt_rdata_ro[13]
  PIN mgmt_rdata_ro[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.960 4.000 523.560 ;
    END
  END mgmt_rdata_ro[14]
  PIN mgmt_rdata_ro[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 528.400 4.000 529.000 ;
    END
  END mgmt_rdata_ro[15]
  PIN mgmt_rdata_ro[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END mgmt_rdata_ro[16]
  PIN mgmt_rdata_ro[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.280 4.000 539.880 ;
    END
  END mgmt_rdata_ro[17]
  PIN mgmt_rdata_ro[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.720 4.000 545.320 ;
    END
  END mgmt_rdata_ro[18]
  PIN mgmt_rdata_ro[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.160 4.000 550.760 ;
    END
  END mgmt_rdata_ro[19]
  PIN mgmt_rdata_ro[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 453.600 4.000 454.200 ;
    END
  END mgmt_rdata_ro[1]
  PIN mgmt_rdata_ro[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 555.600 4.000 556.200 ;
    END
  END mgmt_rdata_ro[20]
  PIN mgmt_rdata_ro[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END mgmt_rdata_ro[21]
  PIN mgmt_rdata_ro[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 566.480 4.000 567.080 ;
    END
  END mgmt_rdata_ro[22]
  PIN mgmt_rdata_ro[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.920 4.000 572.520 ;
    END
  END mgmt_rdata_ro[23]
  PIN mgmt_rdata_ro[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 576.680 4.000 577.280 ;
    END
  END mgmt_rdata_ro[24]
  PIN mgmt_rdata_ro[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END mgmt_rdata_ro[25]
  PIN mgmt_rdata_ro[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 587.560 4.000 588.160 ;
    END
  END mgmt_rdata_ro[26]
  PIN mgmt_rdata_ro[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.000 4.000 593.600 ;
    END
  END mgmt_rdata_ro[27]
  PIN mgmt_rdata_ro[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END mgmt_rdata_ro[28]
  PIN mgmt_rdata_ro[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.880 4.000 604.480 ;
    END
  END mgmt_rdata_ro[29]
  PIN mgmt_rdata_ro[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END mgmt_rdata_ro[2]
  PIN mgmt_rdata_ro[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 609.320 4.000 609.920 ;
    END
  END mgmt_rdata_ro[30]
  PIN mgmt_rdata_ro[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.760 4.000 615.360 ;
    END
  END mgmt_rdata_ro[31]
  PIN mgmt_rdata_ro[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END mgmt_rdata_ro[3]
  PIN mgmt_rdata_ro[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END mgmt_rdata_ro[4]
  PIN mgmt_rdata_ro[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END mgmt_rdata_ro[5]
  PIN mgmt_rdata_ro[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END mgmt_rdata_ro[6]
  PIN mgmt_rdata_ro[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END mgmt_rdata_ro[7]
  PIN mgmt_rdata_ro[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END mgmt_rdata_ro[8]
  PIN mgmt_rdata_ro[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END mgmt_rdata_ro[9]
  PIN mgmt_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.200 4.000 620.800 ;
    END
  END mgmt_wdata[0]
  PIN mgmt_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.920 4.000 674.520 ;
    END
  END mgmt_wdata[10]
  PIN mgmt_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 679.360 4.000 679.960 ;
    END
  END mgmt_wdata[11]
  PIN mgmt_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.800 4.000 685.400 ;
    END
  END mgmt_wdata[12]
  PIN mgmt_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.240 4.000 690.840 ;
    END
  END mgmt_wdata[13]
  PIN mgmt_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.000 4.000 695.600 ;
    END
  END mgmt_wdata[14]
  PIN mgmt_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END mgmt_wdata[15]
  PIN mgmt_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 4.000 706.480 ;
    END
  END mgmt_wdata[16]
  PIN mgmt_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 711.320 4.000 711.920 ;
    END
  END mgmt_wdata[17]
  PIN mgmt_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.760 4.000 717.360 ;
    END
  END mgmt_wdata[18]
  PIN mgmt_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.200 4.000 722.800 ;
    END
  END mgmt_wdata[19]
  PIN mgmt_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END mgmt_wdata[1]
  PIN mgmt_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END mgmt_wdata[20]
  PIN mgmt_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 733.080 4.000 733.680 ;
    END
  END mgmt_wdata[21]
  PIN mgmt_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 738.520 4.000 739.120 ;
    END
  END mgmt_wdata[22]
  PIN mgmt_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.960 4.000 744.560 ;
    END
  END mgmt_wdata[23]
  PIN mgmt_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.720 4.000 749.320 ;
    END
  END mgmt_wdata[24]
  PIN mgmt_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.160 4.000 754.760 ;
    END
  END mgmt_wdata[25]
  PIN mgmt_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 759.600 4.000 760.200 ;
    END
  END mgmt_wdata[26]
  PIN mgmt_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END mgmt_wdata[27]
  PIN mgmt_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 770.480 4.000 771.080 ;
    END
  END mgmt_wdata[28]
  PIN mgmt_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.920 4.000 776.520 ;
    END
  END mgmt_wdata[29]
  PIN mgmt_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.080 4.000 631.680 ;
    END
  END mgmt_wdata[2]
  PIN mgmt_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 781.360 4.000 781.960 ;
    END
  END mgmt_wdata[30]
  PIN mgmt_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 786.800 4.000 787.400 ;
    END
  END mgmt_wdata[31]
  PIN mgmt_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END mgmt_wdata[3]
  PIN mgmt_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 641.280 4.000 641.880 ;
    END
  END mgmt_wdata[4]
  PIN mgmt_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.720 4.000 647.320 ;
    END
  END mgmt_wdata[5]
  PIN mgmt_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.160 4.000 652.760 ;
    END
  END mgmt_wdata[6]
  PIN mgmt_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 657.600 4.000 658.200 ;
    END
  END mgmt_wdata[7]
  PIN mgmt_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END mgmt_wdata[8]
  PIN mgmt_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 668.480 4.000 669.080 ;
    END
  END mgmt_wdata[9]
  PIN mgmt_wen[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.240 4.000 792.840 ;
    END
  END mgmt_wen[0]
  PIN mgmt_wen[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.680 4.000 798.280 ;
    END
  END mgmt_wen[1]
  PIN mgmt_wen_mask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 803.120 4.000 803.720 ;
    END
  END mgmt_wen_mask[0]
  PIN mgmt_wen_mask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.880 4.000 808.480 ;
    END
  END mgmt_wen_mask[1]
  PIN mgmt_wen_mask[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 813.320 4.000 813.920 ;
    END
  END mgmt_wen_mask[2]
  PIN mgmt_wen_mask[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 818.760 4.000 819.360 ;
    END
  END mgmt_wen_mask[3]
  PIN mgmt_wen_mask[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 824.200 4.000 824.800 ;
    END
  END mgmt_wen_mask[4]
  PIN mgmt_wen_mask[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END mgmt_wen_mask[5]
  PIN mgmt_wen_mask[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 835.080 4.000 835.680 ;
    END
  END mgmt_wen_mask[6]
  PIN mgmt_wen_mask[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 840.520 4.000 841.120 ;
    END
  END mgmt_wen_mask[7]
  PIN mprj2_vcc_pwrgood
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2102.750 856.000 2103.030 860.000 ;
    END
  END mprj2_vcc_pwrgood
  PIN mprj2_vdd_pwrgood
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2105.970 856.000 2106.250 860.000 ;
    END
  END mprj2_vdd_pwrgood
  PIN mprj_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 856.000 102.030 860.000 ;
    END
  END mprj_ack_i
  PIN mprj_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 856.000 313.170 860.000 ;
    END
  END mprj_adr_o[0]
  PIN mprj_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 856.000 345.830 860.000 ;
    END
  END mprj_adr_o[10]
  PIN mprj_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 856.000 349.050 860.000 ;
    END
  END mprj_adr_o[11]
  PIN mprj_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 856.000 352.270 860.000 ;
    END
  END mprj_adr_o[12]
  PIN mprj_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 856.000 355.490 860.000 ;
    END
  END mprj_adr_o[13]
  PIN mprj_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 856.000 358.710 860.000 ;
    END
  END mprj_adr_o[14]
  PIN mprj_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 856.000 361.930 860.000 ;
    END
  END mprj_adr_o[15]
  PIN mprj_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 856.000 365.150 860.000 ;
    END
  END mprj_adr_o[16]
  PIN mprj_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 856.000 368.370 860.000 ;
    END
  END mprj_adr_o[17]
  PIN mprj_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 856.000 371.590 860.000 ;
    END
  END mprj_adr_o[18]
  PIN mprj_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 856.000 374.810 860.000 ;
    END
  END mprj_adr_o[19]
  PIN mprj_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 856.000 316.390 860.000 ;
    END
  END mprj_adr_o[1]
  PIN mprj_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 856.000 378.490 860.000 ;
    END
  END mprj_adr_o[20]
  PIN mprj_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 856.000 381.710 860.000 ;
    END
  END mprj_adr_o[21]
  PIN mprj_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 856.000 384.930 860.000 ;
    END
  END mprj_adr_o[22]
  PIN mprj_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 856.000 388.150 860.000 ;
    END
  END mprj_adr_o[23]
  PIN mprj_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 856.000 391.370 860.000 ;
    END
  END mprj_adr_o[24]
  PIN mprj_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 856.000 394.590 860.000 ;
    END
  END mprj_adr_o[25]
  PIN mprj_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 856.000 397.810 860.000 ;
    END
  END mprj_adr_o[26]
  PIN mprj_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.750 856.000 401.030 860.000 ;
    END
  END mprj_adr_o[27]
  PIN mprj_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 856.000 404.250 860.000 ;
    END
  END mprj_adr_o[28]
  PIN mprj_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 856.000 407.470 860.000 ;
    END
  END mprj_adr_o[29]
  PIN mprj_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 856.000 319.610 860.000 ;
    END
  END mprj_adr_o[2]
  PIN mprj_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 856.000 410.690 860.000 ;
    END
  END mprj_adr_o[30]
  PIN mprj_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 856.000 413.910 860.000 ;
    END
  END mprj_adr_o[31]
  PIN mprj_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 856.000 322.830 860.000 ;
    END
  END mprj_adr_o[3]
  PIN mprj_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 856.000 326.510 860.000 ;
    END
  END mprj_adr_o[4]
  PIN mprj_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 856.000 329.730 860.000 ;
    END
  END mprj_adr_o[5]
  PIN mprj_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 856.000 332.950 860.000 ;
    END
  END mprj_adr_o[6]
  PIN mprj_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 856.000 336.170 860.000 ;
    END
  END mprj_adr_o[7]
  PIN mprj_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 856.000 339.390 860.000 ;
    END
  END mprj_adr_o[8]
  PIN mprj_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 856.000 342.610 860.000 ;
    END
  END mprj_adr_o[9]
  PIN mprj_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 856.000 433.690 860.000 ;
    END
  END mprj_cyc_o
  PIN mprj_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 856.000 105.250 860.000 ;
    END
  END mprj_dat_i[0]
  PIN mprj_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 856.000 137.910 860.000 ;
    END
  END mprj_dat_i[10]
  PIN mprj_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 856.000 141.130 860.000 ;
    END
  END mprj_dat_i[11]
  PIN mprj_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 856.000 144.350 860.000 ;
    END
  END mprj_dat_i[12]
  PIN mprj_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 856.000 147.570 860.000 ;
    END
  END mprj_dat_i[13]
  PIN mprj_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 856.000 150.790 860.000 ;
    END
  END mprj_dat_i[14]
  PIN mprj_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 856.000 154.010 860.000 ;
    END
  END mprj_dat_i[15]
  PIN mprj_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 856.000 157.230 860.000 ;
    END
  END mprj_dat_i[16]
  PIN mprj_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 856.000 160.450 860.000 ;
    END
  END mprj_dat_i[17]
  PIN mprj_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 856.000 164.130 860.000 ;
    END
  END mprj_dat_i[18]
  PIN mprj_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 856.000 167.350 860.000 ;
    END
  END mprj_dat_i[19]
  PIN mprj_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 856.000 108.470 860.000 ;
    END
  END mprj_dat_i[1]
  PIN mprj_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 856.000 170.570 860.000 ;
    END
  END mprj_dat_i[20]
  PIN mprj_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 856.000 173.790 860.000 ;
    END
  END mprj_dat_i[21]
  PIN mprj_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 856.000 177.010 860.000 ;
    END
  END mprj_dat_i[22]
  PIN mprj_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 856.000 180.230 860.000 ;
    END
  END mprj_dat_i[23]
  PIN mprj_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 856.000 183.450 860.000 ;
    END
  END mprj_dat_i[24]
  PIN mprj_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 856.000 186.670 860.000 ;
    END
  END mprj_dat_i[25]
  PIN mprj_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 856.000 189.890 860.000 ;
    END
  END mprj_dat_i[26]
  PIN mprj_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 856.000 193.110 860.000 ;
    END
  END mprj_dat_i[27]
  PIN mprj_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 856.000 196.330 860.000 ;
    END
  END mprj_dat_i[28]
  PIN mprj_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 856.000 199.550 860.000 ;
    END
  END mprj_dat_i[29]
  PIN mprj_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 856.000 112.150 860.000 ;
    END
  END mprj_dat_i[2]
  PIN mprj_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 856.000 202.770 860.000 ;
    END
  END mprj_dat_i[30]
  PIN mprj_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 856.000 205.990 860.000 ;
    END
  END mprj_dat_i[31]
  PIN mprj_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 856.000 115.370 860.000 ;
    END
  END mprj_dat_i[3]
  PIN mprj_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 856.000 118.590 860.000 ;
    END
  END mprj_dat_i[4]
  PIN mprj_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 856.000 121.810 860.000 ;
    END
  END mprj_dat_i[5]
  PIN mprj_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 856.000 125.030 860.000 ;
    END
  END mprj_dat_i[6]
  PIN mprj_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 856.000 128.250 860.000 ;
    END
  END mprj_dat_i[7]
  PIN mprj_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 856.000 131.470 860.000 ;
    END
  END mprj_dat_i[8]
  PIN mprj_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 856.000 134.690 860.000 ;
    END
  END mprj_dat_i[9]
  PIN mprj_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 856.000 209.210 860.000 ;
    END
  END mprj_dat_o[0]
  PIN mprj_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 856.000 241.870 860.000 ;
    END
  END mprj_dat_o[10]
  PIN mprj_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 856.000 245.090 860.000 ;
    END
  END mprj_dat_o[11]
  PIN mprj_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 856.000 248.310 860.000 ;
    END
  END mprj_dat_o[12]
  PIN mprj_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 856.000 251.530 860.000 ;
    END
  END mprj_dat_o[13]
  PIN mprj_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 856.000 254.750 860.000 ;
    END
  END mprj_dat_o[14]
  PIN mprj_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 856.000 257.970 860.000 ;
    END
  END mprj_dat_o[15]
  PIN mprj_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 856.000 261.190 860.000 ;
    END
  END mprj_dat_o[16]
  PIN mprj_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 856.000 264.410 860.000 ;
    END
  END mprj_dat_o[17]
  PIN mprj_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 856.000 267.630 860.000 ;
    END
  END mprj_dat_o[18]
  PIN mprj_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 856.000 271.310 860.000 ;
    END
  END mprj_dat_o[19]
  PIN mprj_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 856.000 212.430 860.000 ;
    END
  END mprj_dat_o[1]
  PIN mprj_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 856.000 274.530 860.000 ;
    END
  END mprj_dat_o[20]
  PIN mprj_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 856.000 277.750 860.000 ;
    END
  END mprj_dat_o[21]
  PIN mprj_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 856.000 280.970 860.000 ;
    END
  END mprj_dat_o[22]
  PIN mprj_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 856.000 284.190 860.000 ;
    END
  END mprj_dat_o[23]
  PIN mprj_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 856.000 287.410 860.000 ;
    END
  END mprj_dat_o[24]
  PIN mprj_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 856.000 290.630 860.000 ;
    END
  END mprj_dat_o[25]
  PIN mprj_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 856.000 293.850 860.000 ;
    END
  END mprj_dat_o[26]
  PIN mprj_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 856.000 297.070 860.000 ;
    END
  END mprj_dat_o[27]
  PIN mprj_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 856.000 300.290 860.000 ;
    END
  END mprj_dat_o[28]
  PIN mprj_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 856.000 303.510 860.000 ;
    END
  END mprj_dat_o[29]
  PIN mprj_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 856.000 215.650 860.000 ;
    END
  END mprj_dat_o[2]
  PIN mprj_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 856.000 306.730 860.000 ;
    END
  END mprj_dat_o[30]
  PIN mprj_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 856.000 309.950 860.000 ;
    END
  END mprj_dat_o[31]
  PIN mprj_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 856.000 219.330 860.000 ;
    END
  END mprj_dat_o[3]
  PIN mprj_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 856.000 222.550 860.000 ;
    END
  END mprj_dat_o[4]
  PIN mprj_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 856.000 225.770 860.000 ;
    END
  END mprj_dat_o[5]
  PIN mprj_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 856.000 228.990 860.000 ;
    END
  END mprj_dat_o[6]
  PIN mprj_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 856.000 232.210 860.000 ;
    END
  END mprj_dat_o[7]
  PIN mprj_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 856.000 235.430 860.000 ;
    END
  END mprj_dat_o[8]
  PIN mprj_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 856.000 238.650 860.000 ;
    END
  END mprj_dat_o[9]
  PIN mprj_io_loader_clock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 352.280 2150.000 352.880 ;
    END
  END mprj_io_loader_clock
  PIN mprj_io_loader_data_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2147.830 856.000 2148.110 860.000 ;
    END
  END mprj_io_loader_data_1
  PIN mprj_io_loader_data_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END mprj_io_loader_data_2
  PIN mprj_io_loader_resetn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 342.760 2150.000 343.360 ;
    END
  END mprj_io_loader_resetn
  PIN mprj_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 856.000 417.130 860.000 ;
    END
  END mprj_sel_o[0]
  PIN mprj_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.070 856.000 420.350 860.000 ;
    END
  END mprj_sel_o[1]
  PIN mprj_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 856.000 423.570 860.000 ;
    END
  END mprj_sel_o[2]
  PIN mprj_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 856.000 426.790 860.000 ;
    END
  END mprj_sel_o[3]
  PIN mprj_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 856.000 430.010 860.000 ;
    END
  END mprj_stb_o
  PIN mprj_vcc_pwrgood
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2109.190 856.000 2109.470 860.000 ;
    END
  END mprj_vcc_pwrgood
  PIN mprj_vdd_pwrgood
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.410 856.000 2112.690 860.000 ;
    END
  END mprj_vdd_pwrgood
  PIN mprj_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 856.000 436.910 860.000 ;
    END
  END mprj_we_o
  PIN porb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 313.520 2150.000 314.120 ;
    END
  END porb
  PIN pwr_ctrl_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2115.630 856.000 2115.910 860.000 ;
    END
  END pwr_ctrl_out[0]
  PIN pwr_ctrl_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.850 856.000 2119.130 860.000 ;
    END
  END pwr_ctrl_out[1]
  PIN pwr_ctrl_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2122.070 856.000 2122.350 860.000 ;
    END
  END pwr_ctrl_out[2]
  PIN pwr_ctrl_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2125.290 856.000 2125.570 860.000 ;
    END
  END pwr_ctrl_out[3]
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END resetb
  PIN sdo_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 361.800 2150.000 362.400 ;
    END
  END sdo_out
  PIN sdo_outenb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2146.000 372.000 2150.000 372.600 ;
    END
  END sdo_outenb
  PIN user_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 856.000 8.190 860.000 ;
    END
  END user_clk
  PIN user_irq[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2128.510 856.000 2128.790 860.000 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2131.730 856.000 2132.010 860.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2134.950 856.000 2135.230 860.000 ;
    END
  END user_irq[2]
  PIN user_irq_ena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2138.170 856.000 2138.450 860.000 ;
    END
  END user_irq_ena[0]
  PIN user_irq_ena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2141.390 856.000 2141.670 860.000 ;
    END
  END user_irq_ena[1]
  PIN user_irq_ena[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2144.610 856.000 2144.890 860.000 ;
    END
  END user_irq_ena[2]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2121.040 10.640 2122.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2071.040 10.640 2072.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2021.040 10.640 2022.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1971.040 821.480 1972.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1921.040 10.640 1922.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1871.040 10.640 1872.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1821.040 10.640 1822.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1771.040 10.640 1772.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1721.040 10.640 1722.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1671.040 10.640 1672.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1621.040 10.640 1622.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1571.040 10.640 1572.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1521.040 10.640 1522.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1471.040 10.640 1472.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1421.040 10.640 1422.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1371.040 10.640 1372.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1321.040 10.640 1322.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1271.040 10.640 1272.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1221.040 10.640 1222.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1171.040 10.640 1172.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1121.040 10.640 1122.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1071.040 10.640 1072.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1021.040 10.640 1022.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 971.040 10.640 972.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 921.040 10.640 922.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 871.040 640.760 872.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 821.040 640.760 822.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 771.040 640.760 772.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 721.040 640.760 722.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 671.040 640.760 672.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 621.040 640.760 622.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 571.040 640.760 572.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 521.040 640.760 522.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 471.040 640.760 472.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 421.040 640.760 422.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 371.040 640.760 372.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 321.040 640.760 322.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 271.040 640.760 272.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 221.040 640.760 222.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 171.040 640.760 172.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 121.040 640.760 122.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 71.040 10.640 72.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 848.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1971.040 10.640 1972.640 726.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 871.040 10.640 872.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 821.040 10.640 822.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 771.040 10.640 772.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 721.040 10.640 722.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 671.040 10.640 672.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 621.040 10.640 622.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 571.040 10.640 572.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 521.040 10.640 522.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 421.040 10.640 422.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 371.040 10.640 372.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 271.040 10.640 272.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 221.040 10.640 222.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 121.040 10.640 122.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 806.490 2144.060 808.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 676.490 2144.060 678.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 546.490 2144.060 548.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 416.490 2144.060 418.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 286.490 2144.060 288.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 156.490 2144.060 158.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 2144.060 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2096.040 10.640 2097.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2046.040 10.640 2047.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1996.040 821.480 1997.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1946.040 821.480 1947.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1896.040 10.640 1897.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1846.040 10.640 1847.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1796.040 10.640 1797.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1746.040 10.640 1747.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1696.040 10.640 1697.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1646.040 10.640 1647.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1596.040 10.640 1597.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1546.040 10.640 1547.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1496.040 10.640 1497.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1446.040 10.640 1447.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1396.040 10.640 1397.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1346.040 10.640 1347.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1296.040 10.640 1297.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1246.040 10.640 1247.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1196.040 10.640 1197.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1146.040 10.640 1147.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1096.040 10.640 1097.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1046.040 10.640 1047.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 996.040 10.640 997.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 946.040 10.640 947.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 896.040 10.640 897.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 846.040 640.760 847.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 796.040 640.760 797.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 746.040 640.760 747.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 696.040 640.760 697.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 646.040 640.760 647.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 596.040 640.760 597.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 546.040 640.760 547.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 496.040 640.760 497.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 446.040 640.760 447.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 396.040 640.760 397.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 346.040 640.760 347.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 296.040 640.760 297.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 246.040 640.760 247.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 196.040 640.760 197.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 146.040 640.760 147.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.040 10.640 97.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 46.040 10.640 47.640 848.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1996.040 10.640 1997.640 726.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1946.040 10.640 1947.640 726.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 846.040 10.640 847.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 796.040 10.640 797.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 746.040 10.640 747.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 696.040 10.640 697.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 646.040 10.640 647.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 596.040 10.640 597.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 546.040 10.640 547.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 496.040 10.640 497.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 446.040 10.640 447.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 396.040 10.640 397.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 346.040 10.640 347.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 296.040 10.640 297.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 246.040 10.640 247.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 196.040 10.640 197.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 146.040 10.640 147.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 741.490 2144.060 743.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 611.490 2144.060 613.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 481.490 2144.060 483.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 351.490 2144.060 353.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 221.490 2144.060 223.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 91.490 2144.060 93.090 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 6.545 2144.835 858.415 ;
      LAYER met1 ;
        RECT 1.450 6.500 2148.130 859.820 ;
      LAYER met2 ;
        RECT 2.030 855.720 4.410 859.850 ;
        RECT 5.250 855.720 7.630 859.850 ;
        RECT 8.470 855.720 10.850 859.850 ;
        RECT 11.690 855.720 14.070 859.850 ;
        RECT 14.910 855.720 17.290 859.850 ;
        RECT 18.130 855.720 20.510 859.850 ;
        RECT 21.350 855.720 23.730 859.850 ;
        RECT 24.570 855.720 26.950 859.850 ;
        RECT 27.790 855.720 30.170 859.850 ;
        RECT 31.010 855.720 33.390 859.850 ;
        RECT 34.230 855.720 36.610 859.850 ;
        RECT 37.450 855.720 39.830 859.850 ;
        RECT 40.670 855.720 43.050 859.850 ;
        RECT 43.890 855.720 46.270 859.850 ;
        RECT 47.110 855.720 49.490 859.850 ;
        RECT 50.330 855.720 52.710 859.850 ;
        RECT 53.550 855.720 56.390 859.850 ;
        RECT 57.230 855.720 59.610 859.850 ;
        RECT 60.450 855.720 62.830 859.850 ;
        RECT 63.670 855.720 66.050 859.850 ;
        RECT 66.890 855.720 69.270 859.850 ;
        RECT 70.110 855.720 72.490 859.850 ;
        RECT 73.330 855.720 75.710 859.850 ;
        RECT 76.550 855.720 78.930 859.850 ;
        RECT 79.770 855.720 82.150 859.850 ;
        RECT 82.990 855.720 85.370 859.850 ;
        RECT 86.210 855.720 88.590 859.850 ;
        RECT 89.430 855.720 91.810 859.850 ;
        RECT 92.650 855.720 95.030 859.850 ;
        RECT 95.870 855.720 98.250 859.850 ;
        RECT 99.090 855.720 101.470 859.850 ;
        RECT 102.310 855.720 104.690 859.850 ;
        RECT 105.530 855.720 107.910 859.850 ;
        RECT 108.750 855.720 111.590 859.850 ;
        RECT 112.430 855.720 114.810 859.850 ;
        RECT 115.650 855.720 118.030 859.850 ;
        RECT 118.870 855.720 121.250 859.850 ;
        RECT 122.090 855.720 124.470 859.850 ;
        RECT 125.310 855.720 127.690 859.850 ;
        RECT 128.530 855.720 130.910 859.850 ;
        RECT 131.750 855.720 134.130 859.850 ;
        RECT 134.970 855.720 137.350 859.850 ;
        RECT 138.190 855.720 140.570 859.850 ;
        RECT 141.410 855.720 143.790 859.850 ;
        RECT 144.630 855.720 147.010 859.850 ;
        RECT 147.850 855.720 150.230 859.850 ;
        RECT 151.070 855.720 153.450 859.850 ;
        RECT 154.290 855.720 156.670 859.850 ;
        RECT 157.510 855.720 159.890 859.850 ;
        RECT 160.730 855.720 163.570 859.850 ;
        RECT 164.410 855.720 166.790 859.850 ;
        RECT 167.630 855.720 170.010 859.850 ;
        RECT 170.850 855.720 173.230 859.850 ;
        RECT 174.070 855.720 176.450 859.850 ;
        RECT 177.290 855.720 179.670 859.850 ;
        RECT 180.510 855.720 182.890 859.850 ;
        RECT 183.730 855.720 186.110 859.850 ;
        RECT 186.950 855.720 189.330 859.850 ;
        RECT 190.170 855.720 192.550 859.850 ;
        RECT 193.390 855.720 195.770 859.850 ;
        RECT 196.610 855.720 198.990 859.850 ;
        RECT 199.830 855.720 202.210 859.850 ;
        RECT 203.050 855.720 205.430 859.850 ;
        RECT 206.270 855.720 208.650 859.850 ;
        RECT 209.490 855.720 211.870 859.850 ;
        RECT 212.710 855.720 215.090 859.850 ;
        RECT 215.930 855.720 218.770 859.850 ;
        RECT 219.610 855.720 221.990 859.850 ;
        RECT 222.830 855.720 225.210 859.850 ;
        RECT 226.050 855.720 228.430 859.850 ;
        RECT 229.270 855.720 231.650 859.850 ;
        RECT 232.490 855.720 234.870 859.850 ;
        RECT 235.710 855.720 238.090 859.850 ;
        RECT 238.930 855.720 241.310 859.850 ;
        RECT 242.150 855.720 244.530 859.850 ;
        RECT 245.370 855.720 247.750 859.850 ;
        RECT 248.590 855.720 250.970 859.850 ;
        RECT 251.810 855.720 254.190 859.850 ;
        RECT 255.030 855.720 257.410 859.850 ;
        RECT 258.250 855.720 260.630 859.850 ;
        RECT 261.470 855.720 263.850 859.850 ;
        RECT 264.690 855.720 267.070 859.850 ;
        RECT 267.910 855.720 270.750 859.850 ;
        RECT 271.590 855.720 273.970 859.850 ;
        RECT 274.810 855.720 277.190 859.850 ;
        RECT 278.030 855.720 280.410 859.850 ;
        RECT 281.250 855.720 283.630 859.850 ;
        RECT 284.470 855.720 286.850 859.850 ;
        RECT 287.690 855.720 290.070 859.850 ;
        RECT 290.910 855.720 293.290 859.850 ;
        RECT 294.130 855.720 296.510 859.850 ;
        RECT 297.350 855.720 299.730 859.850 ;
        RECT 300.570 855.720 302.950 859.850 ;
        RECT 303.790 855.720 306.170 859.850 ;
        RECT 307.010 855.720 309.390 859.850 ;
        RECT 310.230 855.720 312.610 859.850 ;
        RECT 313.450 855.720 315.830 859.850 ;
        RECT 316.670 855.720 319.050 859.850 ;
        RECT 319.890 855.720 322.270 859.850 ;
        RECT 323.110 855.720 325.950 859.850 ;
        RECT 326.790 855.720 329.170 859.850 ;
        RECT 330.010 855.720 332.390 859.850 ;
        RECT 333.230 855.720 335.610 859.850 ;
        RECT 336.450 855.720 338.830 859.850 ;
        RECT 339.670 855.720 342.050 859.850 ;
        RECT 342.890 855.720 345.270 859.850 ;
        RECT 346.110 855.720 348.490 859.850 ;
        RECT 349.330 855.720 351.710 859.850 ;
        RECT 352.550 855.720 354.930 859.850 ;
        RECT 355.770 855.720 358.150 859.850 ;
        RECT 358.990 855.720 361.370 859.850 ;
        RECT 362.210 855.720 364.590 859.850 ;
        RECT 365.430 855.720 367.810 859.850 ;
        RECT 368.650 855.720 371.030 859.850 ;
        RECT 371.870 855.720 374.250 859.850 ;
        RECT 375.090 855.720 377.930 859.850 ;
        RECT 378.770 855.720 381.150 859.850 ;
        RECT 381.990 855.720 384.370 859.850 ;
        RECT 385.210 855.720 387.590 859.850 ;
        RECT 388.430 855.720 390.810 859.850 ;
        RECT 391.650 855.720 394.030 859.850 ;
        RECT 394.870 855.720 397.250 859.850 ;
        RECT 398.090 855.720 400.470 859.850 ;
        RECT 401.310 855.720 403.690 859.850 ;
        RECT 404.530 855.720 406.910 859.850 ;
        RECT 407.750 855.720 410.130 859.850 ;
        RECT 410.970 855.720 413.350 859.850 ;
        RECT 414.190 855.720 416.570 859.850 ;
        RECT 417.410 855.720 419.790 859.850 ;
        RECT 420.630 855.720 423.010 859.850 ;
        RECT 423.850 855.720 426.230 859.850 ;
        RECT 427.070 855.720 429.450 859.850 ;
        RECT 430.290 855.720 433.130 859.850 ;
        RECT 433.970 855.720 436.350 859.850 ;
        RECT 437.190 855.720 439.570 859.850 ;
        RECT 440.410 855.720 442.790 859.850 ;
        RECT 443.630 855.720 446.010 859.850 ;
        RECT 446.850 855.720 449.230 859.850 ;
        RECT 450.070 855.720 452.450 859.850 ;
        RECT 453.290 855.720 455.670 859.850 ;
        RECT 456.510 855.720 458.890 859.850 ;
        RECT 459.730 855.720 462.110 859.850 ;
        RECT 462.950 855.720 465.330 859.850 ;
        RECT 466.170 855.720 468.550 859.850 ;
        RECT 469.390 855.720 471.770 859.850 ;
        RECT 472.610 855.720 474.990 859.850 ;
        RECT 475.830 855.720 478.210 859.850 ;
        RECT 479.050 855.720 481.430 859.850 ;
        RECT 482.270 855.720 485.110 859.850 ;
        RECT 485.950 855.720 488.330 859.850 ;
        RECT 489.170 855.720 491.550 859.850 ;
        RECT 492.390 855.720 494.770 859.850 ;
        RECT 495.610 855.720 497.990 859.850 ;
        RECT 498.830 855.720 501.210 859.850 ;
        RECT 502.050 855.720 504.430 859.850 ;
        RECT 505.270 855.720 507.650 859.850 ;
        RECT 508.490 855.720 510.870 859.850 ;
        RECT 511.710 855.720 514.090 859.850 ;
        RECT 514.930 855.720 517.310 859.850 ;
        RECT 518.150 855.720 520.530 859.850 ;
        RECT 521.370 855.720 523.750 859.850 ;
        RECT 524.590 855.720 526.970 859.850 ;
        RECT 527.810 855.720 530.190 859.850 ;
        RECT 531.030 855.720 533.410 859.850 ;
        RECT 534.250 855.720 536.630 859.850 ;
        RECT 537.470 855.720 540.310 859.850 ;
        RECT 541.150 855.720 543.530 859.850 ;
        RECT 544.370 855.720 546.750 859.850 ;
        RECT 547.590 855.720 549.970 859.850 ;
        RECT 550.810 855.720 553.190 859.850 ;
        RECT 554.030 855.720 556.410 859.850 ;
        RECT 557.250 855.720 559.630 859.850 ;
        RECT 560.470 855.720 562.850 859.850 ;
        RECT 563.690 855.720 566.070 859.850 ;
        RECT 566.910 855.720 569.290 859.850 ;
        RECT 570.130 855.720 572.510 859.850 ;
        RECT 573.350 855.720 575.730 859.850 ;
        RECT 576.570 855.720 578.950 859.850 ;
        RECT 579.790 855.720 582.170 859.850 ;
        RECT 583.010 855.720 585.390 859.850 ;
        RECT 586.230 855.720 588.610 859.850 ;
        RECT 589.450 855.720 591.830 859.850 ;
        RECT 592.670 855.720 595.510 859.850 ;
        RECT 596.350 855.720 598.730 859.850 ;
        RECT 599.570 855.720 601.950 859.850 ;
        RECT 602.790 855.720 605.170 859.850 ;
        RECT 606.010 855.720 608.390 859.850 ;
        RECT 609.230 855.720 611.610 859.850 ;
        RECT 612.450 855.720 614.830 859.850 ;
        RECT 615.670 855.720 618.050 859.850 ;
        RECT 618.890 855.720 621.270 859.850 ;
        RECT 622.110 855.720 624.490 859.850 ;
        RECT 625.330 855.720 627.710 859.850 ;
        RECT 628.550 855.720 630.930 859.850 ;
        RECT 631.770 855.720 634.150 859.850 ;
        RECT 634.990 855.720 637.370 859.850 ;
        RECT 638.210 855.720 640.590 859.850 ;
        RECT 641.430 855.720 643.810 859.850 ;
        RECT 644.650 855.720 647.490 859.850 ;
        RECT 648.330 855.720 650.710 859.850 ;
        RECT 651.550 855.720 653.930 859.850 ;
        RECT 654.770 855.720 657.150 859.850 ;
        RECT 657.990 855.720 660.370 859.850 ;
        RECT 661.210 855.720 663.590 859.850 ;
        RECT 664.430 855.720 666.810 859.850 ;
        RECT 667.650 855.720 670.030 859.850 ;
        RECT 670.870 855.720 673.250 859.850 ;
        RECT 674.090 855.720 676.470 859.850 ;
        RECT 677.310 855.720 679.690 859.850 ;
        RECT 680.530 855.720 682.910 859.850 ;
        RECT 683.750 855.720 686.130 859.850 ;
        RECT 686.970 855.720 689.350 859.850 ;
        RECT 690.190 855.720 692.570 859.850 ;
        RECT 693.410 855.720 695.790 859.850 ;
        RECT 696.630 855.720 699.010 859.850 ;
        RECT 699.850 855.720 702.690 859.850 ;
        RECT 703.530 855.720 705.910 859.850 ;
        RECT 706.750 855.720 709.130 859.850 ;
        RECT 709.970 855.720 712.350 859.850 ;
        RECT 713.190 855.720 715.570 859.850 ;
        RECT 716.410 855.720 718.790 859.850 ;
        RECT 719.630 855.720 722.010 859.850 ;
        RECT 722.850 855.720 725.230 859.850 ;
        RECT 726.070 855.720 728.450 859.850 ;
        RECT 729.290 855.720 731.670 859.850 ;
        RECT 732.510 855.720 734.890 859.850 ;
        RECT 735.730 855.720 738.110 859.850 ;
        RECT 738.950 855.720 741.330 859.850 ;
        RECT 742.170 855.720 744.550 859.850 ;
        RECT 745.390 855.720 747.770 859.850 ;
        RECT 748.610 855.720 750.990 859.850 ;
        RECT 751.830 855.720 754.670 859.850 ;
        RECT 755.510 855.720 757.890 859.850 ;
        RECT 758.730 855.720 761.110 859.850 ;
        RECT 761.950 855.720 764.330 859.850 ;
        RECT 765.170 855.720 767.550 859.850 ;
        RECT 768.390 855.720 770.770 859.850 ;
        RECT 771.610 855.720 773.990 859.850 ;
        RECT 774.830 855.720 777.210 859.850 ;
        RECT 778.050 855.720 780.430 859.850 ;
        RECT 781.270 855.720 783.650 859.850 ;
        RECT 784.490 855.720 786.870 859.850 ;
        RECT 787.710 855.720 790.090 859.850 ;
        RECT 790.930 855.720 793.310 859.850 ;
        RECT 794.150 855.720 796.530 859.850 ;
        RECT 797.370 855.720 799.750 859.850 ;
        RECT 800.590 855.720 802.970 859.850 ;
        RECT 803.810 855.720 806.190 859.850 ;
        RECT 807.030 855.720 809.870 859.850 ;
        RECT 810.710 855.720 813.090 859.850 ;
        RECT 813.930 855.720 816.310 859.850 ;
        RECT 817.150 855.720 819.530 859.850 ;
        RECT 820.370 855.720 822.750 859.850 ;
        RECT 823.590 855.720 825.970 859.850 ;
        RECT 826.810 855.720 829.190 859.850 ;
        RECT 830.030 855.720 832.410 859.850 ;
        RECT 833.250 855.720 835.630 859.850 ;
        RECT 836.470 855.720 838.850 859.850 ;
        RECT 839.690 855.720 842.070 859.850 ;
        RECT 842.910 855.720 845.290 859.850 ;
        RECT 846.130 855.720 848.510 859.850 ;
        RECT 849.350 855.720 851.730 859.850 ;
        RECT 852.570 855.720 854.950 859.850 ;
        RECT 855.790 855.720 858.170 859.850 ;
        RECT 859.010 855.720 861.850 859.850 ;
        RECT 862.690 855.720 865.070 859.850 ;
        RECT 865.910 855.720 868.290 859.850 ;
        RECT 869.130 855.720 871.510 859.850 ;
        RECT 872.350 855.720 874.730 859.850 ;
        RECT 875.570 855.720 877.950 859.850 ;
        RECT 878.790 855.720 881.170 859.850 ;
        RECT 882.010 855.720 884.390 859.850 ;
        RECT 885.230 855.720 887.610 859.850 ;
        RECT 888.450 855.720 890.830 859.850 ;
        RECT 891.670 855.720 894.050 859.850 ;
        RECT 894.890 855.720 897.270 859.850 ;
        RECT 898.110 855.720 900.490 859.850 ;
        RECT 901.330 855.720 903.710 859.850 ;
        RECT 904.550 855.720 906.930 859.850 ;
        RECT 907.770 855.720 910.150 859.850 ;
        RECT 910.990 855.720 913.370 859.850 ;
        RECT 914.210 855.720 917.050 859.850 ;
        RECT 917.890 855.720 920.270 859.850 ;
        RECT 921.110 855.720 923.490 859.850 ;
        RECT 924.330 855.720 926.710 859.850 ;
        RECT 927.550 855.720 929.930 859.850 ;
        RECT 930.770 855.720 933.150 859.850 ;
        RECT 933.990 855.720 936.370 859.850 ;
        RECT 937.210 855.720 939.590 859.850 ;
        RECT 940.430 855.720 942.810 859.850 ;
        RECT 943.650 855.720 946.030 859.850 ;
        RECT 946.870 855.720 949.250 859.850 ;
        RECT 950.090 855.720 952.470 859.850 ;
        RECT 953.310 855.720 955.690 859.850 ;
        RECT 956.530 855.720 958.910 859.850 ;
        RECT 959.750 855.720 962.130 859.850 ;
        RECT 962.970 855.720 965.350 859.850 ;
        RECT 966.190 855.720 969.030 859.850 ;
        RECT 969.870 855.720 972.250 859.850 ;
        RECT 973.090 855.720 975.470 859.850 ;
        RECT 976.310 855.720 978.690 859.850 ;
        RECT 979.530 855.720 981.910 859.850 ;
        RECT 982.750 855.720 985.130 859.850 ;
        RECT 985.970 855.720 988.350 859.850 ;
        RECT 989.190 855.720 991.570 859.850 ;
        RECT 992.410 855.720 994.790 859.850 ;
        RECT 995.630 855.720 998.010 859.850 ;
        RECT 998.850 855.720 1001.230 859.850 ;
        RECT 1002.070 855.720 1004.450 859.850 ;
        RECT 1005.290 855.720 1007.670 859.850 ;
        RECT 1008.510 855.720 1010.890 859.850 ;
        RECT 1011.730 855.720 1014.110 859.850 ;
        RECT 1014.950 855.720 1017.330 859.850 ;
        RECT 1018.170 855.720 1020.550 859.850 ;
        RECT 1021.390 855.720 1024.230 859.850 ;
        RECT 1025.070 855.720 1027.450 859.850 ;
        RECT 1028.290 855.720 1030.670 859.850 ;
        RECT 1031.510 855.720 1033.890 859.850 ;
        RECT 1034.730 855.720 1037.110 859.850 ;
        RECT 1037.950 855.720 1040.330 859.850 ;
        RECT 1041.170 855.720 1043.550 859.850 ;
        RECT 1044.390 855.720 1046.770 859.850 ;
        RECT 1047.610 855.720 1049.990 859.850 ;
        RECT 1050.830 855.720 1053.210 859.850 ;
        RECT 1054.050 855.720 1056.430 859.850 ;
        RECT 1057.270 855.720 1059.650 859.850 ;
        RECT 1060.490 855.720 1062.870 859.850 ;
        RECT 1063.710 855.720 1066.090 859.850 ;
        RECT 1066.930 855.720 1069.310 859.850 ;
        RECT 1070.150 855.720 1072.530 859.850 ;
        RECT 1073.370 855.720 1076.210 859.850 ;
        RECT 1077.050 855.720 1079.430 859.850 ;
        RECT 1080.270 855.720 1082.650 859.850 ;
        RECT 1083.490 855.720 1085.870 859.850 ;
        RECT 1086.710 855.720 1089.090 859.850 ;
        RECT 1089.930 855.720 1092.310 859.850 ;
        RECT 1093.150 855.720 1095.530 859.850 ;
        RECT 1096.370 855.720 1098.750 859.850 ;
        RECT 1099.590 855.720 1101.970 859.850 ;
        RECT 1102.810 855.720 1105.190 859.850 ;
        RECT 1106.030 855.720 1108.410 859.850 ;
        RECT 1109.250 855.720 1111.630 859.850 ;
        RECT 1112.470 855.720 1114.850 859.850 ;
        RECT 1115.690 855.720 1118.070 859.850 ;
        RECT 1118.910 855.720 1121.290 859.850 ;
        RECT 1122.130 855.720 1124.510 859.850 ;
        RECT 1125.350 855.720 1127.730 859.850 ;
        RECT 1128.570 855.720 1131.410 859.850 ;
        RECT 1132.250 855.720 1134.630 859.850 ;
        RECT 1135.470 855.720 1137.850 859.850 ;
        RECT 1138.690 855.720 1141.070 859.850 ;
        RECT 1141.910 855.720 1144.290 859.850 ;
        RECT 1145.130 855.720 1147.510 859.850 ;
        RECT 1148.350 855.720 1150.730 859.850 ;
        RECT 1151.570 855.720 1153.950 859.850 ;
        RECT 1154.790 855.720 1157.170 859.850 ;
        RECT 1158.010 855.720 1160.390 859.850 ;
        RECT 1161.230 855.720 1163.610 859.850 ;
        RECT 1164.450 855.720 1166.830 859.850 ;
        RECT 1167.670 855.720 1170.050 859.850 ;
        RECT 1170.890 855.720 1173.270 859.850 ;
        RECT 1174.110 855.720 1176.490 859.850 ;
        RECT 1177.330 855.720 1179.710 859.850 ;
        RECT 1180.550 855.720 1182.930 859.850 ;
        RECT 1183.770 855.720 1186.610 859.850 ;
        RECT 1187.450 855.720 1189.830 859.850 ;
        RECT 1190.670 855.720 1193.050 859.850 ;
        RECT 1193.890 855.720 1196.270 859.850 ;
        RECT 1197.110 855.720 1199.490 859.850 ;
        RECT 1200.330 855.720 1202.710 859.850 ;
        RECT 1203.550 855.720 1205.930 859.850 ;
        RECT 1206.770 855.720 1209.150 859.850 ;
        RECT 1209.990 855.720 1212.370 859.850 ;
        RECT 1213.210 855.720 1215.590 859.850 ;
        RECT 1216.430 855.720 1218.810 859.850 ;
        RECT 1219.650 855.720 1222.030 859.850 ;
        RECT 1222.870 855.720 1225.250 859.850 ;
        RECT 1226.090 855.720 1228.470 859.850 ;
        RECT 1229.310 855.720 1231.690 859.850 ;
        RECT 1232.530 855.720 1234.910 859.850 ;
        RECT 1235.750 855.720 1238.590 859.850 ;
        RECT 1239.430 855.720 1241.810 859.850 ;
        RECT 1242.650 855.720 1245.030 859.850 ;
        RECT 1245.870 855.720 1248.250 859.850 ;
        RECT 1249.090 855.720 1251.470 859.850 ;
        RECT 1252.310 855.720 1254.690 859.850 ;
        RECT 1255.530 855.720 1257.910 859.850 ;
        RECT 1258.750 855.720 1261.130 859.850 ;
        RECT 1261.970 855.720 1264.350 859.850 ;
        RECT 1265.190 855.720 1267.570 859.850 ;
        RECT 1268.410 855.720 1270.790 859.850 ;
        RECT 1271.630 855.720 1274.010 859.850 ;
        RECT 1274.850 855.720 1277.230 859.850 ;
        RECT 1278.070 855.720 1280.450 859.850 ;
        RECT 1281.290 855.720 1283.670 859.850 ;
        RECT 1284.510 855.720 1286.890 859.850 ;
        RECT 1287.730 855.720 1290.110 859.850 ;
        RECT 1290.950 855.720 1293.790 859.850 ;
        RECT 1294.630 855.720 1297.010 859.850 ;
        RECT 1297.850 855.720 1300.230 859.850 ;
        RECT 1301.070 855.720 1303.450 859.850 ;
        RECT 1304.290 855.720 1306.670 859.850 ;
        RECT 1307.510 855.720 1309.890 859.850 ;
        RECT 1310.730 855.720 1313.110 859.850 ;
        RECT 1313.950 855.720 1316.330 859.850 ;
        RECT 1317.170 855.720 1319.550 859.850 ;
        RECT 1320.390 855.720 1322.770 859.850 ;
        RECT 1323.610 855.720 1325.990 859.850 ;
        RECT 1326.830 855.720 1329.210 859.850 ;
        RECT 1330.050 855.720 1332.430 859.850 ;
        RECT 1333.270 855.720 1335.650 859.850 ;
        RECT 1336.490 855.720 1338.870 859.850 ;
        RECT 1339.710 855.720 1342.090 859.850 ;
        RECT 1342.930 855.720 1345.770 859.850 ;
        RECT 1346.610 855.720 1348.990 859.850 ;
        RECT 1349.830 855.720 1352.210 859.850 ;
        RECT 1353.050 855.720 1355.430 859.850 ;
        RECT 1356.270 855.720 1358.650 859.850 ;
        RECT 1359.490 855.720 1361.870 859.850 ;
        RECT 1362.710 855.720 1365.090 859.850 ;
        RECT 1365.930 855.720 1368.310 859.850 ;
        RECT 1369.150 855.720 1371.530 859.850 ;
        RECT 1372.370 855.720 1374.750 859.850 ;
        RECT 1375.590 855.720 1377.970 859.850 ;
        RECT 1378.810 855.720 1381.190 859.850 ;
        RECT 1382.030 855.720 1384.410 859.850 ;
        RECT 1385.250 855.720 1387.630 859.850 ;
        RECT 1388.470 855.720 1390.850 859.850 ;
        RECT 1391.690 855.720 1394.070 859.850 ;
        RECT 1394.910 855.720 1397.290 859.850 ;
        RECT 1398.130 855.720 1400.970 859.850 ;
        RECT 1401.810 855.720 1404.190 859.850 ;
        RECT 1405.030 855.720 1407.410 859.850 ;
        RECT 1408.250 855.720 1410.630 859.850 ;
        RECT 1411.470 855.720 1413.850 859.850 ;
        RECT 1414.690 855.720 1417.070 859.850 ;
        RECT 1417.910 855.720 1420.290 859.850 ;
        RECT 1421.130 855.720 1423.510 859.850 ;
        RECT 1424.350 855.720 1426.730 859.850 ;
        RECT 1427.570 855.720 1429.950 859.850 ;
        RECT 1430.790 855.720 1433.170 859.850 ;
        RECT 1434.010 855.720 1436.390 859.850 ;
        RECT 1437.230 855.720 1439.610 859.850 ;
        RECT 1440.450 855.720 1442.830 859.850 ;
        RECT 1443.670 855.720 1446.050 859.850 ;
        RECT 1446.890 855.720 1449.270 859.850 ;
        RECT 1450.110 855.720 1452.950 859.850 ;
        RECT 1453.790 855.720 1456.170 859.850 ;
        RECT 1457.010 855.720 1459.390 859.850 ;
        RECT 1460.230 855.720 1462.610 859.850 ;
        RECT 1463.450 855.720 1465.830 859.850 ;
        RECT 1466.670 855.720 1469.050 859.850 ;
        RECT 1469.890 855.720 1472.270 859.850 ;
        RECT 1473.110 855.720 1475.490 859.850 ;
        RECT 1476.330 855.720 1478.710 859.850 ;
        RECT 1479.550 855.720 1481.930 859.850 ;
        RECT 1482.770 855.720 1485.150 859.850 ;
        RECT 1485.990 855.720 1488.370 859.850 ;
        RECT 1489.210 855.720 1491.590 859.850 ;
        RECT 1492.430 855.720 1494.810 859.850 ;
        RECT 1495.650 855.720 1498.030 859.850 ;
        RECT 1498.870 855.720 1501.250 859.850 ;
        RECT 1502.090 855.720 1504.470 859.850 ;
        RECT 1505.310 855.720 1508.150 859.850 ;
        RECT 1508.990 855.720 1511.370 859.850 ;
        RECT 1512.210 855.720 1514.590 859.850 ;
        RECT 1515.430 855.720 1517.810 859.850 ;
        RECT 1518.650 855.720 1521.030 859.850 ;
        RECT 1521.870 855.720 1524.250 859.850 ;
        RECT 1525.090 855.720 1527.470 859.850 ;
        RECT 1528.310 855.720 1530.690 859.850 ;
        RECT 1531.530 855.720 1533.910 859.850 ;
        RECT 1534.750 855.720 1537.130 859.850 ;
        RECT 1537.970 855.720 1540.350 859.850 ;
        RECT 1541.190 855.720 1543.570 859.850 ;
        RECT 1544.410 855.720 1546.790 859.850 ;
        RECT 1547.630 855.720 1550.010 859.850 ;
        RECT 1550.850 855.720 1553.230 859.850 ;
        RECT 1554.070 855.720 1556.450 859.850 ;
        RECT 1557.290 855.720 1560.130 859.850 ;
        RECT 1560.970 855.720 1563.350 859.850 ;
        RECT 1564.190 855.720 1566.570 859.850 ;
        RECT 1567.410 855.720 1569.790 859.850 ;
        RECT 1570.630 855.720 1573.010 859.850 ;
        RECT 1573.850 855.720 1576.230 859.850 ;
        RECT 1577.070 855.720 1579.450 859.850 ;
        RECT 1580.290 855.720 1582.670 859.850 ;
        RECT 1583.510 855.720 1585.890 859.850 ;
        RECT 1586.730 855.720 1589.110 859.850 ;
        RECT 1589.950 855.720 1592.330 859.850 ;
        RECT 1593.170 855.720 1595.550 859.850 ;
        RECT 1596.390 855.720 1598.770 859.850 ;
        RECT 1599.610 855.720 1601.990 859.850 ;
        RECT 1602.830 855.720 1605.210 859.850 ;
        RECT 1606.050 855.720 1608.430 859.850 ;
        RECT 1609.270 855.720 1611.650 859.850 ;
        RECT 1612.490 855.720 1615.330 859.850 ;
        RECT 1616.170 855.720 1618.550 859.850 ;
        RECT 1619.390 855.720 1621.770 859.850 ;
        RECT 1622.610 855.720 1624.990 859.850 ;
        RECT 1625.830 855.720 1628.210 859.850 ;
        RECT 1629.050 855.720 1631.430 859.850 ;
        RECT 1632.270 855.720 1634.650 859.850 ;
        RECT 1635.490 855.720 1637.870 859.850 ;
        RECT 1638.710 855.720 1641.090 859.850 ;
        RECT 1641.930 855.720 1644.310 859.850 ;
        RECT 1645.150 855.720 1647.530 859.850 ;
        RECT 1648.370 855.720 1650.750 859.850 ;
        RECT 1651.590 855.720 1653.970 859.850 ;
        RECT 1654.810 855.720 1657.190 859.850 ;
        RECT 1658.030 855.720 1660.410 859.850 ;
        RECT 1661.250 855.720 1663.630 859.850 ;
        RECT 1664.470 855.720 1666.850 859.850 ;
        RECT 1667.690 855.720 1670.530 859.850 ;
        RECT 1671.370 855.720 1673.750 859.850 ;
        RECT 1674.590 855.720 1676.970 859.850 ;
        RECT 1677.810 855.720 1680.190 859.850 ;
        RECT 1681.030 855.720 1683.410 859.850 ;
        RECT 1684.250 855.720 1686.630 859.850 ;
        RECT 1687.470 855.720 1689.850 859.850 ;
        RECT 1690.690 855.720 1693.070 859.850 ;
        RECT 1693.910 855.720 1696.290 859.850 ;
        RECT 1697.130 855.720 1699.510 859.850 ;
        RECT 1700.350 855.720 1702.730 859.850 ;
        RECT 1703.570 855.720 1705.950 859.850 ;
        RECT 1706.790 855.720 1709.170 859.850 ;
        RECT 1710.010 855.720 1712.390 859.850 ;
        RECT 1713.230 855.720 1715.610 859.850 ;
        RECT 1716.450 855.720 1718.830 859.850 ;
        RECT 1719.670 855.720 1722.510 859.850 ;
        RECT 1723.350 855.720 1725.730 859.850 ;
        RECT 1726.570 855.720 1728.950 859.850 ;
        RECT 1729.790 855.720 1732.170 859.850 ;
        RECT 1733.010 855.720 1735.390 859.850 ;
        RECT 1736.230 855.720 1738.610 859.850 ;
        RECT 1739.450 855.720 1741.830 859.850 ;
        RECT 1742.670 855.720 1745.050 859.850 ;
        RECT 1745.890 855.720 1748.270 859.850 ;
        RECT 1749.110 855.720 1751.490 859.850 ;
        RECT 1752.330 855.720 1754.710 859.850 ;
        RECT 1755.550 855.720 1757.930 859.850 ;
        RECT 1758.770 855.720 1761.150 859.850 ;
        RECT 1761.990 855.720 1764.370 859.850 ;
        RECT 1765.210 855.720 1767.590 859.850 ;
        RECT 1768.430 855.720 1770.810 859.850 ;
        RECT 1771.650 855.720 1774.030 859.850 ;
        RECT 1774.870 855.720 1777.710 859.850 ;
        RECT 1778.550 855.720 1780.930 859.850 ;
        RECT 1781.770 855.720 1784.150 859.850 ;
        RECT 1784.990 855.720 1787.370 859.850 ;
        RECT 1788.210 855.720 1790.590 859.850 ;
        RECT 1791.430 855.720 1793.810 859.850 ;
        RECT 1794.650 855.720 1797.030 859.850 ;
        RECT 1797.870 855.720 1800.250 859.850 ;
        RECT 1801.090 855.720 1803.470 859.850 ;
        RECT 1804.310 855.720 1806.690 859.850 ;
        RECT 1807.530 855.720 1809.910 859.850 ;
        RECT 1810.750 855.720 1813.130 859.850 ;
        RECT 1813.970 855.720 1816.350 859.850 ;
        RECT 1817.190 855.720 1819.570 859.850 ;
        RECT 1820.410 855.720 1822.790 859.850 ;
        RECT 1823.630 855.720 1826.010 859.850 ;
        RECT 1826.850 855.720 1829.690 859.850 ;
        RECT 1830.530 855.720 1832.910 859.850 ;
        RECT 1833.750 855.720 1836.130 859.850 ;
        RECT 1836.970 855.720 1839.350 859.850 ;
        RECT 1840.190 855.720 1842.570 859.850 ;
        RECT 1843.410 855.720 1845.790 859.850 ;
        RECT 1846.630 855.720 1849.010 859.850 ;
        RECT 1849.850 855.720 1852.230 859.850 ;
        RECT 1853.070 855.720 1855.450 859.850 ;
        RECT 1856.290 855.720 1858.670 859.850 ;
        RECT 1859.510 855.720 1861.890 859.850 ;
        RECT 1862.730 855.720 1865.110 859.850 ;
        RECT 1865.950 855.720 1868.330 859.850 ;
        RECT 1869.170 855.720 1871.550 859.850 ;
        RECT 1872.390 855.720 1874.770 859.850 ;
        RECT 1875.610 855.720 1877.990 859.850 ;
        RECT 1878.830 855.720 1881.210 859.850 ;
        RECT 1882.050 855.720 1884.890 859.850 ;
        RECT 1885.730 855.720 1888.110 859.850 ;
        RECT 1888.950 855.720 1891.330 859.850 ;
        RECT 1892.170 855.720 1894.550 859.850 ;
        RECT 1895.390 855.720 1897.770 859.850 ;
        RECT 1898.610 855.720 1900.990 859.850 ;
        RECT 1901.830 855.720 1904.210 859.850 ;
        RECT 1905.050 855.720 1907.430 859.850 ;
        RECT 1908.270 855.720 1910.650 859.850 ;
        RECT 1911.490 855.720 1913.870 859.850 ;
        RECT 1914.710 855.720 1917.090 859.850 ;
        RECT 1917.930 855.720 1920.310 859.850 ;
        RECT 1921.150 855.720 1923.530 859.850 ;
        RECT 1924.370 855.720 1926.750 859.850 ;
        RECT 1927.590 855.720 1929.970 859.850 ;
        RECT 1930.810 855.720 1933.190 859.850 ;
        RECT 1934.030 855.720 1936.870 859.850 ;
        RECT 1937.710 855.720 1940.090 859.850 ;
        RECT 1940.930 855.720 1943.310 859.850 ;
        RECT 1944.150 855.720 1946.530 859.850 ;
        RECT 1947.370 855.720 1949.750 859.850 ;
        RECT 1950.590 855.720 1952.970 859.850 ;
        RECT 1953.810 855.720 1956.190 859.850 ;
        RECT 1957.030 855.720 1959.410 859.850 ;
        RECT 1960.250 855.720 1962.630 859.850 ;
        RECT 1963.470 855.720 1965.850 859.850 ;
        RECT 1966.690 855.720 1969.070 859.850 ;
        RECT 1969.910 855.720 1972.290 859.850 ;
        RECT 1973.130 855.720 1975.510 859.850 ;
        RECT 1976.350 855.720 1978.730 859.850 ;
        RECT 1979.570 855.720 1981.950 859.850 ;
        RECT 1982.790 855.720 1985.170 859.850 ;
        RECT 1986.010 855.720 1988.390 859.850 ;
        RECT 1989.230 855.720 1992.070 859.850 ;
        RECT 1992.910 855.720 1995.290 859.850 ;
        RECT 1996.130 855.720 1998.510 859.850 ;
        RECT 1999.350 855.720 2001.730 859.850 ;
        RECT 2002.570 855.720 2004.950 859.850 ;
        RECT 2005.790 855.720 2008.170 859.850 ;
        RECT 2009.010 855.720 2011.390 859.850 ;
        RECT 2012.230 855.720 2014.610 859.850 ;
        RECT 2015.450 855.720 2017.830 859.850 ;
        RECT 2018.670 855.720 2021.050 859.850 ;
        RECT 2021.890 855.720 2024.270 859.850 ;
        RECT 2025.110 855.720 2027.490 859.850 ;
        RECT 2028.330 855.720 2030.710 859.850 ;
        RECT 2031.550 855.720 2033.930 859.850 ;
        RECT 2034.770 855.720 2037.150 859.850 ;
        RECT 2037.990 855.720 2040.370 859.850 ;
        RECT 2041.210 855.720 2044.050 859.850 ;
        RECT 2044.890 855.720 2047.270 859.850 ;
        RECT 2048.110 855.720 2050.490 859.850 ;
        RECT 2051.330 855.720 2053.710 859.850 ;
        RECT 2054.550 855.720 2056.930 859.850 ;
        RECT 2057.770 855.720 2060.150 859.850 ;
        RECT 2060.990 855.720 2063.370 859.850 ;
        RECT 2064.210 855.720 2066.590 859.850 ;
        RECT 2067.430 855.720 2069.810 859.850 ;
        RECT 2070.650 855.720 2073.030 859.850 ;
        RECT 2073.870 855.720 2076.250 859.850 ;
        RECT 2077.090 855.720 2079.470 859.850 ;
        RECT 2080.310 855.720 2082.690 859.850 ;
        RECT 2083.530 855.720 2085.910 859.850 ;
        RECT 2086.750 855.720 2089.130 859.850 ;
        RECT 2089.970 855.720 2092.350 859.850 ;
        RECT 2093.190 855.720 2095.570 859.850 ;
        RECT 2096.410 855.720 2099.250 859.850 ;
        RECT 2100.090 855.720 2102.470 859.850 ;
        RECT 2103.310 855.720 2105.690 859.850 ;
        RECT 2106.530 855.720 2108.910 859.850 ;
        RECT 2109.750 855.720 2112.130 859.850 ;
        RECT 2112.970 855.720 2115.350 859.850 ;
        RECT 2116.190 855.720 2118.570 859.850 ;
        RECT 2119.410 855.720 2121.790 859.850 ;
        RECT 2122.630 855.720 2125.010 859.850 ;
        RECT 2125.850 855.720 2128.230 859.850 ;
        RECT 2129.070 855.720 2131.450 859.850 ;
        RECT 2132.290 855.720 2134.670 859.850 ;
        RECT 2135.510 855.720 2137.890 859.850 ;
        RECT 2138.730 855.720 2141.110 859.850 ;
        RECT 2141.950 855.720 2144.330 859.850 ;
        RECT 2145.170 855.720 2147.550 859.850 ;
        RECT 1.480 4.280 2148.100 855.720 ;
        RECT 1.480 2.195 48.570 4.280 ;
        RECT 49.410 2.195 146.090 4.280 ;
        RECT 146.930 2.195 243.610 4.280 ;
        RECT 244.450 2.195 341.590 4.280 ;
        RECT 342.430 2.195 439.110 4.280 ;
        RECT 439.950 2.195 537.090 4.280 ;
        RECT 537.930 2.195 634.610 4.280 ;
        RECT 635.450 2.195 732.590 4.280 ;
        RECT 733.430 2.195 830.110 4.280 ;
        RECT 830.950 2.195 928.090 4.280 ;
        RECT 928.930 2.195 1025.610 4.280 ;
        RECT 1026.450 2.195 1123.590 4.280 ;
        RECT 1124.430 2.195 1221.110 4.280 ;
        RECT 1221.950 2.195 1318.630 4.280 ;
        RECT 1319.470 2.195 1416.610 4.280 ;
        RECT 1417.450 2.195 1514.130 4.280 ;
        RECT 1514.970 2.195 1612.110 4.280 ;
        RECT 1612.950 2.195 1709.630 4.280 ;
        RECT 1710.470 2.195 1807.610 4.280 ;
        RECT 1808.450 2.195 1905.130 4.280 ;
        RECT 1905.970 2.195 2003.110 4.280 ;
        RECT 2003.950 2.195 2100.630 4.280 ;
        RECT 2101.470 2.195 2148.100 4.280 ;
      LAYER met3 ;
        RECT 4.400 856.440 2146.000 857.305 ;
        RECT 4.000 855.800 2146.000 856.440 ;
        RECT 4.000 854.400 2145.600 855.800 ;
        RECT 4.000 852.400 2146.000 854.400 ;
        RECT 4.400 851.000 2146.000 852.400 ;
        RECT 4.000 846.960 2146.000 851.000 ;
        RECT 4.400 846.280 2146.000 846.960 ;
        RECT 4.400 845.560 2145.600 846.280 ;
        RECT 4.000 844.880 2145.600 845.560 ;
        RECT 4.000 841.520 2146.000 844.880 ;
        RECT 4.400 840.120 2146.000 841.520 ;
        RECT 4.000 836.760 2146.000 840.120 ;
        RECT 4.000 836.080 2145.600 836.760 ;
        RECT 4.400 835.360 2145.600 836.080 ;
        RECT 4.400 834.680 2146.000 835.360 ;
        RECT 4.000 830.640 2146.000 834.680 ;
        RECT 4.400 829.240 2146.000 830.640 ;
        RECT 4.000 827.240 2146.000 829.240 ;
        RECT 4.000 825.840 2145.600 827.240 ;
        RECT 4.000 825.200 2146.000 825.840 ;
        RECT 4.400 823.800 2146.000 825.200 ;
        RECT 4.000 819.760 2146.000 823.800 ;
        RECT 4.400 818.360 2146.000 819.760 ;
        RECT 4.000 817.040 2146.000 818.360 ;
        RECT 4.000 815.640 2145.600 817.040 ;
        RECT 4.000 814.320 2146.000 815.640 ;
        RECT 4.400 812.920 2146.000 814.320 ;
        RECT 4.000 808.880 2146.000 812.920 ;
        RECT 4.400 807.520 2146.000 808.880 ;
        RECT 4.400 807.480 2145.600 807.520 ;
        RECT 4.000 806.120 2145.600 807.480 ;
        RECT 4.000 804.120 2146.000 806.120 ;
        RECT 4.400 802.720 2146.000 804.120 ;
        RECT 4.000 798.680 2146.000 802.720 ;
        RECT 4.400 798.000 2146.000 798.680 ;
        RECT 4.400 797.280 2145.600 798.000 ;
        RECT 4.000 796.600 2145.600 797.280 ;
        RECT 4.000 793.240 2146.000 796.600 ;
        RECT 4.400 791.840 2146.000 793.240 ;
        RECT 4.000 788.480 2146.000 791.840 ;
        RECT 4.000 787.800 2145.600 788.480 ;
        RECT 4.400 787.080 2145.600 787.800 ;
        RECT 4.400 786.400 2146.000 787.080 ;
        RECT 4.000 782.360 2146.000 786.400 ;
        RECT 4.400 780.960 2146.000 782.360 ;
        RECT 4.000 778.960 2146.000 780.960 ;
        RECT 4.000 777.560 2145.600 778.960 ;
        RECT 4.000 776.920 2146.000 777.560 ;
        RECT 4.400 775.520 2146.000 776.920 ;
        RECT 4.000 771.480 2146.000 775.520 ;
        RECT 4.400 770.080 2146.000 771.480 ;
        RECT 4.000 768.760 2146.000 770.080 ;
        RECT 4.000 767.360 2145.600 768.760 ;
        RECT 4.000 766.040 2146.000 767.360 ;
        RECT 4.400 764.640 2146.000 766.040 ;
        RECT 4.000 760.600 2146.000 764.640 ;
        RECT 4.400 759.240 2146.000 760.600 ;
        RECT 4.400 759.200 2145.600 759.240 ;
        RECT 4.000 757.840 2145.600 759.200 ;
        RECT 4.000 755.160 2146.000 757.840 ;
        RECT 4.400 753.760 2146.000 755.160 ;
        RECT 4.000 749.720 2146.000 753.760 ;
        RECT 4.400 748.320 2145.600 749.720 ;
        RECT 4.000 744.960 2146.000 748.320 ;
        RECT 4.400 743.560 2146.000 744.960 ;
        RECT 4.000 740.200 2146.000 743.560 ;
        RECT 4.000 739.520 2145.600 740.200 ;
        RECT 4.400 738.800 2145.600 739.520 ;
        RECT 4.400 738.120 2146.000 738.800 ;
        RECT 4.000 734.080 2146.000 738.120 ;
        RECT 4.400 732.680 2146.000 734.080 ;
        RECT 4.000 730.680 2146.000 732.680 ;
        RECT 4.000 729.280 2145.600 730.680 ;
        RECT 4.000 728.640 2146.000 729.280 ;
        RECT 4.400 727.240 2146.000 728.640 ;
        RECT 4.000 723.200 2146.000 727.240 ;
        RECT 4.400 721.800 2146.000 723.200 ;
        RECT 4.000 720.480 2146.000 721.800 ;
        RECT 4.000 719.080 2145.600 720.480 ;
        RECT 4.000 717.760 2146.000 719.080 ;
        RECT 4.400 716.360 2146.000 717.760 ;
        RECT 4.000 712.320 2146.000 716.360 ;
        RECT 4.400 710.960 2146.000 712.320 ;
        RECT 4.400 710.920 2145.600 710.960 ;
        RECT 4.000 709.560 2145.600 710.920 ;
        RECT 4.000 706.880 2146.000 709.560 ;
        RECT 4.400 705.480 2146.000 706.880 ;
        RECT 4.000 701.440 2146.000 705.480 ;
        RECT 4.400 700.040 2145.600 701.440 ;
        RECT 4.000 696.000 2146.000 700.040 ;
        RECT 4.400 694.600 2146.000 696.000 ;
        RECT 4.000 691.920 2146.000 694.600 ;
        RECT 4.000 691.240 2145.600 691.920 ;
        RECT 4.400 690.520 2145.600 691.240 ;
        RECT 4.400 689.840 2146.000 690.520 ;
        RECT 4.000 685.800 2146.000 689.840 ;
        RECT 4.400 684.400 2146.000 685.800 ;
        RECT 4.000 681.720 2146.000 684.400 ;
        RECT 4.000 680.360 2145.600 681.720 ;
        RECT 4.400 680.320 2145.600 680.360 ;
        RECT 4.400 678.960 2146.000 680.320 ;
        RECT 4.000 674.920 2146.000 678.960 ;
        RECT 4.400 673.520 2146.000 674.920 ;
        RECT 4.000 672.200 2146.000 673.520 ;
        RECT 4.000 670.800 2145.600 672.200 ;
        RECT 4.000 669.480 2146.000 670.800 ;
        RECT 4.400 668.080 2146.000 669.480 ;
        RECT 4.000 664.040 2146.000 668.080 ;
        RECT 4.400 662.680 2146.000 664.040 ;
        RECT 4.400 662.640 2145.600 662.680 ;
        RECT 4.000 661.280 2145.600 662.640 ;
        RECT 4.000 658.600 2146.000 661.280 ;
        RECT 4.400 657.200 2146.000 658.600 ;
        RECT 4.000 653.160 2146.000 657.200 ;
        RECT 4.400 651.760 2145.600 653.160 ;
        RECT 4.000 647.720 2146.000 651.760 ;
        RECT 4.400 646.320 2146.000 647.720 ;
        RECT 4.000 643.640 2146.000 646.320 ;
        RECT 4.000 642.280 2145.600 643.640 ;
        RECT 4.400 642.240 2145.600 642.280 ;
        RECT 4.400 640.880 2146.000 642.240 ;
        RECT 4.000 636.840 2146.000 640.880 ;
        RECT 4.400 635.440 2146.000 636.840 ;
        RECT 4.000 633.440 2146.000 635.440 ;
        RECT 4.000 632.080 2145.600 633.440 ;
        RECT 4.400 632.040 2145.600 632.080 ;
        RECT 4.400 630.680 2146.000 632.040 ;
        RECT 4.000 626.640 2146.000 630.680 ;
        RECT 4.400 625.240 2146.000 626.640 ;
        RECT 4.000 623.920 2146.000 625.240 ;
        RECT 4.000 622.520 2145.600 623.920 ;
        RECT 4.000 621.200 2146.000 622.520 ;
        RECT 4.400 619.800 2146.000 621.200 ;
        RECT 4.000 615.760 2146.000 619.800 ;
        RECT 4.400 614.400 2146.000 615.760 ;
        RECT 4.400 614.360 2145.600 614.400 ;
        RECT 4.000 613.000 2145.600 614.360 ;
        RECT 4.000 610.320 2146.000 613.000 ;
        RECT 4.400 608.920 2146.000 610.320 ;
        RECT 4.000 604.880 2146.000 608.920 ;
        RECT 4.400 603.480 2145.600 604.880 ;
        RECT 4.000 599.440 2146.000 603.480 ;
        RECT 4.400 598.040 2146.000 599.440 ;
        RECT 4.000 595.360 2146.000 598.040 ;
        RECT 4.000 594.000 2145.600 595.360 ;
        RECT 4.400 593.960 2145.600 594.000 ;
        RECT 4.400 592.600 2146.000 593.960 ;
        RECT 4.000 588.560 2146.000 592.600 ;
        RECT 4.400 587.160 2146.000 588.560 ;
        RECT 4.000 585.160 2146.000 587.160 ;
        RECT 4.000 583.760 2145.600 585.160 ;
        RECT 4.000 583.120 2146.000 583.760 ;
        RECT 4.400 581.720 2146.000 583.120 ;
        RECT 4.000 577.680 2146.000 581.720 ;
        RECT 4.400 576.280 2146.000 577.680 ;
        RECT 4.000 575.640 2146.000 576.280 ;
        RECT 4.000 574.240 2145.600 575.640 ;
        RECT 4.000 572.920 2146.000 574.240 ;
        RECT 4.400 571.520 2146.000 572.920 ;
        RECT 4.000 567.480 2146.000 571.520 ;
        RECT 4.400 566.120 2146.000 567.480 ;
        RECT 4.400 566.080 2145.600 566.120 ;
        RECT 4.000 564.720 2145.600 566.080 ;
        RECT 4.000 562.040 2146.000 564.720 ;
        RECT 4.400 560.640 2146.000 562.040 ;
        RECT 4.000 556.600 2146.000 560.640 ;
        RECT 4.400 555.200 2145.600 556.600 ;
        RECT 4.000 551.160 2146.000 555.200 ;
        RECT 4.400 549.760 2146.000 551.160 ;
        RECT 4.000 546.400 2146.000 549.760 ;
        RECT 4.000 545.720 2145.600 546.400 ;
        RECT 4.400 545.000 2145.600 545.720 ;
        RECT 4.400 544.320 2146.000 545.000 ;
        RECT 4.000 540.280 2146.000 544.320 ;
        RECT 4.400 538.880 2146.000 540.280 ;
        RECT 4.000 536.880 2146.000 538.880 ;
        RECT 4.000 535.480 2145.600 536.880 ;
        RECT 4.000 534.840 2146.000 535.480 ;
        RECT 4.400 533.440 2146.000 534.840 ;
        RECT 4.000 529.400 2146.000 533.440 ;
        RECT 4.400 528.000 2146.000 529.400 ;
        RECT 4.000 527.360 2146.000 528.000 ;
        RECT 4.000 525.960 2145.600 527.360 ;
        RECT 4.000 523.960 2146.000 525.960 ;
        RECT 4.400 522.560 2146.000 523.960 ;
        RECT 4.000 519.200 2146.000 522.560 ;
        RECT 4.400 517.840 2146.000 519.200 ;
        RECT 4.400 517.800 2145.600 517.840 ;
        RECT 4.000 516.440 2145.600 517.800 ;
        RECT 4.000 513.760 2146.000 516.440 ;
        RECT 4.400 512.360 2146.000 513.760 ;
        RECT 4.000 508.320 2146.000 512.360 ;
        RECT 4.400 506.920 2145.600 508.320 ;
        RECT 4.000 502.880 2146.000 506.920 ;
        RECT 4.400 501.480 2146.000 502.880 ;
        RECT 4.000 498.120 2146.000 501.480 ;
        RECT 4.000 497.440 2145.600 498.120 ;
        RECT 4.400 496.720 2145.600 497.440 ;
        RECT 4.400 496.040 2146.000 496.720 ;
        RECT 4.000 492.000 2146.000 496.040 ;
        RECT 4.400 490.600 2146.000 492.000 ;
        RECT 4.000 488.600 2146.000 490.600 ;
        RECT 4.000 487.200 2145.600 488.600 ;
        RECT 4.000 486.560 2146.000 487.200 ;
        RECT 4.400 485.160 2146.000 486.560 ;
        RECT 4.000 481.120 2146.000 485.160 ;
        RECT 4.400 479.720 2146.000 481.120 ;
        RECT 4.000 479.080 2146.000 479.720 ;
        RECT 4.000 477.680 2145.600 479.080 ;
        RECT 4.000 475.680 2146.000 477.680 ;
        RECT 4.400 474.280 2146.000 475.680 ;
        RECT 4.000 470.240 2146.000 474.280 ;
        RECT 4.400 469.560 2146.000 470.240 ;
        RECT 4.400 468.840 2145.600 469.560 ;
        RECT 4.000 468.160 2145.600 468.840 ;
        RECT 4.000 464.800 2146.000 468.160 ;
        RECT 4.400 463.400 2146.000 464.800 ;
        RECT 4.000 460.040 2146.000 463.400 ;
        RECT 4.400 458.640 2145.600 460.040 ;
        RECT 4.000 454.600 2146.000 458.640 ;
        RECT 4.400 453.200 2146.000 454.600 ;
        RECT 4.000 449.840 2146.000 453.200 ;
        RECT 4.000 449.160 2145.600 449.840 ;
        RECT 4.400 448.440 2145.600 449.160 ;
        RECT 4.400 447.760 2146.000 448.440 ;
        RECT 4.000 443.720 2146.000 447.760 ;
        RECT 4.400 442.320 2146.000 443.720 ;
        RECT 4.000 440.320 2146.000 442.320 ;
        RECT 4.000 438.920 2145.600 440.320 ;
        RECT 4.000 438.280 2146.000 438.920 ;
        RECT 4.400 436.880 2146.000 438.280 ;
        RECT 4.000 432.840 2146.000 436.880 ;
        RECT 4.400 431.440 2146.000 432.840 ;
        RECT 4.000 430.800 2146.000 431.440 ;
        RECT 4.000 429.400 2145.600 430.800 ;
        RECT 4.000 427.400 2146.000 429.400 ;
        RECT 4.400 426.000 2146.000 427.400 ;
        RECT 4.000 421.960 2146.000 426.000 ;
        RECT 4.400 421.280 2146.000 421.960 ;
        RECT 4.400 420.560 2145.600 421.280 ;
        RECT 4.000 419.880 2145.600 420.560 ;
        RECT 4.000 416.520 2146.000 419.880 ;
        RECT 4.400 415.120 2146.000 416.520 ;
        RECT 4.000 411.080 2146.000 415.120 ;
        RECT 4.400 409.680 2145.600 411.080 ;
        RECT 4.000 405.640 2146.000 409.680 ;
        RECT 4.400 404.240 2146.000 405.640 ;
        RECT 4.000 401.560 2146.000 404.240 ;
        RECT 4.000 400.880 2145.600 401.560 ;
        RECT 4.400 400.160 2145.600 400.880 ;
        RECT 4.400 399.480 2146.000 400.160 ;
        RECT 4.000 395.440 2146.000 399.480 ;
        RECT 4.400 394.040 2146.000 395.440 ;
        RECT 4.000 392.040 2146.000 394.040 ;
        RECT 4.000 390.640 2145.600 392.040 ;
        RECT 4.000 390.000 2146.000 390.640 ;
        RECT 4.400 388.600 2146.000 390.000 ;
        RECT 4.000 384.560 2146.000 388.600 ;
        RECT 4.400 383.160 2146.000 384.560 ;
        RECT 4.000 382.520 2146.000 383.160 ;
        RECT 4.000 381.120 2145.600 382.520 ;
        RECT 4.000 379.120 2146.000 381.120 ;
        RECT 4.400 377.720 2146.000 379.120 ;
        RECT 4.000 373.680 2146.000 377.720 ;
        RECT 4.400 373.000 2146.000 373.680 ;
        RECT 4.400 372.280 2145.600 373.000 ;
        RECT 4.000 371.600 2145.600 372.280 ;
        RECT 4.000 368.240 2146.000 371.600 ;
        RECT 4.400 366.840 2146.000 368.240 ;
        RECT 4.000 362.800 2146.000 366.840 ;
        RECT 4.400 361.400 2145.600 362.800 ;
        RECT 4.000 357.360 2146.000 361.400 ;
        RECT 4.400 355.960 2146.000 357.360 ;
        RECT 4.000 353.280 2146.000 355.960 ;
        RECT 4.000 351.920 2145.600 353.280 ;
        RECT 4.400 351.880 2145.600 351.920 ;
        RECT 4.400 350.520 2146.000 351.880 ;
        RECT 4.000 347.160 2146.000 350.520 ;
        RECT 4.400 345.760 2146.000 347.160 ;
        RECT 4.000 343.760 2146.000 345.760 ;
        RECT 4.000 342.360 2145.600 343.760 ;
        RECT 4.000 341.720 2146.000 342.360 ;
        RECT 4.400 340.320 2146.000 341.720 ;
        RECT 4.000 336.280 2146.000 340.320 ;
        RECT 4.400 334.880 2146.000 336.280 ;
        RECT 4.000 334.240 2146.000 334.880 ;
        RECT 4.000 332.840 2145.600 334.240 ;
        RECT 4.000 330.840 2146.000 332.840 ;
        RECT 4.400 329.440 2146.000 330.840 ;
        RECT 4.000 325.400 2146.000 329.440 ;
        RECT 4.400 324.720 2146.000 325.400 ;
        RECT 4.400 324.000 2145.600 324.720 ;
        RECT 4.000 323.320 2145.600 324.000 ;
        RECT 4.000 319.960 2146.000 323.320 ;
        RECT 4.400 318.560 2146.000 319.960 ;
        RECT 4.000 314.520 2146.000 318.560 ;
        RECT 4.400 313.120 2145.600 314.520 ;
        RECT 4.000 309.080 2146.000 313.120 ;
        RECT 4.400 307.680 2146.000 309.080 ;
        RECT 4.000 305.000 2146.000 307.680 ;
        RECT 4.000 303.640 2145.600 305.000 ;
        RECT 4.400 303.600 2145.600 303.640 ;
        RECT 4.400 302.240 2146.000 303.600 ;
        RECT 4.000 298.200 2146.000 302.240 ;
        RECT 4.400 296.800 2146.000 298.200 ;
        RECT 4.000 295.480 2146.000 296.800 ;
        RECT 4.000 294.080 2145.600 295.480 ;
        RECT 4.000 292.760 2146.000 294.080 ;
        RECT 4.400 291.360 2146.000 292.760 ;
        RECT 4.000 288.000 2146.000 291.360 ;
        RECT 4.400 286.600 2146.000 288.000 ;
        RECT 4.000 285.960 2146.000 286.600 ;
        RECT 4.000 284.560 2145.600 285.960 ;
        RECT 4.000 282.560 2146.000 284.560 ;
        RECT 4.400 281.160 2146.000 282.560 ;
        RECT 4.000 277.120 2146.000 281.160 ;
        RECT 4.400 275.760 2146.000 277.120 ;
        RECT 4.400 275.720 2145.600 275.760 ;
        RECT 4.000 274.360 2145.600 275.720 ;
        RECT 4.000 271.680 2146.000 274.360 ;
        RECT 4.400 270.280 2146.000 271.680 ;
        RECT 4.000 266.240 2146.000 270.280 ;
        RECT 4.400 264.840 2145.600 266.240 ;
        RECT 4.000 260.800 2146.000 264.840 ;
        RECT 4.400 259.400 2146.000 260.800 ;
        RECT 4.000 256.720 2146.000 259.400 ;
        RECT 4.000 255.360 2145.600 256.720 ;
        RECT 4.400 255.320 2145.600 255.360 ;
        RECT 4.400 253.960 2146.000 255.320 ;
        RECT 4.000 249.920 2146.000 253.960 ;
        RECT 4.400 248.520 2146.000 249.920 ;
        RECT 4.000 247.200 2146.000 248.520 ;
        RECT 4.000 245.800 2145.600 247.200 ;
        RECT 4.000 244.480 2146.000 245.800 ;
        RECT 4.400 243.080 2146.000 244.480 ;
        RECT 4.000 239.040 2146.000 243.080 ;
        RECT 4.400 237.680 2146.000 239.040 ;
        RECT 4.400 237.640 2145.600 237.680 ;
        RECT 4.000 236.280 2145.600 237.640 ;
        RECT 4.000 233.600 2146.000 236.280 ;
        RECT 4.400 232.200 2146.000 233.600 ;
        RECT 4.000 228.840 2146.000 232.200 ;
        RECT 4.400 227.480 2146.000 228.840 ;
        RECT 4.400 227.440 2145.600 227.480 ;
        RECT 4.000 226.080 2145.600 227.440 ;
        RECT 4.000 223.400 2146.000 226.080 ;
        RECT 4.400 222.000 2146.000 223.400 ;
        RECT 4.000 217.960 2146.000 222.000 ;
        RECT 4.400 216.560 2145.600 217.960 ;
        RECT 4.000 212.520 2146.000 216.560 ;
        RECT 4.400 211.120 2146.000 212.520 ;
        RECT 4.000 208.440 2146.000 211.120 ;
        RECT 4.000 207.080 2145.600 208.440 ;
        RECT 4.400 207.040 2145.600 207.080 ;
        RECT 4.400 205.680 2146.000 207.040 ;
        RECT 4.000 201.640 2146.000 205.680 ;
        RECT 4.400 200.240 2146.000 201.640 ;
        RECT 4.000 198.920 2146.000 200.240 ;
        RECT 4.000 197.520 2145.600 198.920 ;
        RECT 4.000 196.200 2146.000 197.520 ;
        RECT 4.400 194.800 2146.000 196.200 ;
        RECT 4.000 190.760 2146.000 194.800 ;
        RECT 4.400 189.400 2146.000 190.760 ;
        RECT 4.400 189.360 2145.600 189.400 ;
        RECT 4.000 188.000 2145.600 189.360 ;
        RECT 4.000 185.320 2146.000 188.000 ;
        RECT 4.400 183.920 2146.000 185.320 ;
        RECT 4.000 179.880 2146.000 183.920 ;
        RECT 4.400 179.200 2146.000 179.880 ;
        RECT 4.400 178.480 2145.600 179.200 ;
        RECT 4.000 177.800 2145.600 178.480 ;
        RECT 4.000 175.120 2146.000 177.800 ;
        RECT 4.400 173.720 2146.000 175.120 ;
        RECT 4.000 169.680 2146.000 173.720 ;
        RECT 4.400 168.280 2145.600 169.680 ;
        RECT 4.000 164.240 2146.000 168.280 ;
        RECT 4.400 162.840 2146.000 164.240 ;
        RECT 4.000 160.160 2146.000 162.840 ;
        RECT 4.000 158.800 2145.600 160.160 ;
        RECT 4.400 158.760 2145.600 158.800 ;
        RECT 4.400 157.400 2146.000 158.760 ;
        RECT 4.000 153.360 2146.000 157.400 ;
        RECT 4.400 151.960 2146.000 153.360 ;
        RECT 4.000 150.640 2146.000 151.960 ;
        RECT 4.000 149.240 2145.600 150.640 ;
        RECT 4.000 147.920 2146.000 149.240 ;
        RECT 4.400 146.520 2146.000 147.920 ;
        RECT 4.000 142.480 2146.000 146.520 ;
        RECT 4.400 141.080 2146.000 142.480 ;
        RECT 4.000 140.440 2146.000 141.080 ;
        RECT 4.000 139.040 2145.600 140.440 ;
        RECT 4.000 137.040 2146.000 139.040 ;
        RECT 4.400 135.640 2146.000 137.040 ;
        RECT 4.000 131.600 2146.000 135.640 ;
        RECT 4.400 130.920 2146.000 131.600 ;
        RECT 4.400 130.200 2145.600 130.920 ;
        RECT 4.000 129.520 2145.600 130.200 ;
        RECT 4.000 126.160 2146.000 129.520 ;
        RECT 4.400 124.760 2146.000 126.160 ;
        RECT 4.000 121.400 2146.000 124.760 ;
        RECT 4.000 120.720 2145.600 121.400 ;
        RECT 4.400 120.000 2145.600 120.720 ;
        RECT 4.400 119.320 2146.000 120.000 ;
        RECT 4.000 115.960 2146.000 119.320 ;
        RECT 4.400 114.560 2146.000 115.960 ;
        RECT 4.000 111.880 2146.000 114.560 ;
        RECT 4.000 110.520 2145.600 111.880 ;
        RECT 4.400 110.480 2145.600 110.520 ;
        RECT 4.400 109.120 2146.000 110.480 ;
        RECT 4.000 105.080 2146.000 109.120 ;
        RECT 4.400 103.680 2146.000 105.080 ;
        RECT 4.000 102.360 2146.000 103.680 ;
        RECT 4.000 100.960 2145.600 102.360 ;
        RECT 4.000 99.640 2146.000 100.960 ;
        RECT 4.400 98.240 2146.000 99.640 ;
        RECT 4.000 94.200 2146.000 98.240 ;
        RECT 4.400 92.800 2146.000 94.200 ;
        RECT 4.000 92.160 2146.000 92.800 ;
        RECT 4.000 90.760 2145.600 92.160 ;
        RECT 4.000 88.760 2146.000 90.760 ;
        RECT 4.400 87.360 2146.000 88.760 ;
        RECT 4.000 83.320 2146.000 87.360 ;
        RECT 4.400 82.640 2146.000 83.320 ;
        RECT 4.400 81.920 2145.600 82.640 ;
        RECT 4.000 81.240 2145.600 81.920 ;
        RECT 4.000 77.880 2146.000 81.240 ;
        RECT 4.400 76.480 2146.000 77.880 ;
        RECT 4.000 73.120 2146.000 76.480 ;
        RECT 4.000 72.440 2145.600 73.120 ;
        RECT 4.400 71.720 2145.600 72.440 ;
        RECT 4.400 71.040 2146.000 71.720 ;
        RECT 4.000 67.000 2146.000 71.040 ;
        RECT 4.400 65.600 2146.000 67.000 ;
        RECT 4.000 63.600 2146.000 65.600 ;
        RECT 4.000 62.200 2145.600 63.600 ;
        RECT 4.000 61.560 2146.000 62.200 ;
        RECT 4.400 60.160 2146.000 61.560 ;
        RECT 4.000 56.800 2146.000 60.160 ;
        RECT 4.400 55.400 2146.000 56.800 ;
        RECT 4.000 54.080 2146.000 55.400 ;
        RECT 4.000 52.680 2145.600 54.080 ;
        RECT 4.000 51.360 2146.000 52.680 ;
        RECT 4.400 49.960 2146.000 51.360 ;
        RECT 4.000 45.920 2146.000 49.960 ;
        RECT 4.400 44.520 2146.000 45.920 ;
        RECT 4.000 43.880 2146.000 44.520 ;
        RECT 4.000 42.480 2145.600 43.880 ;
        RECT 4.000 40.480 2146.000 42.480 ;
        RECT 4.400 39.080 2146.000 40.480 ;
        RECT 4.000 35.040 2146.000 39.080 ;
        RECT 4.400 34.360 2146.000 35.040 ;
        RECT 4.400 33.640 2145.600 34.360 ;
        RECT 4.000 32.960 2145.600 33.640 ;
        RECT 4.000 29.600 2146.000 32.960 ;
        RECT 4.400 28.200 2146.000 29.600 ;
        RECT 4.000 24.840 2146.000 28.200 ;
        RECT 4.000 24.160 2145.600 24.840 ;
        RECT 4.400 23.440 2145.600 24.160 ;
        RECT 4.400 22.760 2146.000 23.440 ;
        RECT 4.000 18.720 2146.000 22.760 ;
        RECT 4.400 17.320 2146.000 18.720 ;
        RECT 4.000 15.320 2146.000 17.320 ;
        RECT 4.000 13.920 2145.600 15.320 ;
        RECT 4.000 13.280 2146.000 13.920 ;
        RECT 4.400 11.880 2146.000 13.280 ;
        RECT 4.000 7.840 2146.000 11.880 ;
        RECT 4.400 6.440 2146.000 7.840 ;
        RECT 4.000 5.800 2146.000 6.440 ;
        RECT 4.000 4.400 2145.600 5.800 ;
        RECT 4.000 3.080 2146.000 4.400 ;
        RECT 4.400 2.215 2146.000 3.080 ;
      LAYER met4 ;
        RECT 8.575 849.280 2132.265 855.945 ;
        RECT 8.575 11.735 20.640 849.280 ;
        RECT 23.040 11.735 45.640 849.280 ;
        RECT 48.040 11.735 70.640 849.280 ;
        RECT 73.040 11.735 95.640 849.280 ;
        RECT 98.040 640.360 120.640 849.280 ;
        RECT 123.040 640.360 145.640 849.280 ;
        RECT 148.040 640.360 170.640 849.280 ;
        RECT 173.040 640.360 195.640 849.280 ;
        RECT 198.040 640.360 220.640 849.280 ;
        RECT 223.040 640.360 245.640 849.280 ;
        RECT 248.040 640.360 270.640 849.280 ;
        RECT 273.040 640.360 295.640 849.280 ;
        RECT 298.040 640.360 320.640 849.280 ;
        RECT 323.040 640.360 345.640 849.280 ;
        RECT 348.040 640.360 370.640 849.280 ;
        RECT 373.040 640.360 395.640 849.280 ;
        RECT 398.040 640.360 420.640 849.280 ;
        RECT 423.040 640.360 445.640 849.280 ;
        RECT 448.040 640.360 470.640 849.280 ;
        RECT 473.040 640.360 495.640 849.280 ;
        RECT 498.040 640.360 520.640 849.280 ;
        RECT 523.040 640.360 545.640 849.280 ;
        RECT 548.040 640.360 570.640 849.280 ;
        RECT 573.040 640.360 595.640 849.280 ;
        RECT 598.040 640.360 620.640 849.280 ;
        RECT 623.040 640.360 645.640 849.280 ;
        RECT 648.040 640.360 670.640 849.280 ;
        RECT 673.040 640.360 695.640 849.280 ;
        RECT 698.040 640.360 720.640 849.280 ;
        RECT 723.040 640.360 745.640 849.280 ;
        RECT 748.040 640.360 770.640 849.280 ;
        RECT 773.040 640.360 795.640 849.280 ;
        RECT 798.040 640.360 820.640 849.280 ;
        RECT 823.040 640.360 845.640 849.280 ;
        RECT 848.040 640.360 870.640 849.280 ;
        RECT 873.040 640.360 895.640 849.280 ;
        RECT 98.040 106.640 895.640 640.360 ;
        RECT 98.040 11.735 120.640 106.640 ;
        RECT 123.040 11.735 145.640 106.640 ;
        RECT 148.040 11.735 170.640 106.640 ;
        RECT 173.040 11.735 195.640 106.640 ;
        RECT 198.040 11.735 220.640 106.640 ;
        RECT 223.040 11.735 245.640 106.640 ;
        RECT 248.040 11.735 270.640 106.640 ;
        RECT 273.040 11.735 295.640 106.640 ;
        RECT 298.040 11.735 320.640 106.640 ;
        RECT 323.040 11.735 345.640 106.640 ;
        RECT 348.040 11.735 370.640 106.640 ;
        RECT 373.040 11.735 395.640 106.640 ;
        RECT 398.040 11.735 420.640 106.640 ;
        RECT 423.040 11.735 445.640 106.640 ;
        RECT 448.040 11.735 470.640 106.640 ;
        RECT 473.040 11.735 495.640 106.640 ;
        RECT 498.040 11.735 520.640 106.640 ;
        RECT 523.040 11.735 545.640 106.640 ;
        RECT 548.040 11.735 570.640 106.640 ;
        RECT 573.040 11.735 595.640 106.640 ;
        RECT 598.040 11.735 620.640 106.640 ;
        RECT 623.040 11.735 645.640 106.640 ;
        RECT 648.040 11.735 670.640 106.640 ;
        RECT 673.040 11.735 695.640 106.640 ;
        RECT 698.040 11.735 720.640 106.640 ;
        RECT 723.040 11.735 745.640 106.640 ;
        RECT 748.040 11.735 770.640 106.640 ;
        RECT 773.040 11.735 795.640 106.640 ;
        RECT 798.040 11.735 820.640 106.640 ;
        RECT 823.040 11.735 845.640 106.640 ;
        RECT 848.040 11.735 870.640 106.640 ;
        RECT 873.040 11.735 895.640 106.640 ;
        RECT 898.040 11.735 920.640 849.280 ;
        RECT 923.040 11.735 945.640 849.280 ;
        RECT 948.040 11.735 970.640 849.280 ;
        RECT 973.040 11.735 995.640 849.280 ;
        RECT 998.040 11.735 1020.640 849.280 ;
        RECT 1023.040 11.735 1045.640 849.280 ;
        RECT 1048.040 11.735 1070.640 849.280 ;
        RECT 1073.040 11.735 1095.640 849.280 ;
        RECT 1098.040 11.735 1120.640 849.280 ;
        RECT 1123.040 11.735 1145.640 849.280 ;
        RECT 1148.040 11.735 1170.640 849.280 ;
        RECT 1173.040 11.735 1195.640 849.280 ;
        RECT 1198.040 11.735 1220.640 849.280 ;
        RECT 1223.040 11.735 1245.640 849.280 ;
        RECT 1248.040 11.735 1270.640 849.280 ;
        RECT 1273.040 11.735 1295.640 849.280 ;
        RECT 1298.040 11.735 1320.640 849.280 ;
        RECT 1323.040 11.735 1345.640 849.280 ;
        RECT 1348.040 11.735 1370.640 849.280 ;
        RECT 1373.040 11.735 1395.640 849.280 ;
        RECT 1398.040 11.735 1420.640 849.280 ;
        RECT 1423.040 11.735 1445.640 849.280 ;
        RECT 1448.040 11.735 1470.640 849.280 ;
        RECT 1473.040 11.735 1495.640 849.280 ;
        RECT 1498.040 11.735 1520.640 849.280 ;
        RECT 1523.040 11.735 1545.640 849.280 ;
        RECT 1548.040 11.735 1570.640 849.280 ;
        RECT 1573.040 11.735 1595.640 849.280 ;
        RECT 1598.040 11.735 1620.640 849.280 ;
        RECT 1623.040 11.735 1645.640 849.280 ;
        RECT 1648.040 11.735 1670.640 849.280 ;
        RECT 1673.040 11.735 1695.640 849.280 ;
        RECT 1698.040 11.735 1720.640 849.280 ;
        RECT 1723.040 11.735 1745.640 849.280 ;
        RECT 1748.040 11.735 1770.640 849.280 ;
        RECT 1773.040 11.735 1795.640 849.280 ;
        RECT 1798.040 11.735 1820.640 849.280 ;
        RECT 1823.040 11.735 1845.640 849.280 ;
        RECT 1848.040 11.735 1870.640 849.280 ;
        RECT 1873.040 11.735 1895.640 849.280 ;
        RECT 1898.040 11.735 1920.640 849.280 ;
        RECT 1923.040 821.080 1945.640 849.280 ;
        RECT 1948.040 821.080 1970.640 849.280 ;
        RECT 1973.040 821.080 1995.640 849.280 ;
        RECT 1998.040 821.080 2020.640 849.280 ;
        RECT 1923.040 727.360 2020.640 821.080 ;
        RECT 1923.040 11.735 1945.640 727.360 ;
        RECT 1948.040 11.735 1970.640 727.360 ;
        RECT 1973.040 11.735 1995.640 727.360 ;
        RECT 1998.040 11.735 2020.640 727.360 ;
        RECT 2023.040 11.735 2045.640 849.280 ;
        RECT 2048.040 11.735 2070.640 849.280 ;
        RECT 2073.040 11.735 2095.640 849.280 ;
        RECT 2098.040 11.735 2120.640 849.280 ;
        RECT 2123.040 11.735 2132.265 849.280 ;
  END
END mgmt_core
END LIBRARY

