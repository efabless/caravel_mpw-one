* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_bs_flash__special_sonosfet_star__tox_slope_spectre = 0.0
.param sky130_fd_bs_flash__special_sonosfet_star__vth0_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_bs_flash__special_sonosfet_star__tox_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_bs_flash__special_sonosfet_star__vth0_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_bs_flash__special_sonosfet_star d g s b
+ 
.param  l = 1 w = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 mult = 1.0
Msky130_fd_bs_flash__special_sonosfet_star d g s b sky130_fd_bs_flash__special_sonosfet_star__model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs}
.model sky130_fd_bs_flash__special_sonosfet_star__model.0 nmos
+ lmin = 2.15e-007 lmax = 2.25e-007 wmin = 4.45e-007 wmax = 4.55e-7
+ level = 49.0
+ 
+ tnom = 30.0
+ version = 3.2
+ tox = {1.54e-008*sky130_fd_bs_flash__special_sonosfet_star__tox_mult}
+ toxm = 1.54e-8
+ xj = 1.5000001e-7
+ nch = 1.3069232e+17
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {6.69e-009+sky130_fd_bs_flash__special_sonosfet_star__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {0+sky130_fd_bs_flash__special_sonosfet_star__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ mobmod = 1.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 0.0
* Diode Parameters
+ 
+ ldif = 0.0
+ hdif = 0.0
+ rd = 0.0
+ rs = 0.0
+ rsc = 0.0
+ rdc = 0.0
+ 
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.15+sky130_fd_bs_flash__special_sonosfet_star__vth0_diff_0}
+ k1 = 0.83177
+ k2 = {-0.10077+sky130_fd_bs_flash__special_sonosfet_star__k2_diff_0}
+ k3 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ nlx = 0.0
+ w0 = 0.0
+ k3b = 0.0
+ ngate = 1.0e+23
+ vfb = -0.5627875
* Mobility Parameters
+ vsat = {61317+sky130_fd_bs_flash__special_sonosfet_star__vsat_diff_0}
+ ua = -9.6244e-10
+ ub = 7.44e-18
+ uc = 3.8609e-10
+ rdsw = {0+sky130_fd_bs_flash__special_sonosfet_star__rdsw_diff_0}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.017157+sky130_fd_bs_flash__special_sonosfet_star__u0_diff_0}
+ a0 = 1.0328
+ keta = -0.046049
+ a1 = 0.0
+ a2 = 0.99
+ ags = 0.1
+ b0 = 0.0
+ b1 = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20477+sky130_fd_bs_flash__special_sonosfet_star__voff_diff_0}
+ nfactor = {2.691+sky130_fd_bs_flash__special_sonosfet_star__nfactor_diff_0}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.057437
+ etab = 0.0
+ dsub = 0.0
* Rout Parameters
+ pclm = 1.62
+ pdiblc1 = 0.0
+ pdiblc2 = 0.016156456
+ pdiblcb = 0.2775065
+ drout = 0.0
+ pscbe1 = 4.188539e+8
+ pscbe2 = 1.0e-20
+ pvag = 0.2728709
+ delta = 0.0038
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Temperature Effects Parameters
+ kt1 = {-0.088351+sky130_fd_bs_flash__special_sonosfet_star__kt1_diff_0}
+ kt2 = -0.09179784
+ at = 52118.0
+ ute = -0.5472
+ ua1 = 1.3719e-9
+ ub1 = -2.7626e-18
+ uc1 = 1.4668e-11
+ kt1l = 0.0
+ prt = 0.0
* Capacitance Parameters
+ cj = {0.0012651*sky130_fd_bs_flash__special_sonosfet_star__ajunction_mult}
+ mj = 0.3608
+ pb = 0.729
+ cjsw = {7.3442e-011*sky130_fd_bs_flash__special_sonosfet_star__pjunction_mult}
+ mjsw = 0.13
+ pbsw = 0.729
+ cjswg = {7.3442e-011*sky130_fd_bs_flash__special_sonosfet_star__pjunction_mult}
+ mjswg = 0.13
+ pbswg = 0.729
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.0
+ tcjsw = 0.0
+ tcjswg = 0.0
+ js = 0.000375
+ jsw = 6.0e-10
+ nj = 1.3574
+ xti = 0.13
+ cgdo = {3.0674e-010*sky130_fd_bs_flash__special_sonosfet_star__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_bs_flash__special_sonosfet_star__overlap_mult}
+ cgbo = 0.0
+ capmod = 3.0
+ nqsmod = 0.0
+ elm = 5.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_bs_flash__special_sonosfet_star__overlap_mult}
+ cgdl = {5e-011*sky130_fd_bs_flash__special_sonosfet_star__overlap_mult}
+ ckappa = 0.6
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_bs_flash__special_sonosfet_star__dlc_diff+sky130_fd_bs_flash__special_sonosfet_star__dlc_rotweak}
+ dwc = {0+sky130_fd_bs_flash__special_sonosfet_star__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
.ends sky130_fd_bs_flash__special_sonosfet_star
